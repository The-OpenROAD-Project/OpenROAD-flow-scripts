VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_128x32
  FOREIGN fakeram45_128x32 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 78.470 BY 42.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.400 0.070 1.470 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.680 0.070 1.750 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.960 0.070 2.030 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.240 0.070 2.310 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.520 0.070 2.590 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.800 0.070 2.870 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.080 0.070 3.150 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.360 0.070 3.430 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.640 0.070 3.710 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.920 0.070 3.990 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.200 0.070 4.270 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.480 0.070 4.550 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.760 0.070 4.830 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.040 0.070 5.110 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.320 0.070 5.390 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.600 0.070 5.670 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.880 0.070 5.950 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.160 0.070 6.230 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.440 0.070 6.510 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.720 0.070 6.790 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.000 0.070 7.070 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.280 0.070 7.350 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.560 0.070 7.630 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.840 0.070 7.910 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.120 0.070 8.190 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.400 0.070 8.470 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.680 0.070 8.750 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.960 0.070 9.030 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.240 0.070 9.310 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.520 0.070 9.590 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.800 0.070 9.870 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.080 0.070 10.150 ;
    END
  END w_mask_in[31]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.460 0.070 12.530 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.740 0.070 12.810 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.020 0.070 13.090 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.300 0.070 13.370 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.580 0.070 13.650 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.860 0.070 13.930 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.140 0.070 14.210 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.420 0.070 14.490 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.700 0.070 14.770 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.980 0.070 15.050 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.260 0.070 15.330 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.540 0.070 15.610 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.820 0.070 15.890 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.100 0.070 16.170 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.380 0.070 16.450 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.660 0.070 16.730 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.940 0.070 17.010 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.220 0.070 17.290 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.500 0.070 17.570 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.780 0.070 17.850 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.060 0.070 18.130 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.340 0.070 18.410 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.620 0.070 18.690 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.900 0.070 18.970 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.180 0.070 19.250 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.460 0.070 19.530 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.740 0.070 19.810 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.020 0.070 20.090 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.300 0.070 20.370 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.580 0.070 20.650 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.860 0.070 20.930 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.140 0.070 21.210 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.520 0.070 23.590 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.800 0.070 23.870 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.080 0.070 24.150 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.360 0.070 24.430 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.640 0.070 24.710 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.920 0.070 24.990 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.200 0.070 25.270 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.480 0.070 25.550 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.760 0.070 25.830 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.040 0.070 26.110 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.320 0.070 26.390 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.600 0.070 26.670 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.880 0.070 26.950 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.160 0.070 27.230 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.440 0.070 27.510 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.720 0.070 27.790 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.000 0.070 28.070 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.280 0.070 28.350 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.560 0.070 28.630 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.840 0.070 28.910 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.120 0.070 29.190 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.400 0.070 29.470 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.680 0.070 29.750 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.960 0.070 30.030 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.240 0.070 30.310 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.520 0.070 30.590 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.800 0.070 30.870 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.080 0.070 31.150 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.360 0.070 31.430 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.640 0.070 31.710 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.920 0.070 31.990 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.200 0.070 32.270 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.580 0.070 34.650 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.860 0.070 34.930 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.140 0.070 35.210 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.420 0.070 35.490 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.700 0.070 35.770 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.980 0.070 36.050 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.260 0.070 36.330 ;
    END
  END addr_in[6]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.640 0.070 38.710 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.920 0.070 38.990 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.200 0.070 39.270 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 40.600 ;
      RECT 3.500 1.400 3.780 40.600 ;
      RECT 5.740 1.400 6.020 40.600 ;
      RECT 7.980 1.400 8.260 40.600 ;
      RECT 10.220 1.400 10.500 40.600 ;
      RECT 12.460 1.400 12.740 40.600 ;
      RECT 14.700 1.400 14.980 40.600 ;
      RECT 16.940 1.400 17.220 40.600 ;
      RECT 19.180 1.400 19.460 40.600 ;
      RECT 21.420 1.400 21.700 40.600 ;
      RECT 23.660 1.400 23.940 40.600 ;
      RECT 25.900 1.400 26.180 40.600 ;
      RECT 28.140 1.400 28.420 40.600 ;
      RECT 30.380 1.400 30.660 40.600 ;
      RECT 32.620 1.400 32.900 40.600 ;
      RECT 34.860 1.400 35.140 40.600 ;
      RECT 37.100 1.400 37.380 40.600 ;
      RECT 39.340 1.400 39.620 40.600 ;
      RECT 41.580 1.400 41.860 40.600 ;
      RECT 43.820 1.400 44.100 40.600 ;
      RECT 46.060 1.400 46.340 40.600 ;
      RECT 48.300 1.400 48.580 40.600 ;
      RECT 50.540 1.400 50.820 40.600 ;
      RECT 52.780 1.400 53.060 40.600 ;
      RECT 55.020 1.400 55.300 40.600 ;
      RECT 57.260 1.400 57.540 40.600 ;
      RECT 59.500 1.400 59.780 40.600 ;
      RECT 61.740 1.400 62.020 40.600 ;
      RECT 63.980 1.400 64.260 40.600 ;
      RECT 66.220 1.400 66.500 40.600 ;
      RECT 68.460 1.400 68.740 40.600 ;
      RECT 70.700 1.400 70.980 40.600 ;
      RECT 72.940 1.400 73.220 40.600 ;
      RECT 75.180 1.400 75.460 40.600 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 40.600 ;
      RECT 4.620 1.400 4.900 40.600 ;
      RECT 6.860 1.400 7.140 40.600 ;
      RECT 9.100 1.400 9.380 40.600 ;
      RECT 11.340 1.400 11.620 40.600 ;
      RECT 13.580 1.400 13.860 40.600 ;
      RECT 15.820 1.400 16.100 40.600 ;
      RECT 18.060 1.400 18.340 40.600 ;
      RECT 20.300 1.400 20.580 40.600 ;
      RECT 22.540 1.400 22.820 40.600 ;
      RECT 24.780 1.400 25.060 40.600 ;
      RECT 27.020 1.400 27.300 40.600 ;
      RECT 29.260 1.400 29.540 40.600 ;
      RECT 31.500 1.400 31.780 40.600 ;
      RECT 33.740 1.400 34.020 40.600 ;
      RECT 35.980 1.400 36.260 40.600 ;
      RECT 38.220 1.400 38.500 40.600 ;
      RECT 40.460 1.400 40.740 40.600 ;
      RECT 42.700 1.400 42.980 40.600 ;
      RECT 44.940 1.400 45.220 40.600 ;
      RECT 47.180 1.400 47.460 40.600 ;
      RECT 49.420 1.400 49.700 40.600 ;
      RECT 51.660 1.400 51.940 40.600 ;
      RECT 53.900 1.400 54.180 40.600 ;
      RECT 56.140 1.400 56.420 40.600 ;
      RECT 58.380 1.400 58.660 40.600 ;
      RECT 60.620 1.400 60.900 40.600 ;
      RECT 62.860 1.400 63.140 40.600 ;
      RECT 65.100 1.400 65.380 40.600 ;
      RECT 67.340 1.400 67.620 40.600 ;
      RECT 69.580 1.400 69.860 40.600 ;
      RECT 71.820 1.400 72.100 40.600 ;
      RECT 74.060 1.400 74.340 40.600 ;
      RECT 76.300 1.400 76.580 40.600 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 78.470 42.000 ;
    LAYER metal2 ;
    RECT 0 0 78.470 42.000 ;
    LAYER metal3 ;
    RECT 0.070 0 78.470 42.000 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 1.645 ;
    RECT 0 1.715 0.070 1.925 ;
    RECT 0 1.995 0.070 2.205 ;
    RECT 0 2.275 0.070 2.485 ;
    RECT 0 2.555 0.070 2.765 ;
    RECT 0 2.835 0.070 3.045 ;
    RECT 0 3.115 0.070 3.325 ;
    RECT 0 3.395 0.070 3.605 ;
    RECT 0 3.675 0.070 3.885 ;
    RECT 0 3.955 0.070 4.165 ;
    RECT 0 4.235 0.070 4.445 ;
    RECT 0 4.515 0.070 4.725 ;
    RECT 0 4.795 0.070 5.005 ;
    RECT 0 5.075 0.070 5.285 ;
    RECT 0 5.355 0.070 5.565 ;
    RECT 0 5.635 0.070 5.845 ;
    RECT 0 5.915 0.070 6.125 ;
    RECT 0 6.195 0.070 6.405 ;
    RECT 0 6.475 0.070 6.685 ;
    RECT 0 6.755 0.070 6.965 ;
    RECT 0 7.035 0.070 7.245 ;
    RECT 0 7.315 0.070 7.525 ;
    RECT 0 7.595 0.070 7.805 ;
    RECT 0 7.875 0.070 8.085 ;
    RECT 0 8.155 0.070 8.365 ;
    RECT 0 8.435 0.070 8.645 ;
    RECT 0 8.715 0.070 8.925 ;
    RECT 0 8.995 0.070 9.205 ;
    RECT 0 9.275 0.070 9.485 ;
    RECT 0 9.555 0.070 9.765 ;
    RECT 0 9.835 0.070 10.045 ;
    RECT 0 10.115 0.070 12.425 ;
    RECT 0 12.495 0.070 12.705 ;
    RECT 0 12.775 0.070 12.985 ;
    RECT 0 13.055 0.070 13.265 ;
    RECT 0 13.335 0.070 13.545 ;
    RECT 0 13.615 0.070 13.825 ;
    RECT 0 13.895 0.070 14.105 ;
    RECT 0 14.175 0.070 14.385 ;
    RECT 0 14.455 0.070 14.665 ;
    RECT 0 14.735 0.070 14.945 ;
    RECT 0 15.015 0.070 15.225 ;
    RECT 0 15.295 0.070 15.505 ;
    RECT 0 15.575 0.070 15.785 ;
    RECT 0 15.855 0.070 16.065 ;
    RECT 0 16.135 0.070 16.345 ;
    RECT 0 16.415 0.070 16.625 ;
    RECT 0 16.695 0.070 16.905 ;
    RECT 0 16.975 0.070 17.185 ;
    RECT 0 17.255 0.070 17.465 ;
    RECT 0 17.535 0.070 17.745 ;
    RECT 0 17.815 0.070 18.025 ;
    RECT 0 18.095 0.070 18.305 ;
    RECT 0 18.375 0.070 18.585 ;
    RECT 0 18.655 0.070 18.865 ;
    RECT 0 18.935 0.070 19.145 ;
    RECT 0 19.215 0.070 19.425 ;
    RECT 0 19.495 0.070 19.705 ;
    RECT 0 19.775 0.070 19.985 ;
    RECT 0 20.055 0.070 20.265 ;
    RECT 0 20.335 0.070 20.545 ;
    RECT 0 20.615 0.070 20.825 ;
    RECT 0 20.895 0.070 21.105 ;
    RECT 0 21.175 0.070 23.485 ;
    RECT 0 23.555 0.070 23.765 ;
    RECT 0 23.835 0.070 24.045 ;
    RECT 0 24.115 0.070 24.325 ;
    RECT 0 24.395 0.070 24.605 ;
    RECT 0 24.675 0.070 24.885 ;
    RECT 0 24.955 0.070 25.165 ;
    RECT 0 25.235 0.070 25.445 ;
    RECT 0 25.515 0.070 25.725 ;
    RECT 0 25.795 0.070 26.005 ;
    RECT 0 26.075 0.070 26.285 ;
    RECT 0 26.355 0.070 26.565 ;
    RECT 0 26.635 0.070 26.845 ;
    RECT 0 26.915 0.070 27.125 ;
    RECT 0 27.195 0.070 27.405 ;
    RECT 0 27.475 0.070 27.685 ;
    RECT 0 27.755 0.070 27.965 ;
    RECT 0 28.035 0.070 28.245 ;
    RECT 0 28.315 0.070 28.525 ;
    RECT 0 28.595 0.070 28.805 ;
    RECT 0 28.875 0.070 29.085 ;
    RECT 0 29.155 0.070 29.365 ;
    RECT 0 29.435 0.070 29.645 ;
    RECT 0 29.715 0.070 29.925 ;
    RECT 0 29.995 0.070 30.205 ;
    RECT 0 30.275 0.070 30.485 ;
    RECT 0 30.555 0.070 30.765 ;
    RECT 0 30.835 0.070 31.045 ;
    RECT 0 31.115 0.070 31.325 ;
    RECT 0 31.395 0.070 31.605 ;
    RECT 0 31.675 0.070 31.885 ;
    RECT 0 31.955 0.070 32.165 ;
    RECT 0 32.235 0.070 34.545 ;
    RECT 0 34.615 0.070 34.825 ;
    RECT 0 34.895 0.070 35.105 ;
    RECT 0 35.175 0.070 35.385 ;
    RECT 0 35.455 0.070 35.665 ;
    RECT 0 35.735 0.070 35.945 ;
    RECT 0 36.015 0.070 36.225 ;
    RECT 0 36.295 0.070 38.605 ;
    RECT 0 38.675 0.070 38.885 ;
    RECT 0 38.955 0.070 39.165 ;
    RECT 0 39.235 0.070 42.000 ;
    LAYER metal4 ;
    RECT 0 0 78.470 1.400 ;
    RECT 0 40.600 78.470 42.000 ;
    RECT 0.000 1.400 1.260 40.600 ;
    RECT 1.540 1.400 2.380 40.600 ;
    RECT 2.660 1.400 3.500 40.600 ;
    RECT 3.780 1.400 4.620 40.600 ;
    RECT 4.900 1.400 5.740 40.600 ;
    RECT 6.020 1.400 6.860 40.600 ;
    RECT 7.140 1.400 7.980 40.600 ;
    RECT 8.260 1.400 9.100 40.600 ;
    RECT 9.380 1.400 10.220 40.600 ;
    RECT 10.500 1.400 11.340 40.600 ;
    RECT 11.620 1.400 12.460 40.600 ;
    RECT 12.740 1.400 13.580 40.600 ;
    RECT 13.860 1.400 14.700 40.600 ;
    RECT 14.980 1.400 15.820 40.600 ;
    RECT 16.100 1.400 16.940 40.600 ;
    RECT 17.220 1.400 18.060 40.600 ;
    RECT 18.340 1.400 19.180 40.600 ;
    RECT 19.460 1.400 20.300 40.600 ;
    RECT 20.580 1.400 21.420 40.600 ;
    RECT 21.700 1.400 22.540 40.600 ;
    RECT 22.820 1.400 23.660 40.600 ;
    RECT 23.940 1.400 24.780 40.600 ;
    RECT 25.060 1.400 25.900 40.600 ;
    RECT 26.180 1.400 27.020 40.600 ;
    RECT 27.300 1.400 28.140 40.600 ;
    RECT 28.420 1.400 29.260 40.600 ;
    RECT 29.540 1.400 30.380 40.600 ;
    RECT 30.660 1.400 31.500 40.600 ;
    RECT 31.780 1.400 32.620 40.600 ;
    RECT 32.900 1.400 33.740 40.600 ;
    RECT 34.020 1.400 34.860 40.600 ;
    RECT 35.140 1.400 35.980 40.600 ;
    RECT 36.260 1.400 37.100 40.600 ;
    RECT 37.380 1.400 38.220 40.600 ;
    RECT 38.500 1.400 39.340 40.600 ;
    RECT 39.620 1.400 40.460 40.600 ;
    RECT 40.740 1.400 41.580 40.600 ;
    RECT 41.860 1.400 42.700 40.600 ;
    RECT 42.980 1.400 43.820 40.600 ;
    RECT 44.100 1.400 44.940 40.600 ;
    RECT 45.220 1.400 46.060 40.600 ;
    RECT 46.340 1.400 47.180 40.600 ;
    RECT 47.460 1.400 48.300 40.600 ;
    RECT 48.580 1.400 49.420 40.600 ;
    RECT 49.700 1.400 50.540 40.600 ;
    RECT 50.820 1.400 51.660 40.600 ;
    RECT 51.940 1.400 52.780 40.600 ;
    RECT 53.060 1.400 53.900 40.600 ;
    RECT 54.180 1.400 55.020 40.600 ;
    RECT 55.300 1.400 56.140 40.600 ;
    RECT 56.420 1.400 57.260 40.600 ;
    RECT 57.540 1.400 58.380 40.600 ;
    RECT 58.660 1.400 59.500 40.600 ;
    RECT 59.780 1.400 60.620 40.600 ;
    RECT 60.900 1.400 61.740 40.600 ;
    RECT 62.020 1.400 62.860 40.600 ;
    RECT 63.140 1.400 63.980 40.600 ;
    RECT 64.260 1.400 65.100 40.600 ;
    RECT 65.380 1.400 66.220 40.600 ;
    RECT 66.500 1.400 67.340 40.600 ;
    RECT 67.620 1.400 68.460 40.600 ;
    RECT 68.740 1.400 69.580 40.600 ;
    RECT 69.860 1.400 70.700 40.600 ;
    RECT 70.980 1.400 71.820 40.600 ;
    RECT 72.100 1.400 72.940 40.600 ;
    RECT 73.220 1.400 74.060 40.600 ;
    RECT 74.340 1.400 75.180 40.600 ;
    RECT 75.460 1.400 76.300 40.600 ;
    RECT 76.580 1.400 78.470 40.600 ;
    LAYER OVERLAP ;
    RECT 0 0 78.470 42.000 ;
  END
END fakeram45_128x32

END LIBRARY
