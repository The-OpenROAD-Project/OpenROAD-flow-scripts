module MuxTest_width_256_inputs_1_outputs_8_pipeline_5( // @[:@3.2]
  input          clock, // @[:@4.4]
  input          reset, // @[:@5.4]
  input  [2:0]   io_operation_0, // @[:@6.4]
  input  [2:0]   io_operation_1, // @[:@6.4]
  input  [2:0]   io_operation_2, // @[:@6.4]
  input  [2:0]   io_operation_3, // @[:@6.4]
  input  [2:0]   io_operation_4, // @[:@6.4]
  input  [2:0]   io_operation_5, // @[:@6.4]
  input  [2:0]   io_operation_6, // @[:@6.4]
  input  [2:0]   io_operation_7, // @[:@6.4]
  input  [255:0] io_inputs_0, // @[:@6.4]
  output [255:0] io_outputs_0, // @[:@6.4]
  output [255:0] io_outputs_1, // @[:@6.4]
  output [255:0] io_outputs_2, // @[:@6.4]
  output [255:0] io_outputs_3, // @[:@6.4]
  output [255:0] io_outputs_4, // @[:@6.4]
  output [255:0] io_outputs_5, // @[:@6.4]
  output [255:0] io_outputs_6, // @[:@6.4]
  output [255:0] io_outputs_7 // @[:@6.4]
);
  wire [256:0] _T_404; // @[MuxTest_width_256_inputs_1_outputs_8_pipeline_5s.scala 32:53:@8.4]
  wire [255:0] _T_405; // @[MuxTest_width_256_inputs_1_outputs_8_pipeline_5s.scala 32:53:@9.4]
  wire [511:0] _T_407; // @[MuxTest_width_256_inputs_1_outputs_8_pipeline_5s.scala 33:58:@10.4]
  wire [255:0] _T_409; // @[MuxTest_width_256_inputs_1_outputs_8_pipeline_5s.scala 34:56:@11.4]
  wire  _T_410; // @[Mux.scala 46:19:@12.4]
  wire [255:0] _T_411; // @[Mux.scala 46:16:@13.4]
  wire  _T_412; // @[Mux.scala 46:19:@14.4]
  wire [511:0] _T_413; // @[Mux.scala 46:16:@15.4]
  wire  _T_414; // @[Mux.scala 46:19:@16.4]
  wire [511:0] _T_415; // @[Mux.scala 46:16:@17.4]
  wire  _T_416; // @[Mux.scala 46:19:@18.4]
  wire  _T_427; // @[Mux.scala 46:19:@24.4]
  wire [255:0] _T_428; // @[Mux.scala 46:16:@25.4]
  wire  _T_429; // @[Mux.scala 46:19:@26.4]
  wire [511:0] _T_430; // @[Mux.scala 46:16:@27.4]
  wire  _T_431; // @[Mux.scala 46:19:@28.4]
  wire [511:0] _T_432; // @[Mux.scala 46:16:@29.4]
  wire  _T_433; // @[Mux.scala 46:19:@30.4]
  wire  _T_444; // @[Mux.scala 46:19:@36.4]
  wire [255:0] _T_445; // @[Mux.scala 46:16:@37.4]
  wire  _T_446; // @[Mux.scala 46:19:@38.4]
  wire [511:0] _T_447; // @[Mux.scala 46:16:@39.4]
  wire  _T_448; // @[Mux.scala 46:19:@40.4]
  wire [511:0] _T_449; // @[Mux.scala 46:16:@41.4]
  wire  _T_450; // @[Mux.scala 46:19:@42.4]
  wire  _T_461; // @[Mux.scala 46:19:@48.4]
  wire [255:0] _T_462; // @[Mux.scala 46:16:@49.4]
  wire  _T_463; // @[Mux.scala 46:19:@50.4]
  wire [511:0] _T_464; // @[Mux.scala 46:16:@51.4]
  wire  _T_465; // @[Mux.scala 46:19:@52.4]
  wire [511:0] _T_466; // @[Mux.scala 46:16:@53.4]
  wire  _T_467; // @[Mux.scala 46:19:@54.4]
  wire  _T_478; // @[Mux.scala 46:19:@60.4]
  wire [255:0] _T_479; // @[Mux.scala 46:16:@61.4]
  wire  _T_480; // @[Mux.scala 46:19:@62.4]
  wire [511:0] _T_481; // @[Mux.scala 46:16:@63.4]
  wire  _T_482; // @[Mux.scala 46:19:@64.4]
  wire [511:0] _T_483; // @[Mux.scala 46:16:@65.4]
  wire  _T_484; // @[Mux.scala 46:19:@66.4]
  wire  _T_495; // @[Mux.scala 46:19:@72.4]
  wire [255:0] _T_496; // @[Mux.scala 46:16:@73.4]
  wire  _T_497; // @[Mux.scala 46:19:@74.4]
  wire [511:0] _T_498; // @[Mux.scala 46:16:@75.4]
  wire  _T_499; // @[Mux.scala 46:19:@76.4]
  wire [511:0] _T_500; // @[Mux.scala 46:16:@77.4]
  wire  _T_501; // @[Mux.scala 46:19:@78.4]
  wire  _T_512; // @[Mux.scala 46:19:@84.4]
  wire [255:0] _T_513; // @[Mux.scala 46:16:@85.4]
  wire  _T_514; // @[Mux.scala 46:19:@86.4]
  wire [511:0] _T_515; // @[Mux.scala 46:16:@87.4]
  wire  _T_516; // @[Mux.scala 46:19:@88.4]
  wire [511:0] _T_517; // @[Mux.scala 46:16:@89.4]
  wire  _T_518; // @[Mux.scala 46:19:@90.4]
  wire  _T_529; // @[Mux.scala 46:19:@96.4]
  wire [255:0] _T_530; // @[Mux.scala 46:16:@97.4]
  wire  _T_531; // @[Mux.scala 46:19:@98.4]
  wire [511:0] _T_532; // @[Mux.scala 46:16:@99.4]
  wire  _T_533; // @[Mux.scala 46:19:@100.4]
  wire [511:0] _T_534; // @[Mux.scala 46:16:@101.4]
  wire  _T_535; // @[Mux.scala 46:19:@102.4]
  reg [511:0] _T_539; // @[Reg.scala 11:16:@104.4]
  reg [511:0] _RAND_0;
  reg [511:0] _T_541; // @[Reg.scala 11:16:@108.4]
  reg [511:0] _RAND_1;
  reg [511:0] _T_543; // @[Reg.scala 11:16:@112.4]
  reg [511:0] _RAND_2;
  reg [511:0] _T_545; // @[Reg.scala 11:16:@116.4]
  reg [511:0] _RAND_3;
  reg [511:0] _T_547; // @[Reg.scala 11:16:@120.4]
  reg [511:0] _RAND_4;
  reg [511:0] _T_550; // @[Reg.scala 11:16:@124.4]
  reg [511:0] _RAND_5;
  reg [511:0] _T_552; // @[Reg.scala 11:16:@128.4]
  reg [511:0] _RAND_6;
  reg [511:0] _T_554; // @[Reg.scala 11:16:@132.4]
  reg [511:0] _RAND_7;
  reg [511:0] _T_556; // @[Reg.scala 11:16:@136.4]
  reg [511:0] _RAND_8;
  reg [511:0] _T_558; // @[Reg.scala 11:16:@140.4]
  reg [511:0] _RAND_9;
  reg [511:0] _T_561; // @[Reg.scala 11:16:@144.4]
  reg [511:0] _RAND_10;
  reg [511:0] _T_563; // @[Reg.scala 11:16:@148.4]
  reg [511:0] _RAND_11;
  reg [511:0] _T_565; // @[Reg.scala 11:16:@152.4]
  reg [511:0] _RAND_12;
  reg [511:0] _T_567; // @[Reg.scala 11:16:@156.4]
  reg [511:0] _RAND_13;
  reg [511:0] _T_569; // @[Reg.scala 11:16:@160.4]
  reg [511:0] _RAND_14;
  reg [511:0] _T_572; // @[Reg.scala 11:16:@164.4]
  reg [511:0] _RAND_15;
  reg [511:0] _T_574; // @[Reg.scala 11:16:@168.4]
  reg [511:0] _RAND_16;
  reg [511:0] _T_576; // @[Reg.scala 11:16:@172.4]
  reg [511:0] _RAND_17;
  reg [511:0] _T_578; // @[Reg.scala 11:16:@176.4]
  reg [511:0] _RAND_18;
  reg [511:0] _T_580; // @[Reg.scala 11:16:@180.4]
  reg [511:0] _RAND_19;
  reg [511:0] _T_583; // @[Reg.scala 11:16:@184.4]
  reg [511:0] _RAND_20;
  reg [511:0] _T_585; // @[Reg.scala 11:16:@188.4]
  reg [511:0] _RAND_21;
  reg [511:0] _T_587; // @[Reg.scala 11:16:@192.4]
  reg [511:0] _RAND_22;
  reg [511:0] _T_589; // @[Reg.scala 11:16:@196.4]
  reg [511:0] _RAND_23;
  reg [511:0] _T_591; // @[Reg.scala 11:16:@200.4]
  reg [511:0] _RAND_24;
  reg [511:0] _T_594; // @[Reg.scala 11:16:@204.4]
  reg [511:0] _RAND_25;
  reg [511:0] _T_596; // @[Reg.scala 11:16:@208.4]
  reg [511:0] _RAND_26;
  reg [511:0] _T_598; // @[Reg.scala 11:16:@212.4]
  reg [511:0] _RAND_27;
  reg [511:0] _T_600; // @[Reg.scala 11:16:@216.4]
  reg [511:0] _RAND_28;
  reg [511:0] _T_602; // @[Reg.scala 11:16:@220.4]
  reg [511:0] _RAND_29;
  reg [511:0] _T_605; // @[Reg.scala 11:16:@224.4]
  reg [511:0] _RAND_30;
  reg [511:0] _T_607; // @[Reg.scala 11:16:@228.4]
  reg [511:0] _RAND_31;
  reg [511:0] _T_609; // @[Reg.scala 11:16:@232.4]
  reg [511:0] _RAND_32;
  reg [511:0] _T_611; // @[Reg.scala 11:16:@236.4]
  reg [511:0] _RAND_33;
  reg [511:0] _T_613; // @[Reg.scala 11:16:@240.4]
  reg [511:0] _RAND_34;
  reg [511:0] _T_616; // @[Reg.scala 11:16:@244.4]
  reg [511:0] _RAND_35;
  reg [511:0] _T_618; // @[Reg.scala 11:16:@248.4]
  reg [511:0] _RAND_36;
  reg [511:0] _T_620; // @[Reg.scala 11:16:@252.4]
  reg [511:0] _RAND_37;
  reg [511:0] _T_622; // @[Reg.scala 11:16:@256.4]
  reg [511:0] _RAND_38;
  reg [511:0] _T_624; // @[Reg.scala 11:16:@260.4]
  reg [511:0] _RAND_39;
  assign _T_404 = io_inputs_0 + io_inputs_0; // @[MuxTest_width_256_inputs_1_outputs_8_pipeline_5s.scala 32:53:@8.4]
  assign _T_405 = io_inputs_0 + io_inputs_0; // @[MuxTest_width_256_inputs_1_outputs_8_pipeline_5s.scala 32:53:@9.4]
  assign _T_407 = io_inputs_0 * io_inputs_0; // @[MuxTest_width_256_inputs_1_outputs_8_pipeline_5s.scala 33:58:@10.4]
  assign _T_409 = io_inputs_0 / io_inputs_0; // @[MuxTest_width_256_inputs_1_outputs_8_pipeline_5s.scala 34:56:@11.4]
  assign _T_410 = 3'h3 == io_operation_0; // @[Mux.scala 46:19:@12.4]
  assign _T_411 = _T_410 ? _T_409 : 256'h0; // @[Mux.scala 46:16:@13.4]
  assign _T_412 = 3'h2 == io_operation_0; // @[Mux.scala 46:19:@14.4]
  assign _T_413 = _T_412 ? _T_407 : {{256'd0}, _T_411}; // @[Mux.scala 46:16:@15.4]
  assign _T_414 = 3'h1 == io_operation_0; // @[Mux.scala 46:19:@16.4]
  assign _T_415 = _T_414 ? {{256'd0}, _T_405} : _T_413; // @[Mux.scala 46:16:@17.4]
  assign _T_416 = 3'h0 == io_operation_0; // @[Mux.scala 46:19:@18.4]
  assign _T_427 = 3'h3 == io_operation_1; // @[Mux.scala 46:19:@24.4]
  assign _T_428 = _T_427 ? _T_409 : 256'h0; // @[Mux.scala 46:16:@25.4]
  assign _T_429 = 3'h2 == io_operation_1; // @[Mux.scala 46:19:@26.4]
  assign _T_430 = _T_429 ? _T_407 : {{256'd0}, _T_428}; // @[Mux.scala 46:16:@27.4]
  assign _T_431 = 3'h1 == io_operation_1; // @[Mux.scala 46:19:@28.4]
  assign _T_432 = _T_431 ? {{256'd0}, _T_405} : _T_430; // @[Mux.scala 46:16:@29.4]
  assign _T_433 = 3'h0 == io_operation_1; // @[Mux.scala 46:19:@30.4]
  assign _T_444 = 3'h3 == io_operation_2; // @[Mux.scala 46:19:@36.4]
  assign _T_445 = _T_444 ? _T_409 : 256'h0; // @[Mux.scala 46:16:@37.4]
  assign _T_446 = 3'h2 == io_operation_2; // @[Mux.scala 46:19:@38.4]
  assign _T_447 = _T_446 ? _T_407 : {{256'd0}, _T_445}; // @[Mux.scala 46:16:@39.4]
  assign _T_448 = 3'h1 == io_operation_2; // @[Mux.scala 46:19:@40.4]
  assign _T_449 = _T_448 ? {{256'd0}, _T_405} : _T_447; // @[Mux.scala 46:16:@41.4]
  assign _T_450 = 3'h0 == io_operation_2; // @[Mux.scala 46:19:@42.4]
  assign _T_461 = 3'h3 == io_operation_3; // @[Mux.scala 46:19:@48.4]
  assign _T_462 = _T_461 ? _T_409 : 256'h0; // @[Mux.scala 46:16:@49.4]
  assign _T_463 = 3'h2 == io_operation_3; // @[Mux.scala 46:19:@50.4]
  assign _T_464 = _T_463 ? _T_407 : {{256'd0}, _T_462}; // @[Mux.scala 46:16:@51.4]
  assign _T_465 = 3'h1 == io_operation_3; // @[Mux.scala 46:19:@52.4]
  assign _T_466 = _T_465 ? {{256'd0}, _T_405} : _T_464; // @[Mux.scala 46:16:@53.4]
  assign _T_467 = 3'h0 == io_operation_3; // @[Mux.scala 46:19:@54.4]
  assign _T_478 = 3'h3 == io_operation_4; // @[Mux.scala 46:19:@60.4]
  assign _T_479 = _T_478 ? _T_409 : 256'h0; // @[Mux.scala 46:16:@61.4]
  assign _T_480 = 3'h2 == io_operation_4; // @[Mux.scala 46:19:@62.4]
  assign _T_481 = _T_480 ? _T_407 : {{256'd0}, _T_479}; // @[Mux.scala 46:16:@63.4]
  assign _T_482 = 3'h1 == io_operation_4; // @[Mux.scala 46:19:@64.4]
  assign _T_483 = _T_482 ? {{256'd0}, _T_405} : _T_481; // @[Mux.scala 46:16:@65.4]
  assign _T_484 = 3'h0 == io_operation_4; // @[Mux.scala 46:19:@66.4]
  assign _T_495 = 3'h3 == io_operation_5; // @[Mux.scala 46:19:@72.4]
  assign _T_496 = _T_495 ? _T_409 : 256'h0; // @[Mux.scala 46:16:@73.4]
  assign _T_497 = 3'h2 == io_operation_5; // @[Mux.scala 46:19:@74.4]
  assign _T_498 = _T_497 ? _T_407 : {{256'd0}, _T_496}; // @[Mux.scala 46:16:@75.4]
  assign _T_499 = 3'h1 == io_operation_5; // @[Mux.scala 46:19:@76.4]
  assign _T_500 = _T_499 ? {{256'd0}, _T_405} : _T_498; // @[Mux.scala 46:16:@77.4]
  assign _T_501 = 3'h0 == io_operation_5; // @[Mux.scala 46:19:@78.4]
  assign _T_512 = 3'h3 == io_operation_6; // @[Mux.scala 46:19:@84.4]
  assign _T_513 = _T_512 ? _T_409 : 256'h0; // @[Mux.scala 46:16:@85.4]
  assign _T_514 = 3'h2 == io_operation_6; // @[Mux.scala 46:19:@86.4]
  assign _T_515 = _T_514 ? _T_407 : {{256'd0}, _T_513}; // @[Mux.scala 46:16:@87.4]
  assign _T_516 = 3'h1 == io_operation_6; // @[Mux.scala 46:19:@88.4]
  assign _T_517 = _T_516 ? {{256'd0}, _T_405} : _T_515; // @[Mux.scala 46:16:@89.4]
  assign _T_518 = 3'h0 == io_operation_6; // @[Mux.scala 46:19:@90.4]
  assign _T_529 = 3'h3 == io_operation_7; // @[Mux.scala 46:19:@96.4]
  assign _T_530 = _T_529 ? _T_409 : 256'h0; // @[Mux.scala 46:16:@97.4]
  assign _T_531 = 3'h2 == io_operation_7; // @[Mux.scala 46:19:@98.4]
  assign _T_532 = _T_531 ? _T_407 : {{256'd0}, _T_530}; // @[Mux.scala 46:16:@99.4]
  assign _T_533 = 3'h1 == io_operation_7; // @[Mux.scala 46:19:@100.4]
  assign _T_534 = _T_533 ? {{256'd0}, _T_405} : _T_532; // @[Mux.scala 46:16:@101.4]
  assign _T_535 = 3'h0 == io_operation_7; // @[Mux.scala 46:19:@102.4]
  assign io_outputs_0 = _T_547[255:0]; // @[MuxTest_width_256_inputs_1_outputs_8_pipeline_5s.scala 23:14:@264.4]
  assign io_outputs_1 = _T_558[255:0]; // @[MuxTest_width_256_inputs_1_outputs_8_pipeline_5s.scala 23:14:@265.4]
  assign io_outputs_2 = _T_569[255:0]; // @[MuxTest_width_256_inputs_1_outputs_8_pipeline_5s.scala 23:14:@266.4]
  assign io_outputs_3 = _T_580[255:0]; // @[MuxTest_width_256_inputs_1_outputs_8_pipeline_5s.scala 23:14:@267.4]
  assign io_outputs_4 = _T_591[255:0]; // @[MuxTest_width_256_inputs_1_outputs_8_pipeline_5s.scala 23:14:@268.4]
  assign io_outputs_5 = _T_602[255:0]; // @[MuxTest_width_256_inputs_1_outputs_8_pipeline_5s.scala 23:14:@269.4]
  assign io_outputs_6 = _T_613[255:0]; // @[MuxTest_width_256_inputs_1_outputs_8_pipeline_5s.scala 23:14:@270.4]
  assign io_outputs_7 = _T_624[255:0]; // @[MuxTest_width_256_inputs_1_outputs_8_pipeline_5s.scala 23:14:@271.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {16{`RANDOM}};
  _T_539 = _RAND_0[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {16{`RANDOM}};
  _T_541 = _RAND_1[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {16{`RANDOM}};
  _T_543 = _RAND_2[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {16{`RANDOM}};
  _T_545 = _RAND_3[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {16{`RANDOM}};
  _T_547 = _RAND_4[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {16{`RANDOM}};
  _T_550 = _RAND_5[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {16{`RANDOM}};
  _T_552 = _RAND_6[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {16{`RANDOM}};
  _T_554 = _RAND_7[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {16{`RANDOM}};
  _T_556 = _RAND_8[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {16{`RANDOM}};
  _T_558 = _RAND_9[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {16{`RANDOM}};
  _T_561 = _RAND_10[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {16{`RANDOM}};
  _T_563 = _RAND_11[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {16{`RANDOM}};
  _T_565 = _RAND_12[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {16{`RANDOM}};
  _T_567 = _RAND_13[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {16{`RANDOM}};
  _T_569 = _RAND_14[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {16{`RANDOM}};
  _T_572 = _RAND_15[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {16{`RANDOM}};
  _T_574 = _RAND_16[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {16{`RANDOM}};
  _T_576 = _RAND_17[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {16{`RANDOM}};
  _T_578 = _RAND_18[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {16{`RANDOM}};
  _T_580 = _RAND_19[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {16{`RANDOM}};
  _T_583 = _RAND_20[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {16{`RANDOM}};
  _T_585 = _RAND_21[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {16{`RANDOM}};
  _T_587 = _RAND_22[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {16{`RANDOM}};
  _T_589 = _RAND_23[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {16{`RANDOM}};
  _T_591 = _RAND_24[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {16{`RANDOM}};
  _T_594 = _RAND_25[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {16{`RANDOM}};
  _T_596 = _RAND_26[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {16{`RANDOM}};
  _T_598 = _RAND_27[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {16{`RANDOM}};
  _T_600 = _RAND_28[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {16{`RANDOM}};
  _T_602 = _RAND_29[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {16{`RANDOM}};
  _T_605 = _RAND_30[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {16{`RANDOM}};
  _T_607 = _RAND_31[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {16{`RANDOM}};
  _T_609 = _RAND_32[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {16{`RANDOM}};
  _T_611 = _RAND_33[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {16{`RANDOM}};
  _T_613 = _RAND_34[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {16{`RANDOM}};
  _T_616 = _RAND_35[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {16{`RANDOM}};
  _T_618 = _RAND_36[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {16{`RANDOM}};
  _T_620 = _RAND_37[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {16{`RANDOM}};
  _T_622 = _RAND_38[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {16{`RANDOM}};
  _T_624 = _RAND_39[511:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_416) begin
      _T_539 <= {{256'd0}, io_inputs_0};
    end else begin
      _T_539 <= _T_415;
    end
    _T_541 <= _T_539;
    _T_543 <= _T_541;
    _T_545 <= _T_543;
    _T_547 <= _T_545;
    if (_T_433) begin
      _T_550 <= {{256'd0}, io_inputs_0};
    end else begin
      _T_550 <= _T_432;
    end
    _T_552 <= _T_550;
    _T_554 <= _T_552;
    _T_556 <= _T_554;
    _T_558 <= _T_556;
    if (_T_450) begin
      _T_561 <= {{256'd0}, io_inputs_0};
    end else begin
      _T_561 <= _T_449;
    end
    _T_563 <= _T_561;
    _T_565 <= _T_563;
    _T_567 <= _T_565;
    _T_569 <= _T_567;
    if (_T_467) begin
      _T_572 <= {{256'd0}, io_inputs_0};
    end else begin
      _T_572 <= _T_466;
    end
    _T_574 <= _T_572;
    _T_576 <= _T_574;
    _T_578 <= _T_576;
    _T_580 <= _T_578;
    if (_T_484) begin
      _T_583 <= {{256'd0}, io_inputs_0};
    end else begin
      _T_583 <= _T_483;
    end
    _T_585 <= _T_583;
    _T_587 <= _T_585;
    _T_589 <= _T_587;
    _T_591 <= _T_589;
    if (_T_501) begin
      _T_594 <= {{256'd0}, io_inputs_0};
    end else begin
      _T_594 <= _T_500;
    end
    _T_596 <= _T_594;
    _T_598 <= _T_596;
    _T_600 <= _T_598;
    _T_602 <= _T_600;
    if (_T_518) begin
      _T_605 <= {{256'd0}, io_inputs_0};
    end else begin
      _T_605 <= _T_517;
    end
    _T_607 <= _T_605;
    _T_609 <= _T_607;
    _T_611 <= _T_609;
    _T_613 <= _T_611;
    if (_T_535) begin
      _T_616 <= {{256'd0}, io_inputs_0};
    end else begin
      _T_616 <= _T_534;
    end
    _T_618 <= _T_616;
    _T_620 <= _T_618;
    _T_622 <= _T_620;
    _T_624 <= _T_622;
  end
endmodule
