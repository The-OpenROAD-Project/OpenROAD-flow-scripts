../../../platforms/nangate45/lef/fakeram45_64x15.lef