module fakeram45_256x32 (
   output reg [31:0] rd_out,
   input logic [7:0] addr_in,
   input logic we_in,
   input logic [31:0] wd_in,
   input logic clk,
   input logic ce_in
);
endmodule
