module MockArray(
  input        clock,
  input        reset,
  input  [7:0] io_insHorizontal_0_0,
  input  [7:0] io_insHorizontal_1_0,
  output [7:0] io_outsHorizontal_0_0,
  output [7:0] io_outsHorizontal_1_0,
  input  [7:0] io_insVertical_0_0,
  input  [7:0] io_insVertical_0_1,
  input  [7:0] io_insVertical_0_2,
  input  [7:0] io_insVertical_0_3,
  input  [7:0] io_insVertical_0_4,
  input  [7:0] io_insVertical_0_5,
  input  [7:0] io_insVertical_0_6,
  input  [7:0] io_insVertical_0_7,
  input  [7:0] io_insVertical_0_8,
  input  [7:0] io_insVertical_0_9,
  input  [7:0] io_insVertical_0_10,
  input  [7:0] io_insVertical_0_11,
  input  [7:0] io_insVertical_0_12,
  input  [7:0] io_insVertical_0_13,
  input  [7:0] io_insVertical_0_14,
  input  [7:0] io_insVertical_0_15,
  input  [7:0] io_insVertical_0_16,
  input  [7:0] io_insVertical_0_17,
  input  [7:0] io_insVertical_0_18,
  input  [7:0] io_insVertical_0_19,
  input  [7:0] io_insVertical_0_20,
  input  [7:0] io_insVertical_0_21,
  input  [7:0] io_insVertical_0_22,
  input  [7:0] io_insVertical_0_23,
  input  [7:0] io_insVertical_0_24,
  input  [7:0] io_insVertical_0_25,
  input  [7:0] io_insVertical_0_26,
  input  [7:0] io_insVertical_0_27,
  input  [7:0] io_insVertical_0_28,
  input  [7:0] io_insVertical_0_29,
  input  [7:0] io_insVertical_0_30,
  input  [7:0] io_insVertical_0_31,
  input  [7:0] io_insVertical_0_32,
  input  [7:0] io_insVertical_0_33,
  input  [7:0] io_insVertical_0_34,
  input  [7:0] io_insVertical_0_35,
  input  [7:0] io_insVertical_0_36,
  input  [7:0] io_insVertical_0_37,
  input  [7:0] io_insVertical_0_38,
  input  [7:0] io_insVertical_0_39,
  input  [7:0] io_insVertical_0_40,
  input  [7:0] io_insVertical_0_41,
  input  [7:0] io_insVertical_0_42,
  input  [7:0] io_insVertical_0_43,
  input  [7:0] io_insVertical_0_44,
  input  [7:0] io_insVertical_0_45,
  input  [7:0] io_insVertical_0_46,
  input  [7:0] io_insVertical_0_47,
  input  [7:0] io_insVertical_0_48,
  input  [7:0] io_insVertical_0_49,
  input  [7:0] io_insVertical_0_50,
  input  [7:0] io_insVertical_0_51,
  input  [7:0] io_insVertical_0_52,
  input  [7:0] io_insVertical_0_53,
  input  [7:0] io_insVertical_0_54,
  input  [7:0] io_insVertical_0_55,
  input  [7:0] io_insVertical_0_56,
  input  [7:0] io_insVertical_0_57,
  input  [7:0] io_insVertical_0_58,
  input  [7:0] io_insVertical_0_59,
  input  [7:0] io_insVertical_0_60,
  input  [7:0] io_insVertical_0_61,
  input  [7:0] io_insVertical_0_62,
  input  [7:0] io_insVertical_0_63,
  input  [7:0] io_insVertical_0_64,
  input  [7:0] io_insVertical_0_65,
  input  [7:0] io_insVertical_0_66,
  input  [7:0] io_insVertical_0_67,
  input  [7:0] io_insVertical_0_68,
  input  [7:0] io_insVertical_0_69,
  input  [7:0] io_insVertical_0_70,
  input  [7:0] io_insVertical_0_71,
  input  [7:0] io_insVertical_0_72,
  input  [7:0] io_insVertical_0_73,
  input  [7:0] io_insVertical_0_74,
  input  [7:0] io_insVertical_0_75,
  input  [7:0] io_insVertical_0_76,
  input  [7:0] io_insVertical_0_77,
  input  [7:0] io_insVertical_0_78,
  input  [7:0] io_insVertical_0_79,
  input  [7:0] io_insVertical_0_80,
  input  [7:0] io_insVertical_0_81,
  input  [7:0] io_insVertical_0_82,
  input  [7:0] io_insVertical_0_83,
  input  [7:0] io_insVertical_0_84,
  input  [7:0] io_insVertical_0_85,
  input  [7:0] io_insVertical_0_86,
  input  [7:0] io_insVertical_0_87,
  input  [7:0] io_insVertical_0_88,
  input  [7:0] io_insVertical_0_89,
  input  [7:0] io_insVertical_0_90,
  input  [7:0] io_insVertical_0_91,
  input  [7:0] io_insVertical_0_92,
  input  [7:0] io_insVertical_0_93,
  input  [7:0] io_insVertical_0_94,
  input  [7:0] io_insVertical_0_95,
  input  [7:0] io_insVertical_0_96,
  input  [7:0] io_insVertical_0_97,
  input  [7:0] io_insVertical_0_98,
  input  [7:0] io_insVertical_0_99,
  input  [7:0] io_insVertical_0_100,
  input  [7:0] io_insVertical_0_101,
  input  [7:0] io_insVertical_0_102,
  input  [7:0] io_insVertical_0_103,
  input  [7:0] io_insVertical_0_104,
  input  [7:0] io_insVertical_0_105,
  input  [7:0] io_insVertical_0_106,
  input  [7:0] io_insVertical_0_107,
  input  [7:0] io_insVertical_0_108,
  input  [7:0] io_insVertical_0_109,
  input  [7:0] io_insVertical_0_110,
  input  [7:0] io_insVertical_0_111,
  input  [7:0] io_insVertical_0_112,
  input  [7:0] io_insVertical_0_113,
  input  [7:0] io_insVertical_0_114,
  input  [7:0] io_insVertical_0_115,
  input  [7:0] io_insVertical_0_116,
  input  [7:0] io_insVertical_0_117,
  input  [7:0] io_insVertical_0_118,
  input  [7:0] io_insVertical_0_119,
  input  [7:0] io_insVertical_0_120,
  input  [7:0] io_insVertical_0_121,
  input  [7:0] io_insVertical_0_122,
  input  [7:0] io_insVertical_0_123,
  input  [7:0] io_insVertical_0_124,
  input  [7:0] io_insVertical_0_125,
  input  [7:0] io_insVertical_0_126,
  input  [7:0] io_insVertical_0_127,
  input  [7:0] io_insVertical_0_128,
  input  [7:0] io_insVertical_0_129,
  input  [7:0] io_insVertical_0_130,
  input  [7:0] io_insVertical_0_131,
  input  [7:0] io_insVertical_0_132,
  input  [7:0] io_insVertical_0_133,
  input  [7:0] io_insVertical_0_134,
  input  [7:0] io_insVertical_0_135,
  input  [7:0] io_insVertical_0_136,
  input  [7:0] io_insVertical_0_137,
  input  [7:0] io_insVertical_0_138,
  input  [7:0] io_insVertical_0_139,
  input  [7:0] io_insVertical_0_140,
  input  [7:0] io_insVertical_0_141,
  input  [7:0] io_insVertical_0_142,
  input  [7:0] io_insVertical_0_143,
  input  [7:0] io_insVertical_0_144,
  input  [7:0] io_insVertical_0_145,
  input  [7:0] io_insVertical_0_146,
  input  [7:0] io_insVertical_0_147,
  input  [7:0] io_insVertical_0_148,
  input  [7:0] io_insVertical_0_149,
  input  [7:0] io_insVertical_0_150,
  input  [7:0] io_insVertical_0_151,
  input  [7:0] io_insVertical_0_152,
  input  [7:0] io_insVertical_0_153,
  input  [7:0] io_insVertical_0_154,
  input  [7:0] io_insVertical_0_155,
  input  [7:0] io_insVertical_0_156,
  input  [7:0] io_insVertical_0_157,
  input  [7:0] io_insVertical_0_158,
  input  [7:0] io_insVertical_0_159,
  input  [7:0] io_insVertical_0_160,
  input  [7:0] io_insVertical_0_161,
  input  [7:0] io_insVertical_0_162,
  input  [7:0] io_insVertical_0_163,
  input  [7:0] io_insVertical_0_164,
  input  [7:0] io_insVertical_0_165,
  input  [7:0] io_insVertical_0_166,
  input  [7:0] io_insVertical_0_167,
  input  [7:0] io_insVertical_0_168,
  input  [7:0] io_insVertical_0_169,
  input  [7:0] io_insVertical_0_170,
  input  [7:0] io_insVertical_0_171,
  input  [7:0] io_insVertical_0_172,
  input  [7:0] io_insVertical_0_173,
  input  [7:0] io_insVertical_0_174,
  input  [7:0] io_insVertical_0_175,
  input  [7:0] io_insVertical_0_176,
  input  [7:0] io_insVertical_0_177,
  input  [7:0] io_insVertical_0_178,
  input  [7:0] io_insVertical_0_179,
  input  [7:0] io_insVertical_0_180,
  input  [7:0] io_insVertical_0_181,
  input  [7:0] io_insVertical_0_182,
  input  [7:0] io_insVertical_0_183,
  input  [7:0] io_insVertical_0_184,
  input  [7:0] io_insVertical_0_185,
  input  [7:0] io_insVertical_0_186,
  input  [7:0] io_insVertical_0_187,
  input  [7:0] io_insVertical_0_188,
  input  [7:0] io_insVertical_0_189,
  input  [7:0] io_insVertical_0_190,
  input  [7:0] io_insVertical_0_191,
  input  [7:0] io_insVertical_0_192,
  input  [7:0] io_insVertical_0_193,
  input  [7:0] io_insVertical_0_194,
  input  [7:0] io_insVertical_0_195,
  input  [7:0] io_insVertical_0_196,
  input  [7:0] io_insVertical_0_197,
  input  [7:0] io_insVertical_0_198,
  input  [7:0] io_insVertical_0_199,
  input  [7:0] io_insVertical_0_200,
  input  [7:0] io_insVertical_0_201,
  input  [7:0] io_insVertical_0_202,
  input  [7:0] io_insVertical_0_203,
  input  [7:0] io_insVertical_0_204,
  input  [7:0] io_insVertical_0_205,
  input  [7:0] io_insVertical_0_206,
  input  [7:0] io_insVertical_0_207,
  input  [7:0] io_insVertical_0_208,
  input  [7:0] io_insVertical_0_209,
  input  [7:0] io_insVertical_0_210,
  input  [7:0] io_insVertical_0_211,
  input  [7:0] io_insVertical_0_212,
  input  [7:0] io_insVertical_0_213,
  input  [7:0] io_insVertical_0_214,
  input  [7:0] io_insVertical_0_215,
  input  [7:0] io_insVertical_0_216,
  input  [7:0] io_insVertical_0_217,
  input  [7:0] io_insVertical_0_218,
  input  [7:0] io_insVertical_0_219,
  input  [7:0] io_insVertical_0_220,
  input  [7:0] io_insVertical_0_221,
  input  [7:0] io_insVertical_0_222,
  input  [7:0] io_insVertical_0_223,
  input  [7:0] io_insVertical_0_224,
  input  [7:0] io_insVertical_0_225,
  input  [7:0] io_insVertical_0_226,
  input  [7:0] io_insVertical_0_227,
  input  [7:0] io_insVertical_0_228,
  input  [7:0] io_insVertical_0_229,
  input  [7:0] io_insVertical_0_230,
  input  [7:0] io_insVertical_0_231,
  input  [7:0] io_insVertical_0_232,
  input  [7:0] io_insVertical_0_233,
  input  [7:0] io_insVertical_0_234,
  input  [7:0] io_insVertical_0_235,
  input  [7:0] io_insVertical_0_236,
  input  [7:0] io_insVertical_0_237,
  input  [7:0] io_insVertical_0_238,
  input  [7:0] io_insVertical_0_239,
  input  [7:0] io_insVertical_0_240,
  input  [7:0] io_insVertical_0_241,
  input  [7:0] io_insVertical_0_242,
  input  [7:0] io_insVertical_0_243,
  input  [7:0] io_insVertical_0_244,
  input  [7:0] io_insVertical_0_245,
  input  [7:0] io_insVertical_0_246,
  input  [7:0] io_insVertical_0_247,
  input  [7:0] io_insVertical_0_248,
  input  [7:0] io_insVertical_0_249,
  input  [7:0] io_insVertical_0_250,
  input  [7:0] io_insVertical_0_251,
  input  [7:0] io_insVertical_0_252,
  input  [7:0] io_insVertical_0_253,
  input  [7:0] io_insVertical_0_254,
  input  [7:0] io_insVertical_0_255,
  input  [7:0] io_insVertical_1_0,
  input  [7:0] io_insVertical_1_1,
  input  [7:0] io_insVertical_1_2,
  input  [7:0] io_insVertical_1_3,
  input  [7:0] io_insVertical_1_4,
  input  [7:0] io_insVertical_1_5,
  input  [7:0] io_insVertical_1_6,
  input  [7:0] io_insVertical_1_7,
  input  [7:0] io_insVertical_1_8,
  input  [7:0] io_insVertical_1_9,
  input  [7:0] io_insVertical_1_10,
  input  [7:0] io_insVertical_1_11,
  input  [7:0] io_insVertical_1_12,
  input  [7:0] io_insVertical_1_13,
  input  [7:0] io_insVertical_1_14,
  input  [7:0] io_insVertical_1_15,
  input  [7:0] io_insVertical_1_16,
  input  [7:0] io_insVertical_1_17,
  input  [7:0] io_insVertical_1_18,
  input  [7:0] io_insVertical_1_19,
  input  [7:0] io_insVertical_1_20,
  input  [7:0] io_insVertical_1_21,
  input  [7:0] io_insVertical_1_22,
  input  [7:0] io_insVertical_1_23,
  input  [7:0] io_insVertical_1_24,
  input  [7:0] io_insVertical_1_25,
  input  [7:0] io_insVertical_1_26,
  input  [7:0] io_insVertical_1_27,
  input  [7:0] io_insVertical_1_28,
  input  [7:0] io_insVertical_1_29,
  input  [7:0] io_insVertical_1_30,
  input  [7:0] io_insVertical_1_31,
  input  [7:0] io_insVertical_1_32,
  input  [7:0] io_insVertical_1_33,
  input  [7:0] io_insVertical_1_34,
  input  [7:0] io_insVertical_1_35,
  input  [7:0] io_insVertical_1_36,
  input  [7:0] io_insVertical_1_37,
  input  [7:0] io_insVertical_1_38,
  input  [7:0] io_insVertical_1_39,
  input  [7:0] io_insVertical_1_40,
  input  [7:0] io_insVertical_1_41,
  input  [7:0] io_insVertical_1_42,
  input  [7:0] io_insVertical_1_43,
  input  [7:0] io_insVertical_1_44,
  input  [7:0] io_insVertical_1_45,
  input  [7:0] io_insVertical_1_46,
  input  [7:0] io_insVertical_1_47,
  input  [7:0] io_insVertical_1_48,
  input  [7:0] io_insVertical_1_49,
  input  [7:0] io_insVertical_1_50,
  input  [7:0] io_insVertical_1_51,
  input  [7:0] io_insVertical_1_52,
  input  [7:0] io_insVertical_1_53,
  input  [7:0] io_insVertical_1_54,
  input  [7:0] io_insVertical_1_55,
  input  [7:0] io_insVertical_1_56,
  input  [7:0] io_insVertical_1_57,
  input  [7:0] io_insVertical_1_58,
  input  [7:0] io_insVertical_1_59,
  input  [7:0] io_insVertical_1_60,
  input  [7:0] io_insVertical_1_61,
  input  [7:0] io_insVertical_1_62,
  input  [7:0] io_insVertical_1_63,
  input  [7:0] io_insVertical_1_64,
  input  [7:0] io_insVertical_1_65,
  input  [7:0] io_insVertical_1_66,
  input  [7:0] io_insVertical_1_67,
  input  [7:0] io_insVertical_1_68,
  input  [7:0] io_insVertical_1_69,
  input  [7:0] io_insVertical_1_70,
  input  [7:0] io_insVertical_1_71,
  input  [7:0] io_insVertical_1_72,
  input  [7:0] io_insVertical_1_73,
  input  [7:0] io_insVertical_1_74,
  input  [7:0] io_insVertical_1_75,
  input  [7:0] io_insVertical_1_76,
  input  [7:0] io_insVertical_1_77,
  input  [7:0] io_insVertical_1_78,
  input  [7:0] io_insVertical_1_79,
  input  [7:0] io_insVertical_1_80,
  input  [7:0] io_insVertical_1_81,
  input  [7:0] io_insVertical_1_82,
  input  [7:0] io_insVertical_1_83,
  input  [7:0] io_insVertical_1_84,
  input  [7:0] io_insVertical_1_85,
  input  [7:0] io_insVertical_1_86,
  input  [7:0] io_insVertical_1_87,
  input  [7:0] io_insVertical_1_88,
  input  [7:0] io_insVertical_1_89,
  input  [7:0] io_insVertical_1_90,
  input  [7:0] io_insVertical_1_91,
  input  [7:0] io_insVertical_1_92,
  input  [7:0] io_insVertical_1_93,
  input  [7:0] io_insVertical_1_94,
  input  [7:0] io_insVertical_1_95,
  input  [7:0] io_insVertical_1_96,
  input  [7:0] io_insVertical_1_97,
  input  [7:0] io_insVertical_1_98,
  input  [7:0] io_insVertical_1_99,
  input  [7:0] io_insVertical_1_100,
  input  [7:0] io_insVertical_1_101,
  input  [7:0] io_insVertical_1_102,
  input  [7:0] io_insVertical_1_103,
  input  [7:0] io_insVertical_1_104,
  input  [7:0] io_insVertical_1_105,
  input  [7:0] io_insVertical_1_106,
  input  [7:0] io_insVertical_1_107,
  input  [7:0] io_insVertical_1_108,
  input  [7:0] io_insVertical_1_109,
  input  [7:0] io_insVertical_1_110,
  input  [7:0] io_insVertical_1_111,
  input  [7:0] io_insVertical_1_112,
  input  [7:0] io_insVertical_1_113,
  input  [7:0] io_insVertical_1_114,
  input  [7:0] io_insVertical_1_115,
  input  [7:0] io_insVertical_1_116,
  input  [7:0] io_insVertical_1_117,
  input  [7:0] io_insVertical_1_118,
  input  [7:0] io_insVertical_1_119,
  input  [7:0] io_insVertical_1_120,
  input  [7:0] io_insVertical_1_121,
  input  [7:0] io_insVertical_1_122,
  input  [7:0] io_insVertical_1_123,
  input  [7:0] io_insVertical_1_124,
  input  [7:0] io_insVertical_1_125,
  input  [7:0] io_insVertical_1_126,
  input  [7:0] io_insVertical_1_127,
  input  [7:0] io_insVertical_1_128,
  input  [7:0] io_insVertical_1_129,
  input  [7:0] io_insVertical_1_130,
  input  [7:0] io_insVertical_1_131,
  input  [7:0] io_insVertical_1_132,
  input  [7:0] io_insVertical_1_133,
  input  [7:0] io_insVertical_1_134,
  input  [7:0] io_insVertical_1_135,
  input  [7:0] io_insVertical_1_136,
  input  [7:0] io_insVertical_1_137,
  input  [7:0] io_insVertical_1_138,
  input  [7:0] io_insVertical_1_139,
  input  [7:0] io_insVertical_1_140,
  input  [7:0] io_insVertical_1_141,
  input  [7:0] io_insVertical_1_142,
  input  [7:0] io_insVertical_1_143,
  input  [7:0] io_insVertical_1_144,
  input  [7:0] io_insVertical_1_145,
  input  [7:0] io_insVertical_1_146,
  input  [7:0] io_insVertical_1_147,
  input  [7:0] io_insVertical_1_148,
  input  [7:0] io_insVertical_1_149,
  input  [7:0] io_insVertical_1_150,
  input  [7:0] io_insVertical_1_151,
  input  [7:0] io_insVertical_1_152,
  input  [7:0] io_insVertical_1_153,
  input  [7:0] io_insVertical_1_154,
  input  [7:0] io_insVertical_1_155,
  input  [7:0] io_insVertical_1_156,
  input  [7:0] io_insVertical_1_157,
  input  [7:0] io_insVertical_1_158,
  input  [7:0] io_insVertical_1_159,
  input  [7:0] io_insVertical_1_160,
  input  [7:0] io_insVertical_1_161,
  input  [7:0] io_insVertical_1_162,
  input  [7:0] io_insVertical_1_163,
  input  [7:0] io_insVertical_1_164,
  input  [7:0] io_insVertical_1_165,
  input  [7:0] io_insVertical_1_166,
  input  [7:0] io_insVertical_1_167,
  input  [7:0] io_insVertical_1_168,
  input  [7:0] io_insVertical_1_169,
  input  [7:0] io_insVertical_1_170,
  input  [7:0] io_insVertical_1_171,
  input  [7:0] io_insVertical_1_172,
  input  [7:0] io_insVertical_1_173,
  input  [7:0] io_insVertical_1_174,
  input  [7:0] io_insVertical_1_175,
  input  [7:0] io_insVertical_1_176,
  input  [7:0] io_insVertical_1_177,
  input  [7:0] io_insVertical_1_178,
  input  [7:0] io_insVertical_1_179,
  input  [7:0] io_insVertical_1_180,
  input  [7:0] io_insVertical_1_181,
  input  [7:0] io_insVertical_1_182,
  input  [7:0] io_insVertical_1_183,
  input  [7:0] io_insVertical_1_184,
  input  [7:0] io_insVertical_1_185,
  input  [7:0] io_insVertical_1_186,
  input  [7:0] io_insVertical_1_187,
  input  [7:0] io_insVertical_1_188,
  input  [7:0] io_insVertical_1_189,
  input  [7:0] io_insVertical_1_190,
  input  [7:0] io_insVertical_1_191,
  input  [7:0] io_insVertical_1_192,
  input  [7:0] io_insVertical_1_193,
  input  [7:0] io_insVertical_1_194,
  input  [7:0] io_insVertical_1_195,
  input  [7:0] io_insVertical_1_196,
  input  [7:0] io_insVertical_1_197,
  input  [7:0] io_insVertical_1_198,
  input  [7:0] io_insVertical_1_199,
  input  [7:0] io_insVertical_1_200,
  input  [7:0] io_insVertical_1_201,
  input  [7:0] io_insVertical_1_202,
  input  [7:0] io_insVertical_1_203,
  input  [7:0] io_insVertical_1_204,
  input  [7:0] io_insVertical_1_205,
  input  [7:0] io_insVertical_1_206,
  input  [7:0] io_insVertical_1_207,
  input  [7:0] io_insVertical_1_208,
  input  [7:0] io_insVertical_1_209,
  input  [7:0] io_insVertical_1_210,
  input  [7:0] io_insVertical_1_211,
  input  [7:0] io_insVertical_1_212,
  input  [7:0] io_insVertical_1_213,
  input  [7:0] io_insVertical_1_214,
  input  [7:0] io_insVertical_1_215,
  input  [7:0] io_insVertical_1_216,
  input  [7:0] io_insVertical_1_217,
  input  [7:0] io_insVertical_1_218,
  input  [7:0] io_insVertical_1_219,
  input  [7:0] io_insVertical_1_220,
  input  [7:0] io_insVertical_1_221,
  input  [7:0] io_insVertical_1_222,
  input  [7:0] io_insVertical_1_223,
  input  [7:0] io_insVertical_1_224,
  input  [7:0] io_insVertical_1_225,
  input  [7:0] io_insVertical_1_226,
  input  [7:0] io_insVertical_1_227,
  input  [7:0] io_insVertical_1_228,
  input  [7:0] io_insVertical_1_229,
  input  [7:0] io_insVertical_1_230,
  input  [7:0] io_insVertical_1_231,
  input  [7:0] io_insVertical_1_232,
  input  [7:0] io_insVertical_1_233,
  input  [7:0] io_insVertical_1_234,
  input  [7:0] io_insVertical_1_235,
  input  [7:0] io_insVertical_1_236,
  input  [7:0] io_insVertical_1_237,
  input  [7:0] io_insVertical_1_238,
  input  [7:0] io_insVertical_1_239,
  input  [7:0] io_insVertical_1_240,
  input  [7:0] io_insVertical_1_241,
  input  [7:0] io_insVertical_1_242,
  input  [7:0] io_insVertical_1_243,
  input  [7:0] io_insVertical_1_244,
  input  [7:0] io_insVertical_1_245,
  input  [7:0] io_insVertical_1_246,
  input  [7:0] io_insVertical_1_247,
  input  [7:0] io_insVertical_1_248,
  input  [7:0] io_insVertical_1_249,
  input  [7:0] io_insVertical_1_250,
  input  [7:0] io_insVertical_1_251,
  input  [7:0] io_insVertical_1_252,
  input  [7:0] io_insVertical_1_253,
  input  [7:0] io_insVertical_1_254,
  input  [7:0] io_insVertical_1_255,
  output [7:0] io_outsVertical_0_0,
  output [7:0] io_outsVertical_0_1,
  output [7:0] io_outsVertical_0_2,
  output [7:0] io_outsVertical_0_3,
  output [7:0] io_outsVertical_0_4,
  output [7:0] io_outsVertical_0_5,
  output [7:0] io_outsVertical_0_6,
  output [7:0] io_outsVertical_0_7,
  output [7:0] io_outsVertical_0_8,
  output [7:0] io_outsVertical_0_9,
  output [7:0] io_outsVertical_0_10,
  output [7:0] io_outsVertical_0_11,
  output [7:0] io_outsVertical_0_12,
  output [7:0] io_outsVertical_0_13,
  output [7:0] io_outsVertical_0_14,
  output [7:0] io_outsVertical_0_15,
  output [7:0] io_outsVertical_0_16,
  output [7:0] io_outsVertical_0_17,
  output [7:0] io_outsVertical_0_18,
  output [7:0] io_outsVertical_0_19,
  output [7:0] io_outsVertical_0_20,
  output [7:0] io_outsVertical_0_21,
  output [7:0] io_outsVertical_0_22,
  output [7:0] io_outsVertical_0_23,
  output [7:0] io_outsVertical_0_24,
  output [7:0] io_outsVertical_0_25,
  output [7:0] io_outsVertical_0_26,
  output [7:0] io_outsVertical_0_27,
  output [7:0] io_outsVertical_0_28,
  output [7:0] io_outsVertical_0_29,
  output [7:0] io_outsVertical_0_30,
  output [7:0] io_outsVertical_0_31,
  output [7:0] io_outsVertical_0_32,
  output [7:0] io_outsVertical_0_33,
  output [7:0] io_outsVertical_0_34,
  output [7:0] io_outsVertical_0_35,
  output [7:0] io_outsVertical_0_36,
  output [7:0] io_outsVertical_0_37,
  output [7:0] io_outsVertical_0_38,
  output [7:0] io_outsVertical_0_39,
  output [7:0] io_outsVertical_0_40,
  output [7:0] io_outsVertical_0_41,
  output [7:0] io_outsVertical_0_42,
  output [7:0] io_outsVertical_0_43,
  output [7:0] io_outsVertical_0_44,
  output [7:0] io_outsVertical_0_45,
  output [7:0] io_outsVertical_0_46,
  output [7:0] io_outsVertical_0_47,
  output [7:0] io_outsVertical_0_48,
  output [7:0] io_outsVertical_0_49,
  output [7:0] io_outsVertical_0_50,
  output [7:0] io_outsVertical_0_51,
  output [7:0] io_outsVertical_0_52,
  output [7:0] io_outsVertical_0_53,
  output [7:0] io_outsVertical_0_54,
  output [7:0] io_outsVertical_0_55,
  output [7:0] io_outsVertical_0_56,
  output [7:0] io_outsVertical_0_57,
  output [7:0] io_outsVertical_0_58,
  output [7:0] io_outsVertical_0_59,
  output [7:0] io_outsVertical_0_60,
  output [7:0] io_outsVertical_0_61,
  output [7:0] io_outsVertical_0_62,
  output [7:0] io_outsVertical_0_63,
  output [7:0] io_outsVertical_0_64,
  output [7:0] io_outsVertical_0_65,
  output [7:0] io_outsVertical_0_66,
  output [7:0] io_outsVertical_0_67,
  output [7:0] io_outsVertical_0_68,
  output [7:0] io_outsVertical_0_69,
  output [7:0] io_outsVertical_0_70,
  output [7:0] io_outsVertical_0_71,
  output [7:0] io_outsVertical_0_72,
  output [7:0] io_outsVertical_0_73,
  output [7:0] io_outsVertical_0_74,
  output [7:0] io_outsVertical_0_75,
  output [7:0] io_outsVertical_0_76,
  output [7:0] io_outsVertical_0_77,
  output [7:0] io_outsVertical_0_78,
  output [7:0] io_outsVertical_0_79,
  output [7:0] io_outsVertical_0_80,
  output [7:0] io_outsVertical_0_81,
  output [7:0] io_outsVertical_0_82,
  output [7:0] io_outsVertical_0_83,
  output [7:0] io_outsVertical_0_84,
  output [7:0] io_outsVertical_0_85,
  output [7:0] io_outsVertical_0_86,
  output [7:0] io_outsVertical_0_87,
  output [7:0] io_outsVertical_0_88,
  output [7:0] io_outsVertical_0_89,
  output [7:0] io_outsVertical_0_90,
  output [7:0] io_outsVertical_0_91,
  output [7:0] io_outsVertical_0_92,
  output [7:0] io_outsVertical_0_93,
  output [7:0] io_outsVertical_0_94,
  output [7:0] io_outsVertical_0_95,
  output [7:0] io_outsVertical_0_96,
  output [7:0] io_outsVertical_0_97,
  output [7:0] io_outsVertical_0_98,
  output [7:0] io_outsVertical_0_99,
  output [7:0] io_outsVertical_0_100,
  output [7:0] io_outsVertical_0_101,
  output [7:0] io_outsVertical_0_102,
  output [7:0] io_outsVertical_0_103,
  output [7:0] io_outsVertical_0_104,
  output [7:0] io_outsVertical_0_105,
  output [7:0] io_outsVertical_0_106,
  output [7:0] io_outsVertical_0_107,
  output [7:0] io_outsVertical_0_108,
  output [7:0] io_outsVertical_0_109,
  output [7:0] io_outsVertical_0_110,
  output [7:0] io_outsVertical_0_111,
  output [7:0] io_outsVertical_0_112,
  output [7:0] io_outsVertical_0_113,
  output [7:0] io_outsVertical_0_114,
  output [7:0] io_outsVertical_0_115,
  output [7:0] io_outsVertical_0_116,
  output [7:0] io_outsVertical_0_117,
  output [7:0] io_outsVertical_0_118,
  output [7:0] io_outsVertical_0_119,
  output [7:0] io_outsVertical_0_120,
  output [7:0] io_outsVertical_0_121,
  output [7:0] io_outsVertical_0_122,
  output [7:0] io_outsVertical_0_123,
  output [7:0] io_outsVertical_0_124,
  output [7:0] io_outsVertical_0_125,
  output [7:0] io_outsVertical_0_126,
  output [7:0] io_outsVertical_0_127,
  output [7:0] io_outsVertical_0_128,
  output [7:0] io_outsVertical_0_129,
  output [7:0] io_outsVertical_0_130,
  output [7:0] io_outsVertical_0_131,
  output [7:0] io_outsVertical_0_132,
  output [7:0] io_outsVertical_0_133,
  output [7:0] io_outsVertical_0_134,
  output [7:0] io_outsVertical_0_135,
  output [7:0] io_outsVertical_0_136,
  output [7:0] io_outsVertical_0_137,
  output [7:0] io_outsVertical_0_138,
  output [7:0] io_outsVertical_0_139,
  output [7:0] io_outsVertical_0_140,
  output [7:0] io_outsVertical_0_141,
  output [7:0] io_outsVertical_0_142,
  output [7:0] io_outsVertical_0_143,
  output [7:0] io_outsVertical_0_144,
  output [7:0] io_outsVertical_0_145,
  output [7:0] io_outsVertical_0_146,
  output [7:0] io_outsVertical_0_147,
  output [7:0] io_outsVertical_0_148,
  output [7:0] io_outsVertical_0_149,
  output [7:0] io_outsVertical_0_150,
  output [7:0] io_outsVertical_0_151,
  output [7:0] io_outsVertical_0_152,
  output [7:0] io_outsVertical_0_153,
  output [7:0] io_outsVertical_0_154,
  output [7:0] io_outsVertical_0_155,
  output [7:0] io_outsVertical_0_156,
  output [7:0] io_outsVertical_0_157,
  output [7:0] io_outsVertical_0_158,
  output [7:0] io_outsVertical_0_159,
  output [7:0] io_outsVertical_0_160,
  output [7:0] io_outsVertical_0_161,
  output [7:0] io_outsVertical_0_162,
  output [7:0] io_outsVertical_0_163,
  output [7:0] io_outsVertical_0_164,
  output [7:0] io_outsVertical_0_165,
  output [7:0] io_outsVertical_0_166,
  output [7:0] io_outsVertical_0_167,
  output [7:0] io_outsVertical_0_168,
  output [7:0] io_outsVertical_0_169,
  output [7:0] io_outsVertical_0_170,
  output [7:0] io_outsVertical_0_171,
  output [7:0] io_outsVertical_0_172,
  output [7:0] io_outsVertical_0_173,
  output [7:0] io_outsVertical_0_174,
  output [7:0] io_outsVertical_0_175,
  output [7:0] io_outsVertical_0_176,
  output [7:0] io_outsVertical_0_177,
  output [7:0] io_outsVertical_0_178,
  output [7:0] io_outsVertical_0_179,
  output [7:0] io_outsVertical_0_180,
  output [7:0] io_outsVertical_0_181,
  output [7:0] io_outsVertical_0_182,
  output [7:0] io_outsVertical_0_183,
  output [7:0] io_outsVertical_0_184,
  output [7:0] io_outsVertical_0_185,
  output [7:0] io_outsVertical_0_186,
  output [7:0] io_outsVertical_0_187,
  output [7:0] io_outsVertical_0_188,
  output [7:0] io_outsVertical_0_189,
  output [7:0] io_outsVertical_0_190,
  output [7:0] io_outsVertical_0_191,
  output [7:0] io_outsVertical_0_192,
  output [7:0] io_outsVertical_0_193,
  output [7:0] io_outsVertical_0_194,
  output [7:0] io_outsVertical_0_195,
  output [7:0] io_outsVertical_0_196,
  output [7:0] io_outsVertical_0_197,
  output [7:0] io_outsVertical_0_198,
  output [7:0] io_outsVertical_0_199,
  output [7:0] io_outsVertical_0_200,
  output [7:0] io_outsVertical_0_201,
  output [7:0] io_outsVertical_0_202,
  output [7:0] io_outsVertical_0_203,
  output [7:0] io_outsVertical_0_204,
  output [7:0] io_outsVertical_0_205,
  output [7:0] io_outsVertical_0_206,
  output [7:0] io_outsVertical_0_207,
  output [7:0] io_outsVertical_0_208,
  output [7:0] io_outsVertical_0_209,
  output [7:0] io_outsVertical_0_210,
  output [7:0] io_outsVertical_0_211,
  output [7:0] io_outsVertical_0_212,
  output [7:0] io_outsVertical_0_213,
  output [7:0] io_outsVertical_0_214,
  output [7:0] io_outsVertical_0_215,
  output [7:0] io_outsVertical_0_216,
  output [7:0] io_outsVertical_0_217,
  output [7:0] io_outsVertical_0_218,
  output [7:0] io_outsVertical_0_219,
  output [7:0] io_outsVertical_0_220,
  output [7:0] io_outsVertical_0_221,
  output [7:0] io_outsVertical_0_222,
  output [7:0] io_outsVertical_0_223,
  output [7:0] io_outsVertical_0_224,
  output [7:0] io_outsVertical_0_225,
  output [7:0] io_outsVertical_0_226,
  output [7:0] io_outsVertical_0_227,
  output [7:0] io_outsVertical_0_228,
  output [7:0] io_outsVertical_0_229,
  output [7:0] io_outsVertical_0_230,
  output [7:0] io_outsVertical_0_231,
  output [7:0] io_outsVertical_0_232,
  output [7:0] io_outsVertical_0_233,
  output [7:0] io_outsVertical_0_234,
  output [7:0] io_outsVertical_0_235,
  output [7:0] io_outsVertical_0_236,
  output [7:0] io_outsVertical_0_237,
  output [7:0] io_outsVertical_0_238,
  output [7:0] io_outsVertical_0_239,
  output [7:0] io_outsVertical_0_240,
  output [7:0] io_outsVertical_0_241,
  output [7:0] io_outsVertical_0_242,
  output [7:0] io_outsVertical_0_243,
  output [7:0] io_outsVertical_0_244,
  output [7:0] io_outsVertical_0_245,
  output [7:0] io_outsVertical_0_246,
  output [7:0] io_outsVertical_0_247,
  output [7:0] io_outsVertical_0_248,
  output [7:0] io_outsVertical_0_249,
  output [7:0] io_outsVertical_0_250,
  output [7:0] io_outsVertical_0_251,
  output [7:0] io_outsVertical_0_252,
  output [7:0] io_outsVertical_0_253,
  output [7:0] io_outsVertical_0_254,
  output [7:0] io_outsVertical_0_255,
  output [7:0] io_outsVertical_1_0,
  output [7:0] io_outsVertical_1_1,
  output [7:0] io_outsVertical_1_2,
  output [7:0] io_outsVertical_1_3,
  output [7:0] io_outsVertical_1_4,
  output [7:0] io_outsVertical_1_5,
  output [7:0] io_outsVertical_1_6,
  output [7:0] io_outsVertical_1_7,
  output [7:0] io_outsVertical_1_8,
  output [7:0] io_outsVertical_1_9,
  output [7:0] io_outsVertical_1_10,
  output [7:0] io_outsVertical_1_11,
  output [7:0] io_outsVertical_1_12,
  output [7:0] io_outsVertical_1_13,
  output [7:0] io_outsVertical_1_14,
  output [7:0] io_outsVertical_1_15,
  output [7:0] io_outsVertical_1_16,
  output [7:0] io_outsVertical_1_17,
  output [7:0] io_outsVertical_1_18,
  output [7:0] io_outsVertical_1_19,
  output [7:0] io_outsVertical_1_20,
  output [7:0] io_outsVertical_1_21,
  output [7:0] io_outsVertical_1_22,
  output [7:0] io_outsVertical_1_23,
  output [7:0] io_outsVertical_1_24,
  output [7:0] io_outsVertical_1_25,
  output [7:0] io_outsVertical_1_26,
  output [7:0] io_outsVertical_1_27,
  output [7:0] io_outsVertical_1_28,
  output [7:0] io_outsVertical_1_29,
  output [7:0] io_outsVertical_1_30,
  output [7:0] io_outsVertical_1_31,
  output [7:0] io_outsVertical_1_32,
  output [7:0] io_outsVertical_1_33,
  output [7:0] io_outsVertical_1_34,
  output [7:0] io_outsVertical_1_35,
  output [7:0] io_outsVertical_1_36,
  output [7:0] io_outsVertical_1_37,
  output [7:0] io_outsVertical_1_38,
  output [7:0] io_outsVertical_1_39,
  output [7:0] io_outsVertical_1_40,
  output [7:0] io_outsVertical_1_41,
  output [7:0] io_outsVertical_1_42,
  output [7:0] io_outsVertical_1_43,
  output [7:0] io_outsVertical_1_44,
  output [7:0] io_outsVertical_1_45,
  output [7:0] io_outsVertical_1_46,
  output [7:0] io_outsVertical_1_47,
  output [7:0] io_outsVertical_1_48,
  output [7:0] io_outsVertical_1_49,
  output [7:0] io_outsVertical_1_50,
  output [7:0] io_outsVertical_1_51,
  output [7:0] io_outsVertical_1_52,
  output [7:0] io_outsVertical_1_53,
  output [7:0] io_outsVertical_1_54,
  output [7:0] io_outsVertical_1_55,
  output [7:0] io_outsVertical_1_56,
  output [7:0] io_outsVertical_1_57,
  output [7:0] io_outsVertical_1_58,
  output [7:0] io_outsVertical_1_59,
  output [7:0] io_outsVertical_1_60,
  output [7:0] io_outsVertical_1_61,
  output [7:0] io_outsVertical_1_62,
  output [7:0] io_outsVertical_1_63,
  output [7:0] io_outsVertical_1_64,
  output [7:0] io_outsVertical_1_65,
  output [7:0] io_outsVertical_1_66,
  output [7:0] io_outsVertical_1_67,
  output [7:0] io_outsVertical_1_68,
  output [7:0] io_outsVertical_1_69,
  output [7:0] io_outsVertical_1_70,
  output [7:0] io_outsVertical_1_71,
  output [7:0] io_outsVertical_1_72,
  output [7:0] io_outsVertical_1_73,
  output [7:0] io_outsVertical_1_74,
  output [7:0] io_outsVertical_1_75,
  output [7:0] io_outsVertical_1_76,
  output [7:0] io_outsVertical_1_77,
  output [7:0] io_outsVertical_1_78,
  output [7:0] io_outsVertical_1_79,
  output [7:0] io_outsVertical_1_80,
  output [7:0] io_outsVertical_1_81,
  output [7:0] io_outsVertical_1_82,
  output [7:0] io_outsVertical_1_83,
  output [7:0] io_outsVertical_1_84,
  output [7:0] io_outsVertical_1_85,
  output [7:0] io_outsVertical_1_86,
  output [7:0] io_outsVertical_1_87,
  output [7:0] io_outsVertical_1_88,
  output [7:0] io_outsVertical_1_89,
  output [7:0] io_outsVertical_1_90,
  output [7:0] io_outsVertical_1_91,
  output [7:0] io_outsVertical_1_92,
  output [7:0] io_outsVertical_1_93,
  output [7:0] io_outsVertical_1_94,
  output [7:0] io_outsVertical_1_95,
  output [7:0] io_outsVertical_1_96,
  output [7:0] io_outsVertical_1_97,
  output [7:0] io_outsVertical_1_98,
  output [7:0] io_outsVertical_1_99,
  output [7:0] io_outsVertical_1_100,
  output [7:0] io_outsVertical_1_101,
  output [7:0] io_outsVertical_1_102,
  output [7:0] io_outsVertical_1_103,
  output [7:0] io_outsVertical_1_104,
  output [7:0] io_outsVertical_1_105,
  output [7:0] io_outsVertical_1_106,
  output [7:0] io_outsVertical_1_107,
  output [7:0] io_outsVertical_1_108,
  output [7:0] io_outsVertical_1_109,
  output [7:0] io_outsVertical_1_110,
  output [7:0] io_outsVertical_1_111,
  output [7:0] io_outsVertical_1_112,
  output [7:0] io_outsVertical_1_113,
  output [7:0] io_outsVertical_1_114,
  output [7:0] io_outsVertical_1_115,
  output [7:0] io_outsVertical_1_116,
  output [7:0] io_outsVertical_1_117,
  output [7:0] io_outsVertical_1_118,
  output [7:0] io_outsVertical_1_119,
  output [7:0] io_outsVertical_1_120,
  output [7:0] io_outsVertical_1_121,
  output [7:0] io_outsVertical_1_122,
  output [7:0] io_outsVertical_1_123,
  output [7:0] io_outsVertical_1_124,
  output [7:0] io_outsVertical_1_125,
  output [7:0] io_outsVertical_1_126,
  output [7:0] io_outsVertical_1_127,
  output [7:0] io_outsVertical_1_128,
  output [7:0] io_outsVertical_1_129,
  output [7:0] io_outsVertical_1_130,
  output [7:0] io_outsVertical_1_131,
  output [7:0] io_outsVertical_1_132,
  output [7:0] io_outsVertical_1_133,
  output [7:0] io_outsVertical_1_134,
  output [7:0] io_outsVertical_1_135,
  output [7:0] io_outsVertical_1_136,
  output [7:0] io_outsVertical_1_137,
  output [7:0] io_outsVertical_1_138,
  output [7:0] io_outsVertical_1_139,
  output [7:0] io_outsVertical_1_140,
  output [7:0] io_outsVertical_1_141,
  output [7:0] io_outsVertical_1_142,
  output [7:0] io_outsVertical_1_143,
  output [7:0] io_outsVertical_1_144,
  output [7:0] io_outsVertical_1_145,
  output [7:0] io_outsVertical_1_146,
  output [7:0] io_outsVertical_1_147,
  output [7:0] io_outsVertical_1_148,
  output [7:0] io_outsVertical_1_149,
  output [7:0] io_outsVertical_1_150,
  output [7:0] io_outsVertical_1_151,
  output [7:0] io_outsVertical_1_152,
  output [7:0] io_outsVertical_1_153,
  output [7:0] io_outsVertical_1_154,
  output [7:0] io_outsVertical_1_155,
  output [7:0] io_outsVertical_1_156,
  output [7:0] io_outsVertical_1_157,
  output [7:0] io_outsVertical_1_158,
  output [7:0] io_outsVertical_1_159,
  output [7:0] io_outsVertical_1_160,
  output [7:0] io_outsVertical_1_161,
  output [7:0] io_outsVertical_1_162,
  output [7:0] io_outsVertical_1_163,
  output [7:0] io_outsVertical_1_164,
  output [7:0] io_outsVertical_1_165,
  output [7:0] io_outsVertical_1_166,
  output [7:0] io_outsVertical_1_167,
  output [7:0] io_outsVertical_1_168,
  output [7:0] io_outsVertical_1_169,
  output [7:0] io_outsVertical_1_170,
  output [7:0] io_outsVertical_1_171,
  output [7:0] io_outsVertical_1_172,
  output [7:0] io_outsVertical_1_173,
  output [7:0] io_outsVertical_1_174,
  output [7:0] io_outsVertical_1_175,
  output [7:0] io_outsVertical_1_176,
  output [7:0] io_outsVertical_1_177,
  output [7:0] io_outsVertical_1_178,
  output [7:0] io_outsVertical_1_179,
  output [7:0] io_outsVertical_1_180,
  output [7:0] io_outsVertical_1_181,
  output [7:0] io_outsVertical_1_182,
  output [7:0] io_outsVertical_1_183,
  output [7:0] io_outsVertical_1_184,
  output [7:0] io_outsVertical_1_185,
  output [7:0] io_outsVertical_1_186,
  output [7:0] io_outsVertical_1_187,
  output [7:0] io_outsVertical_1_188,
  output [7:0] io_outsVertical_1_189,
  output [7:0] io_outsVertical_1_190,
  output [7:0] io_outsVertical_1_191,
  output [7:0] io_outsVertical_1_192,
  output [7:0] io_outsVertical_1_193,
  output [7:0] io_outsVertical_1_194,
  output [7:0] io_outsVertical_1_195,
  output [7:0] io_outsVertical_1_196,
  output [7:0] io_outsVertical_1_197,
  output [7:0] io_outsVertical_1_198,
  output [7:0] io_outsVertical_1_199,
  output [7:0] io_outsVertical_1_200,
  output [7:0] io_outsVertical_1_201,
  output [7:0] io_outsVertical_1_202,
  output [7:0] io_outsVertical_1_203,
  output [7:0] io_outsVertical_1_204,
  output [7:0] io_outsVertical_1_205,
  output [7:0] io_outsVertical_1_206,
  output [7:0] io_outsVertical_1_207,
  output [7:0] io_outsVertical_1_208,
  output [7:0] io_outsVertical_1_209,
  output [7:0] io_outsVertical_1_210,
  output [7:0] io_outsVertical_1_211,
  output [7:0] io_outsVertical_1_212,
  output [7:0] io_outsVertical_1_213,
  output [7:0] io_outsVertical_1_214,
  output [7:0] io_outsVertical_1_215,
  output [7:0] io_outsVertical_1_216,
  output [7:0] io_outsVertical_1_217,
  output [7:0] io_outsVertical_1_218,
  output [7:0] io_outsVertical_1_219,
  output [7:0] io_outsVertical_1_220,
  output [7:0] io_outsVertical_1_221,
  output [7:0] io_outsVertical_1_222,
  output [7:0] io_outsVertical_1_223,
  output [7:0] io_outsVertical_1_224,
  output [7:0] io_outsVertical_1_225,
  output [7:0] io_outsVertical_1_226,
  output [7:0] io_outsVertical_1_227,
  output [7:0] io_outsVertical_1_228,
  output [7:0] io_outsVertical_1_229,
  output [7:0] io_outsVertical_1_230,
  output [7:0] io_outsVertical_1_231,
  output [7:0] io_outsVertical_1_232,
  output [7:0] io_outsVertical_1_233,
  output [7:0] io_outsVertical_1_234,
  output [7:0] io_outsVertical_1_235,
  output [7:0] io_outsVertical_1_236,
  output [7:0] io_outsVertical_1_237,
  output [7:0] io_outsVertical_1_238,
  output [7:0] io_outsVertical_1_239,
  output [7:0] io_outsVertical_1_240,
  output [7:0] io_outsVertical_1_241,
  output [7:0] io_outsVertical_1_242,
  output [7:0] io_outsVertical_1_243,
  output [7:0] io_outsVertical_1_244,
  output [7:0] io_outsVertical_1_245,
  output [7:0] io_outsVertical_1_246,
  output [7:0] io_outsVertical_1_247,
  output [7:0] io_outsVertical_1_248,
  output [7:0] io_outsVertical_1_249,
  output [7:0] io_outsVertical_1_250,
  output [7:0] io_outsVertical_1_251,
  output [7:0] io_outsVertical_1_252,
  output [7:0] io_outsVertical_1_253,
  output [7:0] io_outsVertical_1_254,
  output [7:0] io_outsVertical_1_255,
  output       io_lsbs_0,
  output       io_lsbs_1,
  output       io_lsbs_2,
  output       io_lsbs_3,
  output       io_lsbs_4,
  output       io_lsbs_5,
  output       io_lsbs_6,
  output       io_lsbs_7,
  output       io_lsbs_8,
  output       io_lsbs_9,
  output       io_lsbs_10,
  output       io_lsbs_11,
  output       io_lsbs_12,
  output       io_lsbs_13,
  output       io_lsbs_14,
  output       io_lsbs_15,
  output       io_lsbs_16,
  output       io_lsbs_17,
  output       io_lsbs_18,
  output       io_lsbs_19,
  output       io_lsbs_20,
  output       io_lsbs_21,
  output       io_lsbs_22,
  output       io_lsbs_23,
  output       io_lsbs_24,
  output       io_lsbs_25,
  output       io_lsbs_26,
  output       io_lsbs_27,
  output       io_lsbs_28,
  output       io_lsbs_29,
  output       io_lsbs_30,
  output       io_lsbs_31,
  output       io_lsbs_32,
  output       io_lsbs_33,
  output       io_lsbs_34,
  output       io_lsbs_35,
  output       io_lsbs_36,
  output       io_lsbs_37,
  output       io_lsbs_38,
  output       io_lsbs_39,
  output       io_lsbs_40,
  output       io_lsbs_41,
  output       io_lsbs_42,
  output       io_lsbs_43,
  output       io_lsbs_44,
  output       io_lsbs_45,
  output       io_lsbs_46,
  output       io_lsbs_47,
  output       io_lsbs_48,
  output       io_lsbs_49,
  output       io_lsbs_50,
  output       io_lsbs_51,
  output       io_lsbs_52,
  output       io_lsbs_53,
  output       io_lsbs_54,
  output       io_lsbs_55,
  output       io_lsbs_56,
  output       io_lsbs_57,
  output       io_lsbs_58,
  output       io_lsbs_59,
  output       io_lsbs_60,
  output       io_lsbs_61,
  output       io_lsbs_62,
  output       io_lsbs_63,
  output       io_lsbs_64,
  output       io_lsbs_65,
  output       io_lsbs_66,
  output       io_lsbs_67,
  output       io_lsbs_68,
  output       io_lsbs_69,
  output       io_lsbs_70,
  output       io_lsbs_71,
  output       io_lsbs_72,
  output       io_lsbs_73,
  output       io_lsbs_74,
  output       io_lsbs_75,
  output       io_lsbs_76,
  output       io_lsbs_77,
  output       io_lsbs_78,
  output       io_lsbs_79,
  output       io_lsbs_80,
  output       io_lsbs_81,
  output       io_lsbs_82,
  output       io_lsbs_83,
  output       io_lsbs_84,
  output       io_lsbs_85,
  output       io_lsbs_86,
  output       io_lsbs_87,
  output       io_lsbs_88,
  output       io_lsbs_89,
  output       io_lsbs_90,
  output       io_lsbs_91,
  output       io_lsbs_92,
  output       io_lsbs_93,
  output       io_lsbs_94,
  output       io_lsbs_95,
  output       io_lsbs_96,
  output       io_lsbs_97,
  output       io_lsbs_98,
  output       io_lsbs_99,
  output       io_lsbs_100,
  output       io_lsbs_101,
  output       io_lsbs_102,
  output       io_lsbs_103,
  output       io_lsbs_104,
  output       io_lsbs_105,
  output       io_lsbs_106,
  output       io_lsbs_107,
  output       io_lsbs_108,
  output       io_lsbs_109,
  output       io_lsbs_110,
  output       io_lsbs_111,
  output       io_lsbs_112,
  output       io_lsbs_113,
  output       io_lsbs_114,
  output       io_lsbs_115,
  output       io_lsbs_116,
  output       io_lsbs_117,
  output       io_lsbs_118,
  output       io_lsbs_119,
  output       io_lsbs_120,
  output       io_lsbs_121,
  output       io_lsbs_122,
  output       io_lsbs_123,
  output       io_lsbs_124,
  output       io_lsbs_125,
  output       io_lsbs_126,
  output       io_lsbs_127,
  output       io_lsbs_128,
  output       io_lsbs_129,
  output       io_lsbs_130,
  output       io_lsbs_131,
  output       io_lsbs_132,
  output       io_lsbs_133,
  output       io_lsbs_134,
  output       io_lsbs_135,
  output       io_lsbs_136,
  output       io_lsbs_137,
  output       io_lsbs_138,
  output       io_lsbs_139,
  output       io_lsbs_140,
  output       io_lsbs_141,
  output       io_lsbs_142,
  output       io_lsbs_143,
  output       io_lsbs_144,
  output       io_lsbs_145,
  output       io_lsbs_146,
  output       io_lsbs_147,
  output       io_lsbs_148,
  output       io_lsbs_149,
  output       io_lsbs_150,
  output       io_lsbs_151,
  output       io_lsbs_152,
  output       io_lsbs_153,
  output       io_lsbs_154,
  output       io_lsbs_155,
  output       io_lsbs_156,
  output       io_lsbs_157,
  output       io_lsbs_158,
  output       io_lsbs_159,
  output       io_lsbs_160,
  output       io_lsbs_161,
  output       io_lsbs_162,
  output       io_lsbs_163,
  output       io_lsbs_164,
  output       io_lsbs_165,
  output       io_lsbs_166,
  output       io_lsbs_167,
  output       io_lsbs_168,
  output       io_lsbs_169,
  output       io_lsbs_170,
  output       io_lsbs_171,
  output       io_lsbs_172,
  output       io_lsbs_173,
  output       io_lsbs_174,
  output       io_lsbs_175,
  output       io_lsbs_176,
  output       io_lsbs_177,
  output       io_lsbs_178,
  output       io_lsbs_179,
  output       io_lsbs_180,
  output       io_lsbs_181,
  output       io_lsbs_182,
  output       io_lsbs_183,
  output       io_lsbs_184,
  output       io_lsbs_185,
  output       io_lsbs_186,
  output       io_lsbs_187,
  output       io_lsbs_188,
  output       io_lsbs_189,
  output       io_lsbs_190,
  output       io_lsbs_191,
  output       io_lsbs_192,
  output       io_lsbs_193,
  output       io_lsbs_194,
  output       io_lsbs_195,
  output       io_lsbs_196,
  output       io_lsbs_197,
  output       io_lsbs_198,
  output       io_lsbs_199,
  output       io_lsbs_200,
  output       io_lsbs_201,
  output       io_lsbs_202,
  output       io_lsbs_203,
  output       io_lsbs_204,
  output       io_lsbs_205,
  output       io_lsbs_206,
  output       io_lsbs_207,
  output       io_lsbs_208,
  output       io_lsbs_209,
  output       io_lsbs_210,
  output       io_lsbs_211,
  output       io_lsbs_212,
  output       io_lsbs_213,
  output       io_lsbs_214,
  output       io_lsbs_215,
  output       io_lsbs_216,
  output       io_lsbs_217,
  output       io_lsbs_218,
  output       io_lsbs_219,
  output       io_lsbs_220,
  output       io_lsbs_221,
  output       io_lsbs_222,
  output       io_lsbs_223,
  output       io_lsbs_224,
  output       io_lsbs_225,
  output       io_lsbs_226,
  output       io_lsbs_227,
  output       io_lsbs_228,
  output       io_lsbs_229,
  output       io_lsbs_230,
  output       io_lsbs_231,
  output       io_lsbs_232,
  output       io_lsbs_233,
  output       io_lsbs_234,
  output       io_lsbs_235,
  output       io_lsbs_236,
  output       io_lsbs_237,
  output       io_lsbs_238,
  output       io_lsbs_239,
  output       io_lsbs_240,
  output       io_lsbs_241,
  output       io_lsbs_242,
  output       io_lsbs_243,
  output       io_lsbs_244,
  output       io_lsbs_245,
  output       io_lsbs_246,
  output       io_lsbs_247,
  output       io_lsbs_248,
  output       io_lsbs_249,
  output       io_lsbs_250,
  output       io_lsbs_251,
  output       io_lsbs_252,
  output       io_lsbs_253,
  output       io_lsbs_254,
  output       io_lsbs_255
);
  wire  ces_0_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_1_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_1_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_1_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_1_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_1_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_1_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_1_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_1_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_2_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_2_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_2_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_2_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_2_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_2_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_2_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_2_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_3_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_3_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_3_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_3_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_3_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_3_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_3_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_3_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_4_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_4_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_4_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_4_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_4_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_4_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_4_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_4_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_5_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_5_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_5_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_5_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_5_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_5_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_5_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_5_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_6_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_6_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_6_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_6_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_6_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_6_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_6_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_6_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_7_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_7_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_7_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_7_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_7_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_7_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_7_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_7_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_8_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_8_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_8_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_8_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_8_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_8_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_8_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_8_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_9_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_9_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_9_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_9_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_9_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_9_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_9_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_9_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_10_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_10_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_10_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_10_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_10_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_10_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_10_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_10_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_11_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_11_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_11_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_11_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_11_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_11_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_11_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_11_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_12_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_12_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_12_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_12_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_12_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_12_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_12_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_12_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_13_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_13_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_13_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_13_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_13_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_13_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_13_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_13_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_14_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_14_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_14_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_14_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_14_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_14_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_14_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_14_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_15_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_15_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_15_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_15_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_15_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_15_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_15_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_15_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_16_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_16_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_16_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_16_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_16_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_16_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_16_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_16_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_17_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_17_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_17_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_17_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_17_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_17_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_17_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_17_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_18_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_18_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_18_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_18_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_18_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_18_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_18_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_18_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_19_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_19_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_19_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_19_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_19_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_19_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_19_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_19_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_20_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_20_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_20_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_20_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_20_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_20_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_20_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_20_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_21_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_21_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_21_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_21_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_21_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_21_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_21_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_21_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_22_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_22_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_22_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_22_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_22_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_22_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_22_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_22_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_23_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_23_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_23_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_23_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_23_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_23_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_23_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_23_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_24_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_24_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_24_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_24_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_24_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_24_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_24_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_24_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_25_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_25_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_25_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_25_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_25_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_25_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_25_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_25_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_26_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_26_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_26_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_26_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_26_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_26_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_26_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_26_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_27_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_27_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_27_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_27_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_27_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_27_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_27_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_27_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_28_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_28_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_28_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_28_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_28_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_28_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_28_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_28_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_29_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_29_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_29_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_29_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_29_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_29_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_29_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_29_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_30_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_30_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_30_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_30_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_30_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_30_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_30_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_30_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_31_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_31_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_31_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_31_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_31_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_31_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_31_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_31_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_32_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_32_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_32_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_32_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_32_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_32_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_32_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_32_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_32_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_33_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_33_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_33_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_33_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_33_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_33_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_33_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_33_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_33_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_34_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_34_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_34_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_34_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_34_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_34_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_34_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_34_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_34_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_35_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_35_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_35_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_35_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_35_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_35_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_35_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_35_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_35_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_36_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_36_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_36_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_36_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_36_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_36_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_36_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_36_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_36_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_37_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_37_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_37_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_37_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_37_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_37_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_37_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_37_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_37_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_38_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_38_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_38_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_38_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_38_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_38_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_38_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_38_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_38_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_39_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_39_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_39_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_39_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_39_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_39_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_39_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_39_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_39_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_40_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_40_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_40_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_40_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_40_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_40_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_40_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_40_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_40_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_41_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_41_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_41_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_41_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_41_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_41_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_41_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_41_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_41_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_42_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_42_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_42_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_42_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_42_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_42_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_42_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_42_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_42_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_43_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_43_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_43_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_43_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_43_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_43_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_43_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_43_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_43_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_44_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_44_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_44_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_44_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_44_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_44_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_44_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_44_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_44_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_45_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_45_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_45_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_45_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_45_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_45_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_45_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_45_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_45_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_46_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_46_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_46_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_46_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_46_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_46_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_46_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_46_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_46_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_47_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_47_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_47_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_47_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_47_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_47_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_47_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_47_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_47_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_48_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_48_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_48_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_48_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_48_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_48_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_48_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_48_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_48_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_49_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_49_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_49_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_49_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_49_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_49_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_49_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_49_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_49_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_50_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_50_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_50_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_50_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_50_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_50_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_50_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_50_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_50_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_51_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_51_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_51_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_51_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_51_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_51_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_51_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_51_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_51_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_52_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_52_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_52_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_52_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_52_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_52_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_52_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_52_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_52_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_53_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_53_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_53_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_53_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_53_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_53_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_53_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_53_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_53_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_54_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_54_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_54_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_54_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_54_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_54_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_54_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_54_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_54_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_55_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_55_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_55_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_55_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_55_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_55_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_55_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_55_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_55_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_56_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_56_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_56_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_56_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_56_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_56_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_56_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_56_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_56_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_57_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_57_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_57_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_57_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_57_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_57_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_57_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_57_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_57_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_58_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_58_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_58_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_58_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_58_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_58_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_58_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_58_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_58_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_59_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_59_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_59_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_59_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_59_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_59_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_59_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_59_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_59_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_60_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_60_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_60_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_60_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_60_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_60_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_60_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_60_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_60_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_61_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_61_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_61_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_61_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_61_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_61_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_61_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_61_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_61_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_62_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_62_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_62_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_62_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_62_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_62_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_62_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_62_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_62_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_63_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_63_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_63_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_63_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_63_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_63_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_63_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_63_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_63_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_64_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_64_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_64_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_64_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_64_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_64_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_64_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_64_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_64_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_65_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_65_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_65_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_65_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_65_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_65_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_65_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_65_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_65_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_66_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_66_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_66_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_66_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_66_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_66_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_66_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_66_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_66_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_67_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_67_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_67_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_67_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_67_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_67_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_67_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_67_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_67_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_68_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_68_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_68_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_68_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_68_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_68_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_68_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_68_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_68_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_69_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_69_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_69_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_69_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_69_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_69_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_69_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_69_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_69_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_70_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_70_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_70_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_70_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_70_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_70_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_70_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_70_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_70_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_71_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_71_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_71_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_71_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_71_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_71_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_71_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_71_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_71_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_72_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_72_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_72_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_72_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_72_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_72_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_72_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_72_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_72_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_73_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_73_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_73_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_73_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_73_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_73_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_73_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_73_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_73_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_74_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_74_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_74_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_74_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_74_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_74_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_74_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_74_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_74_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_75_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_75_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_75_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_75_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_75_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_75_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_75_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_75_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_75_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_76_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_76_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_76_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_76_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_76_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_76_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_76_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_76_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_76_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_77_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_77_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_77_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_77_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_77_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_77_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_77_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_77_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_77_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_78_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_78_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_78_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_78_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_78_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_78_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_78_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_78_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_78_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_79_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_79_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_79_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_79_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_79_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_79_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_79_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_79_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_79_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_80_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_80_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_80_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_80_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_80_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_80_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_80_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_80_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_80_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_81_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_81_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_81_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_81_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_81_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_81_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_81_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_81_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_81_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_82_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_82_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_82_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_82_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_82_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_82_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_82_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_82_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_82_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_83_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_83_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_83_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_83_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_83_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_83_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_83_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_83_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_83_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_84_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_84_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_84_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_84_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_84_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_84_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_84_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_84_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_84_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_85_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_85_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_85_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_85_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_85_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_85_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_85_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_85_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_85_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_86_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_86_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_86_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_86_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_86_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_86_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_86_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_86_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_86_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_87_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_87_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_87_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_87_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_87_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_87_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_87_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_87_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_87_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_88_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_88_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_88_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_88_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_88_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_88_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_88_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_88_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_88_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_89_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_89_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_89_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_89_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_89_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_89_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_89_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_89_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_89_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_90_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_90_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_90_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_90_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_90_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_90_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_90_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_90_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_90_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_91_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_91_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_91_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_91_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_91_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_91_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_91_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_91_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_91_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_92_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_92_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_92_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_92_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_92_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_92_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_92_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_92_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_92_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_93_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_93_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_93_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_93_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_93_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_93_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_93_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_93_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_93_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_94_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_94_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_94_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_94_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_94_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_94_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_94_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_94_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_94_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_95_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_95_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_95_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_95_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_95_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_95_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_95_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_95_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_95_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_96_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_96_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_96_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_96_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_96_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_96_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_96_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_96_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_96_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_97_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_97_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_97_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_97_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_97_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_97_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_97_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_97_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_97_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_98_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_98_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_98_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_98_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_98_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_98_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_98_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_98_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_98_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_99_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_99_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_99_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_99_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_99_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_99_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_99_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_99_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_99_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_100_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_100_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_100_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_100_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_100_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_100_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_100_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_100_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_100_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_101_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_101_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_101_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_101_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_101_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_101_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_101_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_101_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_101_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_102_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_102_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_102_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_102_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_102_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_102_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_102_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_102_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_102_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_103_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_103_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_103_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_103_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_103_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_103_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_103_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_103_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_103_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_104_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_104_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_104_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_104_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_104_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_104_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_104_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_104_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_104_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_105_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_105_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_105_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_105_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_105_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_105_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_105_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_105_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_105_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_106_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_106_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_106_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_106_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_106_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_106_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_106_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_106_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_106_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_107_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_107_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_107_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_107_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_107_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_107_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_107_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_107_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_107_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_108_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_108_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_108_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_108_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_108_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_108_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_108_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_108_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_108_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_109_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_109_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_109_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_109_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_109_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_109_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_109_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_109_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_109_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_110_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_110_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_110_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_110_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_110_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_110_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_110_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_110_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_110_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_111_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_111_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_111_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_111_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_111_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_111_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_111_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_111_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_111_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_112_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_112_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_112_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_112_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_112_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_112_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_112_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_112_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_112_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_113_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_113_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_113_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_113_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_113_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_113_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_113_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_113_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_113_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_114_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_114_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_114_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_114_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_114_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_114_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_114_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_114_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_114_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_115_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_115_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_115_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_115_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_115_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_115_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_115_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_115_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_115_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_116_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_116_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_116_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_116_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_116_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_116_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_116_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_116_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_116_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_117_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_117_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_117_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_117_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_117_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_117_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_117_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_117_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_117_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_118_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_118_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_118_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_118_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_118_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_118_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_118_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_118_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_118_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_119_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_119_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_119_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_119_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_119_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_119_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_119_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_119_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_119_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_120_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_120_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_120_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_120_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_120_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_120_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_120_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_120_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_120_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_121_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_121_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_121_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_121_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_121_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_121_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_121_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_121_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_121_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_122_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_122_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_122_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_122_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_122_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_122_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_122_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_122_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_122_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_123_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_123_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_123_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_123_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_123_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_123_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_123_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_123_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_123_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_124_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_124_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_124_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_124_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_124_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_124_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_124_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_124_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_124_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_125_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_125_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_125_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_125_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_125_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_125_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_125_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_125_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_125_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_126_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_126_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_126_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_126_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_126_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_126_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_126_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_126_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_126_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_127_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_127_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_127_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_127_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_127_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_127_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_127_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_127_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_127_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_128_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_128_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_128_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_128_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_128_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_128_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_128_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_128_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_128_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_129_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_129_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_129_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_129_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_129_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_129_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_129_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_129_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_129_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_130_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_130_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_130_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_130_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_130_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_130_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_130_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_130_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_130_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_131_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_131_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_131_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_131_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_131_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_131_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_131_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_131_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_131_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_132_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_132_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_132_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_132_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_132_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_132_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_132_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_132_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_132_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_133_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_133_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_133_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_133_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_133_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_133_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_133_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_133_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_133_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_134_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_134_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_134_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_134_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_134_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_134_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_134_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_134_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_134_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_135_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_135_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_135_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_135_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_135_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_135_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_135_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_135_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_135_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_136_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_136_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_136_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_136_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_136_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_136_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_136_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_136_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_136_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_137_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_137_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_137_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_137_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_137_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_137_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_137_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_137_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_137_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_138_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_138_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_138_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_138_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_138_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_138_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_138_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_138_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_138_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_139_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_139_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_139_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_139_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_139_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_139_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_139_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_139_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_139_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_140_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_140_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_140_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_140_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_140_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_140_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_140_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_140_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_140_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_141_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_141_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_141_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_141_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_141_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_141_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_141_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_141_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_141_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_142_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_142_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_142_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_142_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_142_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_142_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_142_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_142_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_142_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_143_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_143_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_143_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_143_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_143_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_143_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_143_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_143_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_143_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_144_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_144_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_144_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_144_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_144_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_144_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_144_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_144_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_144_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_145_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_145_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_145_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_145_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_145_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_145_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_145_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_145_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_145_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_146_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_146_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_146_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_146_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_146_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_146_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_146_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_146_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_146_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_147_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_147_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_147_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_147_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_147_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_147_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_147_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_147_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_147_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_148_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_148_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_148_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_148_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_148_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_148_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_148_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_148_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_148_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_149_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_149_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_149_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_149_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_149_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_149_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_149_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_149_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_149_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_150_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_150_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_150_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_150_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_150_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_150_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_150_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_150_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_150_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_151_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_151_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_151_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_151_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_151_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_151_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_151_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_151_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_151_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_152_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_152_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_152_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_152_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_152_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_152_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_152_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_152_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_152_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_153_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_153_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_153_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_153_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_153_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_153_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_153_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_153_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_153_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_154_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_154_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_154_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_154_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_154_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_154_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_154_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_154_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_154_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_155_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_155_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_155_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_155_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_155_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_155_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_155_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_155_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_155_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_156_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_156_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_156_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_156_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_156_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_156_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_156_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_156_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_156_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_157_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_157_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_157_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_157_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_157_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_157_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_157_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_157_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_157_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_158_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_158_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_158_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_158_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_158_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_158_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_158_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_158_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_158_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_159_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_159_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_159_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_159_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_159_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_159_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_159_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_159_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_159_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_160_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_160_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_160_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_160_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_160_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_160_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_160_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_160_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_160_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_161_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_161_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_161_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_161_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_161_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_161_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_161_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_161_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_161_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_162_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_162_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_162_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_162_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_162_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_162_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_162_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_162_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_162_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_163_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_163_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_163_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_163_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_163_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_163_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_163_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_163_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_163_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_164_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_164_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_164_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_164_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_164_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_164_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_164_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_164_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_164_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_165_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_165_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_165_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_165_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_165_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_165_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_165_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_165_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_165_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_166_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_166_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_166_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_166_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_166_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_166_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_166_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_166_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_166_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_167_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_167_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_167_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_167_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_167_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_167_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_167_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_167_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_167_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_168_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_168_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_168_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_168_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_168_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_168_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_168_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_168_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_168_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_169_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_169_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_169_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_169_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_169_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_169_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_169_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_169_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_169_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_170_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_170_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_170_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_170_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_170_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_170_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_170_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_170_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_170_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_171_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_171_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_171_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_171_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_171_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_171_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_171_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_171_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_171_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_172_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_172_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_172_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_172_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_172_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_172_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_172_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_172_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_172_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_173_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_173_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_173_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_173_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_173_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_173_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_173_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_173_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_173_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_174_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_174_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_174_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_174_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_174_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_174_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_174_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_174_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_174_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_175_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_175_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_175_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_175_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_175_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_175_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_175_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_175_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_175_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_176_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_176_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_176_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_176_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_176_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_176_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_176_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_176_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_176_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_177_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_177_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_177_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_177_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_177_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_177_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_177_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_177_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_177_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_178_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_178_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_178_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_178_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_178_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_178_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_178_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_178_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_178_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_179_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_179_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_179_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_179_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_179_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_179_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_179_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_179_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_179_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_180_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_180_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_180_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_180_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_180_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_180_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_180_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_180_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_180_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_181_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_181_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_181_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_181_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_181_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_181_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_181_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_181_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_181_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_182_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_182_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_182_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_182_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_182_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_182_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_182_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_182_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_182_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_183_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_183_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_183_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_183_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_183_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_183_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_183_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_183_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_183_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_184_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_184_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_184_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_184_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_184_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_184_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_184_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_184_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_184_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_185_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_185_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_185_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_185_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_185_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_185_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_185_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_185_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_185_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_186_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_186_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_186_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_186_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_186_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_186_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_186_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_186_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_186_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_187_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_187_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_187_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_187_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_187_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_187_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_187_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_187_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_187_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_188_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_188_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_188_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_188_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_188_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_188_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_188_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_188_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_188_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_189_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_189_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_189_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_189_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_189_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_189_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_189_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_189_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_189_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_190_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_190_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_190_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_190_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_190_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_190_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_190_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_190_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_190_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_191_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_191_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_191_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_191_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_191_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_191_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_191_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_191_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_191_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_192_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_192_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_192_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_192_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_192_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_192_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_192_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_192_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_192_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_193_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_193_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_193_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_193_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_193_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_193_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_193_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_193_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_193_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_194_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_194_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_194_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_194_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_194_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_194_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_194_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_194_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_194_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_195_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_195_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_195_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_195_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_195_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_195_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_195_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_195_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_195_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_196_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_196_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_196_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_196_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_196_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_196_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_196_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_196_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_196_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_197_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_197_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_197_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_197_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_197_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_197_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_197_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_197_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_197_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_198_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_198_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_198_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_198_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_198_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_198_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_198_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_198_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_198_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_199_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_199_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_199_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_199_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_199_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_199_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_199_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_199_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_199_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_200_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_200_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_200_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_200_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_200_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_200_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_200_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_200_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_200_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_201_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_201_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_201_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_201_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_201_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_201_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_201_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_201_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_201_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_202_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_202_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_202_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_202_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_202_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_202_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_202_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_202_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_202_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_203_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_203_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_203_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_203_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_203_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_203_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_203_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_203_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_203_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_204_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_204_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_204_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_204_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_204_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_204_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_204_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_204_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_204_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_205_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_205_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_205_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_205_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_205_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_205_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_205_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_205_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_205_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_206_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_206_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_206_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_206_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_206_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_206_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_206_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_206_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_206_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_207_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_207_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_207_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_207_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_207_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_207_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_207_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_207_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_207_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_208_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_208_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_208_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_208_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_208_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_208_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_208_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_208_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_208_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_209_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_209_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_209_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_209_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_209_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_209_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_209_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_209_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_209_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_210_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_210_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_210_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_210_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_210_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_210_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_210_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_210_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_210_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_211_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_211_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_211_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_211_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_211_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_211_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_211_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_211_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_211_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_212_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_212_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_212_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_212_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_212_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_212_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_212_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_212_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_212_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_213_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_213_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_213_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_213_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_213_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_213_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_213_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_213_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_213_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_214_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_214_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_214_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_214_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_214_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_214_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_214_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_214_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_214_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_215_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_215_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_215_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_215_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_215_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_215_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_215_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_215_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_215_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_216_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_216_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_216_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_216_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_216_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_216_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_216_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_216_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_216_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_217_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_217_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_217_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_217_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_217_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_217_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_217_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_217_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_217_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_218_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_218_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_218_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_218_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_218_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_218_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_218_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_218_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_218_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_219_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_219_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_219_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_219_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_219_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_219_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_219_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_219_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_219_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_220_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_220_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_220_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_220_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_220_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_220_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_220_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_220_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_220_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_221_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_221_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_221_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_221_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_221_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_221_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_221_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_221_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_221_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_222_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_222_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_222_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_222_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_222_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_222_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_222_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_222_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_222_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_223_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_223_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_223_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_223_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_223_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_223_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_223_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_223_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_223_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_224_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_224_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_224_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_224_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_224_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_224_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_224_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_224_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_224_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_225_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_225_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_225_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_225_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_225_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_225_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_225_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_225_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_225_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_226_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_226_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_226_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_226_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_226_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_226_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_226_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_226_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_226_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_227_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_227_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_227_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_227_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_227_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_227_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_227_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_227_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_227_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_228_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_228_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_228_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_228_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_228_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_228_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_228_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_228_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_228_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_229_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_229_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_229_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_229_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_229_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_229_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_229_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_229_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_229_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_230_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_230_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_230_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_230_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_230_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_230_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_230_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_230_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_230_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_231_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_231_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_231_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_231_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_231_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_231_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_231_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_231_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_231_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_232_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_232_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_232_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_232_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_232_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_232_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_232_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_232_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_232_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_233_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_233_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_233_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_233_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_233_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_233_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_233_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_233_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_233_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_234_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_234_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_234_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_234_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_234_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_234_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_234_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_234_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_234_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_235_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_235_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_235_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_235_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_235_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_235_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_235_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_235_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_235_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_236_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_236_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_236_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_236_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_236_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_236_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_236_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_236_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_236_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_237_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_237_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_237_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_237_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_237_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_237_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_237_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_237_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_237_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_238_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_238_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_238_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_238_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_238_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_238_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_238_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_238_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_238_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_239_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_239_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_239_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_239_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_239_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_239_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_239_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_239_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_239_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_240_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_240_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_240_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_240_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_240_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_240_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_240_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_240_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_240_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_241_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_241_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_241_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_241_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_241_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_241_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_241_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_241_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_241_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_242_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_242_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_242_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_242_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_242_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_242_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_242_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_242_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_242_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_243_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_243_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_243_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_243_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_243_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_243_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_243_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_243_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_243_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_244_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_244_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_244_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_244_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_244_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_244_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_244_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_244_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_244_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_245_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_245_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_245_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_245_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_245_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_245_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_245_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_245_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_245_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_246_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_246_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_246_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_246_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_246_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_246_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_246_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_246_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_246_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_247_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_247_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_247_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_247_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_247_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_247_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_247_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_247_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_247_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_248_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_248_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_248_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_248_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_248_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_248_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_248_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_248_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_248_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_249_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_249_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_249_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_249_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_249_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_249_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_249_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_249_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_249_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_250_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_250_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_250_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_250_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_250_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_250_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_250_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_250_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_250_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_251_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_251_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_251_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_251_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_251_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_251_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_251_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_251_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_251_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_252_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_252_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_252_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_252_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_252_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_252_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_252_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_252_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_252_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_253_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_253_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_253_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_253_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_253_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_253_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_253_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_253_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_253_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_254_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_254_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_254_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_254_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_254_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_254_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_254_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_254_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_254_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_255_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_255_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_255_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_255_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_255_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_255_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_255_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_255_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_255_0_io_outs_3; // @[MockArray.scala 36:52]
  Element ces_0_0 ( // @[MockArray.scala 36:52]
    .clock(ces_0_0_clock),
    .io_ins_0(ces_0_0_io_ins_0),
    .io_ins_1(ces_0_0_io_ins_1),
    .io_ins_2(ces_0_0_io_ins_2),
    .io_ins_3(ces_0_0_io_ins_3),
    .io_outs_0(ces_0_0_io_outs_0),
    .io_outs_1(ces_0_0_io_outs_1),
    .io_outs_2(ces_0_0_io_outs_2),
    .io_outs_3(ces_0_0_io_outs_3)
  );
  Element ces_1_0 ( // @[MockArray.scala 36:52]
    .clock(ces_1_0_clock),
    .io_ins_0(ces_1_0_io_ins_0),
    .io_ins_1(ces_1_0_io_ins_1),
    .io_ins_2(ces_1_0_io_ins_2),
    .io_ins_3(ces_1_0_io_ins_3),
    .io_outs_0(ces_1_0_io_outs_0),
    .io_outs_1(ces_1_0_io_outs_1),
    .io_outs_2(ces_1_0_io_outs_2),
    .io_outs_3(ces_1_0_io_outs_3)
  );
  Element ces_2_0 ( // @[MockArray.scala 36:52]
    .clock(ces_2_0_clock),
    .io_ins_0(ces_2_0_io_ins_0),
    .io_ins_1(ces_2_0_io_ins_1),
    .io_ins_2(ces_2_0_io_ins_2),
    .io_ins_3(ces_2_0_io_ins_3),
    .io_outs_0(ces_2_0_io_outs_0),
    .io_outs_1(ces_2_0_io_outs_1),
    .io_outs_2(ces_2_0_io_outs_2),
    .io_outs_3(ces_2_0_io_outs_3)
  );
  Element ces_3_0 ( // @[MockArray.scala 36:52]
    .clock(ces_3_0_clock),
    .io_ins_0(ces_3_0_io_ins_0),
    .io_ins_1(ces_3_0_io_ins_1),
    .io_ins_2(ces_3_0_io_ins_2),
    .io_ins_3(ces_3_0_io_ins_3),
    .io_outs_0(ces_3_0_io_outs_0),
    .io_outs_1(ces_3_0_io_outs_1),
    .io_outs_2(ces_3_0_io_outs_2),
    .io_outs_3(ces_3_0_io_outs_3)
  );
  Element ces_4_0 ( // @[MockArray.scala 36:52]
    .clock(ces_4_0_clock),
    .io_ins_0(ces_4_0_io_ins_0),
    .io_ins_1(ces_4_0_io_ins_1),
    .io_ins_2(ces_4_0_io_ins_2),
    .io_ins_3(ces_4_0_io_ins_3),
    .io_outs_0(ces_4_0_io_outs_0),
    .io_outs_1(ces_4_0_io_outs_1),
    .io_outs_2(ces_4_0_io_outs_2),
    .io_outs_3(ces_4_0_io_outs_3)
  );
  Element ces_5_0 ( // @[MockArray.scala 36:52]
    .clock(ces_5_0_clock),
    .io_ins_0(ces_5_0_io_ins_0),
    .io_ins_1(ces_5_0_io_ins_1),
    .io_ins_2(ces_5_0_io_ins_2),
    .io_ins_3(ces_5_0_io_ins_3),
    .io_outs_0(ces_5_0_io_outs_0),
    .io_outs_1(ces_5_0_io_outs_1),
    .io_outs_2(ces_5_0_io_outs_2),
    .io_outs_3(ces_5_0_io_outs_3)
  );
  Element ces_6_0 ( // @[MockArray.scala 36:52]
    .clock(ces_6_0_clock),
    .io_ins_0(ces_6_0_io_ins_0),
    .io_ins_1(ces_6_0_io_ins_1),
    .io_ins_2(ces_6_0_io_ins_2),
    .io_ins_3(ces_6_0_io_ins_3),
    .io_outs_0(ces_6_0_io_outs_0),
    .io_outs_1(ces_6_0_io_outs_1),
    .io_outs_2(ces_6_0_io_outs_2),
    .io_outs_3(ces_6_0_io_outs_3)
  );
  Element ces_7_0 ( // @[MockArray.scala 36:52]
    .clock(ces_7_0_clock),
    .io_ins_0(ces_7_0_io_ins_0),
    .io_ins_1(ces_7_0_io_ins_1),
    .io_ins_2(ces_7_0_io_ins_2),
    .io_ins_3(ces_7_0_io_ins_3),
    .io_outs_0(ces_7_0_io_outs_0),
    .io_outs_1(ces_7_0_io_outs_1),
    .io_outs_2(ces_7_0_io_outs_2),
    .io_outs_3(ces_7_0_io_outs_3)
  );
  Element ces_8_0 ( // @[MockArray.scala 36:52]
    .clock(ces_8_0_clock),
    .io_ins_0(ces_8_0_io_ins_0),
    .io_ins_1(ces_8_0_io_ins_1),
    .io_ins_2(ces_8_0_io_ins_2),
    .io_ins_3(ces_8_0_io_ins_3),
    .io_outs_0(ces_8_0_io_outs_0),
    .io_outs_1(ces_8_0_io_outs_1),
    .io_outs_2(ces_8_0_io_outs_2),
    .io_outs_3(ces_8_0_io_outs_3)
  );
  Element ces_9_0 ( // @[MockArray.scala 36:52]
    .clock(ces_9_0_clock),
    .io_ins_0(ces_9_0_io_ins_0),
    .io_ins_1(ces_9_0_io_ins_1),
    .io_ins_2(ces_9_0_io_ins_2),
    .io_ins_3(ces_9_0_io_ins_3),
    .io_outs_0(ces_9_0_io_outs_0),
    .io_outs_1(ces_9_0_io_outs_1),
    .io_outs_2(ces_9_0_io_outs_2),
    .io_outs_3(ces_9_0_io_outs_3)
  );
  Element ces_10_0 ( // @[MockArray.scala 36:52]
    .clock(ces_10_0_clock),
    .io_ins_0(ces_10_0_io_ins_0),
    .io_ins_1(ces_10_0_io_ins_1),
    .io_ins_2(ces_10_0_io_ins_2),
    .io_ins_3(ces_10_0_io_ins_3),
    .io_outs_0(ces_10_0_io_outs_0),
    .io_outs_1(ces_10_0_io_outs_1),
    .io_outs_2(ces_10_0_io_outs_2),
    .io_outs_3(ces_10_0_io_outs_3)
  );
  Element ces_11_0 ( // @[MockArray.scala 36:52]
    .clock(ces_11_0_clock),
    .io_ins_0(ces_11_0_io_ins_0),
    .io_ins_1(ces_11_0_io_ins_1),
    .io_ins_2(ces_11_0_io_ins_2),
    .io_ins_3(ces_11_0_io_ins_3),
    .io_outs_0(ces_11_0_io_outs_0),
    .io_outs_1(ces_11_0_io_outs_1),
    .io_outs_2(ces_11_0_io_outs_2),
    .io_outs_3(ces_11_0_io_outs_3)
  );
  Element ces_12_0 ( // @[MockArray.scala 36:52]
    .clock(ces_12_0_clock),
    .io_ins_0(ces_12_0_io_ins_0),
    .io_ins_1(ces_12_0_io_ins_1),
    .io_ins_2(ces_12_0_io_ins_2),
    .io_ins_3(ces_12_0_io_ins_3),
    .io_outs_0(ces_12_0_io_outs_0),
    .io_outs_1(ces_12_0_io_outs_1),
    .io_outs_2(ces_12_0_io_outs_2),
    .io_outs_3(ces_12_0_io_outs_3)
  );
  Element ces_13_0 ( // @[MockArray.scala 36:52]
    .clock(ces_13_0_clock),
    .io_ins_0(ces_13_0_io_ins_0),
    .io_ins_1(ces_13_0_io_ins_1),
    .io_ins_2(ces_13_0_io_ins_2),
    .io_ins_3(ces_13_0_io_ins_3),
    .io_outs_0(ces_13_0_io_outs_0),
    .io_outs_1(ces_13_0_io_outs_1),
    .io_outs_2(ces_13_0_io_outs_2),
    .io_outs_3(ces_13_0_io_outs_3)
  );
  Element ces_14_0 ( // @[MockArray.scala 36:52]
    .clock(ces_14_0_clock),
    .io_ins_0(ces_14_0_io_ins_0),
    .io_ins_1(ces_14_0_io_ins_1),
    .io_ins_2(ces_14_0_io_ins_2),
    .io_ins_3(ces_14_0_io_ins_3),
    .io_outs_0(ces_14_0_io_outs_0),
    .io_outs_1(ces_14_0_io_outs_1),
    .io_outs_2(ces_14_0_io_outs_2),
    .io_outs_3(ces_14_0_io_outs_3)
  );
  Element ces_15_0 ( // @[MockArray.scala 36:52]
    .clock(ces_15_0_clock),
    .io_ins_0(ces_15_0_io_ins_0),
    .io_ins_1(ces_15_0_io_ins_1),
    .io_ins_2(ces_15_0_io_ins_2),
    .io_ins_3(ces_15_0_io_ins_3),
    .io_outs_0(ces_15_0_io_outs_0),
    .io_outs_1(ces_15_0_io_outs_1),
    .io_outs_2(ces_15_0_io_outs_2),
    .io_outs_3(ces_15_0_io_outs_3)
  );
  Element ces_16_0 ( // @[MockArray.scala 36:52]
    .clock(ces_16_0_clock),
    .io_ins_0(ces_16_0_io_ins_0),
    .io_ins_1(ces_16_0_io_ins_1),
    .io_ins_2(ces_16_0_io_ins_2),
    .io_ins_3(ces_16_0_io_ins_3),
    .io_outs_0(ces_16_0_io_outs_0),
    .io_outs_1(ces_16_0_io_outs_1),
    .io_outs_2(ces_16_0_io_outs_2),
    .io_outs_3(ces_16_0_io_outs_3)
  );
  Element ces_17_0 ( // @[MockArray.scala 36:52]
    .clock(ces_17_0_clock),
    .io_ins_0(ces_17_0_io_ins_0),
    .io_ins_1(ces_17_0_io_ins_1),
    .io_ins_2(ces_17_0_io_ins_2),
    .io_ins_3(ces_17_0_io_ins_3),
    .io_outs_0(ces_17_0_io_outs_0),
    .io_outs_1(ces_17_0_io_outs_1),
    .io_outs_2(ces_17_0_io_outs_2),
    .io_outs_3(ces_17_0_io_outs_3)
  );
  Element ces_18_0 ( // @[MockArray.scala 36:52]
    .clock(ces_18_0_clock),
    .io_ins_0(ces_18_0_io_ins_0),
    .io_ins_1(ces_18_0_io_ins_1),
    .io_ins_2(ces_18_0_io_ins_2),
    .io_ins_3(ces_18_0_io_ins_3),
    .io_outs_0(ces_18_0_io_outs_0),
    .io_outs_1(ces_18_0_io_outs_1),
    .io_outs_2(ces_18_0_io_outs_2),
    .io_outs_3(ces_18_0_io_outs_3)
  );
  Element ces_19_0 ( // @[MockArray.scala 36:52]
    .clock(ces_19_0_clock),
    .io_ins_0(ces_19_0_io_ins_0),
    .io_ins_1(ces_19_0_io_ins_1),
    .io_ins_2(ces_19_0_io_ins_2),
    .io_ins_3(ces_19_0_io_ins_3),
    .io_outs_0(ces_19_0_io_outs_0),
    .io_outs_1(ces_19_0_io_outs_1),
    .io_outs_2(ces_19_0_io_outs_2),
    .io_outs_3(ces_19_0_io_outs_3)
  );
  Element ces_20_0 ( // @[MockArray.scala 36:52]
    .clock(ces_20_0_clock),
    .io_ins_0(ces_20_0_io_ins_0),
    .io_ins_1(ces_20_0_io_ins_1),
    .io_ins_2(ces_20_0_io_ins_2),
    .io_ins_3(ces_20_0_io_ins_3),
    .io_outs_0(ces_20_0_io_outs_0),
    .io_outs_1(ces_20_0_io_outs_1),
    .io_outs_2(ces_20_0_io_outs_2),
    .io_outs_3(ces_20_0_io_outs_3)
  );
  Element ces_21_0 ( // @[MockArray.scala 36:52]
    .clock(ces_21_0_clock),
    .io_ins_0(ces_21_0_io_ins_0),
    .io_ins_1(ces_21_0_io_ins_1),
    .io_ins_2(ces_21_0_io_ins_2),
    .io_ins_3(ces_21_0_io_ins_3),
    .io_outs_0(ces_21_0_io_outs_0),
    .io_outs_1(ces_21_0_io_outs_1),
    .io_outs_2(ces_21_0_io_outs_2),
    .io_outs_3(ces_21_0_io_outs_3)
  );
  Element ces_22_0 ( // @[MockArray.scala 36:52]
    .clock(ces_22_0_clock),
    .io_ins_0(ces_22_0_io_ins_0),
    .io_ins_1(ces_22_0_io_ins_1),
    .io_ins_2(ces_22_0_io_ins_2),
    .io_ins_3(ces_22_0_io_ins_3),
    .io_outs_0(ces_22_0_io_outs_0),
    .io_outs_1(ces_22_0_io_outs_1),
    .io_outs_2(ces_22_0_io_outs_2),
    .io_outs_3(ces_22_0_io_outs_3)
  );
  Element ces_23_0 ( // @[MockArray.scala 36:52]
    .clock(ces_23_0_clock),
    .io_ins_0(ces_23_0_io_ins_0),
    .io_ins_1(ces_23_0_io_ins_1),
    .io_ins_2(ces_23_0_io_ins_2),
    .io_ins_3(ces_23_0_io_ins_3),
    .io_outs_0(ces_23_0_io_outs_0),
    .io_outs_1(ces_23_0_io_outs_1),
    .io_outs_2(ces_23_0_io_outs_2),
    .io_outs_3(ces_23_0_io_outs_3)
  );
  Element ces_24_0 ( // @[MockArray.scala 36:52]
    .clock(ces_24_0_clock),
    .io_ins_0(ces_24_0_io_ins_0),
    .io_ins_1(ces_24_0_io_ins_1),
    .io_ins_2(ces_24_0_io_ins_2),
    .io_ins_3(ces_24_0_io_ins_3),
    .io_outs_0(ces_24_0_io_outs_0),
    .io_outs_1(ces_24_0_io_outs_1),
    .io_outs_2(ces_24_0_io_outs_2),
    .io_outs_3(ces_24_0_io_outs_3)
  );
  Element ces_25_0 ( // @[MockArray.scala 36:52]
    .clock(ces_25_0_clock),
    .io_ins_0(ces_25_0_io_ins_0),
    .io_ins_1(ces_25_0_io_ins_1),
    .io_ins_2(ces_25_0_io_ins_2),
    .io_ins_3(ces_25_0_io_ins_3),
    .io_outs_0(ces_25_0_io_outs_0),
    .io_outs_1(ces_25_0_io_outs_1),
    .io_outs_2(ces_25_0_io_outs_2),
    .io_outs_3(ces_25_0_io_outs_3)
  );
  Element ces_26_0 ( // @[MockArray.scala 36:52]
    .clock(ces_26_0_clock),
    .io_ins_0(ces_26_0_io_ins_0),
    .io_ins_1(ces_26_0_io_ins_1),
    .io_ins_2(ces_26_0_io_ins_2),
    .io_ins_3(ces_26_0_io_ins_3),
    .io_outs_0(ces_26_0_io_outs_0),
    .io_outs_1(ces_26_0_io_outs_1),
    .io_outs_2(ces_26_0_io_outs_2),
    .io_outs_3(ces_26_0_io_outs_3)
  );
  Element ces_27_0 ( // @[MockArray.scala 36:52]
    .clock(ces_27_0_clock),
    .io_ins_0(ces_27_0_io_ins_0),
    .io_ins_1(ces_27_0_io_ins_1),
    .io_ins_2(ces_27_0_io_ins_2),
    .io_ins_3(ces_27_0_io_ins_3),
    .io_outs_0(ces_27_0_io_outs_0),
    .io_outs_1(ces_27_0_io_outs_1),
    .io_outs_2(ces_27_0_io_outs_2),
    .io_outs_3(ces_27_0_io_outs_3)
  );
  Element ces_28_0 ( // @[MockArray.scala 36:52]
    .clock(ces_28_0_clock),
    .io_ins_0(ces_28_0_io_ins_0),
    .io_ins_1(ces_28_0_io_ins_1),
    .io_ins_2(ces_28_0_io_ins_2),
    .io_ins_3(ces_28_0_io_ins_3),
    .io_outs_0(ces_28_0_io_outs_0),
    .io_outs_1(ces_28_0_io_outs_1),
    .io_outs_2(ces_28_0_io_outs_2),
    .io_outs_3(ces_28_0_io_outs_3)
  );
  Element ces_29_0 ( // @[MockArray.scala 36:52]
    .clock(ces_29_0_clock),
    .io_ins_0(ces_29_0_io_ins_0),
    .io_ins_1(ces_29_0_io_ins_1),
    .io_ins_2(ces_29_0_io_ins_2),
    .io_ins_3(ces_29_0_io_ins_3),
    .io_outs_0(ces_29_0_io_outs_0),
    .io_outs_1(ces_29_0_io_outs_1),
    .io_outs_2(ces_29_0_io_outs_2),
    .io_outs_3(ces_29_0_io_outs_3)
  );
  Element ces_30_0 ( // @[MockArray.scala 36:52]
    .clock(ces_30_0_clock),
    .io_ins_0(ces_30_0_io_ins_0),
    .io_ins_1(ces_30_0_io_ins_1),
    .io_ins_2(ces_30_0_io_ins_2),
    .io_ins_3(ces_30_0_io_ins_3),
    .io_outs_0(ces_30_0_io_outs_0),
    .io_outs_1(ces_30_0_io_outs_1),
    .io_outs_2(ces_30_0_io_outs_2),
    .io_outs_3(ces_30_0_io_outs_3)
  );
  Element ces_31_0 ( // @[MockArray.scala 36:52]
    .clock(ces_31_0_clock),
    .io_ins_0(ces_31_0_io_ins_0),
    .io_ins_1(ces_31_0_io_ins_1),
    .io_ins_2(ces_31_0_io_ins_2),
    .io_ins_3(ces_31_0_io_ins_3),
    .io_outs_0(ces_31_0_io_outs_0),
    .io_outs_1(ces_31_0_io_outs_1),
    .io_outs_2(ces_31_0_io_outs_2),
    .io_outs_3(ces_31_0_io_outs_3)
  );
  Element ces_32_0 ( // @[MockArray.scala 36:52]
    .clock(ces_32_0_clock),
    .io_ins_0(ces_32_0_io_ins_0),
    .io_ins_1(ces_32_0_io_ins_1),
    .io_ins_2(ces_32_0_io_ins_2),
    .io_ins_3(ces_32_0_io_ins_3),
    .io_outs_0(ces_32_0_io_outs_0),
    .io_outs_1(ces_32_0_io_outs_1),
    .io_outs_2(ces_32_0_io_outs_2),
    .io_outs_3(ces_32_0_io_outs_3)
  );
  Element ces_33_0 ( // @[MockArray.scala 36:52]
    .clock(ces_33_0_clock),
    .io_ins_0(ces_33_0_io_ins_0),
    .io_ins_1(ces_33_0_io_ins_1),
    .io_ins_2(ces_33_0_io_ins_2),
    .io_ins_3(ces_33_0_io_ins_3),
    .io_outs_0(ces_33_0_io_outs_0),
    .io_outs_1(ces_33_0_io_outs_1),
    .io_outs_2(ces_33_0_io_outs_2),
    .io_outs_3(ces_33_0_io_outs_3)
  );
  Element ces_34_0 ( // @[MockArray.scala 36:52]
    .clock(ces_34_0_clock),
    .io_ins_0(ces_34_0_io_ins_0),
    .io_ins_1(ces_34_0_io_ins_1),
    .io_ins_2(ces_34_0_io_ins_2),
    .io_ins_3(ces_34_0_io_ins_3),
    .io_outs_0(ces_34_0_io_outs_0),
    .io_outs_1(ces_34_0_io_outs_1),
    .io_outs_2(ces_34_0_io_outs_2),
    .io_outs_3(ces_34_0_io_outs_3)
  );
  Element ces_35_0 ( // @[MockArray.scala 36:52]
    .clock(ces_35_0_clock),
    .io_ins_0(ces_35_0_io_ins_0),
    .io_ins_1(ces_35_0_io_ins_1),
    .io_ins_2(ces_35_0_io_ins_2),
    .io_ins_3(ces_35_0_io_ins_3),
    .io_outs_0(ces_35_0_io_outs_0),
    .io_outs_1(ces_35_0_io_outs_1),
    .io_outs_2(ces_35_0_io_outs_2),
    .io_outs_3(ces_35_0_io_outs_3)
  );
  Element ces_36_0 ( // @[MockArray.scala 36:52]
    .clock(ces_36_0_clock),
    .io_ins_0(ces_36_0_io_ins_0),
    .io_ins_1(ces_36_0_io_ins_1),
    .io_ins_2(ces_36_0_io_ins_2),
    .io_ins_3(ces_36_0_io_ins_3),
    .io_outs_0(ces_36_0_io_outs_0),
    .io_outs_1(ces_36_0_io_outs_1),
    .io_outs_2(ces_36_0_io_outs_2),
    .io_outs_3(ces_36_0_io_outs_3)
  );
  Element ces_37_0 ( // @[MockArray.scala 36:52]
    .clock(ces_37_0_clock),
    .io_ins_0(ces_37_0_io_ins_0),
    .io_ins_1(ces_37_0_io_ins_1),
    .io_ins_2(ces_37_0_io_ins_2),
    .io_ins_3(ces_37_0_io_ins_3),
    .io_outs_0(ces_37_0_io_outs_0),
    .io_outs_1(ces_37_0_io_outs_1),
    .io_outs_2(ces_37_0_io_outs_2),
    .io_outs_3(ces_37_0_io_outs_3)
  );
  Element ces_38_0 ( // @[MockArray.scala 36:52]
    .clock(ces_38_0_clock),
    .io_ins_0(ces_38_0_io_ins_0),
    .io_ins_1(ces_38_0_io_ins_1),
    .io_ins_2(ces_38_0_io_ins_2),
    .io_ins_3(ces_38_0_io_ins_3),
    .io_outs_0(ces_38_0_io_outs_0),
    .io_outs_1(ces_38_0_io_outs_1),
    .io_outs_2(ces_38_0_io_outs_2),
    .io_outs_3(ces_38_0_io_outs_3)
  );
  Element ces_39_0 ( // @[MockArray.scala 36:52]
    .clock(ces_39_0_clock),
    .io_ins_0(ces_39_0_io_ins_0),
    .io_ins_1(ces_39_0_io_ins_1),
    .io_ins_2(ces_39_0_io_ins_2),
    .io_ins_3(ces_39_0_io_ins_3),
    .io_outs_0(ces_39_0_io_outs_0),
    .io_outs_1(ces_39_0_io_outs_1),
    .io_outs_2(ces_39_0_io_outs_2),
    .io_outs_3(ces_39_0_io_outs_3)
  );
  Element ces_40_0 ( // @[MockArray.scala 36:52]
    .clock(ces_40_0_clock),
    .io_ins_0(ces_40_0_io_ins_0),
    .io_ins_1(ces_40_0_io_ins_1),
    .io_ins_2(ces_40_0_io_ins_2),
    .io_ins_3(ces_40_0_io_ins_3),
    .io_outs_0(ces_40_0_io_outs_0),
    .io_outs_1(ces_40_0_io_outs_1),
    .io_outs_2(ces_40_0_io_outs_2),
    .io_outs_3(ces_40_0_io_outs_3)
  );
  Element ces_41_0 ( // @[MockArray.scala 36:52]
    .clock(ces_41_0_clock),
    .io_ins_0(ces_41_0_io_ins_0),
    .io_ins_1(ces_41_0_io_ins_1),
    .io_ins_2(ces_41_0_io_ins_2),
    .io_ins_3(ces_41_0_io_ins_3),
    .io_outs_0(ces_41_0_io_outs_0),
    .io_outs_1(ces_41_0_io_outs_1),
    .io_outs_2(ces_41_0_io_outs_2),
    .io_outs_3(ces_41_0_io_outs_3)
  );
  Element ces_42_0 ( // @[MockArray.scala 36:52]
    .clock(ces_42_0_clock),
    .io_ins_0(ces_42_0_io_ins_0),
    .io_ins_1(ces_42_0_io_ins_1),
    .io_ins_2(ces_42_0_io_ins_2),
    .io_ins_3(ces_42_0_io_ins_3),
    .io_outs_0(ces_42_0_io_outs_0),
    .io_outs_1(ces_42_0_io_outs_1),
    .io_outs_2(ces_42_0_io_outs_2),
    .io_outs_3(ces_42_0_io_outs_3)
  );
  Element ces_43_0 ( // @[MockArray.scala 36:52]
    .clock(ces_43_0_clock),
    .io_ins_0(ces_43_0_io_ins_0),
    .io_ins_1(ces_43_0_io_ins_1),
    .io_ins_2(ces_43_0_io_ins_2),
    .io_ins_3(ces_43_0_io_ins_3),
    .io_outs_0(ces_43_0_io_outs_0),
    .io_outs_1(ces_43_0_io_outs_1),
    .io_outs_2(ces_43_0_io_outs_2),
    .io_outs_3(ces_43_0_io_outs_3)
  );
  Element ces_44_0 ( // @[MockArray.scala 36:52]
    .clock(ces_44_0_clock),
    .io_ins_0(ces_44_0_io_ins_0),
    .io_ins_1(ces_44_0_io_ins_1),
    .io_ins_2(ces_44_0_io_ins_2),
    .io_ins_3(ces_44_0_io_ins_3),
    .io_outs_0(ces_44_0_io_outs_0),
    .io_outs_1(ces_44_0_io_outs_1),
    .io_outs_2(ces_44_0_io_outs_2),
    .io_outs_3(ces_44_0_io_outs_3)
  );
  Element ces_45_0 ( // @[MockArray.scala 36:52]
    .clock(ces_45_0_clock),
    .io_ins_0(ces_45_0_io_ins_0),
    .io_ins_1(ces_45_0_io_ins_1),
    .io_ins_2(ces_45_0_io_ins_2),
    .io_ins_3(ces_45_0_io_ins_3),
    .io_outs_0(ces_45_0_io_outs_0),
    .io_outs_1(ces_45_0_io_outs_1),
    .io_outs_2(ces_45_0_io_outs_2),
    .io_outs_3(ces_45_0_io_outs_3)
  );
  Element ces_46_0 ( // @[MockArray.scala 36:52]
    .clock(ces_46_0_clock),
    .io_ins_0(ces_46_0_io_ins_0),
    .io_ins_1(ces_46_0_io_ins_1),
    .io_ins_2(ces_46_0_io_ins_2),
    .io_ins_3(ces_46_0_io_ins_3),
    .io_outs_0(ces_46_0_io_outs_0),
    .io_outs_1(ces_46_0_io_outs_1),
    .io_outs_2(ces_46_0_io_outs_2),
    .io_outs_3(ces_46_0_io_outs_3)
  );
  Element ces_47_0 ( // @[MockArray.scala 36:52]
    .clock(ces_47_0_clock),
    .io_ins_0(ces_47_0_io_ins_0),
    .io_ins_1(ces_47_0_io_ins_1),
    .io_ins_2(ces_47_0_io_ins_2),
    .io_ins_3(ces_47_0_io_ins_3),
    .io_outs_0(ces_47_0_io_outs_0),
    .io_outs_1(ces_47_0_io_outs_1),
    .io_outs_2(ces_47_0_io_outs_2),
    .io_outs_3(ces_47_0_io_outs_3)
  );
  Element ces_48_0 ( // @[MockArray.scala 36:52]
    .clock(ces_48_0_clock),
    .io_ins_0(ces_48_0_io_ins_0),
    .io_ins_1(ces_48_0_io_ins_1),
    .io_ins_2(ces_48_0_io_ins_2),
    .io_ins_3(ces_48_0_io_ins_3),
    .io_outs_0(ces_48_0_io_outs_0),
    .io_outs_1(ces_48_0_io_outs_1),
    .io_outs_2(ces_48_0_io_outs_2),
    .io_outs_3(ces_48_0_io_outs_3)
  );
  Element ces_49_0 ( // @[MockArray.scala 36:52]
    .clock(ces_49_0_clock),
    .io_ins_0(ces_49_0_io_ins_0),
    .io_ins_1(ces_49_0_io_ins_1),
    .io_ins_2(ces_49_0_io_ins_2),
    .io_ins_3(ces_49_0_io_ins_3),
    .io_outs_0(ces_49_0_io_outs_0),
    .io_outs_1(ces_49_0_io_outs_1),
    .io_outs_2(ces_49_0_io_outs_2),
    .io_outs_3(ces_49_0_io_outs_3)
  );
  Element ces_50_0 ( // @[MockArray.scala 36:52]
    .clock(ces_50_0_clock),
    .io_ins_0(ces_50_0_io_ins_0),
    .io_ins_1(ces_50_0_io_ins_1),
    .io_ins_2(ces_50_0_io_ins_2),
    .io_ins_3(ces_50_0_io_ins_3),
    .io_outs_0(ces_50_0_io_outs_0),
    .io_outs_1(ces_50_0_io_outs_1),
    .io_outs_2(ces_50_0_io_outs_2),
    .io_outs_3(ces_50_0_io_outs_3)
  );
  Element ces_51_0 ( // @[MockArray.scala 36:52]
    .clock(ces_51_0_clock),
    .io_ins_0(ces_51_0_io_ins_0),
    .io_ins_1(ces_51_0_io_ins_1),
    .io_ins_2(ces_51_0_io_ins_2),
    .io_ins_3(ces_51_0_io_ins_3),
    .io_outs_0(ces_51_0_io_outs_0),
    .io_outs_1(ces_51_0_io_outs_1),
    .io_outs_2(ces_51_0_io_outs_2),
    .io_outs_3(ces_51_0_io_outs_3)
  );
  Element ces_52_0 ( // @[MockArray.scala 36:52]
    .clock(ces_52_0_clock),
    .io_ins_0(ces_52_0_io_ins_0),
    .io_ins_1(ces_52_0_io_ins_1),
    .io_ins_2(ces_52_0_io_ins_2),
    .io_ins_3(ces_52_0_io_ins_3),
    .io_outs_0(ces_52_0_io_outs_0),
    .io_outs_1(ces_52_0_io_outs_1),
    .io_outs_2(ces_52_0_io_outs_2),
    .io_outs_3(ces_52_0_io_outs_3)
  );
  Element ces_53_0 ( // @[MockArray.scala 36:52]
    .clock(ces_53_0_clock),
    .io_ins_0(ces_53_0_io_ins_0),
    .io_ins_1(ces_53_0_io_ins_1),
    .io_ins_2(ces_53_0_io_ins_2),
    .io_ins_3(ces_53_0_io_ins_3),
    .io_outs_0(ces_53_0_io_outs_0),
    .io_outs_1(ces_53_0_io_outs_1),
    .io_outs_2(ces_53_0_io_outs_2),
    .io_outs_3(ces_53_0_io_outs_3)
  );
  Element ces_54_0 ( // @[MockArray.scala 36:52]
    .clock(ces_54_0_clock),
    .io_ins_0(ces_54_0_io_ins_0),
    .io_ins_1(ces_54_0_io_ins_1),
    .io_ins_2(ces_54_0_io_ins_2),
    .io_ins_3(ces_54_0_io_ins_3),
    .io_outs_0(ces_54_0_io_outs_0),
    .io_outs_1(ces_54_0_io_outs_1),
    .io_outs_2(ces_54_0_io_outs_2),
    .io_outs_3(ces_54_0_io_outs_3)
  );
  Element ces_55_0 ( // @[MockArray.scala 36:52]
    .clock(ces_55_0_clock),
    .io_ins_0(ces_55_0_io_ins_0),
    .io_ins_1(ces_55_0_io_ins_1),
    .io_ins_2(ces_55_0_io_ins_2),
    .io_ins_3(ces_55_0_io_ins_3),
    .io_outs_0(ces_55_0_io_outs_0),
    .io_outs_1(ces_55_0_io_outs_1),
    .io_outs_2(ces_55_0_io_outs_2),
    .io_outs_3(ces_55_0_io_outs_3)
  );
  Element ces_56_0 ( // @[MockArray.scala 36:52]
    .clock(ces_56_0_clock),
    .io_ins_0(ces_56_0_io_ins_0),
    .io_ins_1(ces_56_0_io_ins_1),
    .io_ins_2(ces_56_0_io_ins_2),
    .io_ins_3(ces_56_0_io_ins_3),
    .io_outs_0(ces_56_0_io_outs_0),
    .io_outs_1(ces_56_0_io_outs_1),
    .io_outs_2(ces_56_0_io_outs_2),
    .io_outs_3(ces_56_0_io_outs_3)
  );
  Element ces_57_0 ( // @[MockArray.scala 36:52]
    .clock(ces_57_0_clock),
    .io_ins_0(ces_57_0_io_ins_0),
    .io_ins_1(ces_57_0_io_ins_1),
    .io_ins_2(ces_57_0_io_ins_2),
    .io_ins_3(ces_57_0_io_ins_3),
    .io_outs_0(ces_57_0_io_outs_0),
    .io_outs_1(ces_57_0_io_outs_1),
    .io_outs_2(ces_57_0_io_outs_2),
    .io_outs_3(ces_57_0_io_outs_3)
  );
  Element ces_58_0 ( // @[MockArray.scala 36:52]
    .clock(ces_58_0_clock),
    .io_ins_0(ces_58_0_io_ins_0),
    .io_ins_1(ces_58_0_io_ins_1),
    .io_ins_2(ces_58_0_io_ins_2),
    .io_ins_3(ces_58_0_io_ins_3),
    .io_outs_0(ces_58_0_io_outs_0),
    .io_outs_1(ces_58_0_io_outs_1),
    .io_outs_2(ces_58_0_io_outs_2),
    .io_outs_3(ces_58_0_io_outs_3)
  );
  Element ces_59_0 ( // @[MockArray.scala 36:52]
    .clock(ces_59_0_clock),
    .io_ins_0(ces_59_0_io_ins_0),
    .io_ins_1(ces_59_0_io_ins_1),
    .io_ins_2(ces_59_0_io_ins_2),
    .io_ins_3(ces_59_0_io_ins_3),
    .io_outs_0(ces_59_0_io_outs_0),
    .io_outs_1(ces_59_0_io_outs_1),
    .io_outs_2(ces_59_0_io_outs_2),
    .io_outs_3(ces_59_0_io_outs_3)
  );
  Element ces_60_0 ( // @[MockArray.scala 36:52]
    .clock(ces_60_0_clock),
    .io_ins_0(ces_60_0_io_ins_0),
    .io_ins_1(ces_60_0_io_ins_1),
    .io_ins_2(ces_60_0_io_ins_2),
    .io_ins_3(ces_60_0_io_ins_3),
    .io_outs_0(ces_60_0_io_outs_0),
    .io_outs_1(ces_60_0_io_outs_1),
    .io_outs_2(ces_60_0_io_outs_2),
    .io_outs_3(ces_60_0_io_outs_3)
  );
  Element ces_61_0 ( // @[MockArray.scala 36:52]
    .clock(ces_61_0_clock),
    .io_ins_0(ces_61_0_io_ins_0),
    .io_ins_1(ces_61_0_io_ins_1),
    .io_ins_2(ces_61_0_io_ins_2),
    .io_ins_3(ces_61_0_io_ins_3),
    .io_outs_0(ces_61_0_io_outs_0),
    .io_outs_1(ces_61_0_io_outs_1),
    .io_outs_2(ces_61_0_io_outs_2),
    .io_outs_3(ces_61_0_io_outs_3)
  );
  Element ces_62_0 ( // @[MockArray.scala 36:52]
    .clock(ces_62_0_clock),
    .io_ins_0(ces_62_0_io_ins_0),
    .io_ins_1(ces_62_0_io_ins_1),
    .io_ins_2(ces_62_0_io_ins_2),
    .io_ins_3(ces_62_0_io_ins_3),
    .io_outs_0(ces_62_0_io_outs_0),
    .io_outs_1(ces_62_0_io_outs_1),
    .io_outs_2(ces_62_0_io_outs_2),
    .io_outs_3(ces_62_0_io_outs_3)
  );
  Element ces_63_0 ( // @[MockArray.scala 36:52]
    .clock(ces_63_0_clock),
    .io_ins_0(ces_63_0_io_ins_0),
    .io_ins_1(ces_63_0_io_ins_1),
    .io_ins_2(ces_63_0_io_ins_2),
    .io_ins_3(ces_63_0_io_ins_3),
    .io_outs_0(ces_63_0_io_outs_0),
    .io_outs_1(ces_63_0_io_outs_1),
    .io_outs_2(ces_63_0_io_outs_2),
    .io_outs_3(ces_63_0_io_outs_3)
  );
  Element ces_64_0 ( // @[MockArray.scala 36:52]
    .clock(ces_64_0_clock),
    .io_ins_0(ces_64_0_io_ins_0),
    .io_ins_1(ces_64_0_io_ins_1),
    .io_ins_2(ces_64_0_io_ins_2),
    .io_ins_3(ces_64_0_io_ins_3),
    .io_outs_0(ces_64_0_io_outs_0),
    .io_outs_1(ces_64_0_io_outs_1),
    .io_outs_2(ces_64_0_io_outs_2),
    .io_outs_3(ces_64_0_io_outs_3)
  );
  Element ces_65_0 ( // @[MockArray.scala 36:52]
    .clock(ces_65_0_clock),
    .io_ins_0(ces_65_0_io_ins_0),
    .io_ins_1(ces_65_0_io_ins_1),
    .io_ins_2(ces_65_0_io_ins_2),
    .io_ins_3(ces_65_0_io_ins_3),
    .io_outs_0(ces_65_0_io_outs_0),
    .io_outs_1(ces_65_0_io_outs_1),
    .io_outs_2(ces_65_0_io_outs_2),
    .io_outs_3(ces_65_0_io_outs_3)
  );
  Element ces_66_0 ( // @[MockArray.scala 36:52]
    .clock(ces_66_0_clock),
    .io_ins_0(ces_66_0_io_ins_0),
    .io_ins_1(ces_66_0_io_ins_1),
    .io_ins_2(ces_66_0_io_ins_2),
    .io_ins_3(ces_66_0_io_ins_3),
    .io_outs_0(ces_66_0_io_outs_0),
    .io_outs_1(ces_66_0_io_outs_1),
    .io_outs_2(ces_66_0_io_outs_2),
    .io_outs_3(ces_66_0_io_outs_3)
  );
  Element ces_67_0 ( // @[MockArray.scala 36:52]
    .clock(ces_67_0_clock),
    .io_ins_0(ces_67_0_io_ins_0),
    .io_ins_1(ces_67_0_io_ins_1),
    .io_ins_2(ces_67_0_io_ins_2),
    .io_ins_3(ces_67_0_io_ins_3),
    .io_outs_0(ces_67_0_io_outs_0),
    .io_outs_1(ces_67_0_io_outs_1),
    .io_outs_2(ces_67_0_io_outs_2),
    .io_outs_3(ces_67_0_io_outs_3)
  );
  Element ces_68_0 ( // @[MockArray.scala 36:52]
    .clock(ces_68_0_clock),
    .io_ins_0(ces_68_0_io_ins_0),
    .io_ins_1(ces_68_0_io_ins_1),
    .io_ins_2(ces_68_0_io_ins_2),
    .io_ins_3(ces_68_0_io_ins_3),
    .io_outs_0(ces_68_0_io_outs_0),
    .io_outs_1(ces_68_0_io_outs_1),
    .io_outs_2(ces_68_0_io_outs_2),
    .io_outs_3(ces_68_0_io_outs_3)
  );
  Element ces_69_0 ( // @[MockArray.scala 36:52]
    .clock(ces_69_0_clock),
    .io_ins_0(ces_69_0_io_ins_0),
    .io_ins_1(ces_69_0_io_ins_1),
    .io_ins_2(ces_69_0_io_ins_2),
    .io_ins_3(ces_69_0_io_ins_3),
    .io_outs_0(ces_69_0_io_outs_0),
    .io_outs_1(ces_69_0_io_outs_1),
    .io_outs_2(ces_69_0_io_outs_2),
    .io_outs_3(ces_69_0_io_outs_3)
  );
  Element ces_70_0 ( // @[MockArray.scala 36:52]
    .clock(ces_70_0_clock),
    .io_ins_0(ces_70_0_io_ins_0),
    .io_ins_1(ces_70_0_io_ins_1),
    .io_ins_2(ces_70_0_io_ins_2),
    .io_ins_3(ces_70_0_io_ins_3),
    .io_outs_0(ces_70_0_io_outs_0),
    .io_outs_1(ces_70_0_io_outs_1),
    .io_outs_2(ces_70_0_io_outs_2),
    .io_outs_3(ces_70_0_io_outs_3)
  );
  Element ces_71_0 ( // @[MockArray.scala 36:52]
    .clock(ces_71_0_clock),
    .io_ins_0(ces_71_0_io_ins_0),
    .io_ins_1(ces_71_0_io_ins_1),
    .io_ins_2(ces_71_0_io_ins_2),
    .io_ins_3(ces_71_0_io_ins_3),
    .io_outs_0(ces_71_0_io_outs_0),
    .io_outs_1(ces_71_0_io_outs_1),
    .io_outs_2(ces_71_0_io_outs_2),
    .io_outs_3(ces_71_0_io_outs_3)
  );
  Element ces_72_0 ( // @[MockArray.scala 36:52]
    .clock(ces_72_0_clock),
    .io_ins_0(ces_72_0_io_ins_0),
    .io_ins_1(ces_72_0_io_ins_1),
    .io_ins_2(ces_72_0_io_ins_2),
    .io_ins_3(ces_72_0_io_ins_3),
    .io_outs_0(ces_72_0_io_outs_0),
    .io_outs_1(ces_72_0_io_outs_1),
    .io_outs_2(ces_72_0_io_outs_2),
    .io_outs_3(ces_72_0_io_outs_3)
  );
  Element ces_73_0 ( // @[MockArray.scala 36:52]
    .clock(ces_73_0_clock),
    .io_ins_0(ces_73_0_io_ins_0),
    .io_ins_1(ces_73_0_io_ins_1),
    .io_ins_2(ces_73_0_io_ins_2),
    .io_ins_3(ces_73_0_io_ins_3),
    .io_outs_0(ces_73_0_io_outs_0),
    .io_outs_1(ces_73_0_io_outs_1),
    .io_outs_2(ces_73_0_io_outs_2),
    .io_outs_3(ces_73_0_io_outs_3)
  );
  Element ces_74_0 ( // @[MockArray.scala 36:52]
    .clock(ces_74_0_clock),
    .io_ins_0(ces_74_0_io_ins_0),
    .io_ins_1(ces_74_0_io_ins_1),
    .io_ins_2(ces_74_0_io_ins_2),
    .io_ins_3(ces_74_0_io_ins_3),
    .io_outs_0(ces_74_0_io_outs_0),
    .io_outs_1(ces_74_0_io_outs_1),
    .io_outs_2(ces_74_0_io_outs_2),
    .io_outs_3(ces_74_0_io_outs_3)
  );
  Element ces_75_0 ( // @[MockArray.scala 36:52]
    .clock(ces_75_0_clock),
    .io_ins_0(ces_75_0_io_ins_0),
    .io_ins_1(ces_75_0_io_ins_1),
    .io_ins_2(ces_75_0_io_ins_2),
    .io_ins_3(ces_75_0_io_ins_3),
    .io_outs_0(ces_75_0_io_outs_0),
    .io_outs_1(ces_75_0_io_outs_1),
    .io_outs_2(ces_75_0_io_outs_2),
    .io_outs_3(ces_75_0_io_outs_3)
  );
  Element ces_76_0 ( // @[MockArray.scala 36:52]
    .clock(ces_76_0_clock),
    .io_ins_0(ces_76_0_io_ins_0),
    .io_ins_1(ces_76_0_io_ins_1),
    .io_ins_2(ces_76_0_io_ins_2),
    .io_ins_3(ces_76_0_io_ins_3),
    .io_outs_0(ces_76_0_io_outs_0),
    .io_outs_1(ces_76_0_io_outs_1),
    .io_outs_2(ces_76_0_io_outs_2),
    .io_outs_3(ces_76_0_io_outs_3)
  );
  Element ces_77_0 ( // @[MockArray.scala 36:52]
    .clock(ces_77_0_clock),
    .io_ins_0(ces_77_0_io_ins_0),
    .io_ins_1(ces_77_0_io_ins_1),
    .io_ins_2(ces_77_0_io_ins_2),
    .io_ins_3(ces_77_0_io_ins_3),
    .io_outs_0(ces_77_0_io_outs_0),
    .io_outs_1(ces_77_0_io_outs_1),
    .io_outs_2(ces_77_0_io_outs_2),
    .io_outs_3(ces_77_0_io_outs_3)
  );
  Element ces_78_0 ( // @[MockArray.scala 36:52]
    .clock(ces_78_0_clock),
    .io_ins_0(ces_78_0_io_ins_0),
    .io_ins_1(ces_78_0_io_ins_1),
    .io_ins_2(ces_78_0_io_ins_2),
    .io_ins_3(ces_78_0_io_ins_3),
    .io_outs_0(ces_78_0_io_outs_0),
    .io_outs_1(ces_78_0_io_outs_1),
    .io_outs_2(ces_78_0_io_outs_2),
    .io_outs_3(ces_78_0_io_outs_3)
  );
  Element ces_79_0 ( // @[MockArray.scala 36:52]
    .clock(ces_79_0_clock),
    .io_ins_0(ces_79_0_io_ins_0),
    .io_ins_1(ces_79_0_io_ins_1),
    .io_ins_2(ces_79_0_io_ins_2),
    .io_ins_3(ces_79_0_io_ins_3),
    .io_outs_0(ces_79_0_io_outs_0),
    .io_outs_1(ces_79_0_io_outs_1),
    .io_outs_2(ces_79_0_io_outs_2),
    .io_outs_3(ces_79_0_io_outs_3)
  );
  Element ces_80_0 ( // @[MockArray.scala 36:52]
    .clock(ces_80_0_clock),
    .io_ins_0(ces_80_0_io_ins_0),
    .io_ins_1(ces_80_0_io_ins_1),
    .io_ins_2(ces_80_0_io_ins_2),
    .io_ins_3(ces_80_0_io_ins_3),
    .io_outs_0(ces_80_0_io_outs_0),
    .io_outs_1(ces_80_0_io_outs_1),
    .io_outs_2(ces_80_0_io_outs_2),
    .io_outs_3(ces_80_0_io_outs_3)
  );
  Element ces_81_0 ( // @[MockArray.scala 36:52]
    .clock(ces_81_0_clock),
    .io_ins_0(ces_81_0_io_ins_0),
    .io_ins_1(ces_81_0_io_ins_1),
    .io_ins_2(ces_81_0_io_ins_2),
    .io_ins_3(ces_81_0_io_ins_3),
    .io_outs_0(ces_81_0_io_outs_0),
    .io_outs_1(ces_81_0_io_outs_1),
    .io_outs_2(ces_81_0_io_outs_2),
    .io_outs_3(ces_81_0_io_outs_3)
  );
  Element ces_82_0 ( // @[MockArray.scala 36:52]
    .clock(ces_82_0_clock),
    .io_ins_0(ces_82_0_io_ins_0),
    .io_ins_1(ces_82_0_io_ins_1),
    .io_ins_2(ces_82_0_io_ins_2),
    .io_ins_3(ces_82_0_io_ins_3),
    .io_outs_0(ces_82_0_io_outs_0),
    .io_outs_1(ces_82_0_io_outs_1),
    .io_outs_2(ces_82_0_io_outs_2),
    .io_outs_3(ces_82_0_io_outs_3)
  );
  Element ces_83_0 ( // @[MockArray.scala 36:52]
    .clock(ces_83_0_clock),
    .io_ins_0(ces_83_0_io_ins_0),
    .io_ins_1(ces_83_0_io_ins_1),
    .io_ins_2(ces_83_0_io_ins_2),
    .io_ins_3(ces_83_0_io_ins_3),
    .io_outs_0(ces_83_0_io_outs_0),
    .io_outs_1(ces_83_0_io_outs_1),
    .io_outs_2(ces_83_0_io_outs_2),
    .io_outs_3(ces_83_0_io_outs_3)
  );
  Element ces_84_0 ( // @[MockArray.scala 36:52]
    .clock(ces_84_0_clock),
    .io_ins_0(ces_84_0_io_ins_0),
    .io_ins_1(ces_84_0_io_ins_1),
    .io_ins_2(ces_84_0_io_ins_2),
    .io_ins_3(ces_84_0_io_ins_3),
    .io_outs_0(ces_84_0_io_outs_0),
    .io_outs_1(ces_84_0_io_outs_1),
    .io_outs_2(ces_84_0_io_outs_2),
    .io_outs_3(ces_84_0_io_outs_3)
  );
  Element ces_85_0 ( // @[MockArray.scala 36:52]
    .clock(ces_85_0_clock),
    .io_ins_0(ces_85_0_io_ins_0),
    .io_ins_1(ces_85_0_io_ins_1),
    .io_ins_2(ces_85_0_io_ins_2),
    .io_ins_3(ces_85_0_io_ins_3),
    .io_outs_0(ces_85_0_io_outs_0),
    .io_outs_1(ces_85_0_io_outs_1),
    .io_outs_2(ces_85_0_io_outs_2),
    .io_outs_3(ces_85_0_io_outs_3)
  );
  Element ces_86_0 ( // @[MockArray.scala 36:52]
    .clock(ces_86_0_clock),
    .io_ins_0(ces_86_0_io_ins_0),
    .io_ins_1(ces_86_0_io_ins_1),
    .io_ins_2(ces_86_0_io_ins_2),
    .io_ins_3(ces_86_0_io_ins_3),
    .io_outs_0(ces_86_0_io_outs_0),
    .io_outs_1(ces_86_0_io_outs_1),
    .io_outs_2(ces_86_0_io_outs_2),
    .io_outs_3(ces_86_0_io_outs_3)
  );
  Element ces_87_0 ( // @[MockArray.scala 36:52]
    .clock(ces_87_0_clock),
    .io_ins_0(ces_87_0_io_ins_0),
    .io_ins_1(ces_87_0_io_ins_1),
    .io_ins_2(ces_87_0_io_ins_2),
    .io_ins_3(ces_87_0_io_ins_3),
    .io_outs_0(ces_87_0_io_outs_0),
    .io_outs_1(ces_87_0_io_outs_1),
    .io_outs_2(ces_87_0_io_outs_2),
    .io_outs_3(ces_87_0_io_outs_3)
  );
  Element ces_88_0 ( // @[MockArray.scala 36:52]
    .clock(ces_88_0_clock),
    .io_ins_0(ces_88_0_io_ins_0),
    .io_ins_1(ces_88_0_io_ins_1),
    .io_ins_2(ces_88_0_io_ins_2),
    .io_ins_3(ces_88_0_io_ins_3),
    .io_outs_0(ces_88_0_io_outs_0),
    .io_outs_1(ces_88_0_io_outs_1),
    .io_outs_2(ces_88_0_io_outs_2),
    .io_outs_3(ces_88_0_io_outs_3)
  );
  Element ces_89_0 ( // @[MockArray.scala 36:52]
    .clock(ces_89_0_clock),
    .io_ins_0(ces_89_0_io_ins_0),
    .io_ins_1(ces_89_0_io_ins_1),
    .io_ins_2(ces_89_0_io_ins_2),
    .io_ins_3(ces_89_0_io_ins_3),
    .io_outs_0(ces_89_0_io_outs_0),
    .io_outs_1(ces_89_0_io_outs_1),
    .io_outs_2(ces_89_0_io_outs_2),
    .io_outs_3(ces_89_0_io_outs_3)
  );
  Element ces_90_0 ( // @[MockArray.scala 36:52]
    .clock(ces_90_0_clock),
    .io_ins_0(ces_90_0_io_ins_0),
    .io_ins_1(ces_90_0_io_ins_1),
    .io_ins_2(ces_90_0_io_ins_2),
    .io_ins_3(ces_90_0_io_ins_3),
    .io_outs_0(ces_90_0_io_outs_0),
    .io_outs_1(ces_90_0_io_outs_1),
    .io_outs_2(ces_90_0_io_outs_2),
    .io_outs_3(ces_90_0_io_outs_3)
  );
  Element ces_91_0 ( // @[MockArray.scala 36:52]
    .clock(ces_91_0_clock),
    .io_ins_0(ces_91_0_io_ins_0),
    .io_ins_1(ces_91_0_io_ins_1),
    .io_ins_2(ces_91_0_io_ins_2),
    .io_ins_3(ces_91_0_io_ins_3),
    .io_outs_0(ces_91_0_io_outs_0),
    .io_outs_1(ces_91_0_io_outs_1),
    .io_outs_2(ces_91_0_io_outs_2),
    .io_outs_3(ces_91_0_io_outs_3)
  );
  Element ces_92_0 ( // @[MockArray.scala 36:52]
    .clock(ces_92_0_clock),
    .io_ins_0(ces_92_0_io_ins_0),
    .io_ins_1(ces_92_0_io_ins_1),
    .io_ins_2(ces_92_0_io_ins_2),
    .io_ins_3(ces_92_0_io_ins_3),
    .io_outs_0(ces_92_0_io_outs_0),
    .io_outs_1(ces_92_0_io_outs_1),
    .io_outs_2(ces_92_0_io_outs_2),
    .io_outs_3(ces_92_0_io_outs_3)
  );
  Element ces_93_0 ( // @[MockArray.scala 36:52]
    .clock(ces_93_0_clock),
    .io_ins_0(ces_93_0_io_ins_0),
    .io_ins_1(ces_93_0_io_ins_1),
    .io_ins_2(ces_93_0_io_ins_2),
    .io_ins_3(ces_93_0_io_ins_3),
    .io_outs_0(ces_93_0_io_outs_0),
    .io_outs_1(ces_93_0_io_outs_1),
    .io_outs_2(ces_93_0_io_outs_2),
    .io_outs_3(ces_93_0_io_outs_3)
  );
  Element ces_94_0 ( // @[MockArray.scala 36:52]
    .clock(ces_94_0_clock),
    .io_ins_0(ces_94_0_io_ins_0),
    .io_ins_1(ces_94_0_io_ins_1),
    .io_ins_2(ces_94_0_io_ins_2),
    .io_ins_3(ces_94_0_io_ins_3),
    .io_outs_0(ces_94_0_io_outs_0),
    .io_outs_1(ces_94_0_io_outs_1),
    .io_outs_2(ces_94_0_io_outs_2),
    .io_outs_3(ces_94_0_io_outs_3)
  );
  Element ces_95_0 ( // @[MockArray.scala 36:52]
    .clock(ces_95_0_clock),
    .io_ins_0(ces_95_0_io_ins_0),
    .io_ins_1(ces_95_0_io_ins_1),
    .io_ins_2(ces_95_0_io_ins_2),
    .io_ins_3(ces_95_0_io_ins_3),
    .io_outs_0(ces_95_0_io_outs_0),
    .io_outs_1(ces_95_0_io_outs_1),
    .io_outs_2(ces_95_0_io_outs_2),
    .io_outs_3(ces_95_0_io_outs_3)
  );
  Element ces_96_0 ( // @[MockArray.scala 36:52]
    .clock(ces_96_0_clock),
    .io_ins_0(ces_96_0_io_ins_0),
    .io_ins_1(ces_96_0_io_ins_1),
    .io_ins_2(ces_96_0_io_ins_2),
    .io_ins_3(ces_96_0_io_ins_3),
    .io_outs_0(ces_96_0_io_outs_0),
    .io_outs_1(ces_96_0_io_outs_1),
    .io_outs_2(ces_96_0_io_outs_2),
    .io_outs_3(ces_96_0_io_outs_3)
  );
  Element ces_97_0 ( // @[MockArray.scala 36:52]
    .clock(ces_97_0_clock),
    .io_ins_0(ces_97_0_io_ins_0),
    .io_ins_1(ces_97_0_io_ins_1),
    .io_ins_2(ces_97_0_io_ins_2),
    .io_ins_3(ces_97_0_io_ins_3),
    .io_outs_0(ces_97_0_io_outs_0),
    .io_outs_1(ces_97_0_io_outs_1),
    .io_outs_2(ces_97_0_io_outs_2),
    .io_outs_3(ces_97_0_io_outs_3)
  );
  Element ces_98_0 ( // @[MockArray.scala 36:52]
    .clock(ces_98_0_clock),
    .io_ins_0(ces_98_0_io_ins_0),
    .io_ins_1(ces_98_0_io_ins_1),
    .io_ins_2(ces_98_0_io_ins_2),
    .io_ins_3(ces_98_0_io_ins_3),
    .io_outs_0(ces_98_0_io_outs_0),
    .io_outs_1(ces_98_0_io_outs_1),
    .io_outs_2(ces_98_0_io_outs_2),
    .io_outs_3(ces_98_0_io_outs_3)
  );
  Element ces_99_0 ( // @[MockArray.scala 36:52]
    .clock(ces_99_0_clock),
    .io_ins_0(ces_99_0_io_ins_0),
    .io_ins_1(ces_99_0_io_ins_1),
    .io_ins_2(ces_99_0_io_ins_2),
    .io_ins_3(ces_99_0_io_ins_3),
    .io_outs_0(ces_99_0_io_outs_0),
    .io_outs_1(ces_99_0_io_outs_1),
    .io_outs_2(ces_99_0_io_outs_2),
    .io_outs_3(ces_99_0_io_outs_3)
  );
  Element ces_100_0 ( // @[MockArray.scala 36:52]
    .clock(ces_100_0_clock),
    .io_ins_0(ces_100_0_io_ins_0),
    .io_ins_1(ces_100_0_io_ins_1),
    .io_ins_2(ces_100_0_io_ins_2),
    .io_ins_3(ces_100_0_io_ins_3),
    .io_outs_0(ces_100_0_io_outs_0),
    .io_outs_1(ces_100_0_io_outs_1),
    .io_outs_2(ces_100_0_io_outs_2),
    .io_outs_3(ces_100_0_io_outs_3)
  );
  Element ces_101_0 ( // @[MockArray.scala 36:52]
    .clock(ces_101_0_clock),
    .io_ins_0(ces_101_0_io_ins_0),
    .io_ins_1(ces_101_0_io_ins_1),
    .io_ins_2(ces_101_0_io_ins_2),
    .io_ins_3(ces_101_0_io_ins_3),
    .io_outs_0(ces_101_0_io_outs_0),
    .io_outs_1(ces_101_0_io_outs_1),
    .io_outs_2(ces_101_0_io_outs_2),
    .io_outs_3(ces_101_0_io_outs_3)
  );
  Element ces_102_0 ( // @[MockArray.scala 36:52]
    .clock(ces_102_0_clock),
    .io_ins_0(ces_102_0_io_ins_0),
    .io_ins_1(ces_102_0_io_ins_1),
    .io_ins_2(ces_102_0_io_ins_2),
    .io_ins_3(ces_102_0_io_ins_3),
    .io_outs_0(ces_102_0_io_outs_0),
    .io_outs_1(ces_102_0_io_outs_1),
    .io_outs_2(ces_102_0_io_outs_2),
    .io_outs_3(ces_102_0_io_outs_3)
  );
  Element ces_103_0 ( // @[MockArray.scala 36:52]
    .clock(ces_103_0_clock),
    .io_ins_0(ces_103_0_io_ins_0),
    .io_ins_1(ces_103_0_io_ins_1),
    .io_ins_2(ces_103_0_io_ins_2),
    .io_ins_3(ces_103_0_io_ins_3),
    .io_outs_0(ces_103_0_io_outs_0),
    .io_outs_1(ces_103_0_io_outs_1),
    .io_outs_2(ces_103_0_io_outs_2),
    .io_outs_3(ces_103_0_io_outs_3)
  );
  Element ces_104_0 ( // @[MockArray.scala 36:52]
    .clock(ces_104_0_clock),
    .io_ins_0(ces_104_0_io_ins_0),
    .io_ins_1(ces_104_0_io_ins_1),
    .io_ins_2(ces_104_0_io_ins_2),
    .io_ins_3(ces_104_0_io_ins_3),
    .io_outs_0(ces_104_0_io_outs_0),
    .io_outs_1(ces_104_0_io_outs_1),
    .io_outs_2(ces_104_0_io_outs_2),
    .io_outs_3(ces_104_0_io_outs_3)
  );
  Element ces_105_0 ( // @[MockArray.scala 36:52]
    .clock(ces_105_0_clock),
    .io_ins_0(ces_105_0_io_ins_0),
    .io_ins_1(ces_105_0_io_ins_1),
    .io_ins_2(ces_105_0_io_ins_2),
    .io_ins_3(ces_105_0_io_ins_3),
    .io_outs_0(ces_105_0_io_outs_0),
    .io_outs_1(ces_105_0_io_outs_1),
    .io_outs_2(ces_105_0_io_outs_2),
    .io_outs_3(ces_105_0_io_outs_3)
  );
  Element ces_106_0 ( // @[MockArray.scala 36:52]
    .clock(ces_106_0_clock),
    .io_ins_0(ces_106_0_io_ins_0),
    .io_ins_1(ces_106_0_io_ins_1),
    .io_ins_2(ces_106_0_io_ins_2),
    .io_ins_3(ces_106_0_io_ins_3),
    .io_outs_0(ces_106_0_io_outs_0),
    .io_outs_1(ces_106_0_io_outs_1),
    .io_outs_2(ces_106_0_io_outs_2),
    .io_outs_3(ces_106_0_io_outs_3)
  );
  Element ces_107_0 ( // @[MockArray.scala 36:52]
    .clock(ces_107_0_clock),
    .io_ins_0(ces_107_0_io_ins_0),
    .io_ins_1(ces_107_0_io_ins_1),
    .io_ins_2(ces_107_0_io_ins_2),
    .io_ins_3(ces_107_0_io_ins_3),
    .io_outs_0(ces_107_0_io_outs_0),
    .io_outs_1(ces_107_0_io_outs_1),
    .io_outs_2(ces_107_0_io_outs_2),
    .io_outs_3(ces_107_0_io_outs_3)
  );
  Element ces_108_0 ( // @[MockArray.scala 36:52]
    .clock(ces_108_0_clock),
    .io_ins_0(ces_108_0_io_ins_0),
    .io_ins_1(ces_108_0_io_ins_1),
    .io_ins_2(ces_108_0_io_ins_2),
    .io_ins_3(ces_108_0_io_ins_3),
    .io_outs_0(ces_108_0_io_outs_0),
    .io_outs_1(ces_108_0_io_outs_1),
    .io_outs_2(ces_108_0_io_outs_2),
    .io_outs_3(ces_108_0_io_outs_3)
  );
  Element ces_109_0 ( // @[MockArray.scala 36:52]
    .clock(ces_109_0_clock),
    .io_ins_0(ces_109_0_io_ins_0),
    .io_ins_1(ces_109_0_io_ins_1),
    .io_ins_2(ces_109_0_io_ins_2),
    .io_ins_3(ces_109_0_io_ins_3),
    .io_outs_0(ces_109_0_io_outs_0),
    .io_outs_1(ces_109_0_io_outs_1),
    .io_outs_2(ces_109_0_io_outs_2),
    .io_outs_3(ces_109_0_io_outs_3)
  );
  Element ces_110_0 ( // @[MockArray.scala 36:52]
    .clock(ces_110_0_clock),
    .io_ins_0(ces_110_0_io_ins_0),
    .io_ins_1(ces_110_0_io_ins_1),
    .io_ins_2(ces_110_0_io_ins_2),
    .io_ins_3(ces_110_0_io_ins_3),
    .io_outs_0(ces_110_0_io_outs_0),
    .io_outs_1(ces_110_0_io_outs_1),
    .io_outs_2(ces_110_0_io_outs_2),
    .io_outs_3(ces_110_0_io_outs_3)
  );
  Element ces_111_0 ( // @[MockArray.scala 36:52]
    .clock(ces_111_0_clock),
    .io_ins_0(ces_111_0_io_ins_0),
    .io_ins_1(ces_111_0_io_ins_1),
    .io_ins_2(ces_111_0_io_ins_2),
    .io_ins_3(ces_111_0_io_ins_3),
    .io_outs_0(ces_111_0_io_outs_0),
    .io_outs_1(ces_111_0_io_outs_1),
    .io_outs_2(ces_111_0_io_outs_2),
    .io_outs_3(ces_111_0_io_outs_3)
  );
  Element ces_112_0 ( // @[MockArray.scala 36:52]
    .clock(ces_112_0_clock),
    .io_ins_0(ces_112_0_io_ins_0),
    .io_ins_1(ces_112_0_io_ins_1),
    .io_ins_2(ces_112_0_io_ins_2),
    .io_ins_3(ces_112_0_io_ins_3),
    .io_outs_0(ces_112_0_io_outs_0),
    .io_outs_1(ces_112_0_io_outs_1),
    .io_outs_2(ces_112_0_io_outs_2),
    .io_outs_3(ces_112_0_io_outs_3)
  );
  Element ces_113_0 ( // @[MockArray.scala 36:52]
    .clock(ces_113_0_clock),
    .io_ins_0(ces_113_0_io_ins_0),
    .io_ins_1(ces_113_0_io_ins_1),
    .io_ins_2(ces_113_0_io_ins_2),
    .io_ins_3(ces_113_0_io_ins_3),
    .io_outs_0(ces_113_0_io_outs_0),
    .io_outs_1(ces_113_0_io_outs_1),
    .io_outs_2(ces_113_0_io_outs_2),
    .io_outs_3(ces_113_0_io_outs_3)
  );
  Element ces_114_0 ( // @[MockArray.scala 36:52]
    .clock(ces_114_0_clock),
    .io_ins_0(ces_114_0_io_ins_0),
    .io_ins_1(ces_114_0_io_ins_1),
    .io_ins_2(ces_114_0_io_ins_2),
    .io_ins_3(ces_114_0_io_ins_3),
    .io_outs_0(ces_114_0_io_outs_0),
    .io_outs_1(ces_114_0_io_outs_1),
    .io_outs_2(ces_114_0_io_outs_2),
    .io_outs_3(ces_114_0_io_outs_3)
  );
  Element ces_115_0 ( // @[MockArray.scala 36:52]
    .clock(ces_115_0_clock),
    .io_ins_0(ces_115_0_io_ins_0),
    .io_ins_1(ces_115_0_io_ins_1),
    .io_ins_2(ces_115_0_io_ins_2),
    .io_ins_3(ces_115_0_io_ins_3),
    .io_outs_0(ces_115_0_io_outs_0),
    .io_outs_1(ces_115_0_io_outs_1),
    .io_outs_2(ces_115_0_io_outs_2),
    .io_outs_3(ces_115_0_io_outs_3)
  );
  Element ces_116_0 ( // @[MockArray.scala 36:52]
    .clock(ces_116_0_clock),
    .io_ins_0(ces_116_0_io_ins_0),
    .io_ins_1(ces_116_0_io_ins_1),
    .io_ins_2(ces_116_0_io_ins_2),
    .io_ins_3(ces_116_0_io_ins_3),
    .io_outs_0(ces_116_0_io_outs_0),
    .io_outs_1(ces_116_0_io_outs_1),
    .io_outs_2(ces_116_0_io_outs_2),
    .io_outs_3(ces_116_0_io_outs_3)
  );
  Element ces_117_0 ( // @[MockArray.scala 36:52]
    .clock(ces_117_0_clock),
    .io_ins_0(ces_117_0_io_ins_0),
    .io_ins_1(ces_117_0_io_ins_1),
    .io_ins_2(ces_117_0_io_ins_2),
    .io_ins_3(ces_117_0_io_ins_3),
    .io_outs_0(ces_117_0_io_outs_0),
    .io_outs_1(ces_117_0_io_outs_1),
    .io_outs_2(ces_117_0_io_outs_2),
    .io_outs_3(ces_117_0_io_outs_3)
  );
  Element ces_118_0 ( // @[MockArray.scala 36:52]
    .clock(ces_118_0_clock),
    .io_ins_0(ces_118_0_io_ins_0),
    .io_ins_1(ces_118_0_io_ins_1),
    .io_ins_2(ces_118_0_io_ins_2),
    .io_ins_3(ces_118_0_io_ins_3),
    .io_outs_0(ces_118_0_io_outs_0),
    .io_outs_1(ces_118_0_io_outs_1),
    .io_outs_2(ces_118_0_io_outs_2),
    .io_outs_3(ces_118_0_io_outs_3)
  );
  Element ces_119_0 ( // @[MockArray.scala 36:52]
    .clock(ces_119_0_clock),
    .io_ins_0(ces_119_0_io_ins_0),
    .io_ins_1(ces_119_0_io_ins_1),
    .io_ins_2(ces_119_0_io_ins_2),
    .io_ins_3(ces_119_0_io_ins_3),
    .io_outs_0(ces_119_0_io_outs_0),
    .io_outs_1(ces_119_0_io_outs_1),
    .io_outs_2(ces_119_0_io_outs_2),
    .io_outs_3(ces_119_0_io_outs_3)
  );
  Element ces_120_0 ( // @[MockArray.scala 36:52]
    .clock(ces_120_0_clock),
    .io_ins_0(ces_120_0_io_ins_0),
    .io_ins_1(ces_120_0_io_ins_1),
    .io_ins_2(ces_120_0_io_ins_2),
    .io_ins_3(ces_120_0_io_ins_3),
    .io_outs_0(ces_120_0_io_outs_0),
    .io_outs_1(ces_120_0_io_outs_1),
    .io_outs_2(ces_120_0_io_outs_2),
    .io_outs_3(ces_120_0_io_outs_3)
  );
  Element ces_121_0 ( // @[MockArray.scala 36:52]
    .clock(ces_121_0_clock),
    .io_ins_0(ces_121_0_io_ins_0),
    .io_ins_1(ces_121_0_io_ins_1),
    .io_ins_2(ces_121_0_io_ins_2),
    .io_ins_3(ces_121_0_io_ins_3),
    .io_outs_0(ces_121_0_io_outs_0),
    .io_outs_1(ces_121_0_io_outs_1),
    .io_outs_2(ces_121_0_io_outs_2),
    .io_outs_3(ces_121_0_io_outs_3)
  );
  Element ces_122_0 ( // @[MockArray.scala 36:52]
    .clock(ces_122_0_clock),
    .io_ins_0(ces_122_0_io_ins_0),
    .io_ins_1(ces_122_0_io_ins_1),
    .io_ins_2(ces_122_0_io_ins_2),
    .io_ins_3(ces_122_0_io_ins_3),
    .io_outs_0(ces_122_0_io_outs_0),
    .io_outs_1(ces_122_0_io_outs_1),
    .io_outs_2(ces_122_0_io_outs_2),
    .io_outs_3(ces_122_0_io_outs_3)
  );
  Element ces_123_0 ( // @[MockArray.scala 36:52]
    .clock(ces_123_0_clock),
    .io_ins_0(ces_123_0_io_ins_0),
    .io_ins_1(ces_123_0_io_ins_1),
    .io_ins_2(ces_123_0_io_ins_2),
    .io_ins_3(ces_123_0_io_ins_3),
    .io_outs_0(ces_123_0_io_outs_0),
    .io_outs_1(ces_123_0_io_outs_1),
    .io_outs_2(ces_123_0_io_outs_2),
    .io_outs_3(ces_123_0_io_outs_3)
  );
  Element ces_124_0 ( // @[MockArray.scala 36:52]
    .clock(ces_124_0_clock),
    .io_ins_0(ces_124_0_io_ins_0),
    .io_ins_1(ces_124_0_io_ins_1),
    .io_ins_2(ces_124_0_io_ins_2),
    .io_ins_3(ces_124_0_io_ins_3),
    .io_outs_0(ces_124_0_io_outs_0),
    .io_outs_1(ces_124_0_io_outs_1),
    .io_outs_2(ces_124_0_io_outs_2),
    .io_outs_3(ces_124_0_io_outs_3)
  );
  Element ces_125_0 ( // @[MockArray.scala 36:52]
    .clock(ces_125_0_clock),
    .io_ins_0(ces_125_0_io_ins_0),
    .io_ins_1(ces_125_0_io_ins_1),
    .io_ins_2(ces_125_0_io_ins_2),
    .io_ins_3(ces_125_0_io_ins_3),
    .io_outs_0(ces_125_0_io_outs_0),
    .io_outs_1(ces_125_0_io_outs_1),
    .io_outs_2(ces_125_0_io_outs_2),
    .io_outs_3(ces_125_0_io_outs_3)
  );
  Element ces_126_0 ( // @[MockArray.scala 36:52]
    .clock(ces_126_0_clock),
    .io_ins_0(ces_126_0_io_ins_0),
    .io_ins_1(ces_126_0_io_ins_1),
    .io_ins_2(ces_126_0_io_ins_2),
    .io_ins_3(ces_126_0_io_ins_3),
    .io_outs_0(ces_126_0_io_outs_0),
    .io_outs_1(ces_126_0_io_outs_1),
    .io_outs_2(ces_126_0_io_outs_2),
    .io_outs_3(ces_126_0_io_outs_3)
  );
  Element ces_127_0 ( // @[MockArray.scala 36:52]
    .clock(ces_127_0_clock),
    .io_ins_0(ces_127_0_io_ins_0),
    .io_ins_1(ces_127_0_io_ins_1),
    .io_ins_2(ces_127_0_io_ins_2),
    .io_ins_3(ces_127_0_io_ins_3),
    .io_outs_0(ces_127_0_io_outs_0),
    .io_outs_1(ces_127_0_io_outs_1),
    .io_outs_2(ces_127_0_io_outs_2),
    .io_outs_3(ces_127_0_io_outs_3)
  );
  Element ces_128_0 ( // @[MockArray.scala 36:52]
    .clock(ces_128_0_clock),
    .io_ins_0(ces_128_0_io_ins_0),
    .io_ins_1(ces_128_0_io_ins_1),
    .io_ins_2(ces_128_0_io_ins_2),
    .io_ins_3(ces_128_0_io_ins_3),
    .io_outs_0(ces_128_0_io_outs_0),
    .io_outs_1(ces_128_0_io_outs_1),
    .io_outs_2(ces_128_0_io_outs_2),
    .io_outs_3(ces_128_0_io_outs_3)
  );
  Element ces_129_0 ( // @[MockArray.scala 36:52]
    .clock(ces_129_0_clock),
    .io_ins_0(ces_129_0_io_ins_0),
    .io_ins_1(ces_129_0_io_ins_1),
    .io_ins_2(ces_129_0_io_ins_2),
    .io_ins_3(ces_129_0_io_ins_3),
    .io_outs_0(ces_129_0_io_outs_0),
    .io_outs_1(ces_129_0_io_outs_1),
    .io_outs_2(ces_129_0_io_outs_2),
    .io_outs_3(ces_129_0_io_outs_3)
  );
  Element ces_130_0 ( // @[MockArray.scala 36:52]
    .clock(ces_130_0_clock),
    .io_ins_0(ces_130_0_io_ins_0),
    .io_ins_1(ces_130_0_io_ins_1),
    .io_ins_2(ces_130_0_io_ins_2),
    .io_ins_3(ces_130_0_io_ins_3),
    .io_outs_0(ces_130_0_io_outs_0),
    .io_outs_1(ces_130_0_io_outs_1),
    .io_outs_2(ces_130_0_io_outs_2),
    .io_outs_3(ces_130_0_io_outs_3)
  );
  Element ces_131_0 ( // @[MockArray.scala 36:52]
    .clock(ces_131_0_clock),
    .io_ins_0(ces_131_0_io_ins_0),
    .io_ins_1(ces_131_0_io_ins_1),
    .io_ins_2(ces_131_0_io_ins_2),
    .io_ins_3(ces_131_0_io_ins_3),
    .io_outs_0(ces_131_0_io_outs_0),
    .io_outs_1(ces_131_0_io_outs_1),
    .io_outs_2(ces_131_0_io_outs_2),
    .io_outs_3(ces_131_0_io_outs_3)
  );
  Element ces_132_0 ( // @[MockArray.scala 36:52]
    .clock(ces_132_0_clock),
    .io_ins_0(ces_132_0_io_ins_0),
    .io_ins_1(ces_132_0_io_ins_1),
    .io_ins_2(ces_132_0_io_ins_2),
    .io_ins_3(ces_132_0_io_ins_3),
    .io_outs_0(ces_132_0_io_outs_0),
    .io_outs_1(ces_132_0_io_outs_1),
    .io_outs_2(ces_132_0_io_outs_2),
    .io_outs_3(ces_132_0_io_outs_3)
  );
  Element ces_133_0 ( // @[MockArray.scala 36:52]
    .clock(ces_133_0_clock),
    .io_ins_0(ces_133_0_io_ins_0),
    .io_ins_1(ces_133_0_io_ins_1),
    .io_ins_2(ces_133_0_io_ins_2),
    .io_ins_3(ces_133_0_io_ins_3),
    .io_outs_0(ces_133_0_io_outs_0),
    .io_outs_1(ces_133_0_io_outs_1),
    .io_outs_2(ces_133_0_io_outs_2),
    .io_outs_3(ces_133_0_io_outs_3)
  );
  Element ces_134_0 ( // @[MockArray.scala 36:52]
    .clock(ces_134_0_clock),
    .io_ins_0(ces_134_0_io_ins_0),
    .io_ins_1(ces_134_0_io_ins_1),
    .io_ins_2(ces_134_0_io_ins_2),
    .io_ins_3(ces_134_0_io_ins_3),
    .io_outs_0(ces_134_0_io_outs_0),
    .io_outs_1(ces_134_0_io_outs_1),
    .io_outs_2(ces_134_0_io_outs_2),
    .io_outs_3(ces_134_0_io_outs_3)
  );
  Element ces_135_0 ( // @[MockArray.scala 36:52]
    .clock(ces_135_0_clock),
    .io_ins_0(ces_135_0_io_ins_0),
    .io_ins_1(ces_135_0_io_ins_1),
    .io_ins_2(ces_135_0_io_ins_2),
    .io_ins_3(ces_135_0_io_ins_3),
    .io_outs_0(ces_135_0_io_outs_0),
    .io_outs_1(ces_135_0_io_outs_1),
    .io_outs_2(ces_135_0_io_outs_2),
    .io_outs_3(ces_135_0_io_outs_3)
  );
  Element ces_136_0 ( // @[MockArray.scala 36:52]
    .clock(ces_136_0_clock),
    .io_ins_0(ces_136_0_io_ins_0),
    .io_ins_1(ces_136_0_io_ins_1),
    .io_ins_2(ces_136_0_io_ins_2),
    .io_ins_3(ces_136_0_io_ins_3),
    .io_outs_0(ces_136_0_io_outs_0),
    .io_outs_1(ces_136_0_io_outs_1),
    .io_outs_2(ces_136_0_io_outs_2),
    .io_outs_3(ces_136_0_io_outs_3)
  );
  Element ces_137_0 ( // @[MockArray.scala 36:52]
    .clock(ces_137_0_clock),
    .io_ins_0(ces_137_0_io_ins_0),
    .io_ins_1(ces_137_0_io_ins_1),
    .io_ins_2(ces_137_0_io_ins_2),
    .io_ins_3(ces_137_0_io_ins_3),
    .io_outs_0(ces_137_0_io_outs_0),
    .io_outs_1(ces_137_0_io_outs_1),
    .io_outs_2(ces_137_0_io_outs_2),
    .io_outs_3(ces_137_0_io_outs_3)
  );
  Element ces_138_0 ( // @[MockArray.scala 36:52]
    .clock(ces_138_0_clock),
    .io_ins_0(ces_138_0_io_ins_0),
    .io_ins_1(ces_138_0_io_ins_1),
    .io_ins_2(ces_138_0_io_ins_2),
    .io_ins_3(ces_138_0_io_ins_3),
    .io_outs_0(ces_138_0_io_outs_0),
    .io_outs_1(ces_138_0_io_outs_1),
    .io_outs_2(ces_138_0_io_outs_2),
    .io_outs_3(ces_138_0_io_outs_3)
  );
  Element ces_139_0 ( // @[MockArray.scala 36:52]
    .clock(ces_139_0_clock),
    .io_ins_0(ces_139_0_io_ins_0),
    .io_ins_1(ces_139_0_io_ins_1),
    .io_ins_2(ces_139_0_io_ins_2),
    .io_ins_3(ces_139_0_io_ins_3),
    .io_outs_0(ces_139_0_io_outs_0),
    .io_outs_1(ces_139_0_io_outs_1),
    .io_outs_2(ces_139_0_io_outs_2),
    .io_outs_3(ces_139_0_io_outs_3)
  );
  Element ces_140_0 ( // @[MockArray.scala 36:52]
    .clock(ces_140_0_clock),
    .io_ins_0(ces_140_0_io_ins_0),
    .io_ins_1(ces_140_0_io_ins_1),
    .io_ins_2(ces_140_0_io_ins_2),
    .io_ins_3(ces_140_0_io_ins_3),
    .io_outs_0(ces_140_0_io_outs_0),
    .io_outs_1(ces_140_0_io_outs_1),
    .io_outs_2(ces_140_0_io_outs_2),
    .io_outs_3(ces_140_0_io_outs_3)
  );
  Element ces_141_0 ( // @[MockArray.scala 36:52]
    .clock(ces_141_0_clock),
    .io_ins_0(ces_141_0_io_ins_0),
    .io_ins_1(ces_141_0_io_ins_1),
    .io_ins_2(ces_141_0_io_ins_2),
    .io_ins_3(ces_141_0_io_ins_3),
    .io_outs_0(ces_141_0_io_outs_0),
    .io_outs_1(ces_141_0_io_outs_1),
    .io_outs_2(ces_141_0_io_outs_2),
    .io_outs_3(ces_141_0_io_outs_3)
  );
  Element ces_142_0 ( // @[MockArray.scala 36:52]
    .clock(ces_142_0_clock),
    .io_ins_0(ces_142_0_io_ins_0),
    .io_ins_1(ces_142_0_io_ins_1),
    .io_ins_2(ces_142_0_io_ins_2),
    .io_ins_3(ces_142_0_io_ins_3),
    .io_outs_0(ces_142_0_io_outs_0),
    .io_outs_1(ces_142_0_io_outs_1),
    .io_outs_2(ces_142_0_io_outs_2),
    .io_outs_3(ces_142_0_io_outs_3)
  );
  Element ces_143_0 ( // @[MockArray.scala 36:52]
    .clock(ces_143_0_clock),
    .io_ins_0(ces_143_0_io_ins_0),
    .io_ins_1(ces_143_0_io_ins_1),
    .io_ins_2(ces_143_0_io_ins_2),
    .io_ins_3(ces_143_0_io_ins_3),
    .io_outs_0(ces_143_0_io_outs_0),
    .io_outs_1(ces_143_0_io_outs_1),
    .io_outs_2(ces_143_0_io_outs_2),
    .io_outs_3(ces_143_0_io_outs_3)
  );
  Element ces_144_0 ( // @[MockArray.scala 36:52]
    .clock(ces_144_0_clock),
    .io_ins_0(ces_144_0_io_ins_0),
    .io_ins_1(ces_144_0_io_ins_1),
    .io_ins_2(ces_144_0_io_ins_2),
    .io_ins_3(ces_144_0_io_ins_3),
    .io_outs_0(ces_144_0_io_outs_0),
    .io_outs_1(ces_144_0_io_outs_1),
    .io_outs_2(ces_144_0_io_outs_2),
    .io_outs_3(ces_144_0_io_outs_3)
  );
  Element ces_145_0 ( // @[MockArray.scala 36:52]
    .clock(ces_145_0_clock),
    .io_ins_0(ces_145_0_io_ins_0),
    .io_ins_1(ces_145_0_io_ins_1),
    .io_ins_2(ces_145_0_io_ins_2),
    .io_ins_3(ces_145_0_io_ins_3),
    .io_outs_0(ces_145_0_io_outs_0),
    .io_outs_1(ces_145_0_io_outs_1),
    .io_outs_2(ces_145_0_io_outs_2),
    .io_outs_3(ces_145_0_io_outs_3)
  );
  Element ces_146_0 ( // @[MockArray.scala 36:52]
    .clock(ces_146_0_clock),
    .io_ins_0(ces_146_0_io_ins_0),
    .io_ins_1(ces_146_0_io_ins_1),
    .io_ins_2(ces_146_0_io_ins_2),
    .io_ins_3(ces_146_0_io_ins_3),
    .io_outs_0(ces_146_0_io_outs_0),
    .io_outs_1(ces_146_0_io_outs_1),
    .io_outs_2(ces_146_0_io_outs_2),
    .io_outs_3(ces_146_0_io_outs_3)
  );
  Element ces_147_0 ( // @[MockArray.scala 36:52]
    .clock(ces_147_0_clock),
    .io_ins_0(ces_147_0_io_ins_0),
    .io_ins_1(ces_147_0_io_ins_1),
    .io_ins_2(ces_147_0_io_ins_2),
    .io_ins_3(ces_147_0_io_ins_3),
    .io_outs_0(ces_147_0_io_outs_0),
    .io_outs_1(ces_147_0_io_outs_1),
    .io_outs_2(ces_147_0_io_outs_2),
    .io_outs_3(ces_147_0_io_outs_3)
  );
  Element ces_148_0 ( // @[MockArray.scala 36:52]
    .clock(ces_148_0_clock),
    .io_ins_0(ces_148_0_io_ins_0),
    .io_ins_1(ces_148_0_io_ins_1),
    .io_ins_2(ces_148_0_io_ins_2),
    .io_ins_3(ces_148_0_io_ins_3),
    .io_outs_0(ces_148_0_io_outs_0),
    .io_outs_1(ces_148_0_io_outs_1),
    .io_outs_2(ces_148_0_io_outs_2),
    .io_outs_3(ces_148_0_io_outs_3)
  );
  Element ces_149_0 ( // @[MockArray.scala 36:52]
    .clock(ces_149_0_clock),
    .io_ins_0(ces_149_0_io_ins_0),
    .io_ins_1(ces_149_0_io_ins_1),
    .io_ins_2(ces_149_0_io_ins_2),
    .io_ins_3(ces_149_0_io_ins_3),
    .io_outs_0(ces_149_0_io_outs_0),
    .io_outs_1(ces_149_0_io_outs_1),
    .io_outs_2(ces_149_0_io_outs_2),
    .io_outs_3(ces_149_0_io_outs_3)
  );
  Element ces_150_0 ( // @[MockArray.scala 36:52]
    .clock(ces_150_0_clock),
    .io_ins_0(ces_150_0_io_ins_0),
    .io_ins_1(ces_150_0_io_ins_1),
    .io_ins_2(ces_150_0_io_ins_2),
    .io_ins_3(ces_150_0_io_ins_3),
    .io_outs_0(ces_150_0_io_outs_0),
    .io_outs_1(ces_150_0_io_outs_1),
    .io_outs_2(ces_150_0_io_outs_2),
    .io_outs_3(ces_150_0_io_outs_3)
  );
  Element ces_151_0 ( // @[MockArray.scala 36:52]
    .clock(ces_151_0_clock),
    .io_ins_0(ces_151_0_io_ins_0),
    .io_ins_1(ces_151_0_io_ins_1),
    .io_ins_2(ces_151_0_io_ins_2),
    .io_ins_3(ces_151_0_io_ins_3),
    .io_outs_0(ces_151_0_io_outs_0),
    .io_outs_1(ces_151_0_io_outs_1),
    .io_outs_2(ces_151_0_io_outs_2),
    .io_outs_3(ces_151_0_io_outs_3)
  );
  Element ces_152_0 ( // @[MockArray.scala 36:52]
    .clock(ces_152_0_clock),
    .io_ins_0(ces_152_0_io_ins_0),
    .io_ins_1(ces_152_0_io_ins_1),
    .io_ins_2(ces_152_0_io_ins_2),
    .io_ins_3(ces_152_0_io_ins_3),
    .io_outs_0(ces_152_0_io_outs_0),
    .io_outs_1(ces_152_0_io_outs_1),
    .io_outs_2(ces_152_0_io_outs_2),
    .io_outs_3(ces_152_0_io_outs_3)
  );
  Element ces_153_0 ( // @[MockArray.scala 36:52]
    .clock(ces_153_0_clock),
    .io_ins_0(ces_153_0_io_ins_0),
    .io_ins_1(ces_153_0_io_ins_1),
    .io_ins_2(ces_153_0_io_ins_2),
    .io_ins_3(ces_153_0_io_ins_3),
    .io_outs_0(ces_153_0_io_outs_0),
    .io_outs_1(ces_153_0_io_outs_1),
    .io_outs_2(ces_153_0_io_outs_2),
    .io_outs_3(ces_153_0_io_outs_3)
  );
  Element ces_154_0 ( // @[MockArray.scala 36:52]
    .clock(ces_154_0_clock),
    .io_ins_0(ces_154_0_io_ins_0),
    .io_ins_1(ces_154_0_io_ins_1),
    .io_ins_2(ces_154_0_io_ins_2),
    .io_ins_3(ces_154_0_io_ins_3),
    .io_outs_0(ces_154_0_io_outs_0),
    .io_outs_1(ces_154_0_io_outs_1),
    .io_outs_2(ces_154_0_io_outs_2),
    .io_outs_3(ces_154_0_io_outs_3)
  );
  Element ces_155_0 ( // @[MockArray.scala 36:52]
    .clock(ces_155_0_clock),
    .io_ins_0(ces_155_0_io_ins_0),
    .io_ins_1(ces_155_0_io_ins_1),
    .io_ins_2(ces_155_0_io_ins_2),
    .io_ins_3(ces_155_0_io_ins_3),
    .io_outs_0(ces_155_0_io_outs_0),
    .io_outs_1(ces_155_0_io_outs_1),
    .io_outs_2(ces_155_0_io_outs_2),
    .io_outs_3(ces_155_0_io_outs_3)
  );
  Element ces_156_0 ( // @[MockArray.scala 36:52]
    .clock(ces_156_0_clock),
    .io_ins_0(ces_156_0_io_ins_0),
    .io_ins_1(ces_156_0_io_ins_1),
    .io_ins_2(ces_156_0_io_ins_2),
    .io_ins_3(ces_156_0_io_ins_3),
    .io_outs_0(ces_156_0_io_outs_0),
    .io_outs_1(ces_156_0_io_outs_1),
    .io_outs_2(ces_156_0_io_outs_2),
    .io_outs_3(ces_156_0_io_outs_3)
  );
  Element ces_157_0 ( // @[MockArray.scala 36:52]
    .clock(ces_157_0_clock),
    .io_ins_0(ces_157_0_io_ins_0),
    .io_ins_1(ces_157_0_io_ins_1),
    .io_ins_2(ces_157_0_io_ins_2),
    .io_ins_3(ces_157_0_io_ins_3),
    .io_outs_0(ces_157_0_io_outs_0),
    .io_outs_1(ces_157_0_io_outs_1),
    .io_outs_2(ces_157_0_io_outs_2),
    .io_outs_3(ces_157_0_io_outs_3)
  );
  Element ces_158_0 ( // @[MockArray.scala 36:52]
    .clock(ces_158_0_clock),
    .io_ins_0(ces_158_0_io_ins_0),
    .io_ins_1(ces_158_0_io_ins_1),
    .io_ins_2(ces_158_0_io_ins_2),
    .io_ins_3(ces_158_0_io_ins_3),
    .io_outs_0(ces_158_0_io_outs_0),
    .io_outs_1(ces_158_0_io_outs_1),
    .io_outs_2(ces_158_0_io_outs_2),
    .io_outs_3(ces_158_0_io_outs_3)
  );
  Element ces_159_0 ( // @[MockArray.scala 36:52]
    .clock(ces_159_0_clock),
    .io_ins_0(ces_159_0_io_ins_0),
    .io_ins_1(ces_159_0_io_ins_1),
    .io_ins_2(ces_159_0_io_ins_2),
    .io_ins_3(ces_159_0_io_ins_3),
    .io_outs_0(ces_159_0_io_outs_0),
    .io_outs_1(ces_159_0_io_outs_1),
    .io_outs_2(ces_159_0_io_outs_2),
    .io_outs_3(ces_159_0_io_outs_3)
  );
  Element ces_160_0 ( // @[MockArray.scala 36:52]
    .clock(ces_160_0_clock),
    .io_ins_0(ces_160_0_io_ins_0),
    .io_ins_1(ces_160_0_io_ins_1),
    .io_ins_2(ces_160_0_io_ins_2),
    .io_ins_3(ces_160_0_io_ins_3),
    .io_outs_0(ces_160_0_io_outs_0),
    .io_outs_1(ces_160_0_io_outs_1),
    .io_outs_2(ces_160_0_io_outs_2),
    .io_outs_3(ces_160_0_io_outs_3)
  );
  Element ces_161_0 ( // @[MockArray.scala 36:52]
    .clock(ces_161_0_clock),
    .io_ins_0(ces_161_0_io_ins_0),
    .io_ins_1(ces_161_0_io_ins_1),
    .io_ins_2(ces_161_0_io_ins_2),
    .io_ins_3(ces_161_0_io_ins_3),
    .io_outs_0(ces_161_0_io_outs_0),
    .io_outs_1(ces_161_0_io_outs_1),
    .io_outs_2(ces_161_0_io_outs_2),
    .io_outs_3(ces_161_0_io_outs_3)
  );
  Element ces_162_0 ( // @[MockArray.scala 36:52]
    .clock(ces_162_0_clock),
    .io_ins_0(ces_162_0_io_ins_0),
    .io_ins_1(ces_162_0_io_ins_1),
    .io_ins_2(ces_162_0_io_ins_2),
    .io_ins_3(ces_162_0_io_ins_3),
    .io_outs_0(ces_162_0_io_outs_0),
    .io_outs_1(ces_162_0_io_outs_1),
    .io_outs_2(ces_162_0_io_outs_2),
    .io_outs_3(ces_162_0_io_outs_3)
  );
  Element ces_163_0 ( // @[MockArray.scala 36:52]
    .clock(ces_163_0_clock),
    .io_ins_0(ces_163_0_io_ins_0),
    .io_ins_1(ces_163_0_io_ins_1),
    .io_ins_2(ces_163_0_io_ins_2),
    .io_ins_3(ces_163_0_io_ins_3),
    .io_outs_0(ces_163_0_io_outs_0),
    .io_outs_1(ces_163_0_io_outs_1),
    .io_outs_2(ces_163_0_io_outs_2),
    .io_outs_3(ces_163_0_io_outs_3)
  );
  Element ces_164_0 ( // @[MockArray.scala 36:52]
    .clock(ces_164_0_clock),
    .io_ins_0(ces_164_0_io_ins_0),
    .io_ins_1(ces_164_0_io_ins_1),
    .io_ins_2(ces_164_0_io_ins_2),
    .io_ins_3(ces_164_0_io_ins_3),
    .io_outs_0(ces_164_0_io_outs_0),
    .io_outs_1(ces_164_0_io_outs_1),
    .io_outs_2(ces_164_0_io_outs_2),
    .io_outs_3(ces_164_0_io_outs_3)
  );
  Element ces_165_0 ( // @[MockArray.scala 36:52]
    .clock(ces_165_0_clock),
    .io_ins_0(ces_165_0_io_ins_0),
    .io_ins_1(ces_165_0_io_ins_1),
    .io_ins_2(ces_165_0_io_ins_2),
    .io_ins_3(ces_165_0_io_ins_3),
    .io_outs_0(ces_165_0_io_outs_0),
    .io_outs_1(ces_165_0_io_outs_1),
    .io_outs_2(ces_165_0_io_outs_2),
    .io_outs_3(ces_165_0_io_outs_3)
  );
  Element ces_166_0 ( // @[MockArray.scala 36:52]
    .clock(ces_166_0_clock),
    .io_ins_0(ces_166_0_io_ins_0),
    .io_ins_1(ces_166_0_io_ins_1),
    .io_ins_2(ces_166_0_io_ins_2),
    .io_ins_3(ces_166_0_io_ins_3),
    .io_outs_0(ces_166_0_io_outs_0),
    .io_outs_1(ces_166_0_io_outs_1),
    .io_outs_2(ces_166_0_io_outs_2),
    .io_outs_3(ces_166_0_io_outs_3)
  );
  Element ces_167_0 ( // @[MockArray.scala 36:52]
    .clock(ces_167_0_clock),
    .io_ins_0(ces_167_0_io_ins_0),
    .io_ins_1(ces_167_0_io_ins_1),
    .io_ins_2(ces_167_0_io_ins_2),
    .io_ins_3(ces_167_0_io_ins_3),
    .io_outs_0(ces_167_0_io_outs_0),
    .io_outs_1(ces_167_0_io_outs_1),
    .io_outs_2(ces_167_0_io_outs_2),
    .io_outs_3(ces_167_0_io_outs_3)
  );
  Element ces_168_0 ( // @[MockArray.scala 36:52]
    .clock(ces_168_0_clock),
    .io_ins_0(ces_168_0_io_ins_0),
    .io_ins_1(ces_168_0_io_ins_1),
    .io_ins_2(ces_168_0_io_ins_2),
    .io_ins_3(ces_168_0_io_ins_3),
    .io_outs_0(ces_168_0_io_outs_0),
    .io_outs_1(ces_168_0_io_outs_1),
    .io_outs_2(ces_168_0_io_outs_2),
    .io_outs_3(ces_168_0_io_outs_3)
  );
  Element ces_169_0 ( // @[MockArray.scala 36:52]
    .clock(ces_169_0_clock),
    .io_ins_0(ces_169_0_io_ins_0),
    .io_ins_1(ces_169_0_io_ins_1),
    .io_ins_2(ces_169_0_io_ins_2),
    .io_ins_3(ces_169_0_io_ins_3),
    .io_outs_0(ces_169_0_io_outs_0),
    .io_outs_1(ces_169_0_io_outs_1),
    .io_outs_2(ces_169_0_io_outs_2),
    .io_outs_3(ces_169_0_io_outs_3)
  );
  Element ces_170_0 ( // @[MockArray.scala 36:52]
    .clock(ces_170_0_clock),
    .io_ins_0(ces_170_0_io_ins_0),
    .io_ins_1(ces_170_0_io_ins_1),
    .io_ins_2(ces_170_0_io_ins_2),
    .io_ins_3(ces_170_0_io_ins_3),
    .io_outs_0(ces_170_0_io_outs_0),
    .io_outs_1(ces_170_0_io_outs_1),
    .io_outs_2(ces_170_0_io_outs_2),
    .io_outs_3(ces_170_0_io_outs_3)
  );
  Element ces_171_0 ( // @[MockArray.scala 36:52]
    .clock(ces_171_0_clock),
    .io_ins_0(ces_171_0_io_ins_0),
    .io_ins_1(ces_171_0_io_ins_1),
    .io_ins_2(ces_171_0_io_ins_2),
    .io_ins_3(ces_171_0_io_ins_3),
    .io_outs_0(ces_171_0_io_outs_0),
    .io_outs_1(ces_171_0_io_outs_1),
    .io_outs_2(ces_171_0_io_outs_2),
    .io_outs_3(ces_171_0_io_outs_3)
  );
  Element ces_172_0 ( // @[MockArray.scala 36:52]
    .clock(ces_172_0_clock),
    .io_ins_0(ces_172_0_io_ins_0),
    .io_ins_1(ces_172_0_io_ins_1),
    .io_ins_2(ces_172_0_io_ins_2),
    .io_ins_3(ces_172_0_io_ins_3),
    .io_outs_0(ces_172_0_io_outs_0),
    .io_outs_1(ces_172_0_io_outs_1),
    .io_outs_2(ces_172_0_io_outs_2),
    .io_outs_3(ces_172_0_io_outs_3)
  );
  Element ces_173_0 ( // @[MockArray.scala 36:52]
    .clock(ces_173_0_clock),
    .io_ins_0(ces_173_0_io_ins_0),
    .io_ins_1(ces_173_0_io_ins_1),
    .io_ins_2(ces_173_0_io_ins_2),
    .io_ins_3(ces_173_0_io_ins_3),
    .io_outs_0(ces_173_0_io_outs_0),
    .io_outs_1(ces_173_0_io_outs_1),
    .io_outs_2(ces_173_0_io_outs_2),
    .io_outs_3(ces_173_0_io_outs_3)
  );
  Element ces_174_0 ( // @[MockArray.scala 36:52]
    .clock(ces_174_0_clock),
    .io_ins_0(ces_174_0_io_ins_0),
    .io_ins_1(ces_174_0_io_ins_1),
    .io_ins_2(ces_174_0_io_ins_2),
    .io_ins_3(ces_174_0_io_ins_3),
    .io_outs_0(ces_174_0_io_outs_0),
    .io_outs_1(ces_174_0_io_outs_1),
    .io_outs_2(ces_174_0_io_outs_2),
    .io_outs_3(ces_174_0_io_outs_3)
  );
  Element ces_175_0 ( // @[MockArray.scala 36:52]
    .clock(ces_175_0_clock),
    .io_ins_0(ces_175_0_io_ins_0),
    .io_ins_1(ces_175_0_io_ins_1),
    .io_ins_2(ces_175_0_io_ins_2),
    .io_ins_3(ces_175_0_io_ins_3),
    .io_outs_0(ces_175_0_io_outs_0),
    .io_outs_1(ces_175_0_io_outs_1),
    .io_outs_2(ces_175_0_io_outs_2),
    .io_outs_3(ces_175_0_io_outs_3)
  );
  Element ces_176_0 ( // @[MockArray.scala 36:52]
    .clock(ces_176_0_clock),
    .io_ins_0(ces_176_0_io_ins_0),
    .io_ins_1(ces_176_0_io_ins_1),
    .io_ins_2(ces_176_0_io_ins_2),
    .io_ins_3(ces_176_0_io_ins_3),
    .io_outs_0(ces_176_0_io_outs_0),
    .io_outs_1(ces_176_0_io_outs_1),
    .io_outs_2(ces_176_0_io_outs_2),
    .io_outs_3(ces_176_0_io_outs_3)
  );
  Element ces_177_0 ( // @[MockArray.scala 36:52]
    .clock(ces_177_0_clock),
    .io_ins_0(ces_177_0_io_ins_0),
    .io_ins_1(ces_177_0_io_ins_1),
    .io_ins_2(ces_177_0_io_ins_2),
    .io_ins_3(ces_177_0_io_ins_3),
    .io_outs_0(ces_177_0_io_outs_0),
    .io_outs_1(ces_177_0_io_outs_1),
    .io_outs_2(ces_177_0_io_outs_2),
    .io_outs_3(ces_177_0_io_outs_3)
  );
  Element ces_178_0 ( // @[MockArray.scala 36:52]
    .clock(ces_178_0_clock),
    .io_ins_0(ces_178_0_io_ins_0),
    .io_ins_1(ces_178_0_io_ins_1),
    .io_ins_2(ces_178_0_io_ins_2),
    .io_ins_3(ces_178_0_io_ins_3),
    .io_outs_0(ces_178_0_io_outs_0),
    .io_outs_1(ces_178_0_io_outs_1),
    .io_outs_2(ces_178_0_io_outs_2),
    .io_outs_3(ces_178_0_io_outs_3)
  );
  Element ces_179_0 ( // @[MockArray.scala 36:52]
    .clock(ces_179_0_clock),
    .io_ins_0(ces_179_0_io_ins_0),
    .io_ins_1(ces_179_0_io_ins_1),
    .io_ins_2(ces_179_0_io_ins_2),
    .io_ins_3(ces_179_0_io_ins_3),
    .io_outs_0(ces_179_0_io_outs_0),
    .io_outs_1(ces_179_0_io_outs_1),
    .io_outs_2(ces_179_0_io_outs_2),
    .io_outs_3(ces_179_0_io_outs_3)
  );
  Element ces_180_0 ( // @[MockArray.scala 36:52]
    .clock(ces_180_0_clock),
    .io_ins_0(ces_180_0_io_ins_0),
    .io_ins_1(ces_180_0_io_ins_1),
    .io_ins_2(ces_180_0_io_ins_2),
    .io_ins_3(ces_180_0_io_ins_3),
    .io_outs_0(ces_180_0_io_outs_0),
    .io_outs_1(ces_180_0_io_outs_1),
    .io_outs_2(ces_180_0_io_outs_2),
    .io_outs_3(ces_180_0_io_outs_3)
  );
  Element ces_181_0 ( // @[MockArray.scala 36:52]
    .clock(ces_181_0_clock),
    .io_ins_0(ces_181_0_io_ins_0),
    .io_ins_1(ces_181_0_io_ins_1),
    .io_ins_2(ces_181_0_io_ins_2),
    .io_ins_3(ces_181_0_io_ins_3),
    .io_outs_0(ces_181_0_io_outs_0),
    .io_outs_1(ces_181_0_io_outs_1),
    .io_outs_2(ces_181_0_io_outs_2),
    .io_outs_3(ces_181_0_io_outs_3)
  );
  Element ces_182_0 ( // @[MockArray.scala 36:52]
    .clock(ces_182_0_clock),
    .io_ins_0(ces_182_0_io_ins_0),
    .io_ins_1(ces_182_0_io_ins_1),
    .io_ins_2(ces_182_0_io_ins_2),
    .io_ins_3(ces_182_0_io_ins_3),
    .io_outs_0(ces_182_0_io_outs_0),
    .io_outs_1(ces_182_0_io_outs_1),
    .io_outs_2(ces_182_0_io_outs_2),
    .io_outs_3(ces_182_0_io_outs_3)
  );
  Element ces_183_0 ( // @[MockArray.scala 36:52]
    .clock(ces_183_0_clock),
    .io_ins_0(ces_183_0_io_ins_0),
    .io_ins_1(ces_183_0_io_ins_1),
    .io_ins_2(ces_183_0_io_ins_2),
    .io_ins_3(ces_183_0_io_ins_3),
    .io_outs_0(ces_183_0_io_outs_0),
    .io_outs_1(ces_183_0_io_outs_1),
    .io_outs_2(ces_183_0_io_outs_2),
    .io_outs_3(ces_183_0_io_outs_3)
  );
  Element ces_184_0 ( // @[MockArray.scala 36:52]
    .clock(ces_184_0_clock),
    .io_ins_0(ces_184_0_io_ins_0),
    .io_ins_1(ces_184_0_io_ins_1),
    .io_ins_2(ces_184_0_io_ins_2),
    .io_ins_3(ces_184_0_io_ins_3),
    .io_outs_0(ces_184_0_io_outs_0),
    .io_outs_1(ces_184_0_io_outs_1),
    .io_outs_2(ces_184_0_io_outs_2),
    .io_outs_3(ces_184_0_io_outs_3)
  );
  Element ces_185_0 ( // @[MockArray.scala 36:52]
    .clock(ces_185_0_clock),
    .io_ins_0(ces_185_0_io_ins_0),
    .io_ins_1(ces_185_0_io_ins_1),
    .io_ins_2(ces_185_0_io_ins_2),
    .io_ins_3(ces_185_0_io_ins_3),
    .io_outs_0(ces_185_0_io_outs_0),
    .io_outs_1(ces_185_0_io_outs_1),
    .io_outs_2(ces_185_0_io_outs_2),
    .io_outs_3(ces_185_0_io_outs_3)
  );
  Element ces_186_0 ( // @[MockArray.scala 36:52]
    .clock(ces_186_0_clock),
    .io_ins_0(ces_186_0_io_ins_0),
    .io_ins_1(ces_186_0_io_ins_1),
    .io_ins_2(ces_186_0_io_ins_2),
    .io_ins_3(ces_186_0_io_ins_3),
    .io_outs_0(ces_186_0_io_outs_0),
    .io_outs_1(ces_186_0_io_outs_1),
    .io_outs_2(ces_186_0_io_outs_2),
    .io_outs_3(ces_186_0_io_outs_3)
  );
  Element ces_187_0 ( // @[MockArray.scala 36:52]
    .clock(ces_187_0_clock),
    .io_ins_0(ces_187_0_io_ins_0),
    .io_ins_1(ces_187_0_io_ins_1),
    .io_ins_2(ces_187_0_io_ins_2),
    .io_ins_3(ces_187_0_io_ins_3),
    .io_outs_0(ces_187_0_io_outs_0),
    .io_outs_1(ces_187_0_io_outs_1),
    .io_outs_2(ces_187_0_io_outs_2),
    .io_outs_3(ces_187_0_io_outs_3)
  );
  Element ces_188_0 ( // @[MockArray.scala 36:52]
    .clock(ces_188_0_clock),
    .io_ins_0(ces_188_0_io_ins_0),
    .io_ins_1(ces_188_0_io_ins_1),
    .io_ins_2(ces_188_0_io_ins_2),
    .io_ins_3(ces_188_0_io_ins_3),
    .io_outs_0(ces_188_0_io_outs_0),
    .io_outs_1(ces_188_0_io_outs_1),
    .io_outs_2(ces_188_0_io_outs_2),
    .io_outs_3(ces_188_0_io_outs_3)
  );
  Element ces_189_0 ( // @[MockArray.scala 36:52]
    .clock(ces_189_0_clock),
    .io_ins_0(ces_189_0_io_ins_0),
    .io_ins_1(ces_189_0_io_ins_1),
    .io_ins_2(ces_189_0_io_ins_2),
    .io_ins_3(ces_189_0_io_ins_3),
    .io_outs_0(ces_189_0_io_outs_0),
    .io_outs_1(ces_189_0_io_outs_1),
    .io_outs_2(ces_189_0_io_outs_2),
    .io_outs_3(ces_189_0_io_outs_3)
  );
  Element ces_190_0 ( // @[MockArray.scala 36:52]
    .clock(ces_190_0_clock),
    .io_ins_0(ces_190_0_io_ins_0),
    .io_ins_1(ces_190_0_io_ins_1),
    .io_ins_2(ces_190_0_io_ins_2),
    .io_ins_3(ces_190_0_io_ins_3),
    .io_outs_0(ces_190_0_io_outs_0),
    .io_outs_1(ces_190_0_io_outs_1),
    .io_outs_2(ces_190_0_io_outs_2),
    .io_outs_3(ces_190_0_io_outs_3)
  );
  Element ces_191_0 ( // @[MockArray.scala 36:52]
    .clock(ces_191_0_clock),
    .io_ins_0(ces_191_0_io_ins_0),
    .io_ins_1(ces_191_0_io_ins_1),
    .io_ins_2(ces_191_0_io_ins_2),
    .io_ins_3(ces_191_0_io_ins_3),
    .io_outs_0(ces_191_0_io_outs_0),
    .io_outs_1(ces_191_0_io_outs_1),
    .io_outs_2(ces_191_0_io_outs_2),
    .io_outs_3(ces_191_0_io_outs_3)
  );
  Element ces_192_0 ( // @[MockArray.scala 36:52]
    .clock(ces_192_0_clock),
    .io_ins_0(ces_192_0_io_ins_0),
    .io_ins_1(ces_192_0_io_ins_1),
    .io_ins_2(ces_192_0_io_ins_2),
    .io_ins_3(ces_192_0_io_ins_3),
    .io_outs_0(ces_192_0_io_outs_0),
    .io_outs_1(ces_192_0_io_outs_1),
    .io_outs_2(ces_192_0_io_outs_2),
    .io_outs_3(ces_192_0_io_outs_3)
  );
  Element ces_193_0 ( // @[MockArray.scala 36:52]
    .clock(ces_193_0_clock),
    .io_ins_0(ces_193_0_io_ins_0),
    .io_ins_1(ces_193_0_io_ins_1),
    .io_ins_2(ces_193_0_io_ins_2),
    .io_ins_3(ces_193_0_io_ins_3),
    .io_outs_0(ces_193_0_io_outs_0),
    .io_outs_1(ces_193_0_io_outs_1),
    .io_outs_2(ces_193_0_io_outs_2),
    .io_outs_3(ces_193_0_io_outs_3)
  );
  Element ces_194_0 ( // @[MockArray.scala 36:52]
    .clock(ces_194_0_clock),
    .io_ins_0(ces_194_0_io_ins_0),
    .io_ins_1(ces_194_0_io_ins_1),
    .io_ins_2(ces_194_0_io_ins_2),
    .io_ins_3(ces_194_0_io_ins_3),
    .io_outs_0(ces_194_0_io_outs_0),
    .io_outs_1(ces_194_0_io_outs_1),
    .io_outs_2(ces_194_0_io_outs_2),
    .io_outs_3(ces_194_0_io_outs_3)
  );
  Element ces_195_0 ( // @[MockArray.scala 36:52]
    .clock(ces_195_0_clock),
    .io_ins_0(ces_195_0_io_ins_0),
    .io_ins_1(ces_195_0_io_ins_1),
    .io_ins_2(ces_195_0_io_ins_2),
    .io_ins_3(ces_195_0_io_ins_3),
    .io_outs_0(ces_195_0_io_outs_0),
    .io_outs_1(ces_195_0_io_outs_1),
    .io_outs_2(ces_195_0_io_outs_2),
    .io_outs_3(ces_195_0_io_outs_3)
  );
  Element ces_196_0 ( // @[MockArray.scala 36:52]
    .clock(ces_196_0_clock),
    .io_ins_0(ces_196_0_io_ins_0),
    .io_ins_1(ces_196_0_io_ins_1),
    .io_ins_2(ces_196_0_io_ins_2),
    .io_ins_3(ces_196_0_io_ins_3),
    .io_outs_0(ces_196_0_io_outs_0),
    .io_outs_1(ces_196_0_io_outs_1),
    .io_outs_2(ces_196_0_io_outs_2),
    .io_outs_3(ces_196_0_io_outs_3)
  );
  Element ces_197_0 ( // @[MockArray.scala 36:52]
    .clock(ces_197_0_clock),
    .io_ins_0(ces_197_0_io_ins_0),
    .io_ins_1(ces_197_0_io_ins_1),
    .io_ins_2(ces_197_0_io_ins_2),
    .io_ins_3(ces_197_0_io_ins_3),
    .io_outs_0(ces_197_0_io_outs_0),
    .io_outs_1(ces_197_0_io_outs_1),
    .io_outs_2(ces_197_0_io_outs_2),
    .io_outs_3(ces_197_0_io_outs_3)
  );
  Element ces_198_0 ( // @[MockArray.scala 36:52]
    .clock(ces_198_0_clock),
    .io_ins_0(ces_198_0_io_ins_0),
    .io_ins_1(ces_198_0_io_ins_1),
    .io_ins_2(ces_198_0_io_ins_2),
    .io_ins_3(ces_198_0_io_ins_3),
    .io_outs_0(ces_198_0_io_outs_0),
    .io_outs_1(ces_198_0_io_outs_1),
    .io_outs_2(ces_198_0_io_outs_2),
    .io_outs_3(ces_198_0_io_outs_3)
  );
  Element ces_199_0 ( // @[MockArray.scala 36:52]
    .clock(ces_199_0_clock),
    .io_ins_0(ces_199_0_io_ins_0),
    .io_ins_1(ces_199_0_io_ins_1),
    .io_ins_2(ces_199_0_io_ins_2),
    .io_ins_3(ces_199_0_io_ins_3),
    .io_outs_0(ces_199_0_io_outs_0),
    .io_outs_1(ces_199_0_io_outs_1),
    .io_outs_2(ces_199_0_io_outs_2),
    .io_outs_3(ces_199_0_io_outs_3)
  );
  Element ces_200_0 ( // @[MockArray.scala 36:52]
    .clock(ces_200_0_clock),
    .io_ins_0(ces_200_0_io_ins_0),
    .io_ins_1(ces_200_0_io_ins_1),
    .io_ins_2(ces_200_0_io_ins_2),
    .io_ins_3(ces_200_0_io_ins_3),
    .io_outs_0(ces_200_0_io_outs_0),
    .io_outs_1(ces_200_0_io_outs_1),
    .io_outs_2(ces_200_0_io_outs_2),
    .io_outs_3(ces_200_0_io_outs_3)
  );
  Element ces_201_0 ( // @[MockArray.scala 36:52]
    .clock(ces_201_0_clock),
    .io_ins_0(ces_201_0_io_ins_0),
    .io_ins_1(ces_201_0_io_ins_1),
    .io_ins_2(ces_201_0_io_ins_2),
    .io_ins_3(ces_201_0_io_ins_3),
    .io_outs_0(ces_201_0_io_outs_0),
    .io_outs_1(ces_201_0_io_outs_1),
    .io_outs_2(ces_201_0_io_outs_2),
    .io_outs_3(ces_201_0_io_outs_3)
  );
  Element ces_202_0 ( // @[MockArray.scala 36:52]
    .clock(ces_202_0_clock),
    .io_ins_0(ces_202_0_io_ins_0),
    .io_ins_1(ces_202_0_io_ins_1),
    .io_ins_2(ces_202_0_io_ins_2),
    .io_ins_3(ces_202_0_io_ins_3),
    .io_outs_0(ces_202_0_io_outs_0),
    .io_outs_1(ces_202_0_io_outs_1),
    .io_outs_2(ces_202_0_io_outs_2),
    .io_outs_3(ces_202_0_io_outs_3)
  );
  Element ces_203_0 ( // @[MockArray.scala 36:52]
    .clock(ces_203_0_clock),
    .io_ins_0(ces_203_0_io_ins_0),
    .io_ins_1(ces_203_0_io_ins_1),
    .io_ins_2(ces_203_0_io_ins_2),
    .io_ins_3(ces_203_0_io_ins_3),
    .io_outs_0(ces_203_0_io_outs_0),
    .io_outs_1(ces_203_0_io_outs_1),
    .io_outs_2(ces_203_0_io_outs_2),
    .io_outs_3(ces_203_0_io_outs_3)
  );
  Element ces_204_0 ( // @[MockArray.scala 36:52]
    .clock(ces_204_0_clock),
    .io_ins_0(ces_204_0_io_ins_0),
    .io_ins_1(ces_204_0_io_ins_1),
    .io_ins_2(ces_204_0_io_ins_2),
    .io_ins_3(ces_204_0_io_ins_3),
    .io_outs_0(ces_204_0_io_outs_0),
    .io_outs_1(ces_204_0_io_outs_1),
    .io_outs_2(ces_204_0_io_outs_2),
    .io_outs_3(ces_204_0_io_outs_3)
  );
  Element ces_205_0 ( // @[MockArray.scala 36:52]
    .clock(ces_205_0_clock),
    .io_ins_0(ces_205_0_io_ins_0),
    .io_ins_1(ces_205_0_io_ins_1),
    .io_ins_2(ces_205_0_io_ins_2),
    .io_ins_3(ces_205_0_io_ins_3),
    .io_outs_0(ces_205_0_io_outs_0),
    .io_outs_1(ces_205_0_io_outs_1),
    .io_outs_2(ces_205_0_io_outs_2),
    .io_outs_3(ces_205_0_io_outs_3)
  );
  Element ces_206_0 ( // @[MockArray.scala 36:52]
    .clock(ces_206_0_clock),
    .io_ins_0(ces_206_0_io_ins_0),
    .io_ins_1(ces_206_0_io_ins_1),
    .io_ins_2(ces_206_0_io_ins_2),
    .io_ins_3(ces_206_0_io_ins_3),
    .io_outs_0(ces_206_0_io_outs_0),
    .io_outs_1(ces_206_0_io_outs_1),
    .io_outs_2(ces_206_0_io_outs_2),
    .io_outs_3(ces_206_0_io_outs_3)
  );
  Element ces_207_0 ( // @[MockArray.scala 36:52]
    .clock(ces_207_0_clock),
    .io_ins_0(ces_207_0_io_ins_0),
    .io_ins_1(ces_207_0_io_ins_1),
    .io_ins_2(ces_207_0_io_ins_2),
    .io_ins_3(ces_207_0_io_ins_3),
    .io_outs_0(ces_207_0_io_outs_0),
    .io_outs_1(ces_207_0_io_outs_1),
    .io_outs_2(ces_207_0_io_outs_2),
    .io_outs_3(ces_207_0_io_outs_3)
  );
  Element ces_208_0 ( // @[MockArray.scala 36:52]
    .clock(ces_208_0_clock),
    .io_ins_0(ces_208_0_io_ins_0),
    .io_ins_1(ces_208_0_io_ins_1),
    .io_ins_2(ces_208_0_io_ins_2),
    .io_ins_3(ces_208_0_io_ins_3),
    .io_outs_0(ces_208_0_io_outs_0),
    .io_outs_1(ces_208_0_io_outs_1),
    .io_outs_2(ces_208_0_io_outs_2),
    .io_outs_3(ces_208_0_io_outs_3)
  );
  Element ces_209_0 ( // @[MockArray.scala 36:52]
    .clock(ces_209_0_clock),
    .io_ins_0(ces_209_0_io_ins_0),
    .io_ins_1(ces_209_0_io_ins_1),
    .io_ins_2(ces_209_0_io_ins_2),
    .io_ins_3(ces_209_0_io_ins_3),
    .io_outs_0(ces_209_0_io_outs_0),
    .io_outs_1(ces_209_0_io_outs_1),
    .io_outs_2(ces_209_0_io_outs_2),
    .io_outs_3(ces_209_0_io_outs_3)
  );
  Element ces_210_0 ( // @[MockArray.scala 36:52]
    .clock(ces_210_0_clock),
    .io_ins_0(ces_210_0_io_ins_0),
    .io_ins_1(ces_210_0_io_ins_1),
    .io_ins_2(ces_210_0_io_ins_2),
    .io_ins_3(ces_210_0_io_ins_3),
    .io_outs_0(ces_210_0_io_outs_0),
    .io_outs_1(ces_210_0_io_outs_1),
    .io_outs_2(ces_210_0_io_outs_2),
    .io_outs_3(ces_210_0_io_outs_3)
  );
  Element ces_211_0 ( // @[MockArray.scala 36:52]
    .clock(ces_211_0_clock),
    .io_ins_0(ces_211_0_io_ins_0),
    .io_ins_1(ces_211_0_io_ins_1),
    .io_ins_2(ces_211_0_io_ins_2),
    .io_ins_3(ces_211_0_io_ins_3),
    .io_outs_0(ces_211_0_io_outs_0),
    .io_outs_1(ces_211_0_io_outs_1),
    .io_outs_2(ces_211_0_io_outs_2),
    .io_outs_3(ces_211_0_io_outs_3)
  );
  Element ces_212_0 ( // @[MockArray.scala 36:52]
    .clock(ces_212_0_clock),
    .io_ins_0(ces_212_0_io_ins_0),
    .io_ins_1(ces_212_0_io_ins_1),
    .io_ins_2(ces_212_0_io_ins_2),
    .io_ins_3(ces_212_0_io_ins_3),
    .io_outs_0(ces_212_0_io_outs_0),
    .io_outs_1(ces_212_0_io_outs_1),
    .io_outs_2(ces_212_0_io_outs_2),
    .io_outs_3(ces_212_0_io_outs_3)
  );
  Element ces_213_0 ( // @[MockArray.scala 36:52]
    .clock(ces_213_0_clock),
    .io_ins_0(ces_213_0_io_ins_0),
    .io_ins_1(ces_213_0_io_ins_1),
    .io_ins_2(ces_213_0_io_ins_2),
    .io_ins_3(ces_213_0_io_ins_3),
    .io_outs_0(ces_213_0_io_outs_0),
    .io_outs_1(ces_213_0_io_outs_1),
    .io_outs_2(ces_213_0_io_outs_2),
    .io_outs_3(ces_213_0_io_outs_3)
  );
  Element ces_214_0 ( // @[MockArray.scala 36:52]
    .clock(ces_214_0_clock),
    .io_ins_0(ces_214_0_io_ins_0),
    .io_ins_1(ces_214_0_io_ins_1),
    .io_ins_2(ces_214_0_io_ins_2),
    .io_ins_3(ces_214_0_io_ins_3),
    .io_outs_0(ces_214_0_io_outs_0),
    .io_outs_1(ces_214_0_io_outs_1),
    .io_outs_2(ces_214_0_io_outs_2),
    .io_outs_3(ces_214_0_io_outs_3)
  );
  Element ces_215_0 ( // @[MockArray.scala 36:52]
    .clock(ces_215_0_clock),
    .io_ins_0(ces_215_0_io_ins_0),
    .io_ins_1(ces_215_0_io_ins_1),
    .io_ins_2(ces_215_0_io_ins_2),
    .io_ins_3(ces_215_0_io_ins_3),
    .io_outs_0(ces_215_0_io_outs_0),
    .io_outs_1(ces_215_0_io_outs_1),
    .io_outs_2(ces_215_0_io_outs_2),
    .io_outs_3(ces_215_0_io_outs_3)
  );
  Element ces_216_0 ( // @[MockArray.scala 36:52]
    .clock(ces_216_0_clock),
    .io_ins_0(ces_216_0_io_ins_0),
    .io_ins_1(ces_216_0_io_ins_1),
    .io_ins_2(ces_216_0_io_ins_2),
    .io_ins_3(ces_216_0_io_ins_3),
    .io_outs_0(ces_216_0_io_outs_0),
    .io_outs_1(ces_216_0_io_outs_1),
    .io_outs_2(ces_216_0_io_outs_2),
    .io_outs_3(ces_216_0_io_outs_3)
  );
  Element ces_217_0 ( // @[MockArray.scala 36:52]
    .clock(ces_217_0_clock),
    .io_ins_0(ces_217_0_io_ins_0),
    .io_ins_1(ces_217_0_io_ins_1),
    .io_ins_2(ces_217_0_io_ins_2),
    .io_ins_3(ces_217_0_io_ins_3),
    .io_outs_0(ces_217_0_io_outs_0),
    .io_outs_1(ces_217_0_io_outs_1),
    .io_outs_2(ces_217_0_io_outs_2),
    .io_outs_3(ces_217_0_io_outs_3)
  );
  Element ces_218_0 ( // @[MockArray.scala 36:52]
    .clock(ces_218_0_clock),
    .io_ins_0(ces_218_0_io_ins_0),
    .io_ins_1(ces_218_0_io_ins_1),
    .io_ins_2(ces_218_0_io_ins_2),
    .io_ins_3(ces_218_0_io_ins_3),
    .io_outs_0(ces_218_0_io_outs_0),
    .io_outs_1(ces_218_0_io_outs_1),
    .io_outs_2(ces_218_0_io_outs_2),
    .io_outs_3(ces_218_0_io_outs_3)
  );
  Element ces_219_0 ( // @[MockArray.scala 36:52]
    .clock(ces_219_0_clock),
    .io_ins_0(ces_219_0_io_ins_0),
    .io_ins_1(ces_219_0_io_ins_1),
    .io_ins_2(ces_219_0_io_ins_2),
    .io_ins_3(ces_219_0_io_ins_3),
    .io_outs_0(ces_219_0_io_outs_0),
    .io_outs_1(ces_219_0_io_outs_1),
    .io_outs_2(ces_219_0_io_outs_2),
    .io_outs_3(ces_219_0_io_outs_3)
  );
  Element ces_220_0 ( // @[MockArray.scala 36:52]
    .clock(ces_220_0_clock),
    .io_ins_0(ces_220_0_io_ins_0),
    .io_ins_1(ces_220_0_io_ins_1),
    .io_ins_2(ces_220_0_io_ins_2),
    .io_ins_3(ces_220_0_io_ins_3),
    .io_outs_0(ces_220_0_io_outs_0),
    .io_outs_1(ces_220_0_io_outs_1),
    .io_outs_2(ces_220_0_io_outs_2),
    .io_outs_3(ces_220_0_io_outs_3)
  );
  Element ces_221_0 ( // @[MockArray.scala 36:52]
    .clock(ces_221_0_clock),
    .io_ins_0(ces_221_0_io_ins_0),
    .io_ins_1(ces_221_0_io_ins_1),
    .io_ins_2(ces_221_0_io_ins_2),
    .io_ins_3(ces_221_0_io_ins_3),
    .io_outs_0(ces_221_0_io_outs_0),
    .io_outs_1(ces_221_0_io_outs_1),
    .io_outs_2(ces_221_0_io_outs_2),
    .io_outs_3(ces_221_0_io_outs_3)
  );
  Element ces_222_0 ( // @[MockArray.scala 36:52]
    .clock(ces_222_0_clock),
    .io_ins_0(ces_222_0_io_ins_0),
    .io_ins_1(ces_222_0_io_ins_1),
    .io_ins_2(ces_222_0_io_ins_2),
    .io_ins_3(ces_222_0_io_ins_3),
    .io_outs_0(ces_222_0_io_outs_0),
    .io_outs_1(ces_222_0_io_outs_1),
    .io_outs_2(ces_222_0_io_outs_2),
    .io_outs_3(ces_222_0_io_outs_3)
  );
  Element ces_223_0 ( // @[MockArray.scala 36:52]
    .clock(ces_223_0_clock),
    .io_ins_0(ces_223_0_io_ins_0),
    .io_ins_1(ces_223_0_io_ins_1),
    .io_ins_2(ces_223_0_io_ins_2),
    .io_ins_3(ces_223_0_io_ins_3),
    .io_outs_0(ces_223_0_io_outs_0),
    .io_outs_1(ces_223_0_io_outs_1),
    .io_outs_2(ces_223_0_io_outs_2),
    .io_outs_3(ces_223_0_io_outs_3)
  );
  Element ces_224_0 ( // @[MockArray.scala 36:52]
    .clock(ces_224_0_clock),
    .io_ins_0(ces_224_0_io_ins_0),
    .io_ins_1(ces_224_0_io_ins_1),
    .io_ins_2(ces_224_0_io_ins_2),
    .io_ins_3(ces_224_0_io_ins_3),
    .io_outs_0(ces_224_0_io_outs_0),
    .io_outs_1(ces_224_0_io_outs_1),
    .io_outs_2(ces_224_0_io_outs_2),
    .io_outs_3(ces_224_0_io_outs_3)
  );
  Element ces_225_0 ( // @[MockArray.scala 36:52]
    .clock(ces_225_0_clock),
    .io_ins_0(ces_225_0_io_ins_0),
    .io_ins_1(ces_225_0_io_ins_1),
    .io_ins_2(ces_225_0_io_ins_2),
    .io_ins_3(ces_225_0_io_ins_3),
    .io_outs_0(ces_225_0_io_outs_0),
    .io_outs_1(ces_225_0_io_outs_1),
    .io_outs_2(ces_225_0_io_outs_2),
    .io_outs_3(ces_225_0_io_outs_3)
  );
  Element ces_226_0 ( // @[MockArray.scala 36:52]
    .clock(ces_226_0_clock),
    .io_ins_0(ces_226_0_io_ins_0),
    .io_ins_1(ces_226_0_io_ins_1),
    .io_ins_2(ces_226_0_io_ins_2),
    .io_ins_3(ces_226_0_io_ins_3),
    .io_outs_0(ces_226_0_io_outs_0),
    .io_outs_1(ces_226_0_io_outs_1),
    .io_outs_2(ces_226_0_io_outs_2),
    .io_outs_3(ces_226_0_io_outs_3)
  );
  Element ces_227_0 ( // @[MockArray.scala 36:52]
    .clock(ces_227_0_clock),
    .io_ins_0(ces_227_0_io_ins_0),
    .io_ins_1(ces_227_0_io_ins_1),
    .io_ins_2(ces_227_0_io_ins_2),
    .io_ins_3(ces_227_0_io_ins_3),
    .io_outs_0(ces_227_0_io_outs_0),
    .io_outs_1(ces_227_0_io_outs_1),
    .io_outs_2(ces_227_0_io_outs_2),
    .io_outs_3(ces_227_0_io_outs_3)
  );
  Element ces_228_0 ( // @[MockArray.scala 36:52]
    .clock(ces_228_0_clock),
    .io_ins_0(ces_228_0_io_ins_0),
    .io_ins_1(ces_228_0_io_ins_1),
    .io_ins_2(ces_228_0_io_ins_2),
    .io_ins_3(ces_228_0_io_ins_3),
    .io_outs_0(ces_228_0_io_outs_0),
    .io_outs_1(ces_228_0_io_outs_1),
    .io_outs_2(ces_228_0_io_outs_2),
    .io_outs_3(ces_228_0_io_outs_3)
  );
  Element ces_229_0 ( // @[MockArray.scala 36:52]
    .clock(ces_229_0_clock),
    .io_ins_0(ces_229_0_io_ins_0),
    .io_ins_1(ces_229_0_io_ins_1),
    .io_ins_2(ces_229_0_io_ins_2),
    .io_ins_3(ces_229_0_io_ins_3),
    .io_outs_0(ces_229_0_io_outs_0),
    .io_outs_1(ces_229_0_io_outs_1),
    .io_outs_2(ces_229_0_io_outs_2),
    .io_outs_3(ces_229_0_io_outs_3)
  );
  Element ces_230_0 ( // @[MockArray.scala 36:52]
    .clock(ces_230_0_clock),
    .io_ins_0(ces_230_0_io_ins_0),
    .io_ins_1(ces_230_0_io_ins_1),
    .io_ins_2(ces_230_0_io_ins_2),
    .io_ins_3(ces_230_0_io_ins_3),
    .io_outs_0(ces_230_0_io_outs_0),
    .io_outs_1(ces_230_0_io_outs_1),
    .io_outs_2(ces_230_0_io_outs_2),
    .io_outs_3(ces_230_0_io_outs_3)
  );
  Element ces_231_0 ( // @[MockArray.scala 36:52]
    .clock(ces_231_0_clock),
    .io_ins_0(ces_231_0_io_ins_0),
    .io_ins_1(ces_231_0_io_ins_1),
    .io_ins_2(ces_231_0_io_ins_2),
    .io_ins_3(ces_231_0_io_ins_3),
    .io_outs_0(ces_231_0_io_outs_0),
    .io_outs_1(ces_231_0_io_outs_1),
    .io_outs_2(ces_231_0_io_outs_2),
    .io_outs_3(ces_231_0_io_outs_3)
  );
  Element ces_232_0 ( // @[MockArray.scala 36:52]
    .clock(ces_232_0_clock),
    .io_ins_0(ces_232_0_io_ins_0),
    .io_ins_1(ces_232_0_io_ins_1),
    .io_ins_2(ces_232_0_io_ins_2),
    .io_ins_3(ces_232_0_io_ins_3),
    .io_outs_0(ces_232_0_io_outs_0),
    .io_outs_1(ces_232_0_io_outs_1),
    .io_outs_2(ces_232_0_io_outs_2),
    .io_outs_3(ces_232_0_io_outs_3)
  );
  Element ces_233_0 ( // @[MockArray.scala 36:52]
    .clock(ces_233_0_clock),
    .io_ins_0(ces_233_0_io_ins_0),
    .io_ins_1(ces_233_0_io_ins_1),
    .io_ins_2(ces_233_0_io_ins_2),
    .io_ins_3(ces_233_0_io_ins_3),
    .io_outs_0(ces_233_0_io_outs_0),
    .io_outs_1(ces_233_0_io_outs_1),
    .io_outs_2(ces_233_0_io_outs_2),
    .io_outs_3(ces_233_0_io_outs_3)
  );
  Element ces_234_0 ( // @[MockArray.scala 36:52]
    .clock(ces_234_0_clock),
    .io_ins_0(ces_234_0_io_ins_0),
    .io_ins_1(ces_234_0_io_ins_1),
    .io_ins_2(ces_234_0_io_ins_2),
    .io_ins_3(ces_234_0_io_ins_3),
    .io_outs_0(ces_234_0_io_outs_0),
    .io_outs_1(ces_234_0_io_outs_1),
    .io_outs_2(ces_234_0_io_outs_2),
    .io_outs_3(ces_234_0_io_outs_3)
  );
  Element ces_235_0 ( // @[MockArray.scala 36:52]
    .clock(ces_235_0_clock),
    .io_ins_0(ces_235_0_io_ins_0),
    .io_ins_1(ces_235_0_io_ins_1),
    .io_ins_2(ces_235_0_io_ins_2),
    .io_ins_3(ces_235_0_io_ins_3),
    .io_outs_0(ces_235_0_io_outs_0),
    .io_outs_1(ces_235_0_io_outs_1),
    .io_outs_2(ces_235_0_io_outs_2),
    .io_outs_3(ces_235_0_io_outs_3)
  );
  Element ces_236_0 ( // @[MockArray.scala 36:52]
    .clock(ces_236_0_clock),
    .io_ins_0(ces_236_0_io_ins_0),
    .io_ins_1(ces_236_0_io_ins_1),
    .io_ins_2(ces_236_0_io_ins_2),
    .io_ins_3(ces_236_0_io_ins_3),
    .io_outs_0(ces_236_0_io_outs_0),
    .io_outs_1(ces_236_0_io_outs_1),
    .io_outs_2(ces_236_0_io_outs_2),
    .io_outs_3(ces_236_0_io_outs_3)
  );
  Element ces_237_0 ( // @[MockArray.scala 36:52]
    .clock(ces_237_0_clock),
    .io_ins_0(ces_237_0_io_ins_0),
    .io_ins_1(ces_237_0_io_ins_1),
    .io_ins_2(ces_237_0_io_ins_2),
    .io_ins_3(ces_237_0_io_ins_3),
    .io_outs_0(ces_237_0_io_outs_0),
    .io_outs_1(ces_237_0_io_outs_1),
    .io_outs_2(ces_237_0_io_outs_2),
    .io_outs_3(ces_237_0_io_outs_3)
  );
  Element ces_238_0 ( // @[MockArray.scala 36:52]
    .clock(ces_238_0_clock),
    .io_ins_0(ces_238_0_io_ins_0),
    .io_ins_1(ces_238_0_io_ins_1),
    .io_ins_2(ces_238_0_io_ins_2),
    .io_ins_3(ces_238_0_io_ins_3),
    .io_outs_0(ces_238_0_io_outs_0),
    .io_outs_1(ces_238_0_io_outs_1),
    .io_outs_2(ces_238_0_io_outs_2),
    .io_outs_3(ces_238_0_io_outs_3)
  );
  Element ces_239_0 ( // @[MockArray.scala 36:52]
    .clock(ces_239_0_clock),
    .io_ins_0(ces_239_0_io_ins_0),
    .io_ins_1(ces_239_0_io_ins_1),
    .io_ins_2(ces_239_0_io_ins_2),
    .io_ins_3(ces_239_0_io_ins_3),
    .io_outs_0(ces_239_0_io_outs_0),
    .io_outs_1(ces_239_0_io_outs_1),
    .io_outs_2(ces_239_0_io_outs_2),
    .io_outs_3(ces_239_0_io_outs_3)
  );
  Element ces_240_0 ( // @[MockArray.scala 36:52]
    .clock(ces_240_0_clock),
    .io_ins_0(ces_240_0_io_ins_0),
    .io_ins_1(ces_240_0_io_ins_1),
    .io_ins_2(ces_240_0_io_ins_2),
    .io_ins_3(ces_240_0_io_ins_3),
    .io_outs_0(ces_240_0_io_outs_0),
    .io_outs_1(ces_240_0_io_outs_1),
    .io_outs_2(ces_240_0_io_outs_2),
    .io_outs_3(ces_240_0_io_outs_3)
  );
  Element ces_241_0 ( // @[MockArray.scala 36:52]
    .clock(ces_241_0_clock),
    .io_ins_0(ces_241_0_io_ins_0),
    .io_ins_1(ces_241_0_io_ins_1),
    .io_ins_2(ces_241_0_io_ins_2),
    .io_ins_3(ces_241_0_io_ins_3),
    .io_outs_0(ces_241_0_io_outs_0),
    .io_outs_1(ces_241_0_io_outs_1),
    .io_outs_2(ces_241_0_io_outs_2),
    .io_outs_3(ces_241_0_io_outs_3)
  );
  Element ces_242_0 ( // @[MockArray.scala 36:52]
    .clock(ces_242_0_clock),
    .io_ins_0(ces_242_0_io_ins_0),
    .io_ins_1(ces_242_0_io_ins_1),
    .io_ins_2(ces_242_0_io_ins_2),
    .io_ins_3(ces_242_0_io_ins_3),
    .io_outs_0(ces_242_0_io_outs_0),
    .io_outs_1(ces_242_0_io_outs_1),
    .io_outs_2(ces_242_0_io_outs_2),
    .io_outs_3(ces_242_0_io_outs_3)
  );
  Element ces_243_0 ( // @[MockArray.scala 36:52]
    .clock(ces_243_0_clock),
    .io_ins_0(ces_243_0_io_ins_0),
    .io_ins_1(ces_243_0_io_ins_1),
    .io_ins_2(ces_243_0_io_ins_2),
    .io_ins_3(ces_243_0_io_ins_3),
    .io_outs_0(ces_243_0_io_outs_0),
    .io_outs_1(ces_243_0_io_outs_1),
    .io_outs_2(ces_243_0_io_outs_2),
    .io_outs_3(ces_243_0_io_outs_3)
  );
  Element ces_244_0 ( // @[MockArray.scala 36:52]
    .clock(ces_244_0_clock),
    .io_ins_0(ces_244_0_io_ins_0),
    .io_ins_1(ces_244_0_io_ins_1),
    .io_ins_2(ces_244_0_io_ins_2),
    .io_ins_3(ces_244_0_io_ins_3),
    .io_outs_0(ces_244_0_io_outs_0),
    .io_outs_1(ces_244_0_io_outs_1),
    .io_outs_2(ces_244_0_io_outs_2),
    .io_outs_3(ces_244_0_io_outs_3)
  );
  Element ces_245_0 ( // @[MockArray.scala 36:52]
    .clock(ces_245_0_clock),
    .io_ins_0(ces_245_0_io_ins_0),
    .io_ins_1(ces_245_0_io_ins_1),
    .io_ins_2(ces_245_0_io_ins_2),
    .io_ins_3(ces_245_0_io_ins_3),
    .io_outs_0(ces_245_0_io_outs_0),
    .io_outs_1(ces_245_0_io_outs_1),
    .io_outs_2(ces_245_0_io_outs_2),
    .io_outs_3(ces_245_0_io_outs_3)
  );
  Element ces_246_0 ( // @[MockArray.scala 36:52]
    .clock(ces_246_0_clock),
    .io_ins_0(ces_246_0_io_ins_0),
    .io_ins_1(ces_246_0_io_ins_1),
    .io_ins_2(ces_246_0_io_ins_2),
    .io_ins_3(ces_246_0_io_ins_3),
    .io_outs_0(ces_246_0_io_outs_0),
    .io_outs_1(ces_246_0_io_outs_1),
    .io_outs_2(ces_246_0_io_outs_2),
    .io_outs_3(ces_246_0_io_outs_3)
  );
  Element ces_247_0 ( // @[MockArray.scala 36:52]
    .clock(ces_247_0_clock),
    .io_ins_0(ces_247_0_io_ins_0),
    .io_ins_1(ces_247_0_io_ins_1),
    .io_ins_2(ces_247_0_io_ins_2),
    .io_ins_3(ces_247_0_io_ins_3),
    .io_outs_0(ces_247_0_io_outs_0),
    .io_outs_1(ces_247_0_io_outs_1),
    .io_outs_2(ces_247_0_io_outs_2),
    .io_outs_3(ces_247_0_io_outs_3)
  );
  Element ces_248_0 ( // @[MockArray.scala 36:52]
    .clock(ces_248_0_clock),
    .io_ins_0(ces_248_0_io_ins_0),
    .io_ins_1(ces_248_0_io_ins_1),
    .io_ins_2(ces_248_0_io_ins_2),
    .io_ins_3(ces_248_0_io_ins_3),
    .io_outs_0(ces_248_0_io_outs_0),
    .io_outs_1(ces_248_0_io_outs_1),
    .io_outs_2(ces_248_0_io_outs_2),
    .io_outs_3(ces_248_0_io_outs_3)
  );
  Element ces_249_0 ( // @[MockArray.scala 36:52]
    .clock(ces_249_0_clock),
    .io_ins_0(ces_249_0_io_ins_0),
    .io_ins_1(ces_249_0_io_ins_1),
    .io_ins_2(ces_249_0_io_ins_2),
    .io_ins_3(ces_249_0_io_ins_3),
    .io_outs_0(ces_249_0_io_outs_0),
    .io_outs_1(ces_249_0_io_outs_1),
    .io_outs_2(ces_249_0_io_outs_2),
    .io_outs_3(ces_249_0_io_outs_3)
  );
  Element ces_250_0 ( // @[MockArray.scala 36:52]
    .clock(ces_250_0_clock),
    .io_ins_0(ces_250_0_io_ins_0),
    .io_ins_1(ces_250_0_io_ins_1),
    .io_ins_2(ces_250_0_io_ins_2),
    .io_ins_3(ces_250_0_io_ins_3),
    .io_outs_0(ces_250_0_io_outs_0),
    .io_outs_1(ces_250_0_io_outs_1),
    .io_outs_2(ces_250_0_io_outs_2),
    .io_outs_3(ces_250_0_io_outs_3)
  );
  Element ces_251_0 ( // @[MockArray.scala 36:52]
    .clock(ces_251_0_clock),
    .io_ins_0(ces_251_0_io_ins_0),
    .io_ins_1(ces_251_0_io_ins_1),
    .io_ins_2(ces_251_0_io_ins_2),
    .io_ins_3(ces_251_0_io_ins_3),
    .io_outs_0(ces_251_0_io_outs_0),
    .io_outs_1(ces_251_0_io_outs_1),
    .io_outs_2(ces_251_0_io_outs_2),
    .io_outs_3(ces_251_0_io_outs_3)
  );
  Element ces_252_0 ( // @[MockArray.scala 36:52]
    .clock(ces_252_0_clock),
    .io_ins_0(ces_252_0_io_ins_0),
    .io_ins_1(ces_252_0_io_ins_1),
    .io_ins_2(ces_252_0_io_ins_2),
    .io_ins_3(ces_252_0_io_ins_3),
    .io_outs_0(ces_252_0_io_outs_0),
    .io_outs_1(ces_252_0_io_outs_1),
    .io_outs_2(ces_252_0_io_outs_2),
    .io_outs_3(ces_252_0_io_outs_3)
  );
  Element ces_253_0 ( // @[MockArray.scala 36:52]
    .clock(ces_253_0_clock),
    .io_ins_0(ces_253_0_io_ins_0),
    .io_ins_1(ces_253_0_io_ins_1),
    .io_ins_2(ces_253_0_io_ins_2),
    .io_ins_3(ces_253_0_io_ins_3),
    .io_outs_0(ces_253_0_io_outs_0),
    .io_outs_1(ces_253_0_io_outs_1),
    .io_outs_2(ces_253_0_io_outs_2),
    .io_outs_3(ces_253_0_io_outs_3)
  );
  Element ces_254_0 ( // @[MockArray.scala 36:52]
    .clock(ces_254_0_clock),
    .io_ins_0(ces_254_0_io_ins_0),
    .io_ins_1(ces_254_0_io_ins_1),
    .io_ins_2(ces_254_0_io_ins_2),
    .io_ins_3(ces_254_0_io_ins_3),
    .io_outs_0(ces_254_0_io_outs_0),
    .io_outs_1(ces_254_0_io_outs_1),
    .io_outs_2(ces_254_0_io_outs_2),
    .io_outs_3(ces_254_0_io_outs_3)
  );
  Element ces_255_0 ( // @[MockArray.scala 36:52]
    .clock(ces_255_0_clock),
    .io_ins_0(ces_255_0_io_ins_0),
    .io_ins_1(ces_255_0_io_ins_1),
    .io_ins_2(ces_255_0_io_ins_2),
    .io_ins_3(ces_255_0_io_ins_3),
    .io_outs_0(ces_255_0_io_outs_0),
    .io_outs_1(ces_255_0_io_outs_1),
    .io_outs_2(ces_255_0_io_outs_2),
    .io_outs_3(ces_255_0_io_outs_3)
  );
  assign io_outsHorizontal_0_0 = ces_0_0_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_1_0 = ces_255_0_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_0 = ces_0_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_1 = ces_1_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_2 = ces_2_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_3 = ces_3_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_4 = ces_4_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_5 = ces_5_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_6 = ces_6_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_7 = ces_7_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_8 = ces_8_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_9 = ces_9_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_10 = ces_10_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_11 = ces_11_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_12 = ces_12_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_13 = ces_13_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_14 = ces_14_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_15 = ces_15_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_16 = ces_16_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_17 = ces_17_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_18 = ces_18_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_19 = ces_19_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_20 = ces_20_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_21 = ces_21_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_22 = ces_22_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_23 = ces_23_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_24 = ces_24_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_25 = ces_25_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_26 = ces_26_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_27 = ces_27_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_28 = ces_28_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_29 = ces_29_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_30 = ces_30_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_31 = ces_31_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_32 = ces_32_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_33 = ces_33_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_34 = ces_34_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_35 = ces_35_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_36 = ces_36_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_37 = ces_37_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_38 = ces_38_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_39 = ces_39_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_40 = ces_40_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_41 = ces_41_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_42 = ces_42_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_43 = ces_43_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_44 = ces_44_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_45 = ces_45_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_46 = ces_46_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_47 = ces_47_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_48 = ces_48_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_49 = ces_49_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_50 = ces_50_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_51 = ces_51_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_52 = ces_52_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_53 = ces_53_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_54 = ces_54_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_55 = ces_55_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_56 = ces_56_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_57 = ces_57_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_58 = ces_58_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_59 = ces_59_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_60 = ces_60_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_61 = ces_61_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_62 = ces_62_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_63 = ces_63_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_64 = ces_64_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_65 = ces_65_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_66 = ces_66_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_67 = ces_67_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_68 = ces_68_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_69 = ces_69_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_70 = ces_70_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_71 = ces_71_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_72 = ces_72_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_73 = ces_73_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_74 = ces_74_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_75 = ces_75_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_76 = ces_76_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_77 = ces_77_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_78 = ces_78_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_79 = ces_79_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_80 = ces_80_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_81 = ces_81_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_82 = ces_82_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_83 = ces_83_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_84 = ces_84_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_85 = ces_85_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_86 = ces_86_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_87 = ces_87_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_88 = ces_88_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_89 = ces_89_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_90 = ces_90_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_91 = ces_91_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_92 = ces_92_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_93 = ces_93_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_94 = ces_94_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_95 = ces_95_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_96 = ces_96_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_97 = ces_97_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_98 = ces_98_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_99 = ces_99_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_100 = ces_100_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_101 = ces_101_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_102 = ces_102_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_103 = ces_103_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_104 = ces_104_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_105 = ces_105_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_106 = ces_106_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_107 = ces_107_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_108 = ces_108_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_109 = ces_109_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_110 = ces_110_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_111 = ces_111_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_112 = ces_112_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_113 = ces_113_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_114 = ces_114_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_115 = ces_115_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_116 = ces_116_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_117 = ces_117_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_118 = ces_118_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_119 = ces_119_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_120 = ces_120_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_121 = ces_121_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_122 = ces_122_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_123 = ces_123_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_124 = ces_124_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_125 = ces_125_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_126 = ces_126_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_127 = ces_127_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_128 = ces_128_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_129 = ces_129_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_130 = ces_130_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_131 = ces_131_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_132 = ces_132_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_133 = ces_133_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_134 = ces_134_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_135 = ces_135_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_136 = ces_136_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_137 = ces_137_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_138 = ces_138_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_139 = ces_139_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_140 = ces_140_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_141 = ces_141_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_142 = ces_142_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_143 = ces_143_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_144 = ces_144_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_145 = ces_145_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_146 = ces_146_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_147 = ces_147_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_148 = ces_148_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_149 = ces_149_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_150 = ces_150_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_151 = ces_151_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_152 = ces_152_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_153 = ces_153_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_154 = ces_154_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_155 = ces_155_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_156 = ces_156_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_157 = ces_157_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_158 = ces_158_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_159 = ces_159_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_160 = ces_160_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_161 = ces_161_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_162 = ces_162_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_163 = ces_163_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_164 = ces_164_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_165 = ces_165_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_166 = ces_166_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_167 = ces_167_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_168 = ces_168_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_169 = ces_169_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_170 = ces_170_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_171 = ces_171_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_172 = ces_172_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_173 = ces_173_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_174 = ces_174_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_175 = ces_175_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_176 = ces_176_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_177 = ces_177_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_178 = ces_178_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_179 = ces_179_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_180 = ces_180_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_181 = ces_181_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_182 = ces_182_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_183 = ces_183_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_184 = ces_184_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_185 = ces_185_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_186 = ces_186_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_187 = ces_187_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_188 = ces_188_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_189 = ces_189_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_190 = ces_190_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_191 = ces_191_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_192 = ces_192_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_193 = ces_193_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_194 = ces_194_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_195 = ces_195_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_196 = ces_196_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_197 = ces_197_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_198 = ces_198_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_199 = ces_199_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_200 = ces_200_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_201 = ces_201_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_202 = ces_202_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_203 = ces_203_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_204 = ces_204_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_205 = ces_205_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_206 = ces_206_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_207 = ces_207_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_208 = ces_208_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_209 = ces_209_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_210 = ces_210_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_211 = ces_211_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_212 = ces_212_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_213 = ces_213_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_214 = ces_214_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_215 = ces_215_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_216 = ces_216_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_217 = ces_217_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_218 = ces_218_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_219 = ces_219_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_220 = ces_220_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_221 = ces_221_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_222 = ces_222_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_223 = ces_223_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_224 = ces_224_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_225 = ces_225_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_226 = ces_226_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_227 = ces_227_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_228 = ces_228_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_229 = ces_229_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_230 = ces_230_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_231 = ces_231_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_232 = ces_232_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_233 = ces_233_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_234 = ces_234_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_235 = ces_235_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_236 = ces_236_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_237 = ces_237_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_238 = ces_238_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_239 = ces_239_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_240 = ces_240_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_241 = ces_241_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_242 = ces_242_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_243 = ces_243_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_244 = ces_244_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_245 = ces_245_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_246 = ces_246_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_247 = ces_247_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_248 = ces_248_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_249 = ces_249_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_250 = ces_250_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_251 = ces_251_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_252 = ces_252_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_253 = ces_253_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_254 = ces_254_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_255 = ces_255_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_1_0 = ces_0_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_1 = ces_1_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_2 = ces_2_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_3 = ces_3_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_4 = ces_4_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_5 = ces_5_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_6 = ces_6_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_7 = ces_7_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_8 = ces_8_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_9 = ces_9_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_10 = ces_10_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_11 = ces_11_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_12 = ces_12_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_13 = ces_13_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_14 = ces_14_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_15 = ces_15_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_16 = ces_16_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_17 = ces_17_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_18 = ces_18_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_19 = ces_19_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_20 = ces_20_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_21 = ces_21_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_22 = ces_22_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_23 = ces_23_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_24 = ces_24_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_25 = ces_25_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_26 = ces_26_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_27 = ces_27_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_28 = ces_28_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_29 = ces_29_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_30 = ces_30_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_31 = ces_31_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_32 = ces_32_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_33 = ces_33_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_34 = ces_34_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_35 = ces_35_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_36 = ces_36_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_37 = ces_37_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_38 = ces_38_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_39 = ces_39_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_40 = ces_40_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_41 = ces_41_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_42 = ces_42_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_43 = ces_43_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_44 = ces_44_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_45 = ces_45_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_46 = ces_46_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_47 = ces_47_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_48 = ces_48_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_49 = ces_49_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_50 = ces_50_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_51 = ces_51_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_52 = ces_52_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_53 = ces_53_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_54 = ces_54_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_55 = ces_55_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_56 = ces_56_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_57 = ces_57_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_58 = ces_58_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_59 = ces_59_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_60 = ces_60_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_61 = ces_61_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_62 = ces_62_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_63 = ces_63_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_64 = ces_64_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_65 = ces_65_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_66 = ces_66_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_67 = ces_67_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_68 = ces_68_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_69 = ces_69_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_70 = ces_70_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_71 = ces_71_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_72 = ces_72_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_73 = ces_73_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_74 = ces_74_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_75 = ces_75_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_76 = ces_76_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_77 = ces_77_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_78 = ces_78_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_79 = ces_79_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_80 = ces_80_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_81 = ces_81_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_82 = ces_82_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_83 = ces_83_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_84 = ces_84_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_85 = ces_85_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_86 = ces_86_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_87 = ces_87_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_88 = ces_88_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_89 = ces_89_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_90 = ces_90_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_91 = ces_91_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_92 = ces_92_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_93 = ces_93_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_94 = ces_94_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_95 = ces_95_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_96 = ces_96_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_97 = ces_97_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_98 = ces_98_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_99 = ces_99_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_100 = ces_100_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_101 = ces_101_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_102 = ces_102_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_103 = ces_103_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_104 = ces_104_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_105 = ces_105_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_106 = ces_106_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_107 = ces_107_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_108 = ces_108_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_109 = ces_109_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_110 = ces_110_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_111 = ces_111_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_112 = ces_112_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_113 = ces_113_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_114 = ces_114_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_115 = ces_115_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_116 = ces_116_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_117 = ces_117_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_118 = ces_118_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_119 = ces_119_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_120 = ces_120_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_121 = ces_121_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_122 = ces_122_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_123 = ces_123_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_124 = ces_124_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_125 = ces_125_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_126 = ces_126_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_127 = ces_127_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_128 = ces_128_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_129 = ces_129_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_130 = ces_130_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_131 = ces_131_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_132 = ces_132_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_133 = ces_133_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_134 = ces_134_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_135 = ces_135_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_136 = ces_136_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_137 = ces_137_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_138 = ces_138_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_139 = ces_139_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_140 = ces_140_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_141 = ces_141_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_142 = ces_142_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_143 = ces_143_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_144 = ces_144_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_145 = ces_145_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_146 = ces_146_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_147 = ces_147_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_148 = ces_148_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_149 = ces_149_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_150 = ces_150_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_151 = ces_151_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_152 = ces_152_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_153 = ces_153_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_154 = ces_154_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_155 = ces_155_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_156 = ces_156_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_157 = ces_157_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_158 = ces_158_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_159 = ces_159_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_160 = ces_160_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_161 = ces_161_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_162 = ces_162_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_163 = ces_163_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_164 = ces_164_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_165 = ces_165_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_166 = ces_166_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_167 = ces_167_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_168 = ces_168_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_169 = ces_169_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_170 = ces_170_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_171 = ces_171_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_172 = ces_172_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_173 = ces_173_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_174 = ces_174_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_175 = ces_175_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_176 = ces_176_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_177 = ces_177_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_178 = ces_178_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_179 = ces_179_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_180 = ces_180_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_181 = ces_181_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_182 = ces_182_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_183 = ces_183_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_184 = ces_184_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_185 = ces_185_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_186 = ces_186_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_187 = ces_187_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_188 = ces_188_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_189 = ces_189_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_190 = ces_190_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_191 = ces_191_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_192 = ces_192_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_193 = ces_193_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_194 = ces_194_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_195 = ces_195_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_196 = ces_196_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_197 = ces_197_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_198 = ces_198_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_199 = ces_199_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_200 = ces_200_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_201 = ces_201_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_202 = ces_202_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_203 = ces_203_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_204 = ces_204_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_205 = ces_205_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_206 = ces_206_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_207 = ces_207_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_208 = ces_208_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_209 = ces_209_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_210 = ces_210_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_211 = ces_211_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_212 = ces_212_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_213 = ces_213_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_214 = ces_214_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_215 = ces_215_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_216 = ces_216_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_217 = ces_217_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_218 = ces_218_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_219 = ces_219_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_220 = ces_220_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_221 = ces_221_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_222 = ces_222_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_223 = ces_223_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_224 = ces_224_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_225 = ces_225_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_226 = ces_226_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_227 = ces_227_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_228 = ces_228_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_229 = ces_229_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_230 = ces_230_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_231 = ces_231_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_232 = ces_232_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_233 = ces_233_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_234 = ces_234_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_235 = ces_235_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_236 = ces_236_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_237 = ces_237_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_238 = ces_238_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_239 = ces_239_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_240 = ces_240_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_241 = ces_241_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_242 = ces_242_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_243 = ces_243_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_244 = ces_244_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_245 = ces_245_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_246 = ces_246_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_247 = ces_247_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_248 = ces_248_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_249 = ces_249_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_250 = ces_250_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_251 = ces_251_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_252 = ces_252_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_253 = ces_253_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_254 = ces_254_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_255 = ces_255_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_lsbs_0 = ces_0_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1 = ces_1_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_2 = ces_2_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_3 = ces_3_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_4 = ces_4_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_5 = ces_5_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_6 = ces_6_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_7 = ces_7_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_8 = ces_8_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_9 = ces_9_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_10 = ces_10_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_11 = ces_11_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_12 = ces_12_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_13 = ces_13_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_14 = ces_14_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_15 = ces_15_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_16 = ces_16_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_17 = ces_17_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_18 = ces_18_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_19 = ces_19_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_20 = ces_20_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_21 = ces_21_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_22 = ces_22_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_23 = ces_23_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_24 = ces_24_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_25 = ces_25_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_26 = ces_26_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_27 = ces_27_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_28 = ces_28_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_29 = ces_29_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_30 = ces_30_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_31 = ces_31_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_32 = ces_32_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_33 = ces_33_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_34 = ces_34_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_35 = ces_35_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_36 = ces_36_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_37 = ces_37_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_38 = ces_38_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_39 = ces_39_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_40 = ces_40_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_41 = ces_41_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_42 = ces_42_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_43 = ces_43_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_44 = ces_44_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_45 = ces_45_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_46 = ces_46_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_47 = ces_47_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_48 = ces_48_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_49 = ces_49_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_50 = ces_50_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_51 = ces_51_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_52 = ces_52_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_53 = ces_53_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_54 = ces_54_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_55 = ces_55_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_56 = ces_56_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_57 = ces_57_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_58 = ces_58_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_59 = ces_59_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_60 = ces_60_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_61 = ces_61_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_62 = ces_62_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_63 = ces_63_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_64 = ces_64_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_65 = ces_65_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_66 = ces_66_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_67 = ces_67_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_68 = ces_68_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_69 = ces_69_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_70 = ces_70_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_71 = ces_71_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_72 = ces_72_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_73 = ces_73_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_74 = ces_74_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_75 = ces_75_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_76 = ces_76_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_77 = ces_77_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_78 = ces_78_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_79 = ces_79_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_80 = ces_80_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_81 = ces_81_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_82 = ces_82_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_83 = ces_83_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_84 = ces_84_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_85 = ces_85_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_86 = ces_86_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_87 = ces_87_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_88 = ces_88_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_89 = ces_89_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_90 = ces_90_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_91 = ces_91_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_92 = ces_92_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_93 = ces_93_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_94 = ces_94_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_95 = ces_95_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_96 = ces_96_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_97 = ces_97_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_98 = ces_98_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_99 = ces_99_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_100 = ces_100_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_101 = ces_101_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_102 = ces_102_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_103 = ces_103_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_104 = ces_104_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_105 = ces_105_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_106 = ces_106_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_107 = ces_107_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_108 = ces_108_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_109 = ces_109_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_110 = ces_110_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_111 = ces_111_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_112 = ces_112_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_113 = ces_113_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_114 = ces_114_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_115 = ces_115_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_116 = ces_116_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_117 = ces_117_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_118 = ces_118_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_119 = ces_119_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_120 = ces_120_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_121 = ces_121_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_122 = ces_122_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_123 = ces_123_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_124 = ces_124_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_125 = ces_125_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_126 = ces_126_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_127 = ces_127_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_128 = ces_128_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_129 = ces_129_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_130 = ces_130_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_131 = ces_131_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_132 = ces_132_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_133 = ces_133_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_134 = ces_134_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_135 = ces_135_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_136 = ces_136_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_137 = ces_137_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_138 = ces_138_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_139 = ces_139_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_140 = ces_140_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_141 = ces_141_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_142 = ces_142_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_143 = ces_143_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_144 = ces_144_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_145 = ces_145_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_146 = ces_146_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_147 = ces_147_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_148 = ces_148_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_149 = ces_149_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_150 = ces_150_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_151 = ces_151_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_152 = ces_152_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_153 = ces_153_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_154 = ces_154_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_155 = ces_155_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_156 = ces_156_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_157 = ces_157_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_158 = ces_158_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_159 = ces_159_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_160 = ces_160_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_161 = ces_161_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_162 = ces_162_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_163 = ces_163_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_164 = ces_164_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_165 = ces_165_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_166 = ces_166_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_167 = ces_167_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_168 = ces_168_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_169 = ces_169_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_170 = ces_170_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_171 = ces_171_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_172 = ces_172_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_173 = ces_173_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_174 = ces_174_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_175 = ces_175_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_176 = ces_176_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_177 = ces_177_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_178 = ces_178_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_179 = ces_179_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_180 = ces_180_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_181 = ces_181_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_182 = ces_182_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_183 = ces_183_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_184 = ces_184_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_185 = ces_185_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_186 = ces_186_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_187 = ces_187_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_188 = ces_188_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_189 = ces_189_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_190 = ces_190_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_191 = ces_191_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_192 = ces_192_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_193 = ces_193_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_194 = ces_194_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_195 = ces_195_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_196 = ces_196_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_197 = ces_197_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_198 = ces_198_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_199 = ces_199_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_200 = ces_200_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_201 = ces_201_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_202 = ces_202_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_203 = ces_203_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_204 = ces_204_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_205 = ces_205_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_206 = ces_206_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_207 = ces_207_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_208 = ces_208_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_209 = ces_209_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_210 = ces_210_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_211 = ces_211_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_212 = ces_212_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_213 = ces_213_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_214 = ces_214_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_215 = ces_215_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_216 = ces_216_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_217 = ces_217_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_218 = ces_218_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_219 = ces_219_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_220 = ces_220_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_221 = ces_221_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_222 = ces_222_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_223 = ces_223_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_224 = ces_224_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_225 = ces_225_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_226 = ces_226_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_227 = ces_227_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_228 = ces_228_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_229 = ces_229_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_230 = ces_230_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_231 = ces_231_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_232 = ces_232_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_233 = ces_233_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_234 = ces_234_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_235 = ces_235_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_236 = ces_236_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_237 = ces_237_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_238 = ces_238_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_239 = ces_239_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_240 = ces_240_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_241 = ces_241_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_242 = ces_242_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_243 = ces_243_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_244 = ces_244_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_245 = ces_245_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_246 = ces_246_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_247 = ces_247_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_248 = ces_248_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_249 = ces_249_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_250 = ces_250_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_251 = ces_251_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_252 = ces_252_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_253 = ces_253_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_254 = ces_254_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_255 = ces_255_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign ces_0_0_clock = clock;
  assign ces_0_0_io_ins_0 = io_insHorizontal_0_0; // @[MockArray.scala 44:87]
  assign ces_0_0_io_ins_1 = io_insVertical_0_0; // @[MockArray.scala 45:87]
  assign ces_0_0_io_ins_2 = ces_1_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_0_io_ins_3 = io_insVertical_1_0; // @[MockArray.scala 47:87]
  assign ces_1_0_clock = clock;
  assign ces_1_0_io_ins_0 = ces_0_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_0_io_ins_1 = io_insVertical_0_1; // @[MockArray.scala 45:87]
  assign ces_1_0_io_ins_2 = ces_2_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_0_io_ins_3 = io_insVertical_1_1; // @[MockArray.scala 47:87]
  assign ces_2_0_clock = clock;
  assign ces_2_0_io_ins_0 = ces_1_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_0_io_ins_1 = io_insVertical_0_2; // @[MockArray.scala 45:87]
  assign ces_2_0_io_ins_2 = ces_3_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_0_io_ins_3 = io_insVertical_1_2; // @[MockArray.scala 47:87]
  assign ces_3_0_clock = clock;
  assign ces_3_0_io_ins_0 = ces_2_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_0_io_ins_1 = io_insVertical_0_3; // @[MockArray.scala 45:87]
  assign ces_3_0_io_ins_2 = ces_4_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_0_io_ins_3 = io_insVertical_1_3; // @[MockArray.scala 47:87]
  assign ces_4_0_clock = clock;
  assign ces_4_0_io_ins_0 = ces_3_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_0_io_ins_1 = io_insVertical_0_4; // @[MockArray.scala 45:87]
  assign ces_4_0_io_ins_2 = ces_5_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_0_io_ins_3 = io_insVertical_1_4; // @[MockArray.scala 47:87]
  assign ces_5_0_clock = clock;
  assign ces_5_0_io_ins_0 = ces_4_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_0_io_ins_1 = io_insVertical_0_5; // @[MockArray.scala 45:87]
  assign ces_5_0_io_ins_2 = ces_6_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_0_io_ins_3 = io_insVertical_1_5; // @[MockArray.scala 47:87]
  assign ces_6_0_clock = clock;
  assign ces_6_0_io_ins_0 = ces_5_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_0_io_ins_1 = io_insVertical_0_6; // @[MockArray.scala 45:87]
  assign ces_6_0_io_ins_2 = ces_7_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_0_io_ins_3 = io_insVertical_1_6; // @[MockArray.scala 47:87]
  assign ces_7_0_clock = clock;
  assign ces_7_0_io_ins_0 = ces_6_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_0_io_ins_1 = io_insVertical_0_7; // @[MockArray.scala 45:87]
  assign ces_7_0_io_ins_2 = ces_8_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_0_io_ins_3 = io_insVertical_1_7; // @[MockArray.scala 47:87]
  assign ces_8_0_clock = clock;
  assign ces_8_0_io_ins_0 = ces_7_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_0_io_ins_1 = io_insVertical_0_8; // @[MockArray.scala 45:87]
  assign ces_8_0_io_ins_2 = ces_9_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_0_io_ins_3 = io_insVertical_1_8; // @[MockArray.scala 47:87]
  assign ces_9_0_clock = clock;
  assign ces_9_0_io_ins_0 = ces_8_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_0_io_ins_1 = io_insVertical_0_9; // @[MockArray.scala 45:87]
  assign ces_9_0_io_ins_2 = ces_10_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_0_io_ins_3 = io_insVertical_1_9; // @[MockArray.scala 47:87]
  assign ces_10_0_clock = clock;
  assign ces_10_0_io_ins_0 = ces_9_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_0_io_ins_1 = io_insVertical_0_10; // @[MockArray.scala 45:87]
  assign ces_10_0_io_ins_2 = ces_11_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_0_io_ins_3 = io_insVertical_1_10; // @[MockArray.scala 47:87]
  assign ces_11_0_clock = clock;
  assign ces_11_0_io_ins_0 = ces_10_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_0_io_ins_1 = io_insVertical_0_11; // @[MockArray.scala 45:87]
  assign ces_11_0_io_ins_2 = ces_12_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_0_io_ins_3 = io_insVertical_1_11; // @[MockArray.scala 47:87]
  assign ces_12_0_clock = clock;
  assign ces_12_0_io_ins_0 = ces_11_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_0_io_ins_1 = io_insVertical_0_12; // @[MockArray.scala 45:87]
  assign ces_12_0_io_ins_2 = ces_13_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_0_io_ins_3 = io_insVertical_1_12; // @[MockArray.scala 47:87]
  assign ces_13_0_clock = clock;
  assign ces_13_0_io_ins_0 = ces_12_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_0_io_ins_1 = io_insVertical_0_13; // @[MockArray.scala 45:87]
  assign ces_13_0_io_ins_2 = ces_14_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_0_io_ins_3 = io_insVertical_1_13; // @[MockArray.scala 47:87]
  assign ces_14_0_clock = clock;
  assign ces_14_0_io_ins_0 = ces_13_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_0_io_ins_1 = io_insVertical_0_14; // @[MockArray.scala 45:87]
  assign ces_14_0_io_ins_2 = ces_15_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_0_io_ins_3 = io_insVertical_1_14; // @[MockArray.scala 47:87]
  assign ces_15_0_clock = clock;
  assign ces_15_0_io_ins_0 = ces_14_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_0_io_ins_1 = io_insVertical_0_15; // @[MockArray.scala 45:87]
  assign ces_15_0_io_ins_2 = ces_16_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_0_io_ins_3 = io_insVertical_1_15; // @[MockArray.scala 47:87]
  assign ces_16_0_clock = clock;
  assign ces_16_0_io_ins_0 = ces_15_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_0_io_ins_1 = io_insVertical_0_16; // @[MockArray.scala 45:87]
  assign ces_16_0_io_ins_2 = ces_17_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_0_io_ins_3 = io_insVertical_1_16; // @[MockArray.scala 47:87]
  assign ces_17_0_clock = clock;
  assign ces_17_0_io_ins_0 = ces_16_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_0_io_ins_1 = io_insVertical_0_17; // @[MockArray.scala 45:87]
  assign ces_17_0_io_ins_2 = ces_18_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_0_io_ins_3 = io_insVertical_1_17; // @[MockArray.scala 47:87]
  assign ces_18_0_clock = clock;
  assign ces_18_0_io_ins_0 = ces_17_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_0_io_ins_1 = io_insVertical_0_18; // @[MockArray.scala 45:87]
  assign ces_18_0_io_ins_2 = ces_19_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_0_io_ins_3 = io_insVertical_1_18; // @[MockArray.scala 47:87]
  assign ces_19_0_clock = clock;
  assign ces_19_0_io_ins_0 = ces_18_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_0_io_ins_1 = io_insVertical_0_19; // @[MockArray.scala 45:87]
  assign ces_19_0_io_ins_2 = ces_20_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_0_io_ins_3 = io_insVertical_1_19; // @[MockArray.scala 47:87]
  assign ces_20_0_clock = clock;
  assign ces_20_0_io_ins_0 = ces_19_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_0_io_ins_1 = io_insVertical_0_20; // @[MockArray.scala 45:87]
  assign ces_20_0_io_ins_2 = ces_21_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_0_io_ins_3 = io_insVertical_1_20; // @[MockArray.scala 47:87]
  assign ces_21_0_clock = clock;
  assign ces_21_0_io_ins_0 = ces_20_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_0_io_ins_1 = io_insVertical_0_21; // @[MockArray.scala 45:87]
  assign ces_21_0_io_ins_2 = ces_22_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_0_io_ins_3 = io_insVertical_1_21; // @[MockArray.scala 47:87]
  assign ces_22_0_clock = clock;
  assign ces_22_0_io_ins_0 = ces_21_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_0_io_ins_1 = io_insVertical_0_22; // @[MockArray.scala 45:87]
  assign ces_22_0_io_ins_2 = ces_23_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_0_io_ins_3 = io_insVertical_1_22; // @[MockArray.scala 47:87]
  assign ces_23_0_clock = clock;
  assign ces_23_0_io_ins_0 = ces_22_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_0_io_ins_1 = io_insVertical_0_23; // @[MockArray.scala 45:87]
  assign ces_23_0_io_ins_2 = ces_24_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_0_io_ins_3 = io_insVertical_1_23; // @[MockArray.scala 47:87]
  assign ces_24_0_clock = clock;
  assign ces_24_0_io_ins_0 = ces_23_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_0_io_ins_1 = io_insVertical_0_24; // @[MockArray.scala 45:87]
  assign ces_24_0_io_ins_2 = ces_25_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_0_io_ins_3 = io_insVertical_1_24; // @[MockArray.scala 47:87]
  assign ces_25_0_clock = clock;
  assign ces_25_0_io_ins_0 = ces_24_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_0_io_ins_1 = io_insVertical_0_25; // @[MockArray.scala 45:87]
  assign ces_25_0_io_ins_2 = ces_26_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_0_io_ins_3 = io_insVertical_1_25; // @[MockArray.scala 47:87]
  assign ces_26_0_clock = clock;
  assign ces_26_0_io_ins_0 = ces_25_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_0_io_ins_1 = io_insVertical_0_26; // @[MockArray.scala 45:87]
  assign ces_26_0_io_ins_2 = ces_27_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_0_io_ins_3 = io_insVertical_1_26; // @[MockArray.scala 47:87]
  assign ces_27_0_clock = clock;
  assign ces_27_0_io_ins_0 = ces_26_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_0_io_ins_1 = io_insVertical_0_27; // @[MockArray.scala 45:87]
  assign ces_27_0_io_ins_2 = ces_28_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_0_io_ins_3 = io_insVertical_1_27; // @[MockArray.scala 47:87]
  assign ces_28_0_clock = clock;
  assign ces_28_0_io_ins_0 = ces_27_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_0_io_ins_1 = io_insVertical_0_28; // @[MockArray.scala 45:87]
  assign ces_28_0_io_ins_2 = ces_29_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_0_io_ins_3 = io_insVertical_1_28; // @[MockArray.scala 47:87]
  assign ces_29_0_clock = clock;
  assign ces_29_0_io_ins_0 = ces_28_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_0_io_ins_1 = io_insVertical_0_29; // @[MockArray.scala 45:87]
  assign ces_29_0_io_ins_2 = ces_30_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_0_io_ins_3 = io_insVertical_1_29; // @[MockArray.scala 47:87]
  assign ces_30_0_clock = clock;
  assign ces_30_0_io_ins_0 = ces_29_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_0_io_ins_1 = io_insVertical_0_30; // @[MockArray.scala 45:87]
  assign ces_30_0_io_ins_2 = ces_31_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_0_io_ins_3 = io_insVertical_1_30; // @[MockArray.scala 47:87]
  assign ces_31_0_clock = clock;
  assign ces_31_0_io_ins_0 = ces_30_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_0_io_ins_1 = io_insVertical_0_31; // @[MockArray.scala 45:87]
  assign ces_31_0_io_ins_2 = ces_32_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_31_0_io_ins_3 = io_insVertical_1_31; // @[MockArray.scala 47:87]
  assign ces_32_0_clock = clock;
  assign ces_32_0_io_ins_0 = ces_31_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_32_0_io_ins_1 = io_insVertical_0_32; // @[MockArray.scala 45:87]
  assign ces_32_0_io_ins_2 = ces_33_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_32_0_io_ins_3 = io_insVertical_1_32; // @[MockArray.scala 47:87]
  assign ces_33_0_clock = clock;
  assign ces_33_0_io_ins_0 = ces_32_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_33_0_io_ins_1 = io_insVertical_0_33; // @[MockArray.scala 45:87]
  assign ces_33_0_io_ins_2 = ces_34_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_33_0_io_ins_3 = io_insVertical_1_33; // @[MockArray.scala 47:87]
  assign ces_34_0_clock = clock;
  assign ces_34_0_io_ins_0 = ces_33_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_34_0_io_ins_1 = io_insVertical_0_34; // @[MockArray.scala 45:87]
  assign ces_34_0_io_ins_2 = ces_35_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_34_0_io_ins_3 = io_insVertical_1_34; // @[MockArray.scala 47:87]
  assign ces_35_0_clock = clock;
  assign ces_35_0_io_ins_0 = ces_34_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_35_0_io_ins_1 = io_insVertical_0_35; // @[MockArray.scala 45:87]
  assign ces_35_0_io_ins_2 = ces_36_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_35_0_io_ins_3 = io_insVertical_1_35; // @[MockArray.scala 47:87]
  assign ces_36_0_clock = clock;
  assign ces_36_0_io_ins_0 = ces_35_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_36_0_io_ins_1 = io_insVertical_0_36; // @[MockArray.scala 45:87]
  assign ces_36_0_io_ins_2 = ces_37_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_36_0_io_ins_3 = io_insVertical_1_36; // @[MockArray.scala 47:87]
  assign ces_37_0_clock = clock;
  assign ces_37_0_io_ins_0 = ces_36_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_37_0_io_ins_1 = io_insVertical_0_37; // @[MockArray.scala 45:87]
  assign ces_37_0_io_ins_2 = ces_38_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_37_0_io_ins_3 = io_insVertical_1_37; // @[MockArray.scala 47:87]
  assign ces_38_0_clock = clock;
  assign ces_38_0_io_ins_0 = ces_37_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_38_0_io_ins_1 = io_insVertical_0_38; // @[MockArray.scala 45:87]
  assign ces_38_0_io_ins_2 = ces_39_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_38_0_io_ins_3 = io_insVertical_1_38; // @[MockArray.scala 47:87]
  assign ces_39_0_clock = clock;
  assign ces_39_0_io_ins_0 = ces_38_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_39_0_io_ins_1 = io_insVertical_0_39; // @[MockArray.scala 45:87]
  assign ces_39_0_io_ins_2 = ces_40_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_39_0_io_ins_3 = io_insVertical_1_39; // @[MockArray.scala 47:87]
  assign ces_40_0_clock = clock;
  assign ces_40_0_io_ins_0 = ces_39_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_40_0_io_ins_1 = io_insVertical_0_40; // @[MockArray.scala 45:87]
  assign ces_40_0_io_ins_2 = ces_41_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_40_0_io_ins_3 = io_insVertical_1_40; // @[MockArray.scala 47:87]
  assign ces_41_0_clock = clock;
  assign ces_41_0_io_ins_0 = ces_40_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_41_0_io_ins_1 = io_insVertical_0_41; // @[MockArray.scala 45:87]
  assign ces_41_0_io_ins_2 = ces_42_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_41_0_io_ins_3 = io_insVertical_1_41; // @[MockArray.scala 47:87]
  assign ces_42_0_clock = clock;
  assign ces_42_0_io_ins_0 = ces_41_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_42_0_io_ins_1 = io_insVertical_0_42; // @[MockArray.scala 45:87]
  assign ces_42_0_io_ins_2 = ces_43_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_42_0_io_ins_3 = io_insVertical_1_42; // @[MockArray.scala 47:87]
  assign ces_43_0_clock = clock;
  assign ces_43_0_io_ins_0 = ces_42_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_43_0_io_ins_1 = io_insVertical_0_43; // @[MockArray.scala 45:87]
  assign ces_43_0_io_ins_2 = ces_44_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_43_0_io_ins_3 = io_insVertical_1_43; // @[MockArray.scala 47:87]
  assign ces_44_0_clock = clock;
  assign ces_44_0_io_ins_0 = ces_43_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_44_0_io_ins_1 = io_insVertical_0_44; // @[MockArray.scala 45:87]
  assign ces_44_0_io_ins_2 = ces_45_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_44_0_io_ins_3 = io_insVertical_1_44; // @[MockArray.scala 47:87]
  assign ces_45_0_clock = clock;
  assign ces_45_0_io_ins_0 = ces_44_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_45_0_io_ins_1 = io_insVertical_0_45; // @[MockArray.scala 45:87]
  assign ces_45_0_io_ins_2 = ces_46_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_45_0_io_ins_3 = io_insVertical_1_45; // @[MockArray.scala 47:87]
  assign ces_46_0_clock = clock;
  assign ces_46_0_io_ins_0 = ces_45_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_46_0_io_ins_1 = io_insVertical_0_46; // @[MockArray.scala 45:87]
  assign ces_46_0_io_ins_2 = ces_47_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_46_0_io_ins_3 = io_insVertical_1_46; // @[MockArray.scala 47:87]
  assign ces_47_0_clock = clock;
  assign ces_47_0_io_ins_0 = ces_46_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_47_0_io_ins_1 = io_insVertical_0_47; // @[MockArray.scala 45:87]
  assign ces_47_0_io_ins_2 = ces_48_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_47_0_io_ins_3 = io_insVertical_1_47; // @[MockArray.scala 47:87]
  assign ces_48_0_clock = clock;
  assign ces_48_0_io_ins_0 = ces_47_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_48_0_io_ins_1 = io_insVertical_0_48; // @[MockArray.scala 45:87]
  assign ces_48_0_io_ins_2 = ces_49_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_48_0_io_ins_3 = io_insVertical_1_48; // @[MockArray.scala 47:87]
  assign ces_49_0_clock = clock;
  assign ces_49_0_io_ins_0 = ces_48_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_49_0_io_ins_1 = io_insVertical_0_49; // @[MockArray.scala 45:87]
  assign ces_49_0_io_ins_2 = ces_50_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_49_0_io_ins_3 = io_insVertical_1_49; // @[MockArray.scala 47:87]
  assign ces_50_0_clock = clock;
  assign ces_50_0_io_ins_0 = ces_49_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_50_0_io_ins_1 = io_insVertical_0_50; // @[MockArray.scala 45:87]
  assign ces_50_0_io_ins_2 = ces_51_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_50_0_io_ins_3 = io_insVertical_1_50; // @[MockArray.scala 47:87]
  assign ces_51_0_clock = clock;
  assign ces_51_0_io_ins_0 = ces_50_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_51_0_io_ins_1 = io_insVertical_0_51; // @[MockArray.scala 45:87]
  assign ces_51_0_io_ins_2 = ces_52_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_51_0_io_ins_3 = io_insVertical_1_51; // @[MockArray.scala 47:87]
  assign ces_52_0_clock = clock;
  assign ces_52_0_io_ins_0 = ces_51_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_52_0_io_ins_1 = io_insVertical_0_52; // @[MockArray.scala 45:87]
  assign ces_52_0_io_ins_2 = ces_53_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_52_0_io_ins_3 = io_insVertical_1_52; // @[MockArray.scala 47:87]
  assign ces_53_0_clock = clock;
  assign ces_53_0_io_ins_0 = ces_52_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_53_0_io_ins_1 = io_insVertical_0_53; // @[MockArray.scala 45:87]
  assign ces_53_0_io_ins_2 = ces_54_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_53_0_io_ins_3 = io_insVertical_1_53; // @[MockArray.scala 47:87]
  assign ces_54_0_clock = clock;
  assign ces_54_0_io_ins_0 = ces_53_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_54_0_io_ins_1 = io_insVertical_0_54; // @[MockArray.scala 45:87]
  assign ces_54_0_io_ins_2 = ces_55_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_54_0_io_ins_3 = io_insVertical_1_54; // @[MockArray.scala 47:87]
  assign ces_55_0_clock = clock;
  assign ces_55_0_io_ins_0 = ces_54_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_55_0_io_ins_1 = io_insVertical_0_55; // @[MockArray.scala 45:87]
  assign ces_55_0_io_ins_2 = ces_56_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_55_0_io_ins_3 = io_insVertical_1_55; // @[MockArray.scala 47:87]
  assign ces_56_0_clock = clock;
  assign ces_56_0_io_ins_0 = ces_55_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_56_0_io_ins_1 = io_insVertical_0_56; // @[MockArray.scala 45:87]
  assign ces_56_0_io_ins_2 = ces_57_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_56_0_io_ins_3 = io_insVertical_1_56; // @[MockArray.scala 47:87]
  assign ces_57_0_clock = clock;
  assign ces_57_0_io_ins_0 = ces_56_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_57_0_io_ins_1 = io_insVertical_0_57; // @[MockArray.scala 45:87]
  assign ces_57_0_io_ins_2 = ces_58_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_57_0_io_ins_3 = io_insVertical_1_57; // @[MockArray.scala 47:87]
  assign ces_58_0_clock = clock;
  assign ces_58_0_io_ins_0 = ces_57_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_58_0_io_ins_1 = io_insVertical_0_58; // @[MockArray.scala 45:87]
  assign ces_58_0_io_ins_2 = ces_59_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_58_0_io_ins_3 = io_insVertical_1_58; // @[MockArray.scala 47:87]
  assign ces_59_0_clock = clock;
  assign ces_59_0_io_ins_0 = ces_58_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_59_0_io_ins_1 = io_insVertical_0_59; // @[MockArray.scala 45:87]
  assign ces_59_0_io_ins_2 = ces_60_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_59_0_io_ins_3 = io_insVertical_1_59; // @[MockArray.scala 47:87]
  assign ces_60_0_clock = clock;
  assign ces_60_0_io_ins_0 = ces_59_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_60_0_io_ins_1 = io_insVertical_0_60; // @[MockArray.scala 45:87]
  assign ces_60_0_io_ins_2 = ces_61_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_60_0_io_ins_3 = io_insVertical_1_60; // @[MockArray.scala 47:87]
  assign ces_61_0_clock = clock;
  assign ces_61_0_io_ins_0 = ces_60_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_61_0_io_ins_1 = io_insVertical_0_61; // @[MockArray.scala 45:87]
  assign ces_61_0_io_ins_2 = ces_62_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_61_0_io_ins_3 = io_insVertical_1_61; // @[MockArray.scala 47:87]
  assign ces_62_0_clock = clock;
  assign ces_62_0_io_ins_0 = ces_61_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_62_0_io_ins_1 = io_insVertical_0_62; // @[MockArray.scala 45:87]
  assign ces_62_0_io_ins_2 = ces_63_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_62_0_io_ins_3 = io_insVertical_1_62; // @[MockArray.scala 47:87]
  assign ces_63_0_clock = clock;
  assign ces_63_0_io_ins_0 = ces_62_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_63_0_io_ins_1 = io_insVertical_0_63; // @[MockArray.scala 45:87]
  assign ces_63_0_io_ins_2 = ces_64_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_63_0_io_ins_3 = io_insVertical_1_63; // @[MockArray.scala 47:87]
  assign ces_64_0_clock = clock;
  assign ces_64_0_io_ins_0 = ces_63_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_64_0_io_ins_1 = io_insVertical_0_64; // @[MockArray.scala 45:87]
  assign ces_64_0_io_ins_2 = ces_65_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_64_0_io_ins_3 = io_insVertical_1_64; // @[MockArray.scala 47:87]
  assign ces_65_0_clock = clock;
  assign ces_65_0_io_ins_0 = ces_64_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_65_0_io_ins_1 = io_insVertical_0_65; // @[MockArray.scala 45:87]
  assign ces_65_0_io_ins_2 = ces_66_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_65_0_io_ins_3 = io_insVertical_1_65; // @[MockArray.scala 47:87]
  assign ces_66_0_clock = clock;
  assign ces_66_0_io_ins_0 = ces_65_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_66_0_io_ins_1 = io_insVertical_0_66; // @[MockArray.scala 45:87]
  assign ces_66_0_io_ins_2 = ces_67_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_66_0_io_ins_3 = io_insVertical_1_66; // @[MockArray.scala 47:87]
  assign ces_67_0_clock = clock;
  assign ces_67_0_io_ins_0 = ces_66_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_67_0_io_ins_1 = io_insVertical_0_67; // @[MockArray.scala 45:87]
  assign ces_67_0_io_ins_2 = ces_68_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_67_0_io_ins_3 = io_insVertical_1_67; // @[MockArray.scala 47:87]
  assign ces_68_0_clock = clock;
  assign ces_68_0_io_ins_0 = ces_67_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_68_0_io_ins_1 = io_insVertical_0_68; // @[MockArray.scala 45:87]
  assign ces_68_0_io_ins_2 = ces_69_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_68_0_io_ins_3 = io_insVertical_1_68; // @[MockArray.scala 47:87]
  assign ces_69_0_clock = clock;
  assign ces_69_0_io_ins_0 = ces_68_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_69_0_io_ins_1 = io_insVertical_0_69; // @[MockArray.scala 45:87]
  assign ces_69_0_io_ins_2 = ces_70_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_69_0_io_ins_3 = io_insVertical_1_69; // @[MockArray.scala 47:87]
  assign ces_70_0_clock = clock;
  assign ces_70_0_io_ins_0 = ces_69_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_70_0_io_ins_1 = io_insVertical_0_70; // @[MockArray.scala 45:87]
  assign ces_70_0_io_ins_2 = ces_71_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_70_0_io_ins_3 = io_insVertical_1_70; // @[MockArray.scala 47:87]
  assign ces_71_0_clock = clock;
  assign ces_71_0_io_ins_0 = ces_70_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_71_0_io_ins_1 = io_insVertical_0_71; // @[MockArray.scala 45:87]
  assign ces_71_0_io_ins_2 = ces_72_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_71_0_io_ins_3 = io_insVertical_1_71; // @[MockArray.scala 47:87]
  assign ces_72_0_clock = clock;
  assign ces_72_0_io_ins_0 = ces_71_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_72_0_io_ins_1 = io_insVertical_0_72; // @[MockArray.scala 45:87]
  assign ces_72_0_io_ins_2 = ces_73_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_72_0_io_ins_3 = io_insVertical_1_72; // @[MockArray.scala 47:87]
  assign ces_73_0_clock = clock;
  assign ces_73_0_io_ins_0 = ces_72_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_73_0_io_ins_1 = io_insVertical_0_73; // @[MockArray.scala 45:87]
  assign ces_73_0_io_ins_2 = ces_74_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_73_0_io_ins_3 = io_insVertical_1_73; // @[MockArray.scala 47:87]
  assign ces_74_0_clock = clock;
  assign ces_74_0_io_ins_0 = ces_73_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_74_0_io_ins_1 = io_insVertical_0_74; // @[MockArray.scala 45:87]
  assign ces_74_0_io_ins_2 = ces_75_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_74_0_io_ins_3 = io_insVertical_1_74; // @[MockArray.scala 47:87]
  assign ces_75_0_clock = clock;
  assign ces_75_0_io_ins_0 = ces_74_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_75_0_io_ins_1 = io_insVertical_0_75; // @[MockArray.scala 45:87]
  assign ces_75_0_io_ins_2 = ces_76_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_75_0_io_ins_3 = io_insVertical_1_75; // @[MockArray.scala 47:87]
  assign ces_76_0_clock = clock;
  assign ces_76_0_io_ins_0 = ces_75_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_76_0_io_ins_1 = io_insVertical_0_76; // @[MockArray.scala 45:87]
  assign ces_76_0_io_ins_2 = ces_77_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_76_0_io_ins_3 = io_insVertical_1_76; // @[MockArray.scala 47:87]
  assign ces_77_0_clock = clock;
  assign ces_77_0_io_ins_0 = ces_76_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_77_0_io_ins_1 = io_insVertical_0_77; // @[MockArray.scala 45:87]
  assign ces_77_0_io_ins_2 = ces_78_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_77_0_io_ins_3 = io_insVertical_1_77; // @[MockArray.scala 47:87]
  assign ces_78_0_clock = clock;
  assign ces_78_0_io_ins_0 = ces_77_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_78_0_io_ins_1 = io_insVertical_0_78; // @[MockArray.scala 45:87]
  assign ces_78_0_io_ins_2 = ces_79_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_78_0_io_ins_3 = io_insVertical_1_78; // @[MockArray.scala 47:87]
  assign ces_79_0_clock = clock;
  assign ces_79_0_io_ins_0 = ces_78_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_79_0_io_ins_1 = io_insVertical_0_79; // @[MockArray.scala 45:87]
  assign ces_79_0_io_ins_2 = ces_80_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_79_0_io_ins_3 = io_insVertical_1_79; // @[MockArray.scala 47:87]
  assign ces_80_0_clock = clock;
  assign ces_80_0_io_ins_0 = ces_79_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_80_0_io_ins_1 = io_insVertical_0_80; // @[MockArray.scala 45:87]
  assign ces_80_0_io_ins_2 = ces_81_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_80_0_io_ins_3 = io_insVertical_1_80; // @[MockArray.scala 47:87]
  assign ces_81_0_clock = clock;
  assign ces_81_0_io_ins_0 = ces_80_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_81_0_io_ins_1 = io_insVertical_0_81; // @[MockArray.scala 45:87]
  assign ces_81_0_io_ins_2 = ces_82_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_81_0_io_ins_3 = io_insVertical_1_81; // @[MockArray.scala 47:87]
  assign ces_82_0_clock = clock;
  assign ces_82_0_io_ins_0 = ces_81_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_82_0_io_ins_1 = io_insVertical_0_82; // @[MockArray.scala 45:87]
  assign ces_82_0_io_ins_2 = ces_83_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_82_0_io_ins_3 = io_insVertical_1_82; // @[MockArray.scala 47:87]
  assign ces_83_0_clock = clock;
  assign ces_83_0_io_ins_0 = ces_82_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_83_0_io_ins_1 = io_insVertical_0_83; // @[MockArray.scala 45:87]
  assign ces_83_0_io_ins_2 = ces_84_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_83_0_io_ins_3 = io_insVertical_1_83; // @[MockArray.scala 47:87]
  assign ces_84_0_clock = clock;
  assign ces_84_0_io_ins_0 = ces_83_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_84_0_io_ins_1 = io_insVertical_0_84; // @[MockArray.scala 45:87]
  assign ces_84_0_io_ins_2 = ces_85_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_84_0_io_ins_3 = io_insVertical_1_84; // @[MockArray.scala 47:87]
  assign ces_85_0_clock = clock;
  assign ces_85_0_io_ins_0 = ces_84_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_85_0_io_ins_1 = io_insVertical_0_85; // @[MockArray.scala 45:87]
  assign ces_85_0_io_ins_2 = ces_86_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_85_0_io_ins_3 = io_insVertical_1_85; // @[MockArray.scala 47:87]
  assign ces_86_0_clock = clock;
  assign ces_86_0_io_ins_0 = ces_85_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_86_0_io_ins_1 = io_insVertical_0_86; // @[MockArray.scala 45:87]
  assign ces_86_0_io_ins_2 = ces_87_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_86_0_io_ins_3 = io_insVertical_1_86; // @[MockArray.scala 47:87]
  assign ces_87_0_clock = clock;
  assign ces_87_0_io_ins_0 = ces_86_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_87_0_io_ins_1 = io_insVertical_0_87; // @[MockArray.scala 45:87]
  assign ces_87_0_io_ins_2 = ces_88_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_87_0_io_ins_3 = io_insVertical_1_87; // @[MockArray.scala 47:87]
  assign ces_88_0_clock = clock;
  assign ces_88_0_io_ins_0 = ces_87_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_88_0_io_ins_1 = io_insVertical_0_88; // @[MockArray.scala 45:87]
  assign ces_88_0_io_ins_2 = ces_89_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_88_0_io_ins_3 = io_insVertical_1_88; // @[MockArray.scala 47:87]
  assign ces_89_0_clock = clock;
  assign ces_89_0_io_ins_0 = ces_88_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_89_0_io_ins_1 = io_insVertical_0_89; // @[MockArray.scala 45:87]
  assign ces_89_0_io_ins_2 = ces_90_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_89_0_io_ins_3 = io_insVertical_1_89; // @[MockArray.scala 47:87]
  assign ces_90_0_clock = clock;
  assign ces_90_0_io_ins_0 = ces_89_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_90_0_io_ins_1 = io_insVertical_0_90; // @[MockArray.scala 45:87]
  assign ces_90_0_io_ins_2 = ces_91_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_90_0_io_ins_3 = io_insVertical_1_90; // @[MockArray.scala 47:87]
  assign ces_91_0_clock = clock;
  assign ces_91_0_io_ins_0 = ces_90_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_91_0_io_ins_1 = io_insVertical_0_91; // @[MockArray.scala 45:87]
  assign ces_91_0_io_ins_2 = ces_92_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_91_0_io_ins_3 = io_insVertical_1_91; // @[MockArray.scala 47:87]
  assign ces_92_0_clock = clock;
  assign ces_92_0_io_ins_0 = ces_91_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_92_0_io_ins_1 = io_insVertical_0_92; // @[MockArray.scala 45:87]
  assign ces_92_0_io_ins_2 = ces_93_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_92_0_io_ins_3 = io_insVertical_1_92; // @[MockArray.scala 47:87]
  assign ces_93_0_clock = clock;
  assign ces_93_0_io_ins_0 = ces_92_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_93_0_io_ins_1 = io_insVertical_0_93; // @[MockArray.scala 45:87]
  assign ces_93_0_io_ins_2 = ces_94_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_93_0_io_ins_3 = io_insVertical_1_93; // @[MockArray.scala 47:87]
  assign ces_94_0_clock = clock;
  assign ces_94_0_io_ins_0 = ces_93_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_94_0_io_ins_1 = io_insVertical_0_94; // @[MockArray.scala 45:87]
  assign ces_94_0_io_ins_2 = ces_95_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_94_0_io_ins_3 = io_insVertical_1_94; // @[MockArray.scala 47:87]
  assign ces_95_0_clock = clock;
  assign ces_95_0_io_ins_0 = ces_94_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_95_0_io_ins_1 = io_insVertical_0_95; // @[MockArray.scala 45:87]
  assign ces_95_0_io_ins_2 = ces_96_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_95_0_io_ins_3 = io_insVertical_1_95; // @[MockArray.scala 47:87]
  assign ces_96_0_clock = clock;
  assign ces_96_0_io_ins_0 = ces_95_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_96_0_io_ins_1 = io_insVertical_0_96; // @[MockArray.scala 45:87]
  assign ces_96_0_io_ins_2 = ces_97_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_96_0_io_ins_3 = io_insVertical_1_96; // @[MockArray.scala 47:87]
  assign ces_97_0_clock = clock;
  assign ces_97_0_io_ins_0 = ces_96_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_97_0_io_ins_1 = io_insVertical_0_97; // @[MockArray.scala 45:87]
  assign ces_97_0_io_ins_2 = ces_98_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_97_0_io_ins_3 = io_insVertical_1_97; // @[MockArray.scala 47:87]
  assign ces_98_0_clock = clock;
  assign ces_98_0_io_ins_0 = ces_97_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_98_0_io_ins_1 = io_insVertical_0_98; // @[MockArray.scala 45:87]
  assign ces_98_0_io_ins_2 = ces_99_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_98_0_io_ins_3 = io_insVertical_1_98; // @[MockArray.scala 47:87]
  assign ces_99_0_clock = clock;
  assign ces_99_0_io_ins_0 = ces_98_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_99_0_io_ins_1 = io_insVertical_0_99; // @[MockArray.scala 45:87]
  assign ces_99_0_io_ins_2 = ces_100_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_99_0_io_ins_3 = io_insVertical_1_99; // @[MockArray.scala 47:87]
  assign ces_100_0_clock = clock;
  assign ces_100_0_io_ins_0 = ces_99_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_100_0_io_ins_1 = io_insVertical_0_100; // @[MockArray.scala 45:87]
  assign ces_100_0_io_ins_2 = ces_101_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_100_0_io_ins_3 = io_insVertical_1_100; // @[MockArray.scala 47:87]
  assign ces_101_0_clock = clock;
  assign ces_101_0_io_ins_0 = ces_100_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_101_0_io_ins_1 = io_insVertical_0_101; // @[MockArray.scala 45:87]
  assign ces_101_0_io_ins_2 = ces_102_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_101_0_io_ins_3 = io_insVertical_1_101; // @[MockArray.scala 47:87]
  assign ces_102_0_clock = clock;
  assign ces_102_0_io_ins_0 = ces_101_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_102_0_io_ins_1 = io_insVertical_0_102; // @[MockArray.scala 45:87]
  assign ces_102_0_io_ins_2 = ces_103_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_102_0_io_ins_3 = io_insVertical_1_102; // @[MockArray.scala 47:87]
  assign ces_103_0_clock = clock;
  assign ces_103_0_io_ins_0 = ces_102_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_103_0_io_ins_1 = io_insVertical_0_103; // @[MockArray.scala 45:87]
  assign ces_103_0_io_ins_2 = ces_104_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_103_0_io_ins_3 = io_insVertical_1_103; // @[MockArray.scala 47:87]
  assign ces_104_0_clock = clock;
  assign ces_104_0_io_ins_0 = ces_103_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_104_0_io_ins_1 = io_insVertical_0_104; // @[MockArray.scala 45:87]
  assign ces_104_0_io_ins_2 = ces_105_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_104_0_io_ins_3 = io_insVertical_1_104; // @[MockArray.scala 47:87]
  assign ces_105_0_clock = clock;
  assign ces_105_0_io_ins_0 = ces_104_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_105_0_io_ins_1 = io_insVertical_0_105; // @[MockArray.scala 45:87]
  assign ces_105_0_io_ins_2 = ces_106_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_105_0_io_ins_3 = io_insVertical_1_105; // @[MockArray.scala 47:87]
  assign ces_106_0_clock = clock;
  assign ces_106_0_io_ins_0 = ces_105_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_106_0_io_ins_1 = io_insVertical_0_106; // @[MockArray.scala 45:87]
  assign ces_106_0_io_ins_2 = ces_107_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_106_0_io_ins_3 = io_insVertical_1_106; // @[MockArray.scala 47:87]
  assign ces_107_0_clock = clock;
  assign ces_107_0_io_ins_0 = ces_106_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_107_0_io_ins_1 = io_insVertical_0_107; // @[MockArray.scala 45:87]
  assign ces_107_0_io_ins_2 = ces_108_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_107_0_io_ins_3 = io_insVertical_1_107; // @[MockArray.scala 47:87]
  assign ces_108_0_clock = clock;
  assign ces_108_0_io_ins_0 = ces_107_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_108_0_io_ins_1 = io_insVertical_0_108; // @[MockArray.scala 45:87]
  assign ces_108_0_io_ins_2 = ces_109_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_108_0_io_ins_3 = io_insVertical_1_108; // @[MockArray.scala 47:87]
  assign ces_109_0_clock = clock;
  assign ces_109_0_io_ins_0 = ces_108_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_109_0_io_ins_1 = io_insVertical_0_109; // @[MockArray.scala 45:87]
  assign ces_109_0_io_ins_2 = ces_110_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_109_0_io_ins_3 = io_insVertical_1_109; // @[MockArray.scala 47:87]
  assign ces_110_0_clock = clock;
  assign ces_110_0_io_ins_0 = ces_109_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_110_0_io_ins_1 = io_insVertical_0_110; // @[MockArray.scala 45:87]
  assign ces_110_0_io_ins_2 = ces_111_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_110_0_io_ins_3 = io_insVertical_1_110; // @[MockArray.scala 47:87]
  assign ces_111_0_clock = clock;
  assign ces_111_0_io_ins_0 = ces_110_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_111_0_io_ins_1 = io_insVertical_0_111; // @[MockArray.scala 45:87]
  assign ces_111_0_io_ins_2 = ces_112_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_111_0_io_ins_3 = io_insVertical_1_111; // @[MockArray.scala 47:87]
  assign ces_112_0_clock = clock;
  assign ces_112_0_io_ins_0 = ces_111_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_112_0_io_ins_1 = io_insVertical_0_112; // @[MockArray.scala 45:87]
  assign ces_112_0_io_ins_2 = ces_113_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_112_0_io_ins_3 = io_insVertical_1_112; // @[MockArray.scala 47:87]
  assign ces_113_0_clock = clock;
  assign ces_113_0_io_ins_0 = ces_112_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_113_0_io_ins_1 = io_insVertical_0_113; // @[MockArray.scala 45:87]
  assign ces_113_0_io_ins_2 = ces_114_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_113_0_io_ins_3 = io_insVertical_1_113; // @[MockArray.scala 47:87]
  assign ces_114_0_clock = clock;
  assign ces_114_0_io_ins_0 = ces_113_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_114_0_io_ins_1 = io_insVertical_0_114; // @[MockArray.scala 45:87]
  assign ces_114_0_io_ins_2 = ces_115_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_114_0_io_ins_3 = io_insVertical_1_114; // @[MockArray.scala 47:87]
  assign ces_115_0_clock = clock;
  assign ces_115_0_io_ins_0 = ces_114_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_115_0_io_ins_1 = io_insVertical_0_115; // @[MockArray.scala 45:87]
  assign ces_115_0_io_ins_2 = ces_116_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_115_0_io_ins_3 = io_insVertical_1_115; // @[MockArray.scala 47:87]
  assign ces_116_0_clock = clock;
  assign ces_116_0_io_ins_0 = ces_115_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_116_0_io_ins_1 = io_insVertical_0_116; // @[MockArray.scala 45:87]
  assign ces_116_0_io_ins_2 = ces_117_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_116_0_io_ins_3 = io_insVertical_1_116; // @[MockArray.scala 47:87]
  assign ces_117_0_clock = clock;
  assign ces_117_0_io_ins_0 = ces_116_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_117_0_io_ins_1 = io_insVertical_0_117; // @[MockArray.scala 45:87]
  assign ces_117_0_io_ins_2 = ces_118_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_117_0_io_ins_3 = io_insVertical_1_117; // @[MockArray.scala 47:87]
  assign ces_118_0_clock = clock;
  assign ces_118_0_io_ins_0 = ces_117_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_118_0_io_ins_1 = io_insVertical_0_118; // @[MockArray.scala 45:87]
  assign ces_118_0_io_ins_2 = ces_119_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_118_0_io_ins_3 = io_insVertical_1_118; // @[MockArray.scala 47:87]
  assign ces_119_0_clock = clock;
  assign ces_119_0_io_ins_0 = ces_118_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_119_0_io_ins_1 = io_insVertical_0_119; // @[MockArray.scala 45:87]
  assign ces_119_0_io_ins_2 = ces_120_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_119_0_io_ins_3 = io_insVertical_1_119; // @[MockArray.scala 47:87]
  assign ces_120_0_clock = clock;
  assign ces_120_0_io_ins_0 = ces_119_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_120_0_io_ins_1 = io_insVertical_0_120; // @[MockArray.scala 45:87]
  assign ces_120_0_io_ins_2 = ces_121_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_120_0_io_ins_3 = io_insVertical_1_120; // @[MockArray.scala 47:87]
  assign ces_121_0_clock = clock;
  assign ces_121_0_io_ins_0 = ces_120_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_121_0_io_ins_1 = io_insVertical_0_121; // @[MockArray.scala 45:87]
  assign ces_121_0_io_ins_2 = ces_122_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_121_0_io_ins_3 = io_insVertical_1_121; // @[MockArray.scala 47:87]
  assign ces_122_0_clock = clock;
  assign ces_122_0_io_ins_0 = ces_121_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_122_0_io_ins_1 = io_insVertical_0_122; // @[MockArray.scala 45:87]
  assign ces_122_0_io_ins_2 = ces_123_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_122_0_io_ins_3 = io_insVertical_1_122; // @[MockArray.scala 47:87]
  assign ces_123_0_clock = clock;
  assign ces_123_0_io_ins_0 = ces_122_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_123_0_io_ins_1 = io_insVertical_0_123; // @[MockArray.scala 45:87]
  assign ces_123_0_io_ins_2 = ces_124_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_123_0_io_ins_3 = io_insVertical_1_123; // @[MockArray.scala 47:87]
  assign ces_124_0_clock = clock;
  assign ces_124_0_io_ins_0 = ces_123_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_124_0_io_ins_1 = io_insVertical_0_124; // @[MockArray.scala 45:87]
  assign ces_124_0_io_ins_2 = ces_125_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_124_0_io_ins_3 = io_insVertical_1_124; // @[MockArray.scala 47:87]
  assign ces_125_0_clock = clock;
  assign ces_125_0_io_ins_0 = ces_124_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_125_0_io_ins_1 = io_insVertical_0_125; // @[MockArray.scala 45:87]
  assign ces_125_0_io_ins_2 = ces_126_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_125_0_io_ins_3 = io_insVertical_1_125; // @[MockArray.scala 47:87]
  assign ces_126_0_clock = clock;
  assign ces_126_0_io_ins_0 = ces_125_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_126_0_io_ins_1 = io_insVertical_0_126; // @[MockArray.scala 45:87]
  assign ces_126_0_io_ins_2 = ces_127_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_126_0_io_ins_3 = io_insVertical_1_126; // @[MockArray.scala 47:87]
  assign ces_127_0_clock = clock;
  assign ces_127_0_io_ins_0 = ces_126_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_127_0_io_ins_1 = io_insVertical_0_127; // @[MockArray.scala 45:87]
  assign ces_127_0_io_ins_2 = ces_128_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_127_0_io_ins_3 = io_insVertical_1_127; // @[MockArray.scala 47:87]
  assign ces_128_0_clock = clock;
  assign ces_128_0_io_ins_0 = ces_127_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_128_0_io_ins_1 = io_insVertical_0_128; // @[MockArray.scala 45:87]
  assign ces_128_0_io_ins_2 = ces_129_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_128_0_io_ins_3 = io_insVertical_1_128; // @[MockArray.scala 47:87]
  assign ces_129_0_clock = clock;
  assign ces_129_0_io_ins_0 = ces_128_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_129_0_io_ins_1 = io_insVertical_0_129; // @[MockArray.scala 45:87]
  assign ces_129_0_io_ins_2 = ces_130_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_129_0_io_ins_3 = io_insVertical_1_129; // @[MockArray.scala 47:87]
  assign ces_130_0_clock = clock;
  assign ces_130_0_io_ins_0 = ces_129_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_130_0_io_ins_1 = io_insVertical_0_130; // @[MockArray.scala 45:87]
  assign ces_130_0_io_ins_2 = ces_131_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_130_0_io_ins_3 = io_insVertical_1_130; // @[MockArray.scala 47:87]
  assign ces_131_0_clock = clock;
  assign ces_131_0_io_ins_0 = ces_130_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_131_0_io_ins_1 = io_insVertical_0_131; // @[MockArray.scala 45:87]
  assign ces_131_0_io_ins_2 = ces_132_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_131_0_io_ins_3 = io_insVertical_1_131; // @[MockArray.scala 47:87]
  assign ces_132_0_clock = clock;
  assign ces_132_0_io_ins_0 = ces_131_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_132_0_io_ins_1 = io_insVertical_0_132; // @[MockArray.scala 45:87]
  assign ces_132_0_io_ins_2 = ces_133_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_132_0_io_ins_3 = io_insVertical_1_132; // @[MockArray.scala 47:87]
  assign ces_133_0_clock = clock;
  assign ces_133_0_io_ins_0 = ces_132_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_133_0_io_ins_1 = io_insVertical_0_133; // @[MockArray.scala 45:87]
  assign ces_133_0_io_ins_2 = ces_134_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_133_0_io_ins_3 = io_insVertical_1_133; // @[MockArray.scala 47:87]
  assign ces_134_0_clock = clock;
  assign ces_134_0_io_ins_0 = ces_133_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_134_0_io_ins_1 = io_insVertical_0_134; // @[MockArray.scala 45:87]
  assign ces_134_0_io_ins_2 = ces_135_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_134_0_io_ins_3 = io_insVertical_1_134; // @[MockArray.scala 47:87]
  assign ces_135_0_clock = clock;
  assign ces_135_0_io_ins_0 = ces_134_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_135_0_io_ins_1 = io_insVertical_0_135; // @[MockArray.scala 45:87]
  assign ces_135_0_io_ins_2 = ces_136_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_135_0_io_ins_3 = io_insVertical_1_135; // @[MockArray.scala 47:87]
  assign ces_136_0_clock = clock;
  assign ces_136_0_io_ins_0 = ces_135_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_136_0_io_ins_1 = io_insVertical_0_136; // @[MockArray.scala 45:87]
  assign ces_136_0_io_ins_2 = ces_137_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_136_0_io_ins_3 = io_insVertical_1_136; // @[MockArray.scala 47:87]
  assign ces_137_0_clock = clock;
  assign ces_137_0_io_ins_0 = ces_136_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_137_0_io_ins_1 = io_insVertical_0_137; // @[MockArray.scala 45:87]
  assign ces_137_0_io_ins_2 = ces_138_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_137_0_io_ins_3 = io_insVertical_1_137; // @[MockArray.scala 47:87]
  assign ces_138_0_clock = clock;
  assign ces_138_0_io_ins_0 = ces_137_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_138_0_io_ins_1 = io_insVertical_0_138; // @[MockArray.scala 45:87]
  assign ces_138_0_io_ins_2 = ces_139_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_138_0_io_ins_3 = io_insVertical_1_138; // @[MockArray.scala 47:87]
  assign ces_139_0_clock = clock;
  assign ces_139_0_io_ins_0 = ces_138_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_139_0_io_ins_1 = io_insVertical_0_139; // @[MockArray.scala 45:87]
  assign ces_139_0_io_ins_2 = ces_140_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_139_0_io_ins_3 = io_insVertical_1_139; // @[MockArray.scala 47:87]
  assign ces_140_0_clock = clock;
  assign ces_140_0_io_ins_0 = ces_139_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_140_0_io_ins_1 = io_insVertical_0_140; // @[MockArray.scala 45:87]
  assign ces_140_0_io_ins_2 = ces_141_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_140_0_io_ins_3 = io_insVertical_1_140; // @[MockArray.scala 47:87]
  assign ces_141_0_clock = clock;
  assign ces_141_0_io_ins_0 = ces_140_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_141_0_io_ins_1 = io_insVertical_0_141; // @[MockArray.scala 45:87]
  assign ces_141_0_io_ins_2 = ces_142_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_141_0_io_ins_3 = io_insVertical_1_141; // @[MockArray.scala 47:87]
  assign ces_142_0_clock = clock;
  assign ces_142_0_io_ins_0 = ces_141_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_142_0_io_ins_1 = io_insVertical_0_142; // @[MockArray.scala 45:87]
  assign ces_142_0_io_ins_2 = ces_143_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_142_0_io_ins_3 = io_insVertical_1_142; // @[MockArray.scala 47:87]
  assign ces_143_0_clock = clock;
  assign ces_143_0_io_ins_0 = ces_142_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_143_0_io_ins_1 = io_insVertical_0_143; // @[MockArray.scala 45:87]
  assign ces_143_0_io_ins_2 = ces_144_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_143_0_io_ins_3 = io_insVertical_1_143; // @[MockArray.scala 47:87]
  assign ces_144_0_clock = clock;
  assign ces_144_0_io_ins_0 = ces_143_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_144_0_io_ins_1 = io_insVertical_0_144; // @[MockArray.scala 45:87]
  assign ces_144_0_io_ins_2 = ces_145_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_144_0_io_ins_3 = io_insVertical_1_144; // @[MockArray.scala 47:87]
  assign ces_145_0_clock = clock;
  assign ces_145_0_io_ins_0 = ces_144_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_145_0_io_ins_1 = io_insVertical_0_145; // @[MockArray.scala 45:87]
  assign ces_145_0_io_ins_2 = ces_146_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_145_0_io_ins_3 = io_insVertical_1_145; // @[MockArray.scala 47:87]
  assign ces_146_0_clock = clock;
  assign ces_146_0_io_ins_0 = ces_145_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_146_0_io_ins_1 = io_insVertical_0_146; // @[MockArray.scala 45:87]
  assign ces_146_0_io_ins_2 = ces_147_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_146_0_io_ins_3 = io_insVertical_1_146; // @[MockArray.scala 47:87]
  assign ces_147_0_clock = clock;
  assign ces_147_0_io_ins_0 = ces_146_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_147_0_io_ins_1 = io_insVertical_0_147; // @[MockArray.scala 45:87]
  assign ces_147_0_io_ins_2 = ces_148_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_147_0_io_ins_3 = io_insVertical_1_147; // @[MockArray.scala 47:87]
  assign ces_148_0_clock = clock;
  assign ces_148_0_io_ins_0 = ces_147_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_148_0_io_ins_1 = io_insVertical_0_148; // @[MockArray.scala 45:87]
  assign ces_148_0_io_ins_2 = ces_149_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_148_0_io_ins_3 = io_insVertical_1_148; // @[MockArray.scala 47:87]
  assign ces_149_0_clock = clock;
  assign ces_149_0_io_ins_0 = ces_148_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_149_0_io_ins_1 = io_insVertical_0_149; // @[MockArray.scala 45:87]
  assign ces_149_0_io_ins_2 = ces_150_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_149_0_io_ins_3 = io_insVertical_1_149; // @[MockArray.scala 47:87]
  assign ces_150_0_clock = clock;
  assign ces_150_0_io_ins_0 = ces_149_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_150_0_io_ins_1 = io_insVertical_0_150; // @[MockArray.scala 45:87]
  assign ces_150_0_io_ins_2 = ces_151_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_150_0_io_ins_3 = io_insVertical_1_150; // @[MockArray.scala 47:87]
  assign ces_151_0_clock = clock;
  assign ces_151_0_io_ins_0 = ces_150_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_151_0_io_ins_1 = io_insVertical_0_151; // @[MockArray.scala 45:87]
  assign ces_151_0_io_ins_2 = ces_152_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_151_0_io_ins_3 = io_insVertical_1_151; // @[MockArray.scala 47:87]
  assign ces_152_0_clock = clock;
  assign ces_152_0_io_ins_0 = ces_151_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_152_0_io_ins_1 = io_insVertical_0_152; // @[MockArray.scala 45:87]
  assign ces_152_0_io_ins_2 = ces_153_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_152_0_io_ins_3 = io_insVertical_1_152; // @[MockArray.scala 47:87]
  assign ces_153_0_clock = clock;
  assign ces_153_0_io_ins_0 = ces_152_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_153_0_io_ins_1 = io_insVertical_0_153; // @[MockArray.scala 45:87]
  assign ces_153_0_io_ins_2 = ces_154_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_153_0_io_ins_3 = io_insVertical_1_153; // @[MockArray.scala 47:87]
  assign ces_154_0_clock = clock;
  assign ces_154_0_io_ins_0 = ces_153_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_154_0_io_ins_1 = io_insVertical_0_154; // @[MockArray.scala 45:87]
  assign ces_154_0_io_ins_2 = ces_155_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_154_0_io_ins_3 = io_insVertical_1_154; // @[MockArray.scala 47:87]
  assign ces_155_0_clock = clock;
  assign ces_155_0_io_ins_0 = ces_154_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_155_0_io_ins_1 = io_insVertical_0_155; // @[MockArray.scala 45:87]
  assign ces_155_0_io_ins_2 = ces_156_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_155_0_io_ins_3 = io_insVertical_1_155; // @[MockArray.scala 47:87]
  assign ces_156_0_clock = clock;
  assign ces_156_0_io_ins_0 = ces_155_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_156_0_io_ins_1 = io_insVertical_0_156; // @[MockArray.scala 45:87]
  assign ces_156_0_io_ins_2 = ces_157_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_156_0_io_ins_3 = io_insVertical_1_156; // @[MockArray.scala 47:87]
  assign ces_157_0_clock = clock;
  assign ces_157_0_io_ins_0 = ces_156_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_157_0_io_ins_1 = io_insVertical_0_157; // @[MockArray.scala 45:87]
  assign ces_157_0_io_ins_2 = ces_158_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_157_0_io_ins_3 = io_insVertical_1_157; // @[MockArray.scala 47:87]
  assign ces_158_0_clock = clock;
  assign ces_158_0_io_ins_0 = ces_157_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_158_0_io_ins_1 = io_insVertical_0_158; // @[MockArray.scala 45:87]
  assign ces_158_0_io_ins_2 = ces_159_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_158_0_io_ins_3 = io_insVertical_1_158; // @[MockArray.scala 47:87]
  assign ces_159_0_clock = clock;
  assign ces_159_0_io_ins_0 = ces_158_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_159_0_io_ins_1 = io_insVertical_0_159; // @[MockArray.scala 45:87]
  assign ces_159_0_io_ins_2 = ces_160_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_159_0_io_ins_3 = io_insVertical_1_159; // @[MockArray.scala 47:87]
  assign ces_160_0_clock = clock;
  assign ces_160_0_io_ins_0 = ces_159_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_160_0_io_ins_1 = io_insVertical_0_160; // @[MockArray.scala 45:87]
  assign ces_160_0_io_ins_2 = ces_161_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_160_0_io_ins_3 = io_insVertical_1_160; // @[MockArray.scala 47:87]
  assign ces_161_0_clock = clock;
  assign ces_161_0_io_ins_0 = ces_160_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_161_0_io_ins_1 = io_insVertical_0_161; // @[MockArray.scala 45:87]
  assign ces_161_0_io_ins_2 = ces_162_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_161_0_io_ins_3 = io_insVertical_1_161; // @[MockArray.scala 47:87]
  assign ces_162_0_clock = clock;
  assign ces_162_0_io_ins_0 = ces_161_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_162_0_io_ins_1 = io_insVertical_0_162; // @[MockArray.scala 45:87]
  assign ces_162_0_io_ins_2 = ces_163_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_162_0_io_ins_3 = io_insVertical_1_162; // @[MockArray.scala 47:87]
  assign ces_163_0_clock = clock;
  assign ces_163_0_io_ins_0 = ces_162_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_163_0_io_ins_1 = io_insVertical_0_163; // @[MockArray.scala 45:87]
  assign ces_163_0_io_ins_2 = ces_164_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_163_0_io_ins_3 = io_insVertical_1_163; // @[MockArray.scala 47:87]
  assign ces_164_0_clock = clock;
  assign ces_164_0_io_ins_0 = ces_163_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_164_0_io_ins_1 = io_insVertical_0_164; // @[MockArray.scala 45:87]
  assign ces_164_0_io_ins_2 = ces_165_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_164_0_io_ins_3 = io_insVertical_1_164; // @[MockArray.scala 47:87]
  assign ces_165_0_clock = clock;
  assign ces_165_0_io_ins_0 = ces_164_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_165_0_io_ins_1 = io_insVertical_0_165; // @[MockArray.scala 45:87]
  assign ces_165_0_io_ins_2 = ces_166_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_165_0_io_ins_3 = io_insVertical_1_165; // @[MockArray.scala 47:87]
  assign ces_166_0_clock = clock;
  assign ces_166_0_io_ins_0 = ces_165_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_166_0_io_ins_1 = io_insVertical_0_166; // @[MockArray.scala 45:87]
  assign ces_166_0_io_ins_2 = ces_167_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_166_0_io_ins_3 = io_insVertical_1_166; // @[MockArray.scala 47:87]
  assign ces_167_0_clock = clock;
  assign ces_167_0_io_ins_0 = ces_166_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_167_0_io_ins_1 = io_insVertical_0_167; // @[MockArray.scala 45:87]
  assign ces_167_0_io_ins_2 = ces_168_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_167_0_io_ins_3 = io_insVertical_1_167; // @[MockArray.scala 47:87]
  assign ces_168_0_clock = clock;
  assign ces_168_0_io_ins_0 = ces_167_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_168_0_io_ins_1 = io_insVertical_0_168; // @[MockArray.scala 45:87]
  assign ces_168_0_io_ins_2 = ces_169_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_168_0_io_ins_3 = io_insVertical_1_168; // @[MockArray.scala 47:87]
  assign ces_169_0_clock = clock;
  assign ces_169_0_io_ins_0 = ces_168_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_169_0_io_ins_1 = io_insVertical_0_169; // @[MockArray.scala 45:87]
  assign ces_169_0_io_ins_2 = ces_170_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_169_0_io_ins_3 = io_insVertical_1_169; // @[MockArray.scala 47:87]
  assign ces_170_0_clock = clock;
  assign ces_170_0_io_ins_0 = ces_169_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_170_0_io_ins_1 = io_insVertical_0_170; // @[MockArray.scala 45:87]
  assign ces_170_0_io_ins_2 = ces_171_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_170_0_io_ins_3 = io_insVertical_1_170; // @[MockArray.scala 47:87]
  assign ces_171_0_clock = clock;
  assign ces_171_0_io_ins_0 = ces_170_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_171_0_io_ins_1 = io_insVertical_0_171; // @[MockArray.scala 45:87]
  assign ces_171_0_io_ins_2 = ces_172_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_171_0_io_ins_3 = io_insVertical_1_171; // @[MockArray.scala 47:87]
  assign ces_172_0_clock = clock;
  assign ces_172_0_io_ins_0 = ces_171_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_172_0_io_ins_1 = io_insVertical_0_172; // @[MockArray.scala 45:87]
  assign ces_172_0_io_ins_2 = ces_173_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_172_0_io_ins_3 = io_insVertical_1_172; // @[MockArray.scala 47:87]
  assign ces_173_0_clock = clock;
  assign ces_173_0_io_ins_0 = ces_172_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_173_0_io_ins_1 = io_insVertical_0_173; // @[MockArray.scala 45:87]
  assign ces_173_0_io_ins_2 = ces_174_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_173_0_io_ins_3 = io_insVertical_1_173; // @[MockArray.scala 47:87]
  assign ces_174_0_clock = clock;
  assign ces_174_0_io_ins_0 = ces_173_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_174_0_io_ins_1 = io_insVertical_0_174; // @[MockArray.scala 45:87]
  assign ces_174_0_io_ins_2 = ces_175_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_174_0_io_ins_3 = io_insVertical_1_174; // @[MockArray.scala 47:87]
  assign ces_175_0_clock = clock;
  assign ces_175_0_io_ins_0 = ces_174_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_175_0_io_ins_1 = io_insVertical_0_175; // @[MockArray.scala 45:87]
  assign ces_175_0_io_ins_2 = ces_176_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_175_0_io_ins_3 = io_insVertical_1_175; // @[MockArray.scala 47:87]
  assign ces_176_0_clock = clock;
  assign ces_176_0_io_ins_0 = ces_175_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_176_0_io_ins_1 = io_insVertical_0_176; // @[MockArray.scala 45:87]
  assign ces_176_0_io_ins_2 = ces_177_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_176_0_io_ins_3 = io_insVertical_1_176; // @[MockArray.scala 47:87]
  assign ces_177_0_clock = clock;
  assign ces_177_0_io_ins_0 = ces_176_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_177_0_io_ins_1 = io_insVertical_0_177; // @[MockArray.scala 45:87]
  assign ces_177_0_io_ins_2 = ces_178_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_177_0_io_ins_3 = io_insVertical_1_177; // @[MockArray.scala 47:87]
  assign ces_178_0_clock = clock;
  assign ces_178_0_io_ins_0 = ces_177_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_178_0_io_ins_1 = io_insVertical_0_178; // @[MockArray.scala 45:87]
  assign ces_178_0_io_ins_2 = ces_179_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_178_0_io_ins_3 = io_insVertical_1_178; // @[MockArray.scala 47:87]
  assign ces_179_0_clock = clock;
  assign ces_179_0_io_ins_0 = ces_178_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_179_0_io_ins_1 = io_insVertical_0_179; // @[MockArray.scala 45:87]
  assign ces_179_0_io_ins_2 = ces_180_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_179_0_io_ins_3 = io_insVertical_1_179; // @[MockArray.scala 47:87]
  assign ces_180_0_clock = clock;
  assign ces_180_0_io_ins_0 = ces_179_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_180_0_io_ins_1 = io_insVertical_0_180; // @[MockArray.scala 45:87]
  assign ces_180_0_io_ins_2 = ces_181_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_180_0_io_ins_3 = io_insVertical_1_180; // @[MockArray.scala 47:87]
  assign ces_181_0_clock = clock;
  assign ces_181_0_io_ins_0 = ces_180_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_181_0_io_ins_1 = io_insVertical_0_181; // @[MockArray.scala 45:87]
  assign ces_181_0_io_ins_2 = ces_182_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_181_0_io_ins_3 = io_insVertical_1_181; // @[MockArray.scala 47:87]
  assign ces_182_0_clock = clock;
  assign ces_182_0_io_ins_0 = ces_181_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_182_0_io_ins_1 = io_insVertical_0_182; // @[MockArray.scala 45:87]
  assign ces_182_0_io_ins_2 = ces_183_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_182_0_io_ins_3 = io_insVertical_1_182; // @[MockArray.scala 47:87]
  assign ces_183_0_clock = clock;
  assign ces_183_0_io_ins_0 = ces_182_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_183_0_io_ins_1 = io_insVertical_0_183; // @[MockArray.scala 45:87]
  assign ces_183_0_io_ins_2 = ces_184_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_183_0_io_ins_3 = io_insVertical_1_183; // @[MockArray.scala 47:87]
  assign ces_184_0_clock = clock;
  assign ces_184_0_io_ins_0 = ces_183_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_184_0_io_ins_1 = io_insVertical_0_184; // @[MockArray.scala 45:87]
  assign ces_184_0_io_ins_2 = ces_185_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_184_0_io_ins_3 = io_insVertical_1_184; // @[MockArray.scala 47:87]
  assign ces_185_0_clock = clock;
  assign ces_185_0_io_ins_0 = ces_184_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_185_0_io_ins_1 = io_insVertical_0_185; // @[MockArray.scala 45:87]
  assign ces_185_0_io_ins_2 = ces_186_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_185_0_io_ins_3 = io_insVertical_1_185; // @[MockArray.scala 47:87]
  assign ces_186_0_clock = clock;
  assign ces_186_0_io_ins_0 = ces_185_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_186_0_io_ins_1 = io_insVertical_0_186; // @[MockArray.scala 45:87]
  assign ces_186_0_io_ins_2 = ces_187_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_186_0_io_ins_3 = io_insVertical_1_186; // @[MockArray.scala 47:87]
  assign ces_187_0_clock = clock;
  assign ces_187_0_io_ins_0 = ces_186_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_187_0_io_ins_1 = io_insVertical_0_187; // @[MockArray.scala 45:87]
  assign ces_187_0_io_ins_2 = ces_188_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_187_0_io_ins_3 = io_insVertical_1_187; // @[MockArray.scala 47:87]
  assign ces_188_0_clock = clock;
  assign ces_188_0_io_ins_0 = ces_187_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_188_0_io_ins_1 = io_insVertical_0_188; // @[MockArray.scala 45:87]
  assign ces_188_0_io_ins_2 = ces_189_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_188_0_io_ins_3 = io_insVertical_1_188; // @[MockArray.scala 47:87]
  assign ces_189_0_clock = clock;
  assign ces_189_0_io_ins_0 = ces_188_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_189_0_io_ins_1 = io_insVertical_0_189; // @[MockArray.scala 45:87]
  assign ces_189_0_io_ins_2 = ces_190_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_189_0_io_ins_3 = io_insVertical_1_189; // @[MockArray.scala 47:87]
  assign ces_190_0_clock = clock;
  assign ces_190_0_io_ins_0 = ces_189_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_190_0_io_ins_1 = io_insVertical_0_190; // @[MockArray.scala 45:87]
  assign ces_190_0_io_ins_2 = ces_191_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_190_0_io_ins_3 = io_insVertical_1_190; // @[MockArray.scala 47:87]
  assign ces_191_0_clock = clock;
  assign ces_191_0_io_ins_0 = ces_190_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_191_0_io_ins_1 = io_insVertical_0_191; // @[MockArray.scala 45:87]
  assign ces_191_0_io_ins_2 = ces_192_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_191_0_io_ins_3 = io_insVertical_1_191; // @[MockArray.scala 47:87]
  assign ces_192_0_clock = clock;
  assign ces_192_0_io_ins_0 = ces_191_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_192_0_io_ins_1 = io_insVertical_0_192; // @[MockArray.scala 45:87]
  assign ces_192_0_io_ins_2 = ces_193_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_192_0_io_ins_3 = io_insVertical_1_192; // @[MockArray.scala 47:87]
  assign ces_193_0_clock = clock;
  assign ces_193_0_io_ins_0 = ces_192_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_193_0_io_ins_1 = io_insVertical_0_193; // @[MockArray.scala 45:87]
  assign ces_193_0_io_ins_2 = ces_194_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_193_0_io_ins_3 = io_insVertical_1_193; // @[MockArray.scala 47:87]
  assign ces_194_0_clock = clock;
  assign ces_194_0_io_ins_0 = ces_193_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_194_0_io_ins_1 = io_insVertical_0_194; // @[MockArray.scala 45:87]
  assign ces_194_0_io_ins_2 = ces_195_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_194_0_io_ins_3 = io_insVertical_1_194; // @[MockArray.scala 47:87]
  assign ces_195_0_clock = clock;
  assign ces_195_0_io_ins_0 = ces_194_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_195_0_io_ins_1 = io_insVertical_0_195; // @[MockArray.scala 45:87]
  assign ces_195_0_io_ins_2 = ces_196_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_195_0_io_ins_3 = io_insVertical_1_195; // @[MockArray.scala 47:87]
  assign ces_196_0_clock = clock;
  assign ces_196_0_io_ins_0 = ces_195_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_196_0_io_ins_1 = io_insVertical_0_196; // @[MockArray.scala 45:87]
  assign ces_196_0_io_ins_2 = ces_197_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_196_0_io_ins_3 = io_insVertical_1_196; // @[MockArray.scala 47:87]
  assign ces_197_0_clock = clock;
  assign ces_197_0_io_ins_0 = ces_196_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_197_0_io_ins_1 = io_insVertical_0_197; // @[MockArray.scala 45:87]
  assign ces_197_0_io_ins_2 = ces_198_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_197_0_io_ins_3 = io_insVertical_1_197; // @[MockArray.scala 47:87]
  assign ces_198_0_clock = clock;
  assign ces_198_0_io_ins_0 = ces_197_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_198_0_io_ins_1 = io_insVertical_0_198; // @[MockArray.scala 45:87]
  assign ces_198_0_io_ins_2 = ces_199_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_198_0_io_ins_3 = io_insVertical_1_198; // @[MockArray.scala 47:87]
  assign ces_199_0_clock = clock;
  assign ces_199_0_io_ins_0 = ces_198_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_199_0_io_ins_1 = io_insVertical_0_199; // @[MockArray.scala 45:87]
  assign ces_199_0_io_ins_2 = ces_200_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_199_0_io_ins_3 = io_insVertical_1_199; // @[MockArray.scala 47:87]
  assign ces_200_0_clock = clock;
  assign ces_200_0_io_ins_0 = ces_199_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_200_0_io_ins_1 = io_insVertical_0_200; // @[MockArray.scala 45:87]
  assign ces_200_0_io_ins_2 = ces_201_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_200_0_io_ins_3 = io_insVertical_1_200; // @[MockArray.scala 47:87]
  assign ces_201_0_clock = clock;
  assign ces_201_0_io_ins_0 = ces_200_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_201_0_io_ins_1 = io_insVertical_0_201; // @[MockArray.scala 45:87]
  assign ces_201_0_io_ins_2 = ces_202_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_201_0_io_ins_3 = io_insVertical_1_201; // @[MockArray.scala 47:87]
  assign ces_202_0_clock = clock;
  assign ces_202_0_io_ins_0 = ces_201_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_202_0_io_ins_1 = io_insVertical_0_202; // @[MockArray.scala 45:87]
  assign ces_202_0_io_ins_2 = ces_203_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_202_0_io_ins_3 = io_insVertical_1_202; // @[MockArray.scala 47:87]
  assign ces_203_0_clock = clock;
  assign ces_203_0_io_ins_0 = ces_202_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_203_0_io_ins_1 = io_insVertical_0_203; // @[MockArray.scala 45:87]
  assign ces_203_0_io_ins_2 = ces_204_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_203_0_io_ins_3 = io_insVertical_1_203; // @[MockArray.scala 47:87]
  assign ces_204_0_clock = clock;
  assign ces_204_0_io_ins_0 = ces_203_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_204_0_io_ins_1 = io_insVertical_0_204; // @[MockArray.scala 45:87]
  assign ces_204_0_io_ins_2 = ces_205_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_204_0_io_ins_3 = io_insVertical_1_204; // @[MockArray.scala 47:87]
  assign ces_205_0_clock = clock;
  assign ces_205_0_io_ins_0 = ces_204_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_205_0_io_ins_1 = io_insVertical_0_205; // @[MockArray.scala 45:87]
  assign ces_205_0_io_ins_2 = ces_206_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_205_0_io_ins_3 = io_insVertical_1_205; // @[MockArray.scala 47:87]
  assign ces_206_0_clock = clock;
  assign ces_206_0_io_ins_0 = ces_205_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_206_0_io_ins_1 = io_insVertical_0_206; // @[MockArray.scala 45:87]
  assign ces_206_0_io_ins_2 = ces_207_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_206_0_io_ins_3 = io_insVertical_1_206; // @[MockArray.scala 47:87]
  assign ces_207_0_clock = clock;
  assign ces_207_0_io_ins_0 = ces_206_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_207_0_io_ins_1 = io_insVertical_0_207; // @[MockArray.scala 45:87]
  assign ces_207_0_io_ins_2 = ces_208_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_207_0_io_ins_3 = io_insVertical_1_207; // @[MockArray.scala 47:87]
  assign ces_208_0_clock = clock;
  assign ces_208_0_io_ins_0 = ces_207_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_208_0_io_ins_1 = io_insVertical_0_208; // @[MockArray.scala 45:87]
  assign ces_208_0_io_ins_2 = ces_209_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_208_0_io_ins_3 = io_insVertical_1_208; // @[MockArray.scala 47:87]
  assign ces_209_0_clock = clock;
  assign ces_209_0_io_ins_0 = ces_208_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_209_0_io_ins_1 = io_insVertical_0_209; // @[MockArray.scala 45:87]
  assign ces_209_0_io_ins_2 = ces_210_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_209_0_io_ins_3 = io_insVertical_1_209; // @[MockArray.scala 47:87]
  assign ces_210_0_clock = clock;
  assign ces_210_0_io_ins_0 = ces_209_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_210_0_io_ins_1 = io_insVertical_0_210; // @[MockArray.scala 45:87]
  assign ces_210_0_io_ins_2 = ces_211_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_210_0_io_ins_3 = io_insVertical_1_210; // @[MockArray.scala 47:87]
  assign ces_211_0_clock = clock;
  assign ces_211_0_io_ins_0 = ces_210_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_211_0_io_ins_1 = io_insVertical_0_211; // @[MockArray.scala 45:87]
  assign ces_211_0_io_ins_2 = ces_212_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_211_0_io_ins_3 = io_insVertical_1_211; // @[MockArray.scala 47:87]
  assign ces_212_0_clock = clock;
  assign ces_212_0_io_ins_0 = ces_211_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_212_0_io_ins_1 = io_insVertical_0_212; // @[MockArray.scala 45:87]
  assign ces_212_0_io_ins_2 = ces_213_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_212_0_io_ins_3 = io_insVertical_1_212; // @[MockArray.scala 47:87]
  assign ces_213_0_clock = clock;
  assign ces_213_0_io_ins_0 = ces_212_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_213_0_io_ins_1 = io_insVertical_0_213; // @[MockArray.scala 45:87]
  assign ces_213_0_io_ins_2 = ces_214_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_213_0_io_ins_3 = io_insVertical_1_213; // @[MockArray.scala 47:87]
  assign ces_214_0_clock = clock;
  assign ces_214_0_io_ins_0 = ces_213_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_214_0_io_ins_1 = io_insVertical_0_214; // @[MockArray.scala 45:87]
  assign ces_214_0_io_ins_2 = ces_215_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_214_0_io_ins_3 = io_insVertical_1_214; // @[MockArray.scala 47:87]
  assign ces_215_0_clock = clock;
  assign ces_215_0_io_ins_0 = ces_214_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_215_0_io_ins_1 = io_insVertical_0_215; // @[MockArray.scala 45:87]
  assign ces_215_0_io_ins_2 = ces_216_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_215_0_io_ins_3 = io_insVertical_1_215; // @[MockArray.scala 47:87]
  assign ces_216_0_clock = clock;
  assign ces_216_0_io_ins_0 = ces_215_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_216_0_io_ins_1 = io_insVertical_0_216; // @[MockArray.scala 45:87]
  assign ces_216_0_io_ins_2 = ces_217_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_216_0_io_ins_3 = io_insVertical_1_216; // @[MockArray.scala 47:87]
  assign ces_217_0_clock = clock;
  assign ces_217_0_io_ins_0 = ces_216_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_217_0_io_ins_1 = io_insVertical_0_217; // @[MockArray.scala 45:87]
  assign ces_217_0_io_ins_2 = ces_218_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_217_0_io_ins_3 = io_insVertical_1_217; // @[MockArray.scala 47:87]
  assign ces_218_0_clock = clock;
  assign ces_218_0_io_ins_0 = ces_217_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_218_0_io_ins_1 = io_insVertical_0_218; // @[MockArray.scala 45:87]
  assign ces_218_0_io_ins_2 = ces_219_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_218_0_io_ins_3 = io_insVertical_1_218; // @[MockArray.scala 47:87]
  assign ces_219_0_clock = clock;
  assign ces_219_0_io_ins_0 = ces_218_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_219_0_io_ins_1 = io_insVertical_0_219; // @[MockArray.scala 45:87]
  assign ces_219_0_io_ins_2 = ces_220_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_219_0_io_ins_3 = io_insVertical_1_219; // @[MockArray.scala 47:87]
  assign ces_220_0_clock = clock;
  assign ces_220_0_io_ins_0 = ces_219_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_220_0_io_ins_1 = io_insVertical_0_220; // @[MockArray.scala 45:87]
  assign ces_220_0_io_ins_2 = ces_221_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_220_0_io_ins_3 = io_insVertical_1_220; // @[MockArray.scala 47:87]
  assign ces_221_0_clock = clock;
  assign ces_221_0_io_ins_0 = ces_220_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_221_0_io_ins_1 = io_insVertical_0_221; // @[MockArray.scala 45:87]
  assign ces_221_0_io_ins_2 = ces_222_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_221_0_io_ins_3 = io_insVertical_1_221; // @[MockArray.scala 47:87]
  assign ces_222_0_clock = clock;
  assign ces_222_0_io_ins_0 = ces_221_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_222_0_io_ins_1 = io_insVertical_0_222; // @[MockArray.scala 45:87]
  assign ces_222_0_io_ins_2 = ces_223_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_222_0_io_ins_3 = io_insVertical_1_222; // @[MockArray.scala 47:87]
  assign ces_223_0_clock = clock;
  assign ces_223_0_io_ins_0 = ces_222_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_223_0_io_ins_1 = io_insVertical_0_223; // @[MockArray.scala 45:87]
  assign ces_223_0_io_ins_2 = ces_224_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_223_0_io_ins_3 = io_insVertical_1_223; // @[MockArray.scala 47:87]
  assign ces_224_0_clock = clock;
  assign ces_224_0_io_ins_0 = ces_223_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_224_0_io_ins_1 = io_insVertical_0_224; // @[MockArray.scala 45:87]
  assign ces_224_0_io_ins_2 = ces_225_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_224_0_io_ins_3 = io_insVertical_1_224; // @[MockArray.scala 47:87]
  assign ces_225_0_clock = clock;
  assign ces_225_0_io_ins_0 = ces_224_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_225_0_io_ins_1 = io_insVertical_0_225; // @[MockArray.scala 45:87]
  assign ces_225_0_io_ins_2 = ces_226_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_225_0_io_ins_3 = io_insVertical_1_225; // @[MockArray.scala 47:87]
  assign ces_226_0_clock = clock;
  assign ces_226_0_io_ins_0 = ces_225_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_226_0_io_ins_1 = io_insVertical_0_226; // @[MockArray.scala 45:87]
  assign ces_226_0_io_ins_2 = ces_227_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_226_0_io_ins_3 = io_insVertical_1_226; // @[MockArray.scala 47:87]
  assign ces_227_0_clock = clock;
  assign ces_227_0_io_ins_0 = ces_226_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_227_0_io_ins_1 = io_insVertical_0_227; // @[MockArray.scala 45:87]
  assign ces_227_0_io_ins_2 = ces_228_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_227_0_io_ins_3 = io_insVertical_1_227; // @[MockArray.scala 47:87]
  assign ces_228_0_clock = clock;
  assign ces_228_0_io_ins_0 = ces_227_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_228_0_io_ins_1 = io_insVertical_0_228; // @[MockArray.scala 45:87]
  assign ces_228_0_io_ins_2 = ces_229_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_228_0_io_ins_3 = io_insVertical_1_228; // @[MockArray.scala 47:87]
  assign ces_229_0_clock = clock;
  assign ces_229_0_io_ins_0 = ces_228_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_229_0_io_ins_1 = io_insVertical_0_229; // @[MockArray.scala 45:87]
  assign ces_229_0_io_ins_2 = ces_230_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_229_0_io_ins_3 = io_insVertical_1_229; // @[MockArray.scala 47:87]
  assign ces_230_0_clock = clock;
  assign ces_230_0_io_ins_0 = ces_229_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_230_0_io_ins_1 = io_insVertical_0_230; // @[MockArray.scala 45:87]
  assign ces_230_0_io_ins_2 = ces_231_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_230_0_io_ins_3 = io_insVertical_1_230; // @[MockArray.scala 47:87]
  assign ces_231_0_clock = clock;
  assign ces_231_0_io_ins_0 = ces_230_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_231_0_io_ins_1 = io_insVertical_0_231; // @[MockArray.scala 45:87]
  assign ces_231_0_io_ins_2 = ces_232_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_231_0_io_ins_3 = io_insVertical_1_231; // @[MockArray.scala 47:87]
  assign ces_232_0_clock = clock;
  assign ces_232_0_io_ins_0 = ces_231_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_232_0_io_ins_1 = io_insVertical_0_232; // @[MockArray.scala 45:87]
  assign ces_232_0_io_ins_2 = ces_233_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_232_0_io_ins_3 = io_insVertical_1_232; // @[MockArray.scala 47:87]
  assign ces_233_0_clock = clock;
  assign ces_233_0_io_ins_0 = ces_232_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_233_0_io_ins_1 = io_insVertical_0_233; // @[MockArray.scala 45:87]
  assign ces_233_0_io_ins_2 = ces_234_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_233_0_io_ins_3 = io_insVertical_1_233; // @[MockArray.scala 47:87]
  assign ces_234_0_clock = clock;
  assign ces_234_0_io_ins_0 = ces_233_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_234_0_io_ins_1 = io_insVertical_0_234; // @[MockArray.scala 45:87]
  assign ces_234_0_io_ins_2 = ces_235_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_234_0_io_ins_3 = io_insVertical_1_234; // @[MockArray.scala 47:87]
  assign ces_235_0_clock = clock;
  assign ces_235_0_io_ins_0 = ces_234_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_235_0_io_ins_1 = io_insVertical_0_235; // @[MockArray.scala 45:87]
  assign ces_235_0_io_ins_2 = ces_236_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_235_0_io_ins_3 = io_insVertical_1_235; // @[MockArray.scala 47:87]
  assign ces_236_0_clock = clock;
  assign ces_236_0_io_ins_0 = ces_235_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_236_0_io_ins_1 = io_insVertical_0_236; // @[MockArray.scala 45:87]
  assign ces_236_0_io_ins_2 = ces_237_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_236_0_io_ins_3 = io_insVertical_1_236; // @[MockArray.scala 47:87]
  assign ces_237_0_clock = clock;
  assign ces_237_0_io_ins_0 = ces_236_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_237_0_io_ins_1 = io_insVertical_0_237; // @[MockArray.scala 45:87]
  assign ces_237_0_io_ins_2 = ces_238_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_237_0_io_ins_3 = io_insVertical_1_237; // @[MockArray.scala 47:87]
  assign ces_238_0_clock = clock;
  assign ces_238_0_io_ins_0 = ces_237_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_238_0_io_ins_1 = io_insVertical_0_238; // @[MockArray.scala 45:87]
  assign ces_238_0_io_ins_2 = ces_239_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_238_0_io_ins_3 = io_insVertical_1_238; // @[MockArray.scala 47:87]
  assign ces_239_0_clock = clock;
  assign ces_239_0_io_ins_0 = ces_238_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_239_0_io_ins_1 = io_insVertical_0_239; // @[MockArray.scala 45:87]
  assign ces_239_0_io_ins_2 = ces_240_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_239_0_io_ins_3 = io_insVertical_1_239; // @[MockArray.scala 47:87]
  assign ces_240_0_clock = clock;
  assign ces_240_0_io_ins_0 = ces_239_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_240_0_io_ins_1 = io_insVertical_0_240; // @[MockArray.scala 45:87]
  assign ces_240_0_io_ins_2 = ces_241_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_240_0_io_ins_3 = io_insVertical_1_240; // @[MockArray.scala 47:87]
  assign ces_241_0_clock = clock;
  assign ces_241_0_io_ins_0 = ces_240_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_241_0_io_ins_1 = io_insVertical_0_241; // @[MockArray.scala 45:87]
  assign ces_241_0_io_ins_2 = ces_242_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_241_0_io_ins_3 = io_insVertical_1_241; // @[MockArray.scala 47:87]
  assign ces_242_0_clock = clock;
  assign ces_242_0_io_ins_0 = ces_241_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_242_0_io_ins_1 = io_insVertical_0_242; // @[MockArray.scala 45:87]
  assign ces_242_0_io_ins_2 = ces_243_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_242_0_io_ins_3 = io_insVertical_1_242; // @[MockArray.scala 47:87]
  assign ces_243_0_clock = clock;
  assign ces_243_0_io_ins_0 = ces_242_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_243_0_io_ins_1 = io_insVertical_0_243; // @[MockArray.scala 45:87]
  assign ces_243_0_io_ins_2 = ces_244_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_243_0_io_ins_3 = io_insVertical_1_243; // @[MockArray.scala 47:87]
  assign ces_244_0_clock = clock;
  assign ces_244_0_io_ins_0 = ces_243_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_244_0_io_ins_1 = io_insVertical_0_244; // @[MockArray.scala 45:87]
  assign ces_244_0_io_ins_2 = ces_245_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_244_0_io_ins_3 = io_insVertical_1_244; // @[MockArray.scala 47:87]
  assign ces_245_0_clock = clock;
  assign ces_245_0_io_ins_0 = ces_244_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_245_0_io_ins_1 = io_insVertical_0_245; // @[MockArray.scala 45:87]
  assign ces_245_0_io_ins_2 = ces_246_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_245_0_io_ins_3 = io_insVertical_1_245; // @[MockArray.scala 47:87]
  assign ces_246_0_clock = clock;
  assign ces_246_0_io_ins_0 = ces_245_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_246_0_io_ins_1 = io_insVertical_0_246; // @[MockArray.scala 45:87]
  assign ces_246_0_io_ins_2 = ces_247_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_246_0_io_ins_3 = io_insVertical_1_246; // @[MockArray.scala 47:87]
  assign ces_247_0_clock = clock;
  assign ces_247_0_io_ins_0 = ces_246_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_247_0_io_ins_1 = io_insVertical_0_247; // @[MockArray.scala 45:87]
  assign ces_247_0_io_ins_2 = ces_248_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_247_0_io_ins_3 = io_insVertical_1_247; // @[MockArray.scala 47:87]
  assign ces_248_0_clock = clock;
  assign ces_248_0_io_ins_0 = ces_247_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_248_0_io_ins_1 = io_insVertical_0_248; // @[MockArray.scala 45:87]
  assign ces_248_0_io_ins_2 = ces_249_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_248_0_io_ins_3 = io_insVertical_1_248; // @[MockArray.scala 47:87]
  assign ces_249_0_clock = clock;
  assign ces_249_0_io_ins_0 = ces_248_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_249_0_io_ins_1 = io_insVertical_0_249; // @[MockArray.scala 45:87]
  assign ces_249_0_io_ins_2 = ces_250_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_249_0_io_ins_3 = io_insVertical_1_249; // @[MockArray.scala 47:87]
  assign ces_250_0_clock = clock;
  assign ces_250_0_io_ins_0 = ces_249_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_250_0_io_ins_1 = io_insVertical_0_250; // @[MockArray.scala 45:87]
  assign ces_250_0_io_ins_2 = ces_251_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_250_0_io_ins_3 = io_insVertical_1_250; // @[MockArray.scala 47:87]
  assign ces_251_0_clock = clock;
  assign ces_251_0_io_ins_0 = ces_250_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_251_0_io_ins_1 = io_insVertical_0_251; // @[MockArray.scala 45:87]
  assign ces_251_0_io_ins_2 = ces_252_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_251_0_io_ins_3 = io_insVertical_1_251; // @[MockArray.scala 47:87]
  assign ces_252_0_clock = clock;
  assign ces_252_0_io_ins_0 = ces_251_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_252_0_io_ins_1 = io_insVertical_0_252; // @[MockArray.scala 45:87]
  assign ces_252_0_io_ins_2 = ces_253_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_252_0_io_ins_3 = io_insVertical_1_252; // @[MockArray.scala 47:87]
  assign ces_253_0_clock = clock;
  assign ces_253_0_io_ins_0 = ces_252_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_253_0_io_ins_1 = io_insVertical_0_253; // @[MockArray.scala 45:87]
  assign ces_253_0_io_ins_2 = ces_254_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_253_0_io_ins_3 = io_insVertical_1_253; // @[MockArray.scala 47:87]
  assign ces_254_0_clock = clock;
  assign ces_254_0_io_ins_0 = ces_253_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_254_0_io_ins_1 = io_insVertical_0_254; // @[MockArray.scala 45:87]
  assign ces_254_0_io_ins_2 = ces_255_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_254_0_io_ins_3 = io_insVertical_1_254; // @[MockArray.scala 47:87]
  assign ces_255_0_clock = clock;
  assign ces_255_0_io_ins_0 = ces_254_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_255_0_io_ins_1 = io_insVertical_0_255; // @[MockArray.scala 45:87]
  assign ces_255_0_io_ins_2 = io_insHorizontal_1_0; // @[MockArray.scala 46:87]
  assign ces_255_0_io_ins_3 = io_insVertical_1_255; // @[MockArray.scala 47:87]
endmodule
