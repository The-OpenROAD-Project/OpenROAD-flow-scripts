../../nangate45/lef/fakeram45_64x32.lef