VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_2048x39
  FOREIGN fakeram45_2048x39 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 206.910 BY 219.800 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.535 0.070 3.605 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.475 0.070 6.545 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.945 0.070 8.015 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.415 0.070 9.485 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.355 0.070 12.425 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.825 0.070 13.895 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.295 0.070 15.365 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.235 0.070 18.305 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.705 0.070 19.775 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.175 0.070 21.245 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.115 0.070 24.185 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.585 0.070 25.655 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.055 0.070 27.125 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.525 0.070 28.595 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.995 0.070 30.065 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.465 0.070 31.535 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.935 0.070 33.005 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.405 0.070 34.475 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.875 0.070 35.945 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.345 0.070 37.415 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.815 0.070 38.885 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.755 0.070 41.825 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.225 0.070 43.295 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.695 0.070 44.765 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.635 0.070 47.705 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.105 0.070 49.175 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.575 0.070 50.645 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.045 0.070 52.115 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.515 0.070 53.585 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.985 0.070 55.055 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.455 0.070 56.525 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.925 0.070 57.995 ;
    END
  END w_mask_in[38]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.595 0.070 63.665 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.065 0.070 65.135 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.535 0.070 66.605 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.005 0.070 68.075 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.475 0.070 69.545 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.945 0.070 71.015 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.415 0.070 72.485 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.885 0.070 73.955 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.355 0.070 75.425 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.825 0.070 76.895 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.295 0.070 78.365 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.765 0.070 79.835 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.235 0.070 81.305 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.705 0.070 82.775 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.175 0.070 84.245 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.645 0.070 85.715 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.115 0.070 87.185 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.585 0.070 88.655 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.055 0.070 90.125 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.525 0.070 91.595 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.995 0.070 93.065 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.465 0.070 94.535 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.935 0.070 96.005 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.405 0.070 97.475 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.875 0.070 98.945 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.345 0.070 100.415 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.815 0.070 101.885 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.285 0.070 103.355 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.755 0.070 104.825 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.225 0.070 106.295 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.695 0.070 107.765 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.165 0.070 109.235 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.635 0.070 110.705 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.105 0.070 112.175 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.575 0.070 113.645 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.045 0.070 115.115 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.515 0.070 116.585 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.985 0.070 118.055 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.455 0.070 119.525 ;
    END
  END rd_out[38]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.125 0.070 125.195 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.595 0.070 126.665 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.065 0.070 128.135 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.535 0.070 129.605 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 131.005 0.070 131.075 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.475 0.070 132.545 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 133.945 0.070 134.015 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 135.415 0.070 135.485 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.885 0.070 136.955 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.355 0.070 138.425 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.825 0.070 139.895 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 141.295 0.070 141.365 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.765 0.070 142.835 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.235 0.070 144.305 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.705 0.070 145.775 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.175 0.070 147.245 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.645 0.070 148.715 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.115 0.070 150.185 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.585 0.070 151.655 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.055 0.070 153.125 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.525 0.070 154.595 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.995 0.070 156.065 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.465 0.070 157.535 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.935 0.070 159.005 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.405 0.070 160.475 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.875 0.070 161.945 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.345 0.070 163.415 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.815 0.070 164.885 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.285 0.070 166.355 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.755 0.070 167.825 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.225 0.070 169.295 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.695 0.070 170.765 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.165 0.070 172.235 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.635 0.070 173.705 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.105 0.070 175.175 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.575 0.070 176.645 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.045 0.070 178.115 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.515 0.070 179.585 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.985 0.070 181.055 ;
    END
  END wd_in[38]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.655 0.070 186.725 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.125 0.070 188.195 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.595 0.070 189.665 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.065 0.070 191.135 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.535 0.070 192.605 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.005 0.070 194.075 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.475 0.070 195.545 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.945 0.070 197.015 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 198.415 0.070 198.485 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 199.885 0.070 199.955 ;
    END
  END addr_in[9]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 201.355 0.070 201.425 ;
    END
  END addr_in[10]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 207.025 0.070 207.095 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 208.495 0.070 208.565 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.965 0.070 210.035 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 217.700 ;
      RECT 5.320 2.100 5.600 217.700 ;
      RECT 8.680 2.100 8.960 217.700 ;
      RECT 12.040 2.100 12.320 217.700 ;
      RECT 15.400 2.100 15.680 217.700 ;
      RECT 18.760 2.100 19.040 217.700 ;
      RECT 22.120 2.100 22.400 217.700 ;
      RECT 25.480 2.100 25.760 217.700 ;
      RECT 28.840 2.100 29.120 217.700 ;
      RECT 32.200 2.100 32.480 217.700 ;
      RECT 35.560 2.100 35.840 217.700 ;
      RECT 38.920 2.100 39.200 217.700 ;
      RECT 42.280 2.100 42.560 217.700 ;
      RECT 45.640 2.100 45.920 217.700 ;
      RECT 49.000 2.100 49.280 217.700 ;
      RECT 52.360 2.100 52.640 217.700 ;
      RECT 55.720 2.100 56.000 217.700 ;
      RECT 59.080 2.100 59.360 217.700 ;
      RECT 62.440 2.100 62.720 217.700 ;
      RECT 65.800 2.100 66.080 217.700 ;
      RECT 69.160 2.100 69.440 217.700 ;
      RECT 72.520 2.100 72.800 217.700 ;
      RECT 75.880 2.100 76.160 217.700 ;
      RECT 79.240 2.100 79.520 217.700 ;
      RECT 82.600 2.100 82.880 217.700 ;
      RECT 85.960 2.100 86.240 217.700 ;
      RECT 89.320 2.100 89.600 217.700 ;
      RECT 92.680 2.100 92.960 217.700 ;
      RECT 96.040 2.100 96.320 217.700 ;
      RECT 99.400 2.100 99.680 217.700 ;
      RECT 102.760 2.100 103.040 217.700 ;
      RECT 106.120 2.100 106.400 217.700 ;
      RECT 109.480 2.100 109.760 217.700 ;
      RECT 112.840 2.100 113.120 217.700 ;
      RECT 116.200 2.100 116.480 217.700 ;
      RECT 119.560 2.100 119.840 217.700 ;
      RECT 122.920 2.100 123.200 217.700 ;
      RECT 126.280 2.100 126.560 217.700 ;
      RECT 129.640 2.100 129.920 217.700 ;
      RECT 133.000 2.100 133.280 217.700 ;
      RECT 136.360 2.100 136.640 217.700 ;
      RECT 139.720 2.100 140.000 217.700 ;
      RECT 143.080 2.100 143.360 217.700 ;
      RECT 146.440 2.100 146.720 217.700 ;
      RECT 149.800 2.100 150.080 217.700 ;
      RECT 153.160 2.100 153.440 217.700 ;
      RECT 156.520 2.100 156.800 217.700 ;
      RECT 159.880 2.100 160.160 217.700 ;
      RECT 163.240 2.100 163.520 217.700 ;
      RECT 166.600 2.100 166.880 217.700 ;
      RECT 169.960 2.100 170.240 217.700 ;
      RECT 173.320 2.100 173.600 217.700 ;
      RECT 176.680 2.100 176.960 217.700 ;
      RECT 180.040 2.100 180.320 217.700 ;
      RECT 183.400 2.100 183.680 217.700 ;
      RECT 186.760 2.100 187.040 217.700 ;
      RECT 190.120 2.100 190.400 217.700 ;
      RECT 193.480 2.100 193.760 217.700 ;
      RECT 196.840 2.100 197.120 217.700 ;
      RECT 200.200 2.100 200.480 217.700 ;
      RECT 203.560 2.100 203.840 217.700 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 217.700 ;
      RECT 7.000 2.100 7.280 217.700 ;
      RECT 10.360 2.100 10.640 217.700 ;
      RECT 13.720 2.100 14.000 217.700 ;
      RECT 17.080 2.100 17.360 217.700 ;
      RECT 20.440 2.100 20.720 217.700 ;
      RECT 23.800 2.100 24.080 217.700 ;
      RECT 27.160 2.100 27.440 217.700 ;
      RECT 30.520 2.100 30.800 217.700 ;
      RECT 33.880 2.100 34.160 217.700 ;
      RECT 37.240 2.100 37.520 217.700 ;
      RECT 40.600 2.100 40.880 217.700 ;
      RECT 43.960 2.100 44.240 217.700 ;
      RECT 47.320 2.100 47.600 217.700 ;
      RECT 50.680 2.100 50.960 217.700 ;
      RECT 54.040 2.100 54.320 217.700 ;
      RECT 57.400 2.100 57.680 217.700 ;
      RECT 60.760 2.100 61.040 217.700 ;
      RECT 64.120 2.100 64.400 217.700 ;
      RECT 67.480 2.100 67.760 217.700 ;
      RECT 70.840 2.100 71.120 217.700 ;
      RECT 74.200 2.100 74.480 217.700 ;
      RECT 77.560 2.100 77.840 217.700 ;
      RECT 80.920 2.100 81.200 217.700 ;
      RECT 84.280 2.100 84.560 217.700 ;
      RECT 87.640 2.100 87.920 217.700 ;
      RECT 91.000 2.100 91.280 217.700 ;
      RECT 94.360 2.100 94.640 217.700 ;
      RECT 97.720 2.100 98.000 217.700 ;
      RECT 101.080 2.100 101.360 217.700 ;
      RECT 104.440 2.100 104.720 217.700 ;
      RECT 107.800 2.100 108.080 217.700 ;
      RECT 111.160 2.100 111.440 217.700 ;
      RECT 114.520 2.100 114.800 217.700 ;
      RECT 117.880 2.100 118.160 217.700 ;
      RECT 121.240 2.100 121.520 217.700 ;
      RECT 124.600 2.100 124.880 217.700 ;
      RECT 127.960 2.100 128.240 217.700 ;
      RECT 131.320 2.100 131.600 217.700 ;
      RECT 134.680 2.100 134.960 217.700 ;
      RECT 138.040 2.100 138.320 217.700 ;
      RECT 141.400 2.100 141.680 217.700 ;
      RECT 144.760 2.100 145.040 217.700 ;
      RECT 148.120 2.100 148.400 217.700 ;
      RECT 151.480 2.100 151.760 217.700 ;
      RECT 154.840 2.100 155.120 217.700 ;
      RECT 158.200 2.100 158.480 217.700 ;
      RECT 161.560 2.100 161.840 217.700 ;
      RECT 164.920 2.100 165.200 217.700 ;
      RECT 168.280 2.100 168.560 217.700 ;
      RECT 171.640 2.100 171.920 217.700 ;
      RECT 175.000 2.100 175.280 217.700 ;
      RECT 178.360 2.100 178.640 217.700 ;
      RECT 181.720 2.100 182.000 217.700 ;
      RECT 185.080 2.100 185.360 217.700 ;
      RECT 188.440 2.100 188.720 217.700 ;
      RECT 191.800 2.100 192.080 217.700 ;
      RECT 195.160 2.100 195.440 217.700 ;
      RECT 198.520 2.100 198.800 217.700 ;
      RECT 201.880 2.100 202.160 217.700 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 206.910 219.800 ;
    LAYER metal2 ;
    RECT 0 0 206.910 219.800 ;
    LAYER metal3 ;
    RECT 0.070 0 206.910 219.800 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 3.535 ;
    RECT 0 3.605 0.070 5.005 ;
    RECT 0 5.075 0.070 6.475 ;
    RECT 0 6.545 0.070 7.945 ;
    RECT 0 8.015 0.070 9.415 ;
    RECT 0 9.485 0.070 10.885 ;
    RECT 0 10.955 0.070 12.355 ;
    RECT 0 12.425 0.070 13.825 ;
    RECT 0 13.895 0.070 15.295 ;
    RECT 0 15.365 0.070 16.765 ;
    RECT 0 16.835 0.070 18.235 ;
    RECT 0 18.305 0.070 19.705 ;
    RECT 0 19.775 0.070 21.175 ;
    RECT 0 21.245 0.070 22.645 ;
    RECT 0 22.715 0.070 24.115 ;
    RECT 0 24.185 0.070 25.585 ;
    RECT 0 25.655 0.070 27.055 ;
    RECT 0 27.125 0.070 28.525 ;
    RECT 0 28.595 0.070 29.995 ;
    RECT 0 30.065 0.070 31.465 ;
    RECT 0 31.535 0.070 32.935 ;
    RECT 0 33.005 0.070 34.405 ;
    RECT 0 34.475 0.070 35.875 ;
    RECT 0 35.945 0.070 37.345 ;
    RECT 0 37.415 0.070 38.815 ;
    RECT 0 38.885 0.070 40.285 ;
    RECT 0 40.355 0.070 41.755 ;
    RECT 0 41.825 0.070 43.225 ;
    RECT 0 43.295 0.070 44.695 ;
    RECT 0 44.765 0.070 46.165 ;
    RECT 0 46.235 0.070 47.635 ;
    RECT 0 47.705 0.070 49.105 ;
    RECT 0 49.175 0.070 50.575 ;
    RECT 0 50.645 0.070 52.045 ;
    RECT 0 52.115 0.070 53.515 ;
    RECT 0 53.585 0.070 54.985 ;
    RECT 0 55.055 0.070 56.455 ;
    RECT 0 56.525 0.070 57.925 ;
    RECT 0 57.995 0.070 63.595 ;
    RECT 0 63.665 0.070 65.065 ;
    RECT 0 65.135 0.070 66.535 ;
    RECT 0 66.605 0.070 68.005 ;
    RECT 0 68.075 0.070 69.475 ;
    RECT 0 69.545 0.070 70.945 ;
    RECT 0 71.015 0.070 72.415 ;
    RECT 0 72.485 0.070 73.885 ;
    RECT 0 73.955 0.070 75.355 ;
    RECT 0 75.425 0.070 76.825 ;
    RECT 0 76.895 0.070 78.295 ;
    RECT 0 78.365 0.070 79.765 ;
    RECT 0 79.835 0.070 81.235 ;
    RECT 0 81.305 0.070 82.705 ;
    RECT 0 82.775 0.070 84.175 ;
    RECT 0 84.245 0.070 85.645 ;
    RECT 0 85.715 0.070 87.115 ;
    RECT 0 87.185 0.070 88.585 ;
    RECT 0 88.655 0.070 90.055 ;
    RECT 0 90.125 0.070 91.525 ;
    RECT 0 91.595 0.070 92.995 ;
    RECT 0 93.065 0.070 94.465 ;
    RECT 0 94.535 0.070 95.935 ;
    RECT 0 96.005 0.070 97.405 ;
    RECT 0 97.475 0.070 98.875 ;
    RECT 0 98.945 0.070 100.345 ;
    RECT 0 100.415 0.070 101.815 ;
    RECT 0 101.885 0.070 103.285 ;
    RECT 0 103.355 0.070 104.755 ;
    RECT 0 104.825 0.070 106.225 ;
    RECT 0 106.295 0.070 107.695 ;
    RECT 0 107.765 0.070 109.165 ;
    RECT 0 109.235 0.070 110.635 ;
    RECT 0 110.705 0.070 112.105 ;
    RECT 0 112.175 0.070 113.575 ;
    RECT 0 113.645 0.070 115.045 ;
    RECT 0 115.115 0.070 116.515 ;
    RECT 0 116.585 0.070 117.985 ;
    RECT 0 118.055 0.070 119.455 ;
    RECT 0 119.525 0.070 125.125 ;
    RECT 0 125.195 0.070 126.595 ;
    RECT 0 126.665 0.070 128.065 ;
    RECT 0 128.135 0.070 129.535 ;
    RECT 0 129.605 0.070 131.005 ;
    RECT 0 131.075 0.070 132.475 ;
    RECT 0 132.545 0.070 133.945 ;
    RECT 0 134.015 0.070 135.415 ;
    RECT 0 135.485 0.070 136.885 ;
    RECT 0 136.955 0.070 138.355 ;
    RECT 0 138.425 0.070 139.825 ;
    RECT 0 139.895 0.070 141.295 ;
    RECT 0 141.365 0.070 142.765 ;
    RECT 0 142.835 0.070 144.235 ;
    RECT 0 144.305 0.070 145.705 ;
    RECT 0 145.775 0.070 147.175 ;
    RECT 0 147.245 0.070 148.645 ;
    RECT 0 148.715 0.070 150.115 ;
    RECT 0 150.185 0.070 151.585 ;
    RECT 0 151.655 0.070 153.055 ;
    RECT 0 153.125 0.070 154.525 ;
    RECT 0 154.595 0.070 155.995 ;
    RECT 0 156.065 0.070 157.465 ;
    RECT 0 157.535 0.070 158.935 ;
    RECT 0 159.005 0.070 160.405 ;
    RECT 0 160.475 0.070 161.875 ;
    RECT 0 161.945 0.070 163.345 ;
    RECT 0 163.415 0.070 164.815 ;
    RECT 0 164.885 0.070 166.285 ;
    RECT 0 166.355 0.070 167.755 ;
    RECT 0 167.825 0.070 169.225 ;
    RECT 0 169.295 0.070 170.695 ;
    RECT 0 170.765 0.070 172.165 ;
    RECT 0 172.235 0.070 173.635 ;
    RECT 0 173.705 0.070 175.105 ;
    RECT 0 175.175 0.070 176.575 ;
    RECT 0 176.645 0.070 178.045 ;
    RECT 0 178.115 0.070 179.515 ;
    RECT 0 179.585 0.070 180.985 ;
    RECT 0 181.055 0.070 186.655 ;
    RECT 0 186.725 0.070 188.125 ;
    RECT 0 188.195 0.070 189.595 ;
    RECT 0 189.665 0.070 191.065 ;
    RECT 0 191.135 0.070 192.535 ;
    RECT 0 192.605 0.070 194.005 ;
    RECT 0 194.075 0.070 195.475 ;
    RECT 0 195.545 0.070 196.945 ;
    RECT 0 197.015 0.070 198.415 ;
    RECT 0 198.485 0.070 199.885 ;
    RECT 0 199.955 0.070 201.355 ;
    RECT 0 201.425 0.070 207.025 ;
    RECT 0 207.095 0.070 208.495 ;
    RECT 0 208.565 0.070 209.965 ;
    RECT 0 210.035 0.070 219.800 ;
    LAYER metal4 ;
    RECT 0 0 206.910 2.100 ;
    RECT 0 217.700 206.910 219.800 ;
    RECT 0.000 2.100 1.960 217.700 ;
    RECT 2.240 2.100 3.640 217.700 ;
    RECT 3.920 2.100 5.320 217.700 ;
    RECT 5.600 2.100 7.000 217.700 ;
    RECT 7.280 2.100 8.680 217.700 ;
    RECT 8.960 2.100 10.360 217.700 ;
    RECT 10.640 2.100 12.040 217.700 ;
    RECT 12.320 2.100 13.720 217.700 ;
    RECT 14.000 2.100 15.400 217.700 ;
    RECT 15.680 2.100 17.080 217.700 ;
    RECT 17.360 2.100 18.760 217.700 ;
    RECT 19.040 2.100 20.440 217.700 ;
    RECT 20.720 2.100 22.120 217.700 ;
    RECT 22.400 2.100 23.800 217.700 ;
    RECT 24.080 2.100 25.480 217.700 ;
    RECT 25.760 2.100 27.160 217.700 ;
    RECT 27.440 2.100 28.840 217.700 ;
    RECT 29.120 2.100 30.520 217.700 ;
    RECT 30.800 2.100 32.200 217.700 ;
    RECT 32.480 2.100 33.880 217.700 ;
    RECT 34.160 2.100 35.560 217.700 ;
    RECT 35.840 2.100 37.240 217.700 ;
    RECT 37.520 2.100 38.920 217.700 ;
    RECT 39.200 2.100 40.600 217.700 ;
    RECT 40.880 2.100 42.280 217.700 ;
    RECT 42.560 2.100 43.960 217.700 ;
    RECT 44.240 2.100 45.640 217.700 ;
    RECT 45.920 2.100 47.320 217.700 ;
    RECT 47.600 2.100 49.000 217.700 ;
    RECT 49.280 2.100 50.680 217.700 ;
    RECT 50.960 2.100 52.360 217.700 ;
    RECT 52.640 2.100 54.040 217.700 ;
    RECT 54.320 2.100 55.720 217.700 ;
    RECT 56.000 2.100 57.400 217.700 ;
    RECT 57.680 2.100 59.080 217.700 ;
    RECT 59.360 2.100 60.760 217.700 ;
    RECT 61.040 2.100 62.440 217.700 ;
    RECT 62.720 2.100 64.120 217.700 ;
    RECT 64.400 2.100 65.800 217.700 ;
    RECT 66.080 2.100 67.480 217.700 ;
    RECT 67.760 2.100 69.160 217.700 ;
    RECT 69.440 2.100 70.840 217.700 ;
    RECT 71.120 2.100 72.520 217.700 ;
    RECT 72.800 2.100 74.200 217.700 ;
    RECT 74.480 2.100 75.880 217.700 ;
    RECT 76.160 2.100 77.560 217.700 ;
    RECT 77.840 2.100 79.240 217.700 ;
    RECT 79.520 2.100 80.920 217.700 ;
    RECT 81.200 2.100 82.600 217.700 ;
    RECT 82.880 2.100 84.280 217.700 ;
    RECT 84.560 2.100 85.960 217.700 ;
    RECT 86.240 2.100 87.640 217.700 ;
    RECT 87.920 2.100 89.320 217.700 ;
    RECT 89.600 2.100 91.000 217.700 ;
    RECT 91.280 2.100 92.680 217.700 ;
    RECT 92.960 2.100 94.360 217.700 ;
    RECT 94.640 2.100 96.040 217.700 ;
    RECT 96.320 2.100 97.720 217.700 ;
    RECT 98.000 2.100 99.400 217.700 ;
    RECT 99.680 2.100 101.080 217.700 ;
    RECT 101.360 2.100 102.760 217.700 ;
    RECT 103.040 2.100 104.440 217.700 ;
    RECT 104.720 2.100 106.120 217.700 ;
    RECT 106.400 2.100 107.800 217.700 ;
    RECT 108.080 2.100 109.480 217.700 ;
    RECT 109.760 2.100 111.160 217.700 ;
    RECT 111.440 2.100 112.840 217.700 ;
    RECT 113.120 2.100 114.520 217.700 ;
    RECT 114.800 2.100 116.200 217.700 ;
    RECT 116.480 2.100 117.880 217.700 ;
    RECT 118.160 2.100 119.560 217.700 ;
    RECT 119.840 2.100 121.240 217.700 ;
    RECT 121.520 2.100 122.920 217.700 ;
    RECT 123.200 2.100 124.600 217.700 ;
    RECT 124.880 2.100 126.280 217.700 ;
    RECT 126.560 2.100 127.960 217.700 ;
    RECT 128.240 2.100 129.640 217.700 ;
    RECT 129.920 2.100 131.320 217.700 ;
    RECT 131.600 2.100 133.000 217.700 ;
    RECT 133.280 2.100 134.680 217.700 ;
    RECT 134.960 2.100 136.360 217.700 ;
    RECT 136.640 2.100 138.040 217.700 ;
    RECT 138.320 2.100 139.720 217.700 ;
    RECT 140.000 2.100 141.400 217.700 ;
    RECT 141.680 2.100 143.080 217.700 ;
    RECT 143.360 2.100 144.760 217.700 ;
    RECT 145.040 2.100 146.440 217.700 ;
    RECT 146.720 2.100 148.120 217.700 ;
    RECT 148.400 2.100 149.800 217.700 ;
    RECT 150.080 2.100 151.480 217.700 ;
    RECT 151.760 2.100 153.160 217.700 ;
    RECT 153.440 2.100 154.840 217.700 ;
    RECT 155.120 2.100 156.520 217.700 ;
    RECT 156.800 2.100 158.200 217.700 ;
    RECT 158.480 2.100 159.880 217.700 ;
    RECT 160.160 2.100 161.560 217.700 ;
    RECT 161.840 2.100 163.240 217.700 ;
    RECT 163.520 2.100 164.920 217.700 ;
    RECT 165.200 2.100 166.600 217.700 ;
    RECT 166.880 2.100 168.280 217.700 ;
    RECT 168.560 2.100 169.960 217.700 ;
    RECT 170.240 2.100 171.640 217.700 ;
    RECT 171.920 2.100 173.320 217.700 ;
    RECT 173.600 2.100 175.000 217.700 ;
    RECT 175.280 2.100 176.680 217.700 ;
    RECT 176.960 2.100 178.360 217.700 ;
    RECT 178.640 2.100 180.040 217.700 ;
    RECT 180.320 2.100 181.720 217.700 ;
    RECT 182.000 2.100 183.400 217.700 ;
    RECT 183.680 2.100 185.080 217.700 ;
    RECT 185.360 2.100 186.760 217.700 ;
    RECT 187.040 2.100 188.440 217.700 ;
    RECT 188.720 2.100 190.120 217.700 ;
    RECT 190.400 2.100 191.800 217.700 ;
    RECT 192.080 2.100 193.480 217.700 ;
    RECT 193.760 2.100 195.160 217.700 ;
    RECT 195.440 2.100 196.840 217.700 ;
    RECT 197.120 2.100 198.520 217.700 ;
    RECT 198.800 2.100 200.200 217.700 ;
    RECT 200.480 2.100 201.880 217.700 ;
    RECT 202.160 2.100 203.560 217.700 ;
    RECT 203.840 2.100 206.910 217.700 ;
    LAYER OVERLAP ;
    RECT 0 0 206.910 219.800 ;
  END
END fakeram45_2048x39

END LIBRARY
