module MuxTest_width_1_inputs_8_outputs_16_pipeline_0( // @[:@3.2]
  input        clock, // @[:@4.4]
  input        reset, // @[:@5.4]
  input  [2:0] io_selects_0_0, // @[:@6.4]
  input  [2:0] io_selects_0_1, // @[:@6.4]
  input  [2:0] io_selects_1_0, // @[:@6.4]
  input  [2:0] io_selects_1_1, // @[:@6.4]
  input  [2:0] io_selects_2_0, // @[:@6.4]
  input  [2:0] io_selects_2_1, // @[:@6.4]
  input  [2:0] io_selects_3_0, // @[:@6.4]
  input  [2:0] io_selects_3_1, // @[:@6.4]
  input  [2:0] io_selects_4_0, // @[:@6.4]
  input  [2:0] io_selects_4_1, // @[:@6.4]
  input  [2:0] io_selects_5_0, // @[:@6.4]
  input  [2:0] io_selects_5_1, // @[:@6.4]
  input  [2:0] io_selects_6_0, // @[:@6.4]
  input  [2:0] io_selects_6_1, // @[:@6.4]
  input  [2:0] io_selects_7_0, // @[:@6.4]
  input  [2:0] io_selects_7_1, // @[:@6.4]
  input  [2:0] io_selects_8_0, // @[:@6.4]
  input  [2:0] io_selects_8_1, // @[:@6.4]
  input  [2:0] io_selects_9_0, // @[:@6.4]
  input  [2:0] io_selects_9_1, // @[:@6.4]
  input  [2:0] io_selects_10_0, // @[:@6.4]
  input  [2:0] io_selects_10_1, // @[:@6.4]
  input  [2:0] io_selects_11_0, // @[:@6.4]
  input  [2:0] io_selects_11_1, // @[:@6.4]
  input  [2:0] io_selects_12_0, // @[:@6.4]
  input  [2:0] io_selects_12_1, // @[:@6.4]
  input  [2:0] io_selects_13_0, // @[:@6.4]
  input  [2:0] io_selects_13_1, // @[:@6.4]
  input  [2:0] io_selects_14_0, // @[:@6.4]
  input  [2:0] io_selects_14_1, // @[:@6.4]
  input  [2:0] io_selects_15_0, // @[:@6.4]
  input  [2:0] io_selects_15_1, // @[:@6.4]
  input  [2:0] io_operation_0, // @[:@6.4]
  input  [2:0] io_operation_1, // @[:@6.4]
  input  [2:0] io_operation_2, // @[:@6.4]
  input  [2:0] io_operation_3, // @[:@6.4]
  input  [2:0] io_operation_4, // @[:@6.4]
  input  [2:0] io_operation_5, // @[:@6.4]
  input  [2:0] io_operation_6, // @[:@6.4]
  input  [2:0] io_operation_7, // @[:@6.4]
  input  [2:0] io_operation_8, // @[:@6.4]
  input  [2:0] io_operation_9, // @[:@6.4]
  input  [2:0] io_operation_10, // @[:@6.4]
  input  [2:0] io_operation_11, // @[:@6.4]
  input  [2:0] io_operation_12, // @[:@6.4]
  input  [2:0] io_operation_13, // @[:@6.4]
  input  [2:0] io_operation_14, // @[:@6.4]
  input  [2:0] io_operation_15, // @[:@6.4]
  input        io_inputs_0, // @[:@6.4]
  input        io_inputs_1, // @[:@6.4]
  input        io_inputs_2, // @[:@6.4]
  input        io_inputs_3, // @[:@6.4]
  input        io_inputs_4, // @[:@6.4]
  input        io_inputs_5, // @[:@6.4]
  input        io_inputs_6, // @[:@6.4]
  input        io_inputs_7, // @[:@6.4]
  output       io_outputs_0, // @[:@6.4]
  output       io_outputs_1, // @[:@6.4]
  output       io_outputs_2, // @[:@6.4]
  output       io_outputs_3, // @[:@6.4]
  output       io_outputs_4, // @[:@6.4]
  output       io_outputs_5, // @[:@6.4]
  output       io_outputs_6, // @[:@6.4]
  output       io_outputs_7, // @[:@6.4]
  output       io_outputs_8, // @[:@6.4]
  output       io_outputs_9, // @[:@6.4]
  output       io_outputs_10, // @[:@6.4]
  output       io_outputs_11, // @[:@6.4]
  output       io_outputs_12, // @[:@6.4]
  output       io_outputs_13, // @[:@6.4]
  output       io_outputs_14, // @[:@6.4]
  output       io_outputs_15 // @[:@6.4]
);
  wire  _GEN_1; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  wire  _GEN_2; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  wire  _GEN_3; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  wire  _GEN_4; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  wire  _GEN_5; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  wire  _GEN_6; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  wire  _GEN_7; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  wire  _GEN_9; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  wire  _GEN_10; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  wire  _GEN_11; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  wire  _GEN_12; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  wire  _GEN_13; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  wire  _GEN_14; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  wire  _GEN_15; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  wire [1:0] _T_706; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  wire  _T_707; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@9.4]
  wire [1:0] _T_709; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@10.4]
  wire  _T_711; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@11.4]
  wire  _T_712; // @[Mux.scala 46:19:@12.4]
  wire  _T_713; // @[Mux.scala 46:16:@13.4]
  wire  _T_714; // @[Mux.scala 46:19:@14.4]
  wire [1:0] _T_715; // @[Mux.scala 46:16:@15.4]
  wire  _T_716; // @[Mux.scala 46:19:@16.4]
  wire [1:0] _T_717; // @[Mux.scala 46:16:@17.4]
  wire  _T_718; // @[Mux.scala 46:19:@18.4]
  wire [1:0] _T_719; // @[Mux.scala 46:16:@19.4]
  wire  _GEN_17; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  wire  _GEN_18; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  wire  _GEN_19; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  wire  _GEN_20; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  wire  _GEN_21; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  wire  _GEN_22; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  wire  _GEN_23; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  wire  _GEN_25; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  wire  _GEN_26; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  wire  _GEN_27; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  wire  _GEN_28; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  wire  _GEN_29; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  wire  _GEN_30; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  wire  _GEN_31; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  wire [1:0] _T_723; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  wire  _T_724; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@21.4]
  wire [1:0] _T_726; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@22.4]
  wire  _T_728; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@23.4]
  wire  _T_729; // @[Mux.scala 46:19:@24.4]
  wire  _T_730; // @[Mux.scala 46:16:@25.4]
  wire  _T_731; // @[Mux.scala 46:19:@26.4]
  wire [1:0] _T_732; // @[Mux.scala 46:16:@27.4]
  wire  _T_733; // @[Mux.scala 46:19:@28.4]
  wire [1:0] _T_734; // @[Mux.scala 46:16:@29.4]
  wire  _T_735; // @[Mux.scala 46:19:@30.4]
  wire [1:0] _T_736; // @[Mux.scala 46:16:@31.4]
  wire  _GEN_33; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  wire  _GEN_34; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  wire  _GEN_35; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  wire  _GEN_36; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  wire  _GEN_37; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  wire  _GEN_38; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  wire  _GEN_39; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  wire  _GEN_41; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  wire  _GEN_42; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  wire  _GEN_43; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  wire  _GEN_44; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  wire  _GEN_45; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  wire  _GEN_46; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  wire  _GEN_47; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  wire [1:0] _T_740; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  wire  _T_741; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@33.4]
  wire [1:0] _T_743; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@34.4]
  wire  _T_745; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@35.4]
  wire  _T_746; // @[Mux.scala 46:19:@36.4]
  wire  _T_747; // @[Mux.scala 46:16:@37.4]
  wire  _T_748; // @[Mux.scala 46:19:@38.4]
  wire [1:0] _T_749; // @[Mux.scala 46:16:@39.4]
  wire  _T_750; // @[Mux.scala 46:19:@40.4]
  wire [1:0] _T_751; // @[Mux.scala 46:16:@41.4]
  wire  _T_752; // @[Mux.scala 46:19:@42.4]
  wire [1:0] _T_753; // @[Mux.scala 46:16:@43.4]
  wire  _GEN_49; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  wire  _GEN_50; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  wire  _GEN_51; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  wire  _GEN_52; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  wire  _GEN_53; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  wire  _GEN_54; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  wire  _GEN_55; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  wire  _GEN_57; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  wire  _GEN_58; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  wire  _GEN_59; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  wire  _GEN_60; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  wire  _GEN_61; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  wire  _GEN_62; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  wire  _GEN_63; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  wire [1:0] _T_757; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  wire  _T_758; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@45.4]
  wire [1:0] _T_760; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@46.4]
  wire  _T_762; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@47.4]
  wire  _T_763; // @[Mux.scala 46:19:@48.4]
  wire  _T_764; // @[Mux.scala 46:16:@49.4]
  wire  _T_765; // @[Mux.scala 46:19:@50.4]
  wire [1:0] _T_766; // @[Mux.scala 46:16:@51.4]
  wire  _T_767; // @[Mux.scala 46:19:@52.4]
  wire [1:0] _T_768; // @[Mux.scala 46:16:@53.4]
  wire  _T_769; // @[Mux.scala 46:19:@54.4]
  wire [1:0] _T_770; // @[Mux.scala 46:16:@55.4]
  wire  _GEN_65; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  wire  _GEN_66; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  wire  _GEN_67; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  wire  _GEN_68; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  wire  _GEN_69; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  wire  _GEN_70; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  wire  _GEN_71; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  wire  _GEN_73; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  wire  _GEN_74; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  wire  _GEN_75; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  wire  _GEN_76; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  wire  _GEN_77; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  wire  _GEN_78; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  wire  _GEN_79; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  wire [1:0] _T_774; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  wire  _T_775; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@57.4]
  wire [1:0] _T_777; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@58.4]
  wire  _T_779; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@59.4]
  wire  _T_780; // @[Mux.scala 46:19:@60.4]
  wire  _T_781; // @[Mux.scala 46:16:@61.4]
  wire  _T_782; // @[Mux.scala 46:19:@62.4]
  wire [1:0] _T_783; // @[Mux.scala 46:16:@63.4]
  wire  _T_784; // @[Mux.scala 46:19:@64.4]
  wire [1:0] _T_785; // @[Mux.scala 46:16:@65.4]
  wire  _T_786; // @[Mux.scala 46:19:@66.4]
  wire [1:0] _T_787; // @[Mux.scala 46:16:@67.4]
  wire  _GEN_81; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  wire  _GEN_82; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  wire  _GEN_83; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  wire  _GEN_84; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  wire  _GEN_85; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  wire  _GEN_86; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  wire  _GEN_87; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  wire  _GEN_89; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  wire  _GEN_90; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  wire  _GEN_91; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  wire  _GEN_92; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  wire  _GEN_93; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  wire  _GEN_94; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  wire  _GEN_95; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  wire [1:0] _T_791; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  wire  _T_792; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@69.4]
  wire [1:0] _T_794; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@70.4]
  wire  _T_796; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@71.4]
  wire  _T_797; // @[Mux.scala 46:19:@72.4]
  wire  _T_798; // @[Mux.scala 46:16:@73.4]
  wire  _T_799; // @[Mux.scala 46:19:@74.4]
  wire [1:0] _T_800; // @[Mux.scala 46:16:@75.4]
  wire  _T_801; // @[Mux.scala 46:19:@76.4]
  wire [1:0] _T_802; // @[Mux.scala 46:16:@77.4]
  wire  _T_803; // @[Mux.scala 46:19:@78.4]
  wire [1:0] _T_804; // @[Mux.scala 46:16:@79.4]
  wire  _GEN_97; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  wire  _GEN_98; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  wire  _GEN_99; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  wire  _GEN_100; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  wire  _GEN_101; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  wire  _GEN_102; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  wire  _GEN_103; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  wire  _GEN_105; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  wire  _GEN_106; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  wire  _GEN_107; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  wire  _GEN_108; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  wire  _GEN_109; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  wire  _GEN_110; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  wire  _GEN_111; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  wire [1:0] _T_808; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  wire  _T_809; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@81.4]
  wire [1:0] _T_811; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@82.4]
  wire  _T_813; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@83.4]
  wire  _T_814; // @[Mux.scala 46:19:@84.4]
  wire  _T_815; // @[Mux.scala 46:16:@85.4]
  wire  _T_816; // @[Mux.scala 46:19:@86.4]
  wire [1:0] _T_817; // @[Mux.scala 46:16:@87.4]
  wire  _T_818; // @[Mux.scala 46:19:@88.4]
  wire [1:0] _T_819; // @[Mux.scala 46:16:@89.4]
  wire  _T_820; // @[Mux.scala 46:19:@90.4]
  wire [1:0] _T_821; // @[Mux.scala 46:16:@91.4]
  wire  _GEN_113; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  wire  _GEN_114; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  wire  _GEN_115; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  wire  _GEN_116; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  wire  _GEN_117; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  wire  _GEN_118; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  wire  _GEN_119; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  wire  _GEN_121; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  wire  _GEN_122; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  wire  _GEN_123; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  wire  _GEN_124; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  wire  _GEN_125; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  wire  _GEN_126; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  wire  _GEN_127; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  wire [1:0] _T_825; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  wire  _T_826; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@93.4]
  wire [1:0] _T_828; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@94.4]
  wire  _T_830; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@95.4]
  wire  _T_831; // @[Mux.scala 46:19:@96.4]
  wire  _T_832; // @[Mux.scala 46:16:@97.4]
  wire  _T_833; // @[Mux.scala 46:19:@98.4]
  wire [1:0] _T_834; // @[Mux.scala 46:16:@99.4]
  wire  _T_835; // @[Mux.scala 46:19:@100.4]
  wire [1:0] _T_836; // @[Mux.scala 46:16:@101.4]
  wire  _T_837; // @[Mux.scala 46:19:@102.4]
  wire [1:0] _T_838; // @[Mux.scala 46:16:@103.4]
  wire  _GEN_129; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  wire  _GEN_130; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  wire  _GEN_131; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  wire  _GEN_132; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  wire  _GEN_133; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  wire  _GEN_134; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  wire  _GEN_135; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  wire  _GEN_137; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  wire  _GEN_138; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  wire  _GEN_139; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  wire  _GEN_140; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  wire  _GEN_141; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  wire  _GEN_142; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  wire  _GEN_143; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  wire [1:0] _T_842; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  wire  _T_843; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@105.4]
  wire [1:0] _T_845; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@106.4]
  wire  _T_847; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@107.4]
  wire  _T_848; // @[Mux.scala 46:19:@108.4]
  wire  _T_849; // @[Mux.scala 46:16:@109.4]
  wire  _T_850; // @[Mux.scala 46:19:@110.4]
  wire [1:0] _T_851; // @[Mux.scala 46:16:@111.4]
  wire  _T_852; // @[Mux.scala 46:19:@112.4]
  wire [1:0] _T_853; // @[Mux.scala 46:16:@113.4]
  wire  _T_854; // @[Mux.scala 46:19:@114.4]
  wire [1:0] _T_855; // @[Mux.scala 46:16:@115.4]
  wire  _GEN_145; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  wire  _GEN_146; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  wire  _GEN_147; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  wire  _GEN_148; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  wire  _GEN_149; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  wire  _GEN_150; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  wire  _GEN_151; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  wire  _GEN_153; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  wire  _GEN_154; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  wire  _GEN_155; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  wire  _GEN_156; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  wire  _GEN_157; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  wire  _GEN_158; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  wire  _GEN_159; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  wire [1:0] _T_859; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  wire  _T_860; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@117.4]
  wire [1:0] _T_862; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@118.4]
  wire  _T_864; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@119.4]
  wire  _T_865; // @[Mux.scala 46:19:@120.4]
  wire  _T_866; // @[Mux.scala 46:16:@121.4]
  wire  _T_867; // @[Mux.scala 46:19:@122.4]
  wire [1:0] _T_868; // @[Mux.scala 46:16:@123.4]
  wire  _T_869; // @[Mux.scala 46:19:@124.4]
  wire [1:0] _T_870; // @[Mux.scala 46:16:@125.4]
  wire  _T_871; // @[Mux.scala 46:19:@126.4]
  wire [1:0] _T_872; // @[Mux.scala 46:16:@127.4]
  wire  _GEN_161; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  wire  _GEN_162; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  wire  _GEN_163; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  wire  _GEN_164; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  wire  _GEN_165; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  wire  _GEN_166; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  wire  _GEN_167; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  wire  _GEN_169; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  wire  _GEN_170; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  wire  _GEN_171; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  wire  _GEN_172; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  wire  _GEN_173; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  wire  _GEN_174; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  wire  _GEN_175; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  wire [1:0] _T_876; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  wire  _T_877; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@129.4]
  wire [1:0] _T_879; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@130.4]
  wire  _T_881; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@131.4]
  wire  _T_882; // @[Mux.scala 46:19:@132.4]
  wire  _T_883; // @[Mux.scala 46:16:@133.4]
  wire  _T_884; // @[Mux.scala 46:19:@134.4]
  wire [1:0] _T_885; // @[Mux.scala 46:16:@135.4]
  wire  _T_886; // @[Mux.scala 46:19:@136.4]
  wire [1:0] _T_887; // @[Mux.scala 46:16:@137.4]
  wire  _T_888; // @[Mux.scala 46:19:@138.4]
  wire [1:0] _T_889; // @[Mux.scala 46:16:@139.4]
  wire  _GEN_177; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  wire  _GEN_178; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  wire  _GEN_179; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  wire  _GEN_180; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  wire  _GEN_181; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  wire  _GEN_182; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  wire  _GEN_183; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  wire  _GEN_185; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  wire  _GEN_186; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  wire  _GEN_187; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  wire  _GEN_188; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  wire  _GEN_189; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  wire  _GEN_190; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  wire  _GEN_191; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  wire [1:0] _T_893; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  wire  _T_894; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@141.4]
  wire [1:0] _T_896; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@142.4]
  wire  _T_898; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@143.4]
  wire  _T_899; // @[Mux.scala 46:19:@144.4]
  wire  _T_900; // @[Mux.scala 46:16:@145.4]
  wire  _T_901; // @[Mux.scala 46:19:@146.4]
  wire [1:0] _T_902; // @[Mux.scala 46:16:@147.4]
  wire  _T_903; // @[Mux.scala 46:19:@148.4]
  wire [1:0] _T_904; // @[Mux.scala 46:16:@149.4]
  wire  _T_905; // @[Mux.scala 46:19:@150.4]
  wire [1:0] _T_906; // @[Mux.scala 46:16:@151.4]
  wire  _GEN_193; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  wire  _GEN_194; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  wire  _GEN_195; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  wire  _GEN_196; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  wire  _GEN_197; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  wire  _GEN_198; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  wire  _GEN_199; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  wire  _GEN_201; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  wire  _GEN_202; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  wire  _GEN_203; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  wire  _GEN_204; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  wire  _GEN_205; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  wire  _GEN_206; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  wire  _GEN_207; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  wire [1:0] _T_910; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  wire  _T_911; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@153.4]
  wire [1:0] _T_913; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@154.4]
  wire  _T_915; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@155.4]
  wire  _T_916; // @[Mux.scala 46:19:@156.4]
  wire  _T_917; // @[Mux.scala 46:16:@157.4]
  wire  _T_918; // @[Mux.scala 46:19:@158.4]
  wire [1:0] _T_919; // @[Mux.scala 46:16:@159.4]
  wire  _T_920; // @[Mux.scala 46:19:@160.4]
  wire [1:0] _T_921; // @[Mux.scala 46:16:@161.4]
  wire  _T_922; // @[Mux.scala 46:19:@162.4]
  wire [1:0] _T_923; // @[Mux.scala 46:16:@163.4]
  wire  _GEN_209; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  wire  _GEN_210; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  wire  _GEN_211; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  wire  _GEN_212; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  wire  _GEN_213; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  wire  _GEN_214; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  wire  _GEN_215; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  wire  _GEN_217; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  wire  _GEN_218; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  wire  _GEN_219; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  wire  _GEN_220; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  wire  _GEN_221; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  wire  _GEN_222; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  wire  _GEN_223; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  wire [1:0] _T_927; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  wire  _T_928; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@165.4]
  wire [1:0] _T_930; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@166.4]
  wire  _T_932; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@167.4]
  wire  _T_933; // @[Mux.scala 46:19:@168.4]
  wire  _T_934; // @[Mux.scala 46:16:@169.4]
  wire  _T_935; // @[Mux.scala 46:19:@170.4]
  wire [1:0] _T_936; // @[Mux.scala 46:16:@171.4]
  wire  _T_937; // @[Mux.scala 46:19:@172.4]
  wire [1:0] _T_938; // @[Mux.scala 46:16:@173.4]
  wire  _T_939; // @[Mux.scala 46:19:@174.4]
  wire [1:0] _T_940; // @[Mux.scala 46:16:@175.4]
  wire  _GEN_225; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  wire  _GEN_226; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  wire  _GEN_227; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  wire  _GEN_228; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  wire  _GEN_229; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  wire  _GEN_230; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  wire  _GEN_231; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  wire  _GEN_233; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  wire  _GEN_234; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  wire  _GEN_235; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  wire  _GEN_236; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  wire  _GEN_237; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  wire  _GEN_238; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  wire  _GEN_239; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  wire [1:0] _T_944; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  wire  _T_945; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@177.4]
  wire [1:0] _T_947; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@178.4]
  wire  _T_949; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@179.4]
  wire  _T_950; // @[Mux.scala 46:19:@180.4]
  wire  _T_951; // @[Mux.scala 46:16:@181.4]
  wire  _T_952; // @[Mux.scala 46:19:@182.4]
  wire [1:0] _T_953; // @[Mux.scala 46:16:@183.4]
  wire  _T_954; // @[Mux.scala 46:19:@184.4]
  wire [1:0] _T_955; // @[Mux.scala 46:16:@185.4]
  wire  _T_956; // @[Mux.scala 46:19:@186.4]
  wire [1:0] _T_957; // @[Mux.scala 46:16:@187.4]
  wire  _GEN_241; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  wire  _GEN_242; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  wire  _GEN_243; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  wire  _GEN_244; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  wire  _GEN_245; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  wire  _GEN_246; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  wire  _GEN_247; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  wire  _GEN_249; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  wire  _GEN_250; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  wire  _GEN_251; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  wire  _GEN_252; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  wire  _GEN_253; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  wire  _GEN_254; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  wire  _GEN_255; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  wire [1:0] _T_961; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  wire  _T_962; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@189.4]
  wire [1:0] _T_964; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@190.4]
  wire  _T_966; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@191.4]
  wire  _T_967; // @[Mux.scala 46:19:@192.4]
  wire  _T_968; // @[Mux.scala 46:16:@193.4]
  wire  _T_969; // @[Mux.scala 46:19:@194.4]
  wire [1:0] _T_970; // @[Mux.scala 46:16:@195.4]
  wire  _T_971; // @[Mux.scala 46:19:@196.4]
  wire [1:0] _T_972; // @[Mux.scala 46:16:@197.4]
  wire  _T_973; // @[Mux.scala 46:19:@198.4]
  wire [1:0] _T_974; // @[Mux.scala 46:16:@199.4]
  assign _GEN_1 = 3'h1 == io_selects_0_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_2 = 3'h2 == io_selects_0_0 ? io_inputs_2 : _GEN_1; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_3 = 3'h3 == io_selects_0_0 ? io_inputs_3 : _GEN_2; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_4 = 3'h4 == io_selects_0_0 ? io_inputs_4 : _GEN_3; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_5 = 3'h5 == io_selects_0_0 ? io_inputs_5 : _GEN_4; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_6 = 3'h6 == io_selects_0_0 ? io_inputs_6 : _GEN_5; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_7 = 3'h7 == io_selects_0_0 ? io_inputs_7 : _GEN_6; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_9 = 3'h1 == io_selects_0_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_10 = 3'h2 == io_selects_0_1 ? io_inputs_2 : _GEN_9; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_11 = 3'h3 == io_selects_0_1 ? io_inputs_3 : _GEN_10; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_12 = 3'h4 == io_selects_0_1 ? io_inputs_4 : _GEN_11; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_13 = 3'h5 == io_selects_0_1 ? io_inputs_5 : _GEN_12; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_14 = 3'h6 == io_selects_0_1 ? io_inputs_6 : _GEN_13; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_15 = 3'h7 == io_selects_0_1 ? io_inputs_7 : _GEN_14; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  assign _T_706 = _GEN_7 + _GEN_15; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@8.4]
  assign _T_707 = _GEN_7 + _GEN_15; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@9.4]
  assign _T_709 = _GEN_7 * _GEN_15; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@10.4]
  assign _T_711 = _GEN_7 / _GEN_15; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@11.4]
  assign _T_712 = 3'h3 == io_operation_0; // @[Mux.scala 46:19:@12.4]
  assign _T_713 = _T_712 ? _T_711 : 1'h0; // @[Mux.scala 46:16:@13.4]
  assign _T_714 = 3'h2 == io_operation_0; // @[Mux.scala 46:19:@14.4]
  assign _T_715 = _T_714 ? _T_709 : {{1'd0}, _T_713}; // @[Mux.scala 46:16:@15.4]
  assign _T_716 = 3'h1 == io_operation_0; // @[Mux.scala 46:19:@16.4]
  assign _T_717 = _T_716 ? {{1'd0}, _T_707} : _T_715; // @[Mux.scala 46:16:@17.4]
  assign _T_718 = 3'h0 == io_operation_0; // @[Mux.scala 46:19:@18.4]
  assign _T_719 = _T_718 ? {{1'd0}, _GEN_7} : _T_717; // @[Mux.scala 46:16:@19.4]
  assign _GEN_17 = 3'h1 == io_selects_1_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_18 = 3'h2 == io_selects_1_0 ? io_inputs_2 : _GEN_17; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_19 = 3'h3 == io_selects_1_0 ? io_inputs_3 : _GEN_18; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_20 = 3'h4 == io_selects_1_0 ? io_inputs_4 : _GEN_19; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_21 = 3'h5 == io_selects_1_0 ? io_inputs_5 : _GEN_20; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_22 = 3'h6 == io_selects_1_0 ? io_inputs_6 : _GEN_21; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_23 = 3'h7 == io_selects_1_0 ? io_inputs_7 : _GEN_22; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_25 = 3'h1 == io_selects_1_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_26 = 3'h2 == io_selects_1_1 ? io_inputs_2 : _GEN_25; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_27 = 3'h3 == io_selects_1_1 ? io_inputs_3 : _GEN_26; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_28 = 3'h4 == io_selects_1_1 ? io_inputs_4 : _GEN_27; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_29 = 3'h5 == io_selects_1_1 ? io_inputs_5 : _GEN_28; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_30 = 3'h6 == io_selects_1_1 ? io_inputs_6 : _GEN_29; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_31 = 3'h7 == io_selects_1_1 ? io_inputs_7 : _GEN_30; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  assign _T_723 = _GEN_23 + _GEN_31; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@20.4]
  assign _T_724 = _GEN_23 + _GEN_31; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@21.4]
  assign _T_726 = _GEN_23 * _GEN_31; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@22.4]
  assign _T_728 = _GEN_23 / _GEN_31; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@23.4]
  assign _T_729 = 3'h3 == io_operation_1; // @[Mux.scala 46:19:@24.4]
  assign _T_730 = _T_729 ? _T_728 : 1'h0; // @[Mux.scala 46:16:@25.4]
  assign _T_731 = 3'h2 == io_operation_1; // @[Mux.scala 46:19:@26.4]
  assign _T_732 = _T_731 ? _T_726 : {{1'd0}, _T_730}; // @[Mux.scala 46:16:@27.4]
  assign _T_733 = 3'h1 == io_operation_1; // @[Mux.scala 46:19:@28.4]
  assign _T_734 = _T_733 ? {{1'd0}, _T_724} : _T_732; // @[Mux.scala 46:16:@29.4]
  assign _T_735 = 3'h0 == io_operation_1; // @[Mux.scala 46:19:@30.4]
  assign _T_736 = _T_735 ? {{1'd0}, _GEN_23} : _T_734; // @[Mux.scala 46:16:@31.4]
  assign _GEN_33 = 3'h1 == io_selects_2_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_34 = 3'h2 == io_selects_2_0 ? io_inputs_2 : _GEN_33; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_35 = 3'h3 == io_selects_2_0 ? io_inputs_3 : _GEN_34; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_36 = 3'h4 == io_selects_2_0 ? io_inputs_4 : _GEN_35; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_37 = 3'h5 == io_selects_2_0 ? io_inputs_5 : _GEN_36; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_38 = 3'h6 == io_selects_2_0 ? io_inputs_6 : _GEN_37; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_39 = 3'h7 == io_selects_2_0 ? io_inputs_7 : _GEN_38; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_41 = 3'h1 == io_selects_2_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_42 = 3'h2 == io_selects_2_1 ? io_inputs_2 : _GEN_41; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_43 = 3'h3 == io_selects_2_1 ? io_inputs_3 : _GEN_42; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_44 = 3'h4 == io_selects_2_1 ? io_inputs_4 : _GEN_43; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_45 = 3'h5 == io_selects_2_1 ? io_inputs_5 : _GEN_44; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_46 = 3'h6 == io_selects_2_1 ? io_inputs_6 : _GEN_45; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_47 = 3'h7 == io_selects_2_1 ? io_inputs_7 : _GEN_46; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  assign _T_740 = _GEN_39 + _GEN_47; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@32.4]
  assign _T_741 = _GEN_39 + _GEN_47; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@33.4]
  assign _T_743 = _GEN_39 * _GEN_47; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@34.4]
  assign _T_745 = _GEN_39 / _GEN_47; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@35.4]
  assign _T_746 = 3'h3 == io_operation_2; // @[Mux.scala 46:19:@36.4]
  assign _T_747 = _T_746 ? _T_745 : 1'h0; // @[Mux.scala 46:16:@37.4]
  assign _T_748 = 3'h2 == io_operation_2; // @[Mux.scala 46:19:@38.4]
  assign _T_749 = _T_748 ? _T_743 : {{1'd0}, _T_747}; // @[Mux.scala 46:16:@39.4]
  assign _T_750 = 3'h1 == io_operation_2; // @[Mux.scala 46:19:@40.4]
  assign _T_751 = _T_750 ? {{1'd0}, _T_741} : _T_749; // @[Mux.scala 46:16:@41.4]
  assign _T_752 = 3'h0 == io_operation_2; // @[Mux.scala 46:19:@42.4]
  assign _T_753 = _T_752 ? {{1'd0}, _GEN_39} : _T_751; // @[Mux.scala 46:16:@43.4]
  assign _GEN_49 = 3'h1 == io_selects_3_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_50 = 3'h2 == io_selects_3_0 ? io_inputs_2 : _GEN_49; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_51 = 3'h3 == io_selects_3_0 ? io_inputs_3 : _GEN_50; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_52 = 3'h4 == io_selects_3_0 ? io_inputs_4 : _GEN_51; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_53 = 3'h5 == io_selects_3_0 ? io_inputs_5 : _GEN_52; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_54 = 3'h6 == io_selects_3_0 ? io_inputs_6 : _GEN_53; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_55 = 3'h7 == io_selects_3_0 ? io_inputs_7 : _GEN_54; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_57 = 3'h1 == io_selects_3_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_58 = 3'h2 == io_selects_3_1 ? io_inputs_2 : _GEN_57; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_59 = 3'h3 == io_selects_3_1 ? io_inputs_3 : _GEN_58; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_60 = 3'h4 == io_selects_3_1 ? io_inputs_4 : _GEN_59; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_61 = 3'h5 == io_selects_3_1 ? io_inputs_5 : _GEN_60; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_62 = 3'h6 == io_selects_3_1 ? io_inputs_6 : _GEN_61; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_63 = 3'h7 == io_selects_3_1 ? io_inputs_7 : _GEN_62; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  assign _T_757 = _GEN_55 + _GEN_63; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@44.4]
  assign _T_758 = _GEN_55 + _GEN_63; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@45.4]
  assign _T_760 = _GEN_55 * _GEN_63; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@46.4]
  assign _T_762 = _GEN_55 / _GEN_63; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@47.4]
  assign _T_763 = 3'h3 == io_operation_3; // @[Mux.scala 46:19:@48.4]
  assign _T_764 = _T_763 ? _T_762 : 1'h0; // @[Mux.scala 46:16:@49.4]
  assign _T_765 = 3'h2 == io_operation_3; // @[Mux.scala 46:19:@50.4]
  assign _T_766 = _T_765 ? _T_760 : {{1'd0}, _T_764}; // @[Mux.scala 46:16:@51.4]
  assign _T_767 = 3'h1 == io_operation_3; // @[Mux.scala 46:19:@52.4]
  assign _T_768 = _T_767 ? {{1'd0}, _T_758} : _T_766; // @[Mux.scala 46:16:@53.4]
  assign _T_769 = 3'h0 == io_operation_3; // @[Mux.scala 46:19:@54.4]
  assign _T_770 = _T_769 ? {{1'd0}, _GEN_55} : _T_768; // @[Mux.scala 46:16:@55.4]
  assign _GEN_65 = 3'h1 == io_selects_4_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_66 = 3'h2 == io_selects_4_0 ? io_inputs_2 : _GEN_65; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_67 = 3'h3 == io_selects_4_0 ? io_inputs_3 : _GEN_66; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_68 = 3'h4 == io_selects_4_0 ? io_inputs_4 : _GEN_67; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_69 = 3'h5 == io_selects_4_0 ? io_inputs_5 : _GEN_68; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_70 = 3'h6 == io_selects_4_0 ? io_inputs_6 : _GEN_69; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_71 = 3'h7 == io_selects_4_0 ? io_inputs_7 : _GEN_70; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_73 = 3'h1 == io_selects_4_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_74 = 3'h2 == io_selects_4_1 ? io_inputs_2 : _GEN_73; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_75 = 3'h3 == io_selects_4_1 ? io_inputs_3 : _GEN_74; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_76 = 3'h4 == io_selects_4_1 ? io_inputs_4 : _GEN_75; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_77 = 3'h5 == io_selects_4_1 ? io_inputs_5 : _GEN_76; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_78 = 3'h6 == io_selects_4_1 ? io_inputs_6 : _GEN_77; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_79 = 3'h7 == io_selects_4_1 ? io_inputs_7 : _GEN_78; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  assign _T_774 = _GEN_71 + _GEN_79; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@56.4]
  assign _T_775 = _GEN_71 + _GEN_79; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@57.4]
  assign _T_777 = _GEN_71 * _GEN_79; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@58.4]
  assign _T_779 = _GEN_71 / _GEN_79; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@59.4]
  assign _T_780 = 3'h3 == io_operation_4; // @[Mux.scala 46:19:@60.4]
  assign _T_781 = _T_780 ? _T_779 : 1'h0; // @[Mux.scala 46:16:@61.4]
  assign _T_782 = 3'h2 == io_operation_4; // @[Mux.scala 46:19:@62.4]
  assign _T_783 = _T_782 ? _T_777 : {{1'd0}, _T_781}; // @[Mux.scala 46:16:@63.4]
  assign _T_784 = 3'h1 == io_operation_4; // @[Mux.scala 46:19:@64.4]
  assign _T_785 = _T_784 ? {{1'd0}, _T_775} : _T_783; // @[Mux.scala 46:16:@65.4]
  assign _T_786 = 3'h0 == io_operation_4; // @[Mux.scala 46:19:@66.4]
  assign _T_787 = _T_786 ? {{1'd0}, _GEN_71} : _T_785; // @[Mux.scala 46:16:@67.4]
  assign _GEN_81 = 3'h1 == io_selects_5_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_82 = 3'h2 == io_selects_5_0 ? io_inputs_2 : _GEN_81; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_83 = 3'h3 == io_selects_5_0 ? io_inputs_3 : _GEN_82; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_84 = 3'h4 == io_selects_5_0 ? io_inputs_4 : _GEN_83; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_85 = 3'h5 == io_selects_5_0 ? io_inputs_5 : _GEN_84; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_86 = 3'h6 == io_selects_5_0 ? io_inputs_6 : _GEN_85; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_87 = 3'h7 == io_selects_5_0 ? io_inputs_7 : _GEN_86; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_89 = 3'h1 == io_selects_5_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_90 = 3'h2 == io_selects_5_1 ? io_inputs_2 : _GEN_89; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_91 = 3'h3 == io_selects_5_1 ? io_inputs_3 : _GEN_90; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_92 = 3'h4 == io_selects_5_1 ? io_inputs_4 : _GEN_91; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_93 = 3'h5 == io_selects_5_1 ? io_inputs_5 : _GEN_92; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_94 = 3'h6 == io_selects_5_1 ? io_inputs_6 : _GEN_93; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_95 = 3'h7 == io_selects_5_1 ? io_inputs_7 : _GEN_94; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  assign _T_791 = _GEN_87 + _GEN_95; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@68.4]
  assign _T_792 = _GEN_87 + _GEN_95; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@69.4]
  assign _T_794 = _GEN_87 * _GEN_95; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@70.4]
  assign _T_796 = _GEN_87 / _GEN_95; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@71.4]
  assign _T_797 = 3'h3 == io_operation_5; // @[Mux.scala 46:19:@72.4]
  assign _T_798 = _T_797 ? _T_796 : 1'h0; // @[Mux.scala 46:16:@73.4]
  assign _T_799 = 3'h2 == io_operation_5; // @[Mux.scala 46:19:@74.4]
  assign _T_800 = _T_799 ? _T_794 : {{1'd0}, _T_798}; // @[Mux.scala 46:16:@75.4]
  assign _T_801 = 3'h1 == io_operation_5; // @[Mux.scala 46:19:@76.4]
  assign _T_802 = _T_801 ? {{1'd0}, _T_792} : _T_800; // @[Mux.scala 46:16:@77.4]
  assign _T_803 = 3'h0 == io_operation_5; // @[Mux.scala 46:19:@78.4]
  assign _T_804 = _T_803 ? {{1'd0}, _GEN_87} : _T_802; // @[Mux.scala 46:16:@79.4]
  assign _GEN_97 = 3'h1 == io_selects_6_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_98 = 3'h2 == io_selects_6_0 ? io_inputs_2 : _GEN_97; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_99 = 3'h3 == io_selects_6_0 ? io_inputs_3 : _GEN_98; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_100 = 3'h4 == io_selects_6_0 ? io_inputs_4 : _GEN_99; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_101 = 3'h5 == io_selects_6_0 ? io_inputs_5 : _GEN_100; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_102 = 3'h6 == io_selects_6_0 ? io_inputs_6 : _GEN_101; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_103 = 3'h7 == io_selects_6_0 ? io_inputs_7 : _GEN_102; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_105 = 3'h1 == io_selects_6_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_106 = 3'h2 == io_selects_6_1 ? io_inputs_2 : _GEN_105; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_107 = 3'h3 == io_selects_6_1 ? io_inputs_3 : _GEN_106; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_108 = 3'h4 == io_selects_6_1 ? io_inputs_4 : _GEN_107; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_109 = 3'h5 == io_selects_6_1 ? io_inputs_5 : _GEN_108; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_110 = 3'h6 == io_selects_6_1 ? io_inputs_6 : _GEN_109; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_111 = 3'h7 == io_selects_6_1 ? io_inputs_7 : _GEN_110; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  assign _T_808 = _GEN_103 + _GEN_111; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@80.4]
  assign _T_809 = _GEN_103 + _GEN_111; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@81.4]
  assign _T_811 = _GEN_103 * _GEN_111; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@82.4]
  assign _T_813 = _GEN_103 / _GEN_111; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@83.4]
  assign _T_814 = 3'h3 == io_operation_6; // @[Mux.scala 46:19:@84.4]
  assign _T_815 = _T_814 ? _T_813 : 1'h0; // @[Mux.scala 46:16:@85.4]
  assign _T_816 = 3'h2 == io_operation_6; // @[Mux.scala 46:19:@86.4]
  assign _T_817 = _T_816 ? _T_811 : {{1'd0}, _T_815}; // @[Mux.scala 46:16:@87.4]
  assign _T_818 = 3'h1 == io_operation_6; // @[Mux.scala 46:19:@88.4]
  assign _T_819 = _T_818 ? {{1'd0}, _T_809} : _T_817; // @[Mux.scala 46:16:@89.4]
  assign _T_820 = 3'h0 == io_operation_6; // @[Mux.scala 46:19:@90.4]
  assign _T_821 = _T_820 ? {{1'd0}, _GEN_103} : _T_819; // @[Mux.scala 46:16:@91.4]
  assign _GEN_113 = 3'h1 == io_selects_7_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_114 = 3'h2 == io_selects_7_0 ? io_inputs_2 : _GEN_113; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_115 = 3'h3 == io_selects_7_0 ? io_inputs_3 : _GEN_114; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_116 = 3'h4 == io_selects_7_0 ? io_inputs_4 : _GEN_115; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_117 = 3'h5 == io_selects_7_0 ? io_inputs_5 : _GEN_116; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_118 = 3'h6 == io_selects_7_0 ? io_inputs_6 : _GEN_117; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_119 = 3'h7 == io_selects_7_0 ? io_inputs_7 : _GEN_118; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_121 = 3'h1 == io_selects_7_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_122 = 3'h2 == io_selects_7_1 ? io_inputs_2 : _GEN_121; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_123 = 3'h3 == io_selects_7_1 ? io_inputs_3 : _GEN_122; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_124 = 3'h4 == io_selects_7_1 ? io_inputs_4 : _GEN_123; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_125 = 3'h5 == io_selects_7_1 ? io_inputs_5 : _GEN_124; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_126 = 3'h6 == io_selects_7_1 ? io_inputs_6 : _GEN_125; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_127 = 3'h7 == io_selects_7_1 ? io_inputs_7 : _GEN_126; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  assign _T_825 = _GEN_119 + _GEN_127; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@92.4]
  assign _T_826 = _GEN_119 + _GEN_127; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@93.4]
  assign _T_828 = _GEN_119 * _GEN_127; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@94.4]
  assign _T_830 = _GEN_119 / _GEN_127; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@95.4]
  assign _T_831 = 3'h3 == io_operation_7; // @[Mux.scala 46:19:@96.4]
  assign _T_832 = _T_831 ? _T_830 : 1'h0; // @[Mux.scala 46:16:@97.4]
  assign _T_833 = 3'h2 == io_operation_7; // @[Mux.scala 46:19:@98.4]
  assign _T_834 = _T_833 ? _T_828 : {{1'd0}, _T_832}; // @[Mux.scala 46:16:@99.4]
  assign _T_835 = 3'h1 == io_operation_7; // @[Mux.scala 46:19:@100.4]
  assign _T_836 = _T_835 ? {{1'd0}, _T_826} : _T_834; // @[Mux.scala 46:16:@101.4]
  assign _T_837 = 3'h0 == io_operation_7; // @[Mux.scala 46:19:@102.4]
  assign _T_838 = _T_837 ? {{1'd0}, _GEN_119} : _T_836; // @[Mux.scala 46:16:@103.4]
  assign _GEN_129 = 3'h1 == io_selects_8_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  assign _GEN_130 = 3'h2 == io_selects_8_0 ? io_inputs_2 : _GEN_129; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  assign _GEN_131 = 3'h3 == io_selects_8_0 ? io_inputs_3 : _GEN_130; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  assign _GEN_132 = 3'h4 == io_selects_8_0 ? io_inputs_4 : _GEN_131; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  assign _GEN_133 = 3'h5 == io_selects_8_0 ? io_inputs_5 : _GEN_132; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  assign _GEN_134 = 3'h6 == io_selects_8_0 ? io_inputs_6 : _GEN_133; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  assign _GEN_135 = 3'h7 == io_selects_8_0 ? io_inputs_7 : _GEN_134; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  assign _GEN_137 = 3'h1 == io_selects_8_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  assign _GEN_138 = 3'h2 == io_selects_8_1 ? io_inputs_2 : _GEN_137; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  assign _GEN_139 = 3'h3 == io_selects_8_1 ? io_inputs_3 : _GEN_138; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  assign _GEN_140 = 3'h4 == io_selects_8_1 ? io_inputs_4 : _GEN_139; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  assign _GEN_141 = 3'h5 == io_selects_8_1 ? io_inputs_5 : _GEN_140; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  assign _GEN_142 = 3'h6 == io_selects_8_1 ? io_inputs_6 : _GEN_141; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  assign _GEN_143 = 3'h7 == io_selects_8_1 ? io_inputs_7 : _GEN_142; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  assign _T_842 = _GEN_135 + _GEN_143; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@104.4]
  assign _T_843 = _GEN_135 + _GEN_143; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@105.4]
  assign _T_845 = _GEN_135 * _GEN_143; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@106.4]
  assign _T_847 = _GEN_135 / _GEN_143; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@107.4]
  assign _T_848 = 3'h3 == io_operation_8; // @[Mux.scala 46:19:@108.4]
  assign _T_849 = _T_848 ? _T_847 : 1'h0; // @[Mux.scala 46:16:@109.4]
  assign _T_850 = 3'h2 == io_operation_8; // @[Mux.scala 46:19:@110.4]
  assign _T_851 = _T_850 ? _T_845 : {{1'd0}, _T_849}; // @[Mux.scala 46:16:@111.4]
  assign _T_852 = 3'h1 == io_operation_8; // @[Mux.scala 46:19:@112.4]
  assign _T_853 = _T_852 ? {{1'd0}, _T_843} : _T_851; // @[Mux.scala 46:16:@113.4]
  assign _T_854 = 3'h0 == io_operation_8; // @[Mux.scala 46:19:@114.4]
  assign _T_855 = _T_854 ? {{1'd0}, _GEN_135} : _T_853; // @[Mux.scala 46:16:@115.4]
  assign _GEN_145 = 3'h1 == io_selects_9_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  assign _GEN_146 = 3'h2 == io_selects_9_0 ? io_inputs_2 : _GEN_145; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  assign _GEN_147 = 3'h3 == io_selects_9_0 ? io_inputs_3 : _GEN_146; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  assign _GEN_148 = 3'h4 == io_selects_9_0 ? io_inputs_4 : _GEN_147; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  assign _GEN_149 = 3'h5 == io_selects_9_0 ? io_inputs_5 : _GEN_148; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  assign _GEN_150 = 3'h6 == io_selects_9_0 ? io_inputs_6 : _GEN_149; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  assign _GEN_151 = 3'h7 == io_selects_9_0 ? io_inputs_7 : _GEN_150; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  assign _GEN_153 = 3'h1 == io_selects_9_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  assign _GEN_154 = 3'h2 == io_selects_9_1 ? io_inputs_2 : _GEN_153; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  assign _GEN_155 = 3'h3 == io_selects_9_1 ? io_inputs_3 : _GEN_154; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  assign _GEN_156 = 3'h4 == io_selects_9_1 ? io_inputs_4 : _GEN_155; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  assign _GEN_157 = 3'h5 == io_selects_9_1 ? io_inputs_5 : _GEN_156; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  assign _GEN_158 = 3'h6 == io_selects_9_1 ? io_inputs_6 : _GEN_157; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  assign _GEN_159 = 3'h7 == io_selects_9_1 ? io_inputs_7 : _GEN_158; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  assign _T_859 = _GEN_151 + _GEN_159; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@116.4]
  assign _T_860 = _GEN_151 + _GEN_159; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@117.4]
  assign _T_862 = _GEN_151 * _GEN_159; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@118.4]
  assign _T_864 = _GEN_151 / _GEN_159; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@119.4]
  assign _T_865 = 3'h3 == io_operation_9; // @[Mux.scala 46:19:@120.4]
  assign _T_866 = _T_865 ? _T_864 : 1'h0; // @[Mux.scala 46:16:@121.4]
  assign _T_867 = 3'h2 == io_operation_9; // @[Mux.scala 46:19:@122.4]
  assign _T_868 = _T_867 ? _T_862 : {{1'd0}, _T_866}; // @[Mux.scala 46:16:@123.4]
  assign _T_869 = 3'h1 == io_operation_9; // @[Mux.scala 46:19:@124.4]
  assign _T_870 = _T_869 ? {{1'd0}, _T_860} : _T_868; // @[Mux.scala 46:16:@125.4]
  assign _T_871 = 3'h0 == io_operation_9; // @[Mux.scala 46:19:@126.4]
  assign _T_872 = _T_871 ? {{1'd0}, _GEN_151} : _T_870; // @[Mux.scala 46:16:@127.4]
  assign _GEN_161 = 3'h1 == io_selects_10_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  assign _GEN_162 = 3'h2 == io_selects_10_0 ? io_inputs_2 : _GEN_161; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  assign _GEN_163 = 3'h3 == io_selects_10_0 ? io_inputs_3 : _GEN_162; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  assign _GEN_164 = 3'h4 == io_selects_10_0 ? io_inputs_4 : _GEN_163; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  assign _GEN_165 = 3'h5 == io_selects_10_0 ? io_inputs_5 : _GEN_164; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  assign _GEN_166 = 3'h6 == io_selects_10_0 ? io_inputs_6 : _GEN_165; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  assign _GEN_167 = 3'h7 == io_selects_10_0 ? io_inputs_7 : _GEN_166; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  assign _GEN_169 = 3'h1 == io_selects_10_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  assign _GEN_170 = 3'h2 == io_selects_10_1 ? io_inputs_2 : _GEN_169; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  assign _GEN_171 = 3'h3 == io_selects_10_1 ? io_inputs_3 : _GEN_170; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  assign _GEN_172 = 3'h4 == io_selects_10_1 ? io_inputs_4 : _GEN_171; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  assign _GEN_173 = 3'h5 == io_selects_10_1 ? io_inputs_5 : _GEN_172; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  assign _GEN_174 = 3'h6 == io_selects_10_1 ? io_inputs_6 : _GEN_173; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  assign _GEN_175 = 3'h7 == io_selects_10_1 ? io_inputs_7 : _GEN_174; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  assign _T_876 = _GEN_167 + _GEN_175; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@128.4]
  assign _T_877 = _GEN_167 + _GEN_175; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@129.4]
  assign _T_879 = _GEN_167 * _GEN_175; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@130.4]
  assign _T_881 = _GEN_167 / _GEN_175; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@131.4]
  assign _T_882 = 3'h3 == io_operation_10; // @[Mux.scala 46:19:@132.4]
  assign _T_883 = _T_882 ? _T_881 : 1'h0; // @[Mux.scala 46:16:@133.4]
  assign _T_884 = 3'h2 == io_operation_10; // @[Mux.scala 46:19:@134.4]
  assign _T_885 = _T_884 ? _T_879 : {{1'd0}, _T_883}; // @[Mux.scala 46:16:@135.4]
  assign _T_886 = 3'h1 == io_operation_10; // @[Mux.scala 46:19:@136.4]
  assign _T_887 = _T_886 ? {{1'd0}, _T_877} : _T_885; // @[Mux.scala 46:16:@137.4]
  assign _T_888 = 3'h0 == io_operation_10; // @[Mux.scala 46:19:@138.4]
  assign _T_889 = _T_888 ? {{1'd0}, _GEN_167} : _T_887; // @[Mux.scala 46:16:@139.4]
  assign _GEN_177 = 3'h1 == io_selects_11_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  assign _GEN_178 = 3'h2 == io_selects_11_0 ? io_inputs_2 : _GEN_177; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  assign _GEN_179 = 3'h3 == io_selects_11_0 ? io_inputs_3 : _GEN_178; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  assign _GEN_180 = 3'h4 == io_selects_11_0 ? io_inputs_4 : _GEN_179; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  assign _GEN_181 = 3'h5 == io_selects_11_0 ? io_inputs_5 : _GEN_180; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  assign _GEN_182 = 3'h6 == io_selects_11_0 ? io_inputs_6 : _GEN_181; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  assign _GEN_183 = 3'h7 == io_selects_11_0 ? io_inputs_7 : _GEN_182; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  assign _GEN_185 = 3'h1 == io_selects_11_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  assign _GEN_186 = 3'h2 == io_selects_11_1 ? io_inputs_2 : _GEN_185; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  assign _GEN_187 = 3'h3 == io_selects_11_1 ? io_inputs_3 : _GEN_186; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  assign _GEN_188 = 3'h4 == io_selects_11_1 ? io_inputs_4 : _GEN_187; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  assign _GEN_189 = 3'h5 == io_selects_11_1 ? io_inputs_5 : _GEN_188; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  assign _GEN_190 = 3'h6 == io_selects_11_1 ? io_inputs_6 : _GEN_189; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  assign _GEN_191 = 3'h7 == io_selects_11_1 ? io_inputs_7 : _GEN_190; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  assign _T_893 = _GEN_183 + _GEN_191; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@140.4]
  assign _T_894 = _GEN_183 + _GEN_191; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@141.4]
  assign _T_896 = _GEN_183 * _GEN_191; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@142.4]
  assign _T_898 = _GEN_183 / _GEN_191; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@143.4]
  assign _T_899 = 3'h3 == io_operation_11; // @[Mux.scala 46:19:@144.4]
  assign _T_900 = _T_899 ? _T_898 : 1'h0; // @[Mux.scala 46:16:@145.4]
  assign _T_901 = 3'h2 == io_operation_11; // @[Mux.scala 46:19:@146.4]
  assign _T_902 = _T_901 ? _T_896 : {{1'd0}, _T_900}; // @[Mux.scala 46:16:@147.4]
  assign _T_903 = 3'h1 == io_operation_11; // @[Mux.scala 46:19:@148.4]
  assign _T_904 = _T_903 ? {{1'd0}, _T_894} : _T_902; // @[Mux.scala 46:16:@149.4]
  assign _T_905 = 3'h0 == io_operation_11; // @[Mux.scala 46:19:@150.4]
  assign _T_906 = _T_905 ? {{1'd0}, _GEN_183} : _T_904; // @[Mux.scala 46:16:@151.4]
  assign _GEN_193 = 3'h1 == io_selects_12_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  assign _GEN_194 = 3'h2 == io_selects_12_0 ? io_inputs_2 : _GEN_193; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  assign _GEN_195 = 3'h3 == io_selects_12_0 ? io_inputs_3 : _GEN_194; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  assign _GEN_196 = 3'h4 == io_selects_12_0 ? io_inputs_4 : _GEN_195; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  assign _GEN_197 = 3'h5 == io_selects_12_0 ? io_inputs_5 : _GEN_196; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  assign _GEN_198 = 3'h6 == io_selects_12_0 ? io_inputs_6 : _GEN_197; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  assign _GEN_199 = 3'h7 == io_selects_12_0 ? io_inputs_7 : _GEN_198; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  assign _GEN_201 = 3'h1 == io_selects_12_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  assign _GEN_202 = 3'h2 == io_selects_12_1 ? io_inputs_2 : _GEN_201; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  assign _GEN_203 = 3'h3 == io_selects_12_1 ? io_inputs_3 : _GEN_202; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  assign _GEN_204 = 3'h4 == io_selects_12_1 ? io_inputs_4 : _GEN_203; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  assign _GEN_205 = 3'h5 == io_selects_12_1 ? io_inputs_5 : _GEN_204; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  assign _GEN_206 = 3'h6 == io_selects_12_1 ? io_inputs_6 : _GEN_205; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  assign _GEN_207 = 3'h7 == io_selects_12_1 ? io_inputs_7 : _GEN_206; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  assign _T_910 = _GEN_199 + _GEN_207; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@152.4]
  assign _T_911 = _GEN_199 + _GEN_207; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@153.4]
  assign _T_913 = _GEN_199 * _GEN_207; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@154.4]
  assign _T_915 = _GEN_199 / _GEN_207; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@155.4]
  assign _T_916 = 3'h3 == io_operation_12; // @[Mux.scala 46:19:@156.4]
  assign _T_917 = _T_916 ? _T_915 : 1'h0; // @[Mux.scala 46:16:@157.4]
  assign _T_918 = 3'h2 == io_operation_12; // @[Mux.scala 46:19:@158.4]
  assign _T_919 = _T_918 ? _T_913 : {{1'd0}, _T_917}; // @[Mux.scala 46:16:@159.4]
  assign _T_920 = 3'h1 == io_operation_12; // @[Mux.scala 46:19:@160.4]
  assign _T_921 = _T_920 ? {{1'd0}, _T_911} : _T_919; // @[Mux.scala 46:16:@161.4]
  assign _T_922 = 3'h0 == io_operation_12; // @[Mux.scala 46:19:@162.4]
  assign _T_923 = _T_922 ? {{1'd0}, _GEN_199} : _T_921; // @[Mux.scala 46:16:@163.4]
  assign _GEN_209 = 3'h1 == io_selects_13_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  assign _GEN_210 = 3'h2 == io_selects_13_0 ? io_inputs_2 : _GEN_209; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  assign _GEN_211 = 3'h3 == io_selects_13_0 ? io_inputs_3 : _GEN_210; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  assign _GEN_212 = 3'h4 == io_selects_13_0 ? io_inputs_4 : _GEN_211; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  assign _GEN_213 = 3'h5 == io_selects_13_0 ? io_inputs_5 : _GEN_212; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  assign _GEN_214 = 3'h6 == io_selects_13_0 ? io_inputs_6 : _GEN_213; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  assign _GEN_215 = 3'h7 == io_selects_13_0 ? io_inputs_7 : _GEN_214; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  assign _GEN_217 = 3'h1 == io_selects_13_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  assign _GEN_218 = 3'h2 == io_selects_13_1 ? io_inputs_2 : _GEN_217; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  assign _GEN_219 = 3'h3 == io_selects_13_1 ? io_inputs_3 : _GEN_218; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  assign _GEN_220 = 3'h4 == io_selects_13_1 ? io_inputs_4 : _GEN_219; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  assign _GEN_221 = 3'h5 == io_selects_13_1 ? io_inputs_5 : _GEN_220; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  assign _GEN_222 = 3'h6 == io_selects_13_1 ? io_inputs_6 : _GEN_221; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  assign _GEN_223 = 3'h7 == io_selects_13_1 ? io_inputs_7 : _GEN_222; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  assign _T_927 = _GEN_215 + _GEN_223; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@164.4]
  assign _T_928 = _GEN_215 + _GEN_223; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@165.4]
  assign _T_930 = _GEN_215 * _GEN_223; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@166.4]
  assign _T_932 = _GEN_215 / _GEN_223; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@167.4]
  assign _T_933 = 3'h3 == io_operation_13; // @[Mux.scala 46:19:@168.4]
  assign _T_934 = _T_933 ? _T_932 : 1'h0; // @[Mux.scala 46:16:@169.4]
  assign _T_935 = 3'h2 == io_operation_13; // @[Mux.scala 46:19:@170.4]
  assign _T_936 = _T_935 ? _T_930 : {{1'd0}, _T_934}; // @[Mux.scala 46:16:@171.4]
  assign _T_937 = 3'h1 == io_operation_13; // @[Mux.scala 46:19:@172.4]
  assign _T_938 = _T_937 ? {{1'd0}, _T_928} : _T_936; // @[Mux.scala 46:16:@173.4]
  assign _T_939 = 3'h0 == io_operation_13; // @[Mux.scala 46:19:@174.4]
  assign _T_940 = _T_939 ? {{1'd0}, _GEN_215} : _T_938; // @[Mux.scala 46:16:@175.4]
  assign _GEN_225 = 3'h1 == io_selects_14_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  assign _GEN_226 = 3'h2 == io_selects_14_0 ? io_inputs_2 : _GEN_225; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  assign _GEN_227 = 3'h3 == io_selects_14_0 ? io_inputs_3 : _GEN_226; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  assign _GEN_228 = 3'h4 == io_selects_14_0 ? io_inputs_4 : _GEN_227; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  assign _GEN_229 = 3'h5 == io_selects_14_0 ? io_inputs_5 : _GEN_228; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  assign _GEN_230 = 3'h6 == io_selects_14_0 ? io_inputs_6 : _GEN_229; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  assign _GEN_231 = 3'h7 == io_selects_14_0 ? io_inputs_7 : _GEN_230; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  assign _GEN_233 = 3'h1 == io_selects_14_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  assign _GEN_234 = 3'h2 == io_selects_14_1 ? io_inputs_2 : _GEN_233; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  assign _GEN_235 = 3'h3 == io_selects_14_1 ? io_inputs_3 : _GEN_234; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  assign _GEN_236 = 3'h4 == io_selects_14_1 ? io_inputs_4 : _GEN_235; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  assign _GEN_237 = 3'h5 == io_selects_14_1 ? io_inputs_5 : _GEN_236; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  assign _GEN_238 = 3'h6 == io_selects_14_1 ? io_inputs_6 : _GEN_237; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  assign _GEN_239 = 3'h7 == io_selects_14_1 ? io_inputs_7 : _GEN_238; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  assign _T_944 = _GEN_231 + _GEN_239; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@176.4]
  assign _T_945 = _GEN_231 + _GEN_239; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@177.4]
  assign _T_947 = _GEN_231 * _GEN_239; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@178.4]
  assign _T_949 = _GEN_231 / _GEN_239; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@179.4]
  assign _T_950 = 3'h3 == io_operation_14; // @[Mux.scala 46:19:@180.4]
  assign _T_951 = _T_950 ? _T_949 : 1'h0; // @[Mux.scala 46:16:@181.4]
  assign _T_952 = 3'h2 == io_operation_14; // @[Mux.scala 46:19:@182.4]
  assign _T_953 = _T_952 ? _T_947 : {{1'd0}, _T_951}; // @[Mux.scala 46:16:@183.4]
  assign _T_954 = 3'h1 == io_operation_14; // @[Mux.scala 46:19:@184.4]
  assign _T_955 = _T_954 ? {{1'd0}, _T_945} : _T_953; // @[Mux.scala 46:16:@185.4]
  assign _T_956 = 3'h0 == io_operation_14; // @[Mux.scala 46:19:@186.4]
  assign _T_957 = _T_956 ? {{1'd0}, _GEN_231} : _T_955; // @[Mux.scala 46:16:@187.4]
  assign _GEN_241 = 3'h1 == io_selects_15_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  assign _GEN_242 = 3'h2 == io_selects_15_0 ? io_inputs_2 : _GEN_241; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  assign _GEN_243 = 3'h3 == io_selects_15_0 ? io_inputs_3 : _GEN_242; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  assign _GEN_244 = 3'h4 == io_selects_15_0 ? io_inputs_4 : _GEN_243; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  assign _GEN_245 = 3'h5 == io_selects_15_0 ? io_inputs_5 : _GEN_244; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  assign _GEN_246 = 3'h6 == io_selects_15_0 ? io_inputs_6 : _GEN_245; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  assign _GEN_247 = 3'h7 == io_selects_15_0 ? io_inputs_7 : _GEN_246; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  assign _GEN_249 = 3'h1 == io_selects_15_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  assign _GEN_250 = 3'h2 == io_selects_15_1 ? io_inputs_2 : _GEN_249; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  assign _GEN_251 = 3'h3 == io_selects_15_1 ? io_inputs_3 : _GEN_250; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  assign _GEN_252 = 3'h4 == io_selects_15_1 ? io_inputs_4 : _GEN_251; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  assign _GEN_253 = 3'h5 == io_selects_15_1 ? io_inputs_5 : _GEN_252; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  assign _GEN_254 = 3'h6 == io_selects_15_1 ? io_inputs_6 : _GEN_253; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  assign _GEN_255 = 3'h7 == io_selects_15_1 ? io_inputs_7 : _GEN_254; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  assign _T_961 = _GEN_247 + _GEN_255; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@188.4]
  assign _T_962 = _GEN_247 + _GEN_255; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 32:53:@189.4]
  assign _T_964 = _GEN_247 * _GEN_255; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 33:58:@190.4]
  assign _T_966 = _GEN_247 / _GEN_255; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 34:56:@191.4]
  assign _T_967 = 3'h3 == io_operation_15; // @[Mux.scala 46:19:@192.4]
  assign _T_968 = _T_967 ? _T_966 : 1'h0; // @[Mux.scala 46:16:@193.4]
  assign _T_969 = 3'h2 == io_operation_15; // @[Mux.scala 46:19:@194.4]
  assign _T_970 = _T_969 ? _T_964 : {{1'd0}, _T_968}; // @[Mux.scala 46:16:@195.4]
  assign _T_971 = 3'h1 == io_operation_15; // @[Mux.scala 46:19:@196.4]
  assign _T_972 = _T_971 ? {{1'd0}, _T_962} : _T_970; // @[Mux.scala 46:16:@197.4]
  assign _T_973 = 3'h0 == io_operation_15; // @[Mux.scala 46:19:@198.4]
  assign _T_974 = _T_973 ? {{1'd0}, _GEN_247} : _T_972; // @[Mux.scala 46:16:@199.4]
  assign io_outputs_0 = _T_719[0]; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 23:14:@200.4]
  assign io_outputs_1 = _T_736[0]; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 23:14:@201.4]
  assign io_outputs_2 = _T_753[0]; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 23:14:@202.4]
  assign io_outputs_3 = _T_770[0]; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 23:14:@203.4]
  assign io_outputs_4 = _T_787[0]; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 23:14:@204.4]
  assign io_outputs_5 = _T_804[0]; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 23:14:@205.4]
  assign io_outputs_6 = _T_821[0]; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 23:14:@206.4]
  assign io_outputs_7 = _T_838[0]; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 23:14:@207.4]
  assign io_outputs_8 = _T_855[0]; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 23:14:@208.4]
  assign io_outputs_9 = _T_872[0]; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 23:14:@209.4]
  assign io_outputs_10 = _T_889[0]; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 23:14:@210.4]
  assign io_outputs_11 = _T_906[0]; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 23:14:@211.4]
  assign io_outputs_12 = _T_923[0]; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 23:14:@212.4]
  assign io_outputs_13 = _T_940[0]; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 23:14:@213.4]
  assign io_outputs_14 = _T_957[0]; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 23:14:@214.4]
  assign io_outputs_15 = _T_974[0]; // @[MuxTest_width_1_inputs_8_outputs_16_pipeline_0s.scala 23:14:@215.4]
endmodule
