VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS
MACRO memory4
  FOREIGN memory4 0 0 ;
  CLASS BLOCK ;
  SIZE 391.95 BY 235.97 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal7 ;
        RECT  2.94 202.7 339.34 204.1 ;
        RECT  2.94 162.7 339.34 164.1 ;
        RECT  2.94 122.7 339.34 124.1 ;
        RECT  2.94 82.7 339.34 84.1 ;
        RECT  2.94 42.7 339.34 44.1 ;
        RECT  2.94 2.7 339.34 4.1 ;
      LAYER metal4 ;
        RECT  339.04 1.33 339.24 233.87 ;
        RECT  283.04 1.33 283.24 233.87 ;
        RECT  227.04 1.33 227.24 233.87 ;
        RECT  171.04 1.33 171.24 233.87 ;
        RECT  115.04 1.33 115.24 233.87 ;
        RECT  59.04 1.33 59.24 233.87 ;
        RECT  3.04 1.33 3.24 233.87 ;
      LAYER metal1 ;
        RECT  1.14 233.75 390.83 233.85 ;
        RECT  1.14 230.95 390.83 231.05 ;
        RECT  1.14 228.15 390.83 228.25 ;
        RECT  1.14 225.35 390.83 225.45 ;
        RECT  1.14 222.55 390.83 222.65 ;
        RECT  1.14 219.75 390.83 219.85 ;
        RECT  1.14 216.95 390.83 217.05 ;
        RECT  1.14 214.15 390.83 214.25 ;
        RECT  1.14 211.35 390.83 211.45 ;
        RECT  1.14 208.55 390.83 208.65 ;
        RECT  1.14 205.75 390.83 205.85 ;
        RECT  1.14 202.95 390.83 203.05 ;
        RECT  1.14 200.15 390.83 200.25 ;
        RECT  1.14 197.35 390.83 197.45 ;
        RECT  1.14 194.55 390.83 194.65 ;
        RECT  1.14 191.75 390.83 191.85 ;
        RECT  1.14 188.95 390.83 189.05 ;
        RECT  1.14 186.15 390.83 186.25 ;
        RECT  1.14 183.35 390.83 183.45 ;
        RECT  1.14 180.55 390.83 180.65 ;
        RECT  1.14 177.75 390.83 177.85 ;
        RECT  1.14 174.95 390.83 175.05 ;
        RECT  1.14 172.15 390.83 172.25 ;
        RECT  1.14 169.35 390.83 169.45 ;
        RECT  1.14 166.55 390.83 166.65 ;
        RECT  1.14 163.75 390.83 163.85 ;
        RECT  1.14 160.95 390.83 161.05 ;
        RECT  1.14 158.15 390.83 158.25 ;
        RECT  1.14 155.35 390.83 155.45 ;
        RECT  1.14 152.55 390.83 152.65 ;
        RECT  1.14 149.75 390.83 149.85 ;
        RECT  1.14 146.95 390.83 147.05 ;
        RECT  1.14 144.15 390.83 144.25 ;
        RECT  1.14 141.35 390.83 141.45 ;
        RECT  1.14 138.55 390.83 138.65 ;
        RECT  1.14 135.75 390.83 135.85 ;
        RECT  1.14 132.95 390.83 133.05 ;
        RECT  1.14 130.15 390.83 130.25 ;
        RECT  1.14 127.35 390.83 127.45 ;
        RECT  1.14 124.55 390.83 124.65 ;
        RECT  1.14 121.75 390.83 121.85 ;
        RECT  1.14 118.95 390.83 119.05 ;
        RECT  1.14 116.15 390.83 116.25 ;
        RECT  1.14 113.35 390.83 113.45 ;
        RECT  1.14 110.55 390.83 110.65 ;
        RECT  1.14 107.75 390.83 107.85 ;
        RECT  1.14 104.95 390.83 105.05 ;
        RECT  1.14 102.15 390.83 102.25 ;
        RECT  1.14 99.35 390.83 99.45 ;
        RECT  1.14 96.55 390.83 96.65 ;
        RECT  1.14 93.75 390.83 93.85 ;
        RECT  1.14 90.95 390.83 91.05 ;
        RECT  1.14 88.15 390.83 88.25 ;
        RECT  1.14 85.35 390.83 85.45 ;
        RECT  1.14 82.55 390.83 82.65 ;
        RECT  1.14 79.75 390.83 79.85 ;
        RECT  1.14 76.95 390.83 77.05 ;
        RECT  1.14 74.15 390.83 74.25 ;
        RECT  1.14 71.35 390.83 71.45 ;
        RECT  1.14 68.55 390.83 68.65 ;
        RECT  1.14 65.75 390.83 65.85 ;
        RECT  1.14 62.95 390.83 63.05 ;
        RECT  1.14 60.15 390.83 60.25 ;
        RECT  1.14 57.35 390.83 57.45 ;
        RECT  1.14 54.55 390.83 54.65 ;
        RECT  1.14 51.75 390.83 51.85 ;
        RECT  1.14 48.95 390.83 49.05 ;
        RECT  1.14 46.15 390.83 46.25 ;
        RECT  1.14 43.35 390.83 43.45 ;
        RECT  1.14 40.55 390.83 40.65 ;
        RECT  1.14 37.75 390.83 37.85 ;
        RECT  1.14 34.95 390.83 35.05 ;
        RECT  1.14 32.15 390.83 32.25 ;
        RECT  1.14 29.35 390.83 29.45 ;
        RECT  1.14 26.55 390.83 26.65 ;
        RECT  1.14 23.75 390.83 23.85 ;
        RECT  1.14 20.95 390.83 21.05 ;
        RECT  1.14 18.15 390.83 18.25 ;
        RECT  1.14 15.35 390.83 15.45 ;
        RECT  1.14 12.55 390.83 12.65 ;
        RECT  1.14 9.75 390.83 9.85 ;
        RECT  1.14 6.95 390.83 7.05 ;
        RECT  1.14 4.15 390.83 4.25 ;
        RECT  1.14 1.35 390.83 1.45 ;
      VIA 339.14 203.4 via6_7_400_2800_4_1_600_600 ;
      VIA 339.14 203.4 via5_6_400_2800_5_1_600_600 ;
      VIA 339.14 203.4 via4_5_400_2800_5_1_600_600 ;
      VIA 339.14 163.4 via6_7_400_2800_4_1_600_600 ;
      VIA 339.14 163.4 via5_6_400_2800_5_1_600_600 ;
      VIA 339.14 163.4 via4_5_400_2800_5_1_600_600 ;
      VIA 339.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 339.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 339.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 339.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 339.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 339.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 339.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 339.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 339.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 339.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 339.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 339.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 203.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 203.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 203.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 163.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 163.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 163.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 203.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 203.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 203.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 163.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 163.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 163.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 203.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 203.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 203.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 163.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 163.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 163.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 203.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 203.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 203.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 163.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 163.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 163.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 203.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 203.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 203.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 163.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 163.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 163.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 203.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 203.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 203.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 163.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 163.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 163.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 339.14 233.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 233.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 233.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 231 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 231 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 231 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 228.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 228.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 228.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 225.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 225.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 225.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 222.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 222.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 222.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 219.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 219.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 219.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 217 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 217 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 217 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 214.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 214.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 214.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 211.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 211.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 211.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 208.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 208.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 208.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 205.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 205.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 205.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 203 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 203 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 203 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 200.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 200.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 200.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 197.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 197.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 197.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 194.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 194.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 194.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 191.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 191.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 191.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 189 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 189 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 189 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 186.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 186.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 186.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 183.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 183.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 183.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 180.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 180.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 180.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 177.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 177.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 177.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 175 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 175 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 175 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 172.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 172.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 172.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 169.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 169.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 169.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 166.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 166.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 166.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 163.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 163.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 163.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 161 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 161 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 161 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 158.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 158.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 158.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 155.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 155.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 155.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 152.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 152.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 152.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 149.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 149.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 149.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 147 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 147 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 147 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 144.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 144.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 144.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 141.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 141.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 141.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 138.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 138.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 138.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 1.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 233.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 233.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 233.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 231 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 231 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 231 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 228.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 228.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 228.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 225.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 225.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 225.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 222.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 222.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 222.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 219.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 219.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 219.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 217 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 217 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 217 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 214.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 214.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 214.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 211.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 211.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 211.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 208.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 208.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 208.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 205.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 205.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 205.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 203 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 203 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 203 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 200.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 200.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 200.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 197.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 197.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 197.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 194.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 194.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 194.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 191.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 191.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 191.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 189 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 189 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 189 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 186.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 186.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 186.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 183.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 183.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 183.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 180.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 180.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 180.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 177.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 177.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 177.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 175 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 175 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 175 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 172.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 172.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 172.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 169.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 169.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 169.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 166.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 166.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 166.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 163.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 163.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 163.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 161 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 161 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 161 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 158.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 158.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 158.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 155.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 155.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 155.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 152.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 152.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 152.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 149.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 149.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 149.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 147 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 147 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 147 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 144.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 144.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 144.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 141.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 141.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 141.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 138.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 138.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 138.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 1.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 233.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 233.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 233.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 231 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 231 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 231 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 228.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 228.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 228.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 225.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 225.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 225.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 222.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 222.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 222.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 219.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 219.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 219.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 217 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 217 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 217 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 214.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 214.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 214.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 211.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 211.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 211.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 208.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 208.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 208.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 205.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 205.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 205.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 203 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 203 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 203 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 200.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 200.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 200.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 197.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 197.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 197.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 194.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 194.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 194.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 191.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 191.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 191.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 189 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 189 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 189 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 186.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 186.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 186.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 183.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 183.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 183.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 180.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 180.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 180.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 177.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 177.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 177.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 175 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 175 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 175 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 172.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 172.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 172.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 169.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 169.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 169.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 166.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 166.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 166.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 163.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 163.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 163.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 161 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 161 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 161 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 158.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 158.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 158.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 155.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 155.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 155.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 152.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 152.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 152.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 149.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 149.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 149.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 147 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 147 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 147 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 144.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 144.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 144.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 141.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 141.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 141.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 138.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 138.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 138.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 1.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 233.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 233.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 233.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 231 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 231 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 231 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 228.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 228.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 228.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 225.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 225.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 225.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 222.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 222.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 222.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 219.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 219.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 219.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 217 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 217 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 217 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 214.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 214.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 214.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 211.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 211.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 211.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 208.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 208.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 208.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 205.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 205.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 205.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 203 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 203 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 203 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 200.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 200.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 200.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 197.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 197.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 197.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 194.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 194.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 194.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 191.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 191.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 191.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 189 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 189 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 189 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 186.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 186.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 186.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 183.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 183.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 183.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 180.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 180.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 180.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 177.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 177.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 177.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 175 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 175 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 175 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 172.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 172.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 172.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 169.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 169.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 169.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 166.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 166.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 166.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 163.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 163.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 163.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 161 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 161 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 161 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 158.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 158.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 158.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 155.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 155.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 155.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 152.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 152.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 152.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 149.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 149.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 149.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 147 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 147 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 147 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 144.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 144.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 144.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 141.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 141.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 141.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 138.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 138.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 138.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 1.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 233.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 233.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 233.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 231 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 231 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 231 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 228.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 228.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 228.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 225.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 225.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 225.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 222.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 222.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 222.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 219.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 219.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 219.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 217 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 217 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 217 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 214.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 214.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 214.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 211.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 211.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 211.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 208.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 208.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 208.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 205.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 205.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 205.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 203 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 203 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 203 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 200.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 200.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 200.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 197.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 197.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 197.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 194.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 194.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 194.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 191.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 191.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 191.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 189 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 189 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 189 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 186.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 186.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 186.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 183.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 183.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 183.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 180.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 180.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 180.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 177.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 177.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 177.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 175 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 175 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 175 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 172.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 172.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 172.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 169.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 169.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 169.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 166.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 166.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 166.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 163.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 163.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 163.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 161 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 161 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 161 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 158.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 158.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 158.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 155.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 155.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 155.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 152.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 152.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 152.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 149.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 149.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 149.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 147 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 147 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 147 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 144.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 144.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 144.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 141.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 141.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 141.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 138.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 138.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 138.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 1.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 233.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 233.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 233.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 231 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 231 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 231 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 228.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 228.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 228.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 225.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 225.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 225.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 222.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 222.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 222.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 219.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 219.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 219.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 217 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 217 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 217 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 214.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 214.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 214.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 211.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 211.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 211.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 208.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 208.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 208.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 205.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 205.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 205.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 203 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 203 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 203 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 200.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 200.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 200.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 197.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 197.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 197.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 194.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 194.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 194.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 191.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 191.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 191.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 189 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 189 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 189 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 186.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 186.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 186.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 183.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 183.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 183.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 180.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 180.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 180.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 177.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 177.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 177.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 175 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 175 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 175 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 172.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 172.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 172.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 169.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 169.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 169.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 166.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 166.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 166.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 163.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 163.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 163.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 161 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 161 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 161 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 158.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 158.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 158.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 155.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 155.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 155.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 152.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 152.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 152.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 149.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 149.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 149.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 147 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 147 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 147 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 144.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 144.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 144.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 141.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 141.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 141.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 138.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 138.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 138.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 1.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 233.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 233.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 233.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 231 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 231 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 231 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 228.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 228.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 228.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 225.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 225.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 225.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 222.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 222.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 222.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 219.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 219.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 219.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 217 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 217 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 217 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 214.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 214.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 214.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 211.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 211.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 211.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 208.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 208.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 208.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 205.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 205.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 205.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 203 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 203 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 203 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 200.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 200.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 200.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 197.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 197.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 197.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 194.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 194.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 194.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 191.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 191.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 191.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 189 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 189 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 189 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 186.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 186.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 186.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 183.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 183.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 183.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 180.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 180.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 180.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 177.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 177.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 177.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 175 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 175 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 175 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 172.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 172.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 172.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 169.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 169.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 169.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 166.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 166.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 166.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 163.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 163.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 163.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 161 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 161 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 161 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 158.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 158.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 158.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 155.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 155.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 155.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 152.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 152.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 152.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 149.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 149.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 149.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 147 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 147 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 147 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 144.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 144.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 144.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 141.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 141.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 141.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 138.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 138.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 138.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 1.4 via1_2_400_200_1_1_300_300 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal7 ;
        RECT  30.94 222.7 367.34 224.1 ;
        RECT  30.94 182.7 367.34 184.1 ;
        RECT  30.94 142.7 367.34 144.1 ;
        RECT  30.94 102.7 367.34 104.1 ;
        RECT  30.94 62.7 367.34 64.1 ;
        RECT  30.94 22.7 367.34 24.1 ;
      LAYER metal4 ;
        RECT  367.04 2.73 367.24 232.47 ;
        RECT  311.04 2.73 311.24 232.47 ;
        RECT  255.04 2.73 255.24 232.47 ;
        RECT  199.04 2.73 199.24 232.47 ;
        RECT  143.04 2.73 143.24 232.47 ;
        RECT  87.04 2.73 87.24 232.47 ;
        RECT  31.04 2.73 31.24 232.47 ;
      LAYER metal1 ;
        RECT  1.14 232.35 390.83 232.45 ;
        RECT  1.14 229.55 390.83 229.65 ;
        RECT  1.14 226.75 390.83 226.85 ;
        RECT  1.14 223.95 390.83 224.05 ;
        RECT  1.14 221.15 390.83 221.25 ;
        RECT  1.14 218.35 390.83 218.45 ;
        RECT  1.14 215.55 390.83 215.65 ;
        RECT  1.14 212.75 390.83 212.85 ;
        RECT  1.14 209.95 390.83 210.05 ;
        RECT  1.14 207.15 390.83 207.25 ;
        RECT  1.14 204.35 390.83 204.45 ;
        RECT  1.14 201.55 390.83 201.65 ;
        RECT  1.14 198.75 390.83 198.85 ;
        RECT  1.14 195.95 390.83 196.05 ;
        RECT  1.14 193.15 390.83 193.25 ;
        RECT  1.14 190.35 390.83 190.45 ;
        RECT  1.14 187.55 390.83 187.65 ;
        RECT  1.14 184.75 390.83 184.85 ;
        RECT  1.14 181.95 390.83 182.05 ;
        RECT  1.14 179.15 390.83 179.25 ;
        RECT  1.14 176.35 390.83 176.45 ;
        RECT  1.14 173.55 390.83 173.65 ;
        RECT  1.14 170.75 390.83 170.85 ;
        RECT  1.14 167.95 390.83 168.05 ;
        RECT  1.14 165.15 390.83 165.25 ;
        RECT  1.14 162.35 390.83 162.45 ;
        RECT  1.14 159.55 390.83 159.65 ;
        RECT  1.14 156.75 390.83 156.85 ;
        RECT  1.14 153.95 390.83 154.05 ;
        RECT  1.14 151.15 390.83 151.25 ;
        RECT  1.14 148.35 390.83 148.45 ;
        RECT  1.14 145.55 390.83 145.65 ;
        RECT  1.14 142.75 390.83 142.85 ;
        RECT  1.14 139.95 390.83 140.05 ;
        RECT  1.14 137.15 390.83 137.25 ;
        RECT  1.14 134.35 390.83 134.45 ;
        RECT  1.14 131.55 390.83 131.65 ;
        RECT  1.14 128.75 390.83 128.85 ;
        RECT  1.14 125.95 390.83 126.05 ;
        RECT  1.14 123.15 390.83 123.25 ;
        RECT  1.14 120.35 390.83 120.45 ;
        RECT  1.14 117.55 390.83 117.65 ;
        RECT  1.14 114.75 390.83 114.85 ;
        RECT  1.14 111.95 390.83 112.05 ;
        RECT  1.14 109.15 390.83 109.25 ;
        RECT  1.14 106.35 390.83 106.45 ;
        RECT  1.14 103.55 390.83 103.65 ;
        RECT  1.14 100.75 390.83 100.85 ;
        RECT  1.14 97.95 390.83 98.05 ;
        RECT  1.14 95.15 390.83 95.25 ;
        RECT  1.14 92.35 390.83 92.45 ;
        RECT  1.14 89.55 390.83 89.65 ;
        RECT  1.14 86.75 390.83 86.85 ;
        RECT  1.14 83.95 390.83 84.05 ;
        RECT  1.14 81.15 390.83 81.25 ;
        RECT  1.14 78.35 390.83 78.45 ;
        RECT  1.14 75.55 390.83 75.65 ;
        RECT  1.14 72.75 390.83 72.85 ;
        RECT  1.14 69.95 390.83 70.05 ;
        RECT  1.14 67.15 390.83 67.25 ;
        RECT  1.14 64.35 390.83 64.45 ;
        RECT  1.14 61.55 390.83 61.65 ;
        RECT  1.14 58.75 390.83 58.85 ;
        RECT  1.14 55.95 390.83 56.05 ;
        RECT  1.14 53.15 390.83 53.25 ;
        RECT  1.14 50.35 390.83 50.45 ;
        RECT  1.14 47.55 390.83 47.65 ;
        RECT  1.14 44.75 390.83 44.85 ;
        RECT  1.14 41.95 390.83 42.05 ;
        RECT  1.14 39.15 390.83 39.25 ;
        RECT  1.14 36.35 390.83 36.45 ;
        RECT  1.14 33.55 390.83 33.65 ;
        RECT  1.14 30.75 390.83 30.85 ;
        RECT  1.14 27.95 390.83 28.05 ;
        RECT  1.14 25.15 390.83 25.25 ;
        RECT  1.14 22.35 390.83 22.45 ;
        RECT  1.14 19.55 390.83 19.65 ;
        RECT  1.14 16.75 390.83 16.85 ;
        RECT  1.14 13.95 390.83 14.05 ;
        RECT  1.14 11.15 390.83 11.25 ;
        RECT  1.14 8.35 390.83 8.45 ;
        RECT  1.14 5.55 390.83 5.65 ;
        RECT  1.14 2.75 390.83 2.85 ;
      VIA 367.14 223.4 via6_7_400_2800_4_1_600_600 ;
      VIA 367.14 223.4 via5_6_400_2800_5_1_600_600 ;
      VIA 367.14 223.4 via4_5_400_2800_5_1_600_600 ;
      VIA 367.14 183.4 via6_7_400_2800_4_1_600_600 ;
      VIA 367.14 183.4 via5_6_400_2800_5_1_600_600 ;
      VIA 367.14 183.4 via4_5_400_2800_5_1_600_600 ;
      VIA 367.14 143.4 via6_7_400_2800_4_1_600_600 ;
      VIA 367.14 143.4 via5_6_400_2800_5_1_600_600 ;
      VIA 367.14 143.4 via4_5_400_2800_5_1_600_600 ;
      VIA 367.14 103.4 via6_7_400_2800_4_1_600_600 ;
      VIA 367.14 103.4 via5_6_400_2800_5_1_600_600 ;
      VIA 367.14 103.4 via4_5_400_2800_5_1_600_600 ;
      VIA 367.14 63.4 via6_7_400_2800_4_1_600_600 ;
      VIA 367.14 63.4 via5_6_400_2800_5_1_600_600 ;
      VIA 367.14 63.4 via4_5_400_2800_5_1_600_600 ;
      VIA 367.14 23.4 via6_7_400_2800_4_1_600_600 ;
      VIA 367.14 23.4 via5_6_400_2800_5_1_600_600 ;
      VIA 367.14 23.4 via4_5_400_2800_5_1_600_600 ;
      VIA 311.14 223.4 via6_7_400_2800_4_1_600_600 ;
      VIA 311.14 223.4 via5_6_400_2800_5_1_600_600 ;
      VIA 311.14 223.4 via4_5_400_2800_5_1_600_600 ;
      VIA 311.14 183.4 via6_7_400_2800_4_1_600_600 ;
      VIA 311.14 183.4 via5_6_400_2800_5_1_600_600 ;
      VIA 311.14 183.4 via4_5_400_2800_5_1_600_600 ;
      VIA 311.14 143.4 via6_7_400_2800_4_1_600_600 ;
      VIA 311.14 143.4 via5_6_400_2800_5_1_600_600 ;
      VIA 311.14 143.4 via4_5_400_2800_5_1_600_600 ;
      VIA 311.14 103.4 via6_7_400_2800_4_1_600_600 ;
      VIA 311.14 103.4 via5_6_400_2800_5_1_600_600 ;
      VIA 311.14 103.4 via4_5_400_2800_5_1_600_600 ;
      VIA 311.14 63.4 via6_7_400_2800_4_1_600_600 ;
      VIA 311.14 63.4 via5_6_400_2800_5_1_600_600 ;
      VIA 311.14 63.4 via4_5_400_2800_5_1_600_600 ;
      VIA 311.14 23.4 via6_7_400_2800_4_1_600_600 ;
      VIA 311.14 23.4 via5_6_400_2800_5_1_600_600 ;
      VIA 311.14 23.4 via4_5_400_2800_5_1_600_600 ;
      VIA 255.14 223.4 via6_7_400_2800_4_1_600_600 ;
      VIA 255.14 223.4 via5_6_400_2800_5_1_600_600 ;
      VIA 255.14 223.4 via4_5_400_2800_5_1_600_600 ;
      VIA 255.14 183.4 via6_7_400_2800_4_1_600_600 ;
      VIA 255.14 183.4 via5_6_400_2800_5_1_600_600 ;
      VIA 255.14 183.4 via4_5_400_2800_5_1_600_600 ;
      VIA 255.14 143.4 via6_7_400_2800_4_1_600_600 ;
      VIA 255.14 143.4 via5_6_400_2800_5_1_600_600 ;
      VIA 255.14 143.4 via4_5_400_2800_5_1_600_600 ;
      VIA 255.14 103.4 via6_7_400_2800_4_1_600_600 ;
      VIA 255.14 103.4 via5_6_400_2800_5_1_600_600 ;
      VIA 255.14 103.4 via4_5_400_2800_5_1_600_600 ;
      VIA 255.14 63.4 via6_7_400_2800_4_1_600_600 ;
      VIA 255.14 63.4 via5_6_400_2800_5_1_600_600 ;
      VIA 255.14 63.4 via4_5_400_2800_5_1_600_600 ;
      VIA 255.14 23.4 via6_7_400_2800_4_1_600_600 ;
      VIA 255.14 23.4 via5_6_400_2800_5_1_600_600 ;
      VIA 255.14 23.4 via4_5_400_2800_5_1_600_600 ;
      VIA 199.14 223.4 via6_7_400_2800_4_1_600_600 ;
      VIA 199.14 223.4 via5_6_400_2800_5_1_600_600 ;
      VIA 199.14 223.4 via4_5_400_2800_5_1_600_600 ;
      VIA 199.14 183.4 via6_7_400_2800_4_1_600_600 ;
      VIA 199.14 183.4 via5_6_400_2800_5_1_600_600 ;
      VIA 199.14 183.4 via4_5_400_2800_5_1_600_600 ;
      VIA 199.14 143.4 via6_7_400_2800_4_1_600_600 ;
      VIA 199.14 143.4 via5_6_400_2800_5_1_600_600 ;
      VIA 199.14 143.4 via4_5_400_2800_5_1_600_600 ;
      VIA 199.14 103.4 via6_7_400_2800_4_1_600_600 ;
      VIA 199.14 103.4 via5_6_400_2800_5_1_600_600 ;
      VIA 199.14 103.4 via4_5_400_2800_5_1_600_600 ;
      VIA 199.14 63.4 via6_7_400_2800_4_1_600_600 ;
      VIA 199.14 63.4 via5_6_400_2800_5_1_600_600 ;
      VIA 199.14 63.4 via4_5_400_2800_5_1_600_600 ;
      VIA 199.14 23.4 via6_7_400_2800_4_1_600_600 ;
      VIA 199.14 23.4 via5_6_400_2800_5_1_600_600 ;
      VIA 199.14 23.4 via4_5_400_2800_5_1_600_600 ;
      VIA 143.14 223.4 via6_7_400_2800_4_1_600_600 ;
      VIA 143.14 223.4 via5_6_400_2800_5_1_600_600 ;
      VIA 143.14 223.4 via4_5_400_2800_5_1_600_600 ;
      VIA 143.14 183.4 via6_7_400_2800_4_1_600_600 ;
      VIA 143.14 183.4 via5_6_400_2800_5_1_600_600 ;
      VIA 143.14 183.4 via4_5_400_2800_5_1_600_600 ;
      VIA 143.14 143.4 via6_7_400_2800_4_1_600_600 ;
      VIA 143.14 143.4 via5_6_400_2800_5_1_600_600 ;
      VIA 143.14 143.4 via4_5_400_2800_5_1_600_600 ;
      VIA 143.14 103.4 via6_7_400_2800_4_1_600_600 ;
      VIA 143.14 103.4 via5_6_400_2800_5_1_600_600 ;
      VIA 143.14 103.4 via4_5_400_2800_5_1_600_600 ;
      VIA 143.14 63.4 via6_7_400_2800_4_1_600_600 ;
      VIA 143.14 63.4 via5_6_400_2800_5_1_600_600 ;
      VIA 143.14 63.4 via4_5_400_2800_5_1_600_600 ;
      VIA 143.14 23.4 via6_7_400_2800_4_1_600_600 ;
      VIA 143.14 23.4 via5_6_400_2800_5_1_600_600 ;
      VIA 143.14 23.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 223.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 223.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 223.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 183.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 183.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 183.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 143.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 143.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 143.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 103.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 103.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 103.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 63.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 63.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 63.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 23.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 23.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 23.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 223.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 223.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 223.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 183.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 183.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 183.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 143.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 143.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 143.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 103.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 103.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 103.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 63.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 63.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 63.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 23.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 23.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 23.4 via4_5_400_2800_5_1_600_600 ;
      VIA 367.14 232.4 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 232.4 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 232.4 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 229.6 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 229.6 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 229.6 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 226.8 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 226.8 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 226.8 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 224 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 224 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 224 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 221.2 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 221.2 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 221.2 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 218.4 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 218.4 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 218.4 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 215.6 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 215.6 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 215.6 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 212.8 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 212.8 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 212.8 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 210 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 210 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 210 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 207.2 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 207.2 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 207.2 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 204.4 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 204.4 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 204.4 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 201.6 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 201.6 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 201.6 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 198.8 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 198.8 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 198.8 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 196 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 196 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 196 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 193.2 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 193.2 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 193.2 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 190.4 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 190.4 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 190.4 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 187.6 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 187.6 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 187.6 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 184.8 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 184.8 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 184.8 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 182 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 182 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 182 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 179.2 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 179.2 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 179.2 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 176.4 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 176.4 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 176.4 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 173.6 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 173.6 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 173.6 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 170.8 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 170.8 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 170.8 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 168 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 168 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 168 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 165.2 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 165.2 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 165.2 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 162.4 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 162.4 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 162.4 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 159.6 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 159.6 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 159.6 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 156.8 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 156.8 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 156.8 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 154 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 154 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 154 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 151.2 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 151.2 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 151.2 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 148.4 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 148.4 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 148.4 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 145.6 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 145.6 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 145.6 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 142.8 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 142.8 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 142.8 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 140 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 140 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 140 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 137.2 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 137.2 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 137.2 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 134.4 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 134.4 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 134.4 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 131.6 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 131.6 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 131.6 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 128.8 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 128.8 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 128.8 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 126 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 126 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 126 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 123.2 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 123.2 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 123.2 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 120.4 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 120.4 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 120.4 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 117.6 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 117.6 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 117.6 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 114.8 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 114.8 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 114.8 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 112 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 112 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 112 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 109.2 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 109.2 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 109.2 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 106.4 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 106.4 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 106.4 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 103.6 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 103.6 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 103.6 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 100.8 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 100.8 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 100.8 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 98 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 98 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 98 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 95.2 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 95.2 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 95.2 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 92.4 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 92.4 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 92.4 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 89.6 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 89.6 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 89.6 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 86.8 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 86.8 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 86.8 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 84 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 84 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 84 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 81.2 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 81.2 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 81.2 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 78.4 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 78.4 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 78.4 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 75.6 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 75.6 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 75.6 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 72.8 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 72.8 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 72.8 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 70 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 70 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 70 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 67.2 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 67.2 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 67.2 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 64.4 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 64.4 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 64.4 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 61.6 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 61.6 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 61.6 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 58.8 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 58.8 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 58.8 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 56 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 56 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 56 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 53.2 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 53.2 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 53.2 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 50.4 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 50.4 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 50.4 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 47.6 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 47.6 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 47.6 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 44.8 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 44.8 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 44.8 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 42 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 42 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 42 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 39.2 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 39.2 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 39.2 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 36.4 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 36.4 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 36.4 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 33.6 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 33.6 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 33.6 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 30.8 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 30.8 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 30.8 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 28 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 28 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 28 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 25.2 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 25.2 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 25.2 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 22.4 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 22.4 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 22.4 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 19.6 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 19.6 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 19.6 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 16.8 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 16.8 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 16.8 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 14 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 14 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 14 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 11.2 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 11.2 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 11.2 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 8.4 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 8.4 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 8.4 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 5.6 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 5.6 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 5.6 via1_2_400_200_1_1_300_300 ;
      VIA 367.14 2.8 via3_4_400_200_1_1_320_320 ;
      VIA 367.14 2.8 via2_3_400_200_1_1_320_320 ;
      VIA 367.14 2.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 232.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 232.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 232.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 229.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 229.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 229.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 226.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 226.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 226.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 224 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 224 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 224 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 221.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 221.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 221.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 218.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 218.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 218.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 215.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 215.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 215.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 212.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 212.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 212.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 210 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 210 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 210 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 207.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 207.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 207.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 204.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 204.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 204.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 201.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 201.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 201.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 198.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 198.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 198.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 196 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 196 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 196 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 193.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 193.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 193.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 190.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 190.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 190.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 187.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 187.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 187.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 184.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 184.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 184.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 182 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 182 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 182 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 179.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 179.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 179.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 176.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 176.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 176.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 173.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 173.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 173.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 170.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 170.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 170.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 168 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 168 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 168 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 165.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 165.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 165.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 162.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 162.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 162.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 159.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 159.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 159.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 156.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 156.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 156.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 154 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 154 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 154 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 151.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 151.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 151.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 148.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 148.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 148.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 145.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 145.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 145.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 142.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 142.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 142.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 140 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 140 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 140 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 137.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 137.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 137.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 134.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 134.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 134.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 131.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 131.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 131.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 128.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 128.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 128.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 126 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 126 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 126 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 123.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 123.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 123.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 120.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 120.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 120.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 117.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 117.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 117.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 114.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 114.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 114.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 112 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 112 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 112 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 109.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 109.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 109.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 106.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 106.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 106.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 103.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 103.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 103.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 100.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 100.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 100.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 98 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 98 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 98 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 95.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 95.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 95.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 92.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 92.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 92.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 89.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 89.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 89.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 86.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 86.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 86.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 84 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 84 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 84 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 81.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 81.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 81.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 78.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 78.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 78.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 75.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 75.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 75.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 72.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 72.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 72.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 70 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 70 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 70 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 67.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 67.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 67.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 64.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 64.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 64.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 61.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 61.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 61.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 58.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 58.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 58.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 56 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 56 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 56 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 53.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 53.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 53.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 50.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 50.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 50.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 47.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 47.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 47.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 44.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 44.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 44.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 42 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 42 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 42 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 39.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 39.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 39.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 36.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 36.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 36.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 33.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 33.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 33.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 30.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 30.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 30.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 28 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 28 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 28 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 25.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 25.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 25.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 22.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 22.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 22.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 19.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 19.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 19.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 16.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 16.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 16.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 14 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 14 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 14 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 11.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 11.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 11.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 8.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 8.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 8.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 5.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 5.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 5.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 2.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 2.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 2.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 232.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 232.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 232.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 229.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 229.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 229.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 226.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 226.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 226.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 224 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 224 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 224 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 221.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 221.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 221.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 218.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 218.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 218.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 215.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 215.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 215.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 212.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 212.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 212.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 210 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 210 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 210 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 207.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 207.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 207.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 204.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 204.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 204.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 201.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 201.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 201.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 198.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 198.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 198.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 196 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 196 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 196 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 193.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 193.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 193.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 190.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 190.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 190.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 187.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 187.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 187.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 184.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 184.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 184.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 182 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 182 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 182 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 179.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 179.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 179.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 176.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 176.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 176.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 173.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 173.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 173.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 170.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 170.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 170.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 168 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 168 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 168 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 165.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 165.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 165.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 162.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 162.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 162.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 159.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 159.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 159.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 156.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 156.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 156.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 154 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 154 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 154 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 151.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 151.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 151.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 148.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 148.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 148.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 145.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 145.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 145.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 142.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 142.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 142.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 140 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 140 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 140 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 137.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 137.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 137.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 134.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 134.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 134.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 131.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 131.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 131.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 128.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 128.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 128.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 126 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 126 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 126 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 123.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 123.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 123.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 120.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 120.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 120.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 117.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 117.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 117.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 114.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 114.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 114.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 112 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 112 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 112 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 109.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 109.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 109.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 106.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 106.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 106.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 103.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 103.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 103.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 100.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 100.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 100.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 98 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 98 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 98 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 95.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 95.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 95.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 92.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 92.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 92.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 89.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 89.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 89.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 86.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 86.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 86.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 84 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 84 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 84 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 81.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 81.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 81.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 78.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 78.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 78.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 75.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 75.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 75.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 72.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 72.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 72.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 70 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 70 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 70 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 67.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 67.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 67.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 64.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 64.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 64.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 61.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 61.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 61.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 58.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 58.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 58.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 56 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 56 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 56 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 53.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 53.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 53.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 50.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 50.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 50.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 47.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 47.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 47.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 44.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 44.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 44.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 42 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 42 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 42 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 39.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 39.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 39.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 36.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 36.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 36.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 33.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 33.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 33.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 30.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 30.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 30.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 28 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 28 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 28 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 25.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 25.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 25.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 22.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 22.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 22.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 19.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 19.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 19.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 16.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 16.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 16.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 14 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 14 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 14 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 11.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 11.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 11.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 8.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 8.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 8.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 5.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 5.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 5.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 2.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 2.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 2.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 232.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 232.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 232.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 229.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 229.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 229.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 226.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 226.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 226.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 224 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 224 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 224 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 221.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 221.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 221.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 218.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 218.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 218.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 215.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 215.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 215.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 212.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 212.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 212.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 210 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 210 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 210 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 207.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 207.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 207.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 204.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 204.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 204.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 201.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 201.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 201.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 198.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 198.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 198.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 196 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 196 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 196 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 193.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 193.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 193.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 190.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 190.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 190.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 187.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 187.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 187.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 184.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 184.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 184.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 182 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 182 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 182 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 179.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 179.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 179.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 176.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 176.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 176.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 173.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 173.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 173.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 170.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 170.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 170.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 168 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 168 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 168 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 165.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 165.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 165.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 162.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 162.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 162.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 159.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 159.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 159.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 156.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 156.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 156.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 154 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 154 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 154 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 151.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 151.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 151.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 148.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 148.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 148.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 145.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 145.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 145.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 142.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 142.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 142.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 140 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 140 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 140 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 137.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 137.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 137.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 134.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 134.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 134.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 131.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 131.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 131.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 128.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 128.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 128.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 126 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 126 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 126 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 123.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 123.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 123.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 120.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 120.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 120.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 117.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 117.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 117.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 114.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 114.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 114.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 112 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 112 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 112 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 109.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 109.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 109.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 106.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 106.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 106.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 103.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 103.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 103.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 100.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 100.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 100.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 98 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 98 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 98 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 95.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 95.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 95.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 92.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 92.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 92.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 89.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 89.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 89.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 86.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 86.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 86.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 84 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 84 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 84 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 81.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 81.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 81.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 78.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 78.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 78.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 75.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 75.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 75.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 72.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 72.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 72.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 70 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 70 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 70 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 67.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 67.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 67.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 64.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 64.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 64.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 61.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 61.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 61.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 58.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 58.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 58.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 56 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 56 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 56 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 53.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 53.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 53.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 50.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 50.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 50.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 47.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 47.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 47.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 44.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 44.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 44.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 42 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 42 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 42 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 39.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 39.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 39.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 36.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 36.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 36.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 33.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 33.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 33.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 30.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 30.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 30.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 28 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 28 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 28 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 25.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 25.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 25.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 22.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 22.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 22.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 19.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 19.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 19.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 16.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 16.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 16.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 14 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 14 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 14 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 11.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 11.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 11.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 8.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 8.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 8.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 5.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 5.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 5.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 2.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 2.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 2.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 232.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 232.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 232.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 229.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 229.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 229.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 226.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 226.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 226.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 224 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 224 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 224 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 221.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 221.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 221.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 218.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 218.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 218.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 215.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 215.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 215.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 212.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 212.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 212.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 210 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 210 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 210 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 207.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 207.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 207.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 204.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 204.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 204.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 201.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 201.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 201.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 198.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 198.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 198.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 196 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 196 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 196 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 193.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 193.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 193.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 190.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 190.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 190.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 187.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 187.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 187.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 184.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 184.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 184.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 182 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 182 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 182 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 179.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 179.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 179.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 176.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 176.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 176.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 173.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 173.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 173.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 170.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 170.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 170.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 168 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 168 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 168 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 165.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 165.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 165.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 162.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 162.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 162.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 159.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 159.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 159.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 156.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 156.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 156.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 154 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 154 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 154 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 151.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 151.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 151.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 148.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 148.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 148.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 145.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 145.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 145.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 142.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 142.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 142.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 140 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 140 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 140 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 137.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 137.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 137.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 134.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 134.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 134.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 131.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 131.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 131.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 128.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 128.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 128.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 126 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 126 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 126 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 123.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 123.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 123.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 120.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 120.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 120.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 117.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 117.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 117.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 114.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 114.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 114.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 112 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 112 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 112 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 109.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 109.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 109.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 106.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 106.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 106.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 103.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 103.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 103.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 100.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 100.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 100.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 98 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 98 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 98 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 95.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 95.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 95.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 92.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 92.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 92.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 89.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 89.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 89.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 86.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 86.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 86.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 84 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 84 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 84 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 81.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 81.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 81.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 78.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 78.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 78.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 75.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 75.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 75.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 72.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 72.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 72.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 70 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 70 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 70 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 67.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 67.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 67.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 64.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 64.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 64.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 61.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 61.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 61.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 58.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 58.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 58.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 56 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 56 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 56 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 53.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 53.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 53.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 50.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 50.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 50.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 47.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 47.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 47.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 44.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 44.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 44.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 42 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 42 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 42 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 39.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 39.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 39.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 36.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 36.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 36.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 33.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 33.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 33.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 30.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 30.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 30.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 28 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 28 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 28 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 25.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 25.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 25.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 22.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 22.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 22.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 19.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 19.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 19.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 16.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 16.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 16.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 14 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 14 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 14 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 11.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 11.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 11.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 8.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 8.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 8.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 5.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 5.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 5.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 2.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 2.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 2.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 232.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 232.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 232.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 229.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 229.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 229.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 226.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 226.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 226.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 224 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 224 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 224 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 221.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 221.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 221.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 218.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 218.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 218.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 215.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 215.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 215.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 212.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 212.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 212.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 210 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 210 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 210 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 207.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 207.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 207.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 204.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 204.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 204.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 201.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 201.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 201.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 198.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 198.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 198.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 196 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 196 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 196 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 193.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 193.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 193.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 190.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 190.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 190.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 187.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 187.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 187.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 184.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 184.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 184.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 182 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 182 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 182 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 179.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 179.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 179.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 176.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 176.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 176.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 173.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 173.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 173.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 170.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 170.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 170.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 168 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 168 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 168 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 165.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 165.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 165.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 162.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 162.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 162.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 159.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 159.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 159.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 156.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 156.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 156.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 154 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 154 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 154 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 151.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 151.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 151.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 148.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 148.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 148.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 145.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 145.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 145.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 142.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 142.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 142.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 140 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 140 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 140 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 137.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 137.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 137.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 134.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 134.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 134.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 131.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 131.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 131.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 128.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 128.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 128.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 126 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 126 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 126 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 123.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 123.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 123.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 120.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 120.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 120.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 117.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 117.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 117.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 114.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 114.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 114.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 112 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 112 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 112 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 109.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 109.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 109.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 106.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 106.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 106.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 103.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 103.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 103.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 100.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 100.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 100.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 98 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 98 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 98 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 95.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 95.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 95.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 92.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 92.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 92.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 89.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 89.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 89.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 86.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 86.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 86.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 84 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 84 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 84 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 81.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 81.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 81.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 78.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 78.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 78.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 75.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 75.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 75.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 72.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 72.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 72.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 70 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 70 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 70 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 67.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 67.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 67.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 64.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 64.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 64.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 61.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 61.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 61.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 58.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 58.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 58.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 56 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 56 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 56 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 53.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 53.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 53.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 50.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 50.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 50.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 47.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 47.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 47.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 44.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 44.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 44.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 42 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 42 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 42 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 39.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 39.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 39.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 36.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 36.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 36.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 33.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 33.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 33.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 30.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 30.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 30.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 28 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 28 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 28 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 25.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 25.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 25.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 22.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 22.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 22.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 19.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 19.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 19.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 16.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 16.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 16.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 14 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 14 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 14 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 11.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 11.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 11.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 8.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 8.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 8.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 5.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 5.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 5.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 2.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 2.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 2.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 232.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 232.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 232.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 229.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 229.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 229.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 226.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 226.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 226.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 224 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 224 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 224 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 221.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 221.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 221.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 218.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 218.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 218.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 215.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 215.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 215.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 212.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 212.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 212.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 210 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 210 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 210 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 207.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 207.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 207.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 204.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 204.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 204.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 201.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 201.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 201.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 198.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 198.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 198.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 196 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 196 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 196 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 193.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 193.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 193.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 190.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 190.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 190.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 187.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 187.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 187.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 184.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 184.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 184.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 182 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 182 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 182 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 179.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 179.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 179.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 176.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 176.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 176.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 173.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 173.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 173.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 170.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 170.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 170.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 168 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 168 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 168 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 165.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 165.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 165.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 162.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 162.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 162.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 159.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 159.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 159.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 156.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 156.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 156.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 154 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 154 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 154 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 151.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 151.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 151.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 148.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 148.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 148.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 145.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 145.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 145.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 142.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 142.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 142.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 140 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 140 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 140 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 137.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 137.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 137.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 134.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 134.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 134.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 131.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 131.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 131.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 128.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 128.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 128.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 126 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 126 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 126 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 123.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 123.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 123.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 120.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 120.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 120.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 117.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 117.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 117.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 114.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 114.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 114.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 112 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 112 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 112 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 109.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 109.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 109.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 106.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 106.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 106.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 103.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 103.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 103.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 100.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 100.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 100.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 98 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 98 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 98 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 95.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 95.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 95.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 92.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 92.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 92.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 89.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 89.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 89.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 86.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 86.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 86.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 84 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 84 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 84 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 81.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 81.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 81.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 78.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 78.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 78.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 75.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 75.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 75.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 72.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 72.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 72.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 70 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 70 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 70 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 67.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 67.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 67.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 64.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 64.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 64.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 61.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 61.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 61.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 58.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 58.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 58.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 56 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 56 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 56 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 53.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 53.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 53.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 50.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 50.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 50.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 47.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 47.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 47.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 44.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 44.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 44.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 42 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 42 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 42 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 39.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 39.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 39.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 36.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 36.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 36.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 33.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 33.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 33.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 30.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 30.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 30.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 28 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 28 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 28 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 25.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 25.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 25.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 22.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 22.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 22.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 19.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 19.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 19.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 16.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 16.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 16.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 14 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 14 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 14 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 11.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 11.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 11.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 8.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 8.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 8.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 5.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 5.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 5.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 2.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 2.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 2.8 via1_2_400_200_1_1_300_300 ;
    END
  END VDD
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  334.345 235.83 334.485 235.97 ;
    END
  END addr[0]
  PIN addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  220.665 235.83 220.805 235.97 ;
    END
  END addr[10]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  391.81 178.64 391.95 178.78 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  391.81 7.84 391.95 7.98 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  163.545 235.83 163.685 235.97 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 227.92 0.14 228.06 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 114.24 0.14 114.38 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  341.625 0 341.765 0.14 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  227.945 0 228.085 0.14 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  0.585 0 0.725 0.14 ;
    END
  END addr[8]
  PIN addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  390.905 235.83 391.045 235.97 ;
    END
  END addr[9]
  PIN ce
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  57.145 0 57.285 0.14 ;
    END
  END ce
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  285.065 0 285.205 0.14 ;
    END
  END clk
  PIN di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  114.265 0 114.405 0.14 ;
    END
  END di[0]
  PIN di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 57.12 0.14 57.26 ;
    END
  END di[1]
  PIN di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  391.81 121.52 391.95 121.66 ;
    END
  END di[2]
  PIN di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  49.865 235.83 50.005 235.97 ;
    END
  END di[3]
  PIN doq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  277.225 235.83 277.365 235.97 ;
    END
  END doq[0]
  PIN doq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  170.825 0 170.965 0.14 ;
    END
  END doq[1]
  PIN doq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 170.8 0.14 170.94 ;
    END
  END doq[2]
  PIN doq[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  106.425 235.83 106.565 235.97 ;
    END
  END doq[3]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  391.81 64.96 391.95 65.1 ;
    END
  END we
  OBS
    LAYER metal1 ;
     RECT  0 0 391.95 235.97 ;
    LAYER metal2 ;
     RECT  0 0 391.95 235.97 ;
    LAYER metal3 ;
     RECT  0 0 391.95 235.97 ;
    LAYER metal4 ;
     RECT  0 0 391.95 235.97 ;
    LAYER metal5 ;
     RECT  0 0 391.95 235.97 ;
    LAYER metal6 ;
     RECT  0 0 391.95 235.97 ;
    LAYER metal7 ;
     RECT  0 0 391.95 235.97 ;
    LAYER metal8 ;
     RECT  0 0 391.95 235.97 ;
    LAYER metal9 ;
     RECT  0 0 391.95 235.97 ;
  END
END memory4
END LIBRARY
