VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS
MACRO or1200_spram2
  FOREIGN or1200_spram2 0 0 ;
  CLASS BLOCK ;
  SIZE 340.72 BY 340.72 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal7 ;
        RECT  2.94 322.7 339.34 324.1 ;
        RECT  2.94 282.7 339.34 284.1 ;
        RECT  2.94 242.7 339.34 244.1 ;
        RECT  2.94 202.7 339.34 204.1 ;
        RECT  2.94 162.7 339.34 164.1 ;
        RECT  2.94 122.7 339.34 124.1 ;
        RECT  2.94 82.7 339.34 84.1 ;
        RECT  2.94 42.7 339.34 44.1 ;
        RECT  2.94 2.7 339.34 4.1 ;
      LAYER metal4 ;
        RECT  339.04 1.33 339.24 337.47 ;
        RECT  283.04 1.33 283.24 337.47 ;
        RECT  227.04 1.33 227.24 337.47 ;
        RECT  171.04 1.33 171.24 337.47 ;
        RECT  115.04 1.33 115.24 337.47 ;
        RECT  59.04 1.33 59.24 337.47 ;
        RECT  3.04 1.33 3.24 337.47 ;
      LAYER metal1 ;
        RECT  1.14 337.35 339.53 337.45 ;
        RECT  1.14 334.55 339.53 334.65 ;
        RECT  1.14 331.75 339.53 331.85 ;
        RECT  1.14 328.95 339.53 329.05 ;
        RECT  1.14 326.15 339.53 326.25 ;
        RECT  1.14 323.35 339.53 323.45 ;
        RECT  1.14 320.55 339.53 320.65 ;
        RECT  1.14 317.75 339.53 317.85 ;
        RECT  1.14 314.95 339.53 315.05 ;
        RECT  1.14 312.15 339.53 312.25 ;
        RECT  1.14 309.35 339.53 309.45 ;
        RECT  1.14 306.55 339.53 306.65 ;
        RECT  1.14 303.75 339.53 303.85 ;
        RECT  1.14 300.95 339.53 301.05 ;
        RECT  1.14 298.15 339.53 298.25 ;
        RECT  1.14 295.35 339.53 295.45 ;
        RECT  1.14 292.55 339.53 292.65 ;
        RECT  1.14 289.75 339.53 289.85 ;
        RECT  1.14 286.95 339.53 287.05 ;
        RECT  1.14 284.15 339.53 284.25 ;
        RECT  1.14 281.35 339.53 281.45 ;
        RECT  1.14 278.55 339.53 278.65 ;
        RECT  1.14 275.75 339.53 275.85 ;
        RECT  1.14 272.95 339.53 273.05 ;
        RECT  1.14 270.15 339.53 270.25 ;
        RECT  1.14 267.35 339.53 267.45 ;
        RECT  1.14 264.55 339.53 264.65 ;
        RECT  1.14 261.75 339.53 261.85 ;
        RECT  1.14 258.95 339.53 259.05 ;
        RECT  1.14 256.15 339.53 256.25 ;
        RECT  1.14 253.35 339.53 253.45 ;
        RECT  1.14 250.55 339.53 250.65 ;
        RECT  1.14 247.75 339.53 247.85 ;
        RECT  1.14 244.95 339.53 245.05 ;
        RECT  1.14 242.15 339.53 242.25 ;
        RECT  1.14 239.35 339.53 239.45 ;
        RECT  1.14 236.55 339.53 236.65 ;
        RECT  1.14 233.75 339.53 233.85 ;
        RECT  1.14 230.95 339.53 231.05 ;
        RECT  1.14 228.15 339.53 228.25 ;
        RECT  1.14 225.35 339.53 225.45 ;
        RECT  1.14 222.55 339.53 222.65 ;
        RECT  1.14 219.75 339.53 219.85 ;
        RECT  1.14 216.95 339.53 217.05 ;
        RECT  1.14 214.15 339.53 214.25 ;
        RECT  1.14 211.35 339.53 211.45 ;
        RECT  1.14 208.55 339.53 208.65 ;
        RECT  1.14 205.75 339.53 205.85 ;
        RECT  1.14 202.95 339.53 203.05 ;
        RECT  1.14 200.15 339.53 200.25 ;
        RECT  1.14 197.35 339.53 197.45 ;
        RECT  1.14 194.55 339.53 194.65 ;
        RECT  1.14 191.75 339.53 191.85 ;
        RECT  1.14 188.95 339.53 189.05 ;
        RECT  1.14 186.15 339.53 186.25 ;
        RECT  1.14 183.35 339.53 183.45 ;
        RECT  1.14 180.55 339.53 180.65 ;
        RECT  1.14 177.75 339.53 177.85 ;
        RECT  1.14 174.95 339.53 175.05 ;
        RECT  1.14 172.15 339.53 172.25 ;
        RECT  1.14 169.35 339.53 169.45 ;
        RECT  1.14 166.55 339.53 166.65 ;
        RECT  1.14 163.75 339.53 163.85 ;
        RECT  1.14 160.95 339.53 161.05 ;
        RECT  1.14 158.15 339.53 158.25 ;
        RECT  1.14 155.35 339.53 155.45 ;
        RECT  1.14 152.55 339.53 152.65 ;
        RECT  1.14 149.75 339.53 149.85 ;
        RECT  1.14 146.95 339.53 147.05 ;
        RECT  1.14 144.15 339.53 144.25 ;
        RECT  1.14 141.35 339.53 141.45 ;
        RECT  1.14 138.55 339.53 138.65 ;
        RECT  1.14 135.75 339.53 135.85 ;
        RECT  1.14 132.95 339.53 133.05 ;
        RECT  1.14 130.15 339.53 130.25 ;
        RECT  1.14 127.35 339.53 127.45 ;
        RECT  1.14 124.55 339.53 124.65 ;
        RECT  1.14 121.75 339.53 121.85 ;
        RECT  1.14 118.95 339.53 119.05 ;
        RECT  1.14 116.15 339.53 116.25 ;
        RECT  1.14 113.35 339.53 113.45 ;
        RECT  1.14 110.55 339.53 110.65 ;
        RECT  1.14 107.75 339.53 107.85 ;
        RECT  1.14 104.95 339.53 105.05 ;
        RECT  1.14 102.15 339.53 102.25 ;
        RECT  1.14 99.35 339.53 99.45 ;
        RECT  1.14 96.55 339.53 96.65 ;
        RECT  1.14 93.75 339.53 93.85 ;
        RECT  1.14 90.95 339.53 91.05 ;
        RECT  1.14 88.15 339.53 88.25 ;
        RECT  1.14 85.35 339.53 85.45 ;
        RECT  1.14 82.55 339.53 82.65 ;
        RECT  1.14 79.75 339.53 79.85 ;
        RECT  1.14 76.95 339.53 77.05 ;
        RECT  1.14 74.15 339.53 74.25 ;
        RECT  1.14 71.35 339.53 71.45 ;
        RECT  1.14 68.55 339.53 68.65 ;
        RECT  1.14 65.75 339.53 65.85 ;
        RECT  1.14 62.95 339.53 63.05 ;
        RECT  1.14 60.15 339.53 60.25 ;
        RECT  1.14 57.35 339.53 57.45 ;
        RECT  1.14 54.55 339.53 54.65 ;
        RECT  1.14 51.75 339.53 51.85 ;
        RECT  1.14 48.95 339.53 49.05 ;
        RECT  1.14 46.15 339.53 46.25 ;
        RECT  1.14 43.35 339.53 43.45 ;
        RECT  1.14 40.55 339.53 40.65 ;
        RECT  1.14 37.75 339.53 37.85 ;
        RECT  1.14 34.95 339.53 35.05 ;
        RECT  1.14 32.15 339.53 32.25 ;
        RECT  1.14 29.35 339.53 29.45 ;
        RECT  1.14 26.55 339.53 26.65 ;
        RECT  1.14 23.75 339.53 23.85 ;
        RECT  1.14 20.95 339.53 21.05 ;
        RECT  1.14 18.15 339.53 18.25 ;
        RECT  1.14 15.35 339.53 15.45 ;
        RECT  1.14 12.55 339.53 12.65 ;
        RECT  1.14 9.75 339.53 9.85 ;
        RECT  1.14 6.95 339.53 7.05 ;
        RECT  1.14 4.15 339.53 4.25 ;
        RECT  1.14 1.35 339.53 1.45 ;
      VIA 339.14 323.4 via6_7_400_2800_4_1_600_600 ;
      VIA 339.14 323.4 via5_6_400_2800_5_1_600_600 ;
      VIA 339.14 323.4 via4_5_400_2800_5_1_600_600 ;
      VIA 339.14 283.4 via6_7_400_2800_4_1_600_600 ;
      VIA 339.14 283.4 via5_6_400_2800_5_1_600_600 ;
      VIA 339.14 283.4 via4_5_400_2800_5_1_600_600 ;
      VIA 339.14 243.4 via6_7_400_2800_4_1_600_600 ;
      VIA 339.14 243.4 via5_6_400_2800_5_1_600_600 ;
      VIA 339.14 243.4 via4_5_400_2800_5_1_600_600 ;
      VIA 339.14 203.4 via6_7_400_2800_4_1_600_600 ;
      VIA 339.14 203.4 via5_6_400_2800_5_1_600_600 ;
      VIA 339.14 203.4 via4_5_400_2800_5_1_600_600 ;
      VIA 339.14 163.4 via6_7_400_2800_4_1_600_600 ;
      VIA 339.14 163.4 via5_6_400_2800_5_1_600_600 ;
      VIA 339.14 163.4 via4_5_400_2800_5_1_600_600 ;
      VIA 339.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 339.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 339.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 339.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 339.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 339.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 339.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 339.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 339.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 339.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 339.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 339.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 323.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 323.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 323.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 283.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 283.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 283.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 243.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 243.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 243.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 203.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 203.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 203.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 163.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 163.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 163.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 323.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 323.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 323.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 283.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 283.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 283.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 243.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 243.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 243.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 203.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 203.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 203.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 163.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 163.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 163.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 323.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 323.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 323.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 283.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 283.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 283.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 243.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 243.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 243.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 203.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 203.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 203.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 163.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 163.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 163.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 323.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 323.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 323.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 283.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 283.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 283.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 243.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 243.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 243.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 203.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 203.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 203.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 163.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 163.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 163.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 323.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 323.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 323.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 283.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 283.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 283.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 243.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 243.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 243.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 203.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 203.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 203.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 163.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 163.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 163.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 323.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 323.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 323.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 283.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 283.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 283.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 243.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 243.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 243.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 203.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 203.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 203.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 163.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 163.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 163.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 339.14 337.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 337.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 337.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 334.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 334.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 334.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 331.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 331.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 331.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 329 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 329 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 329 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 326.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 326.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 326.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 323.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 323.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 323.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 320.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 320.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 320.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 317.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 317.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 317.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 315 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 315 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 315 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 312.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 312.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 312.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 309.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 309.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 309.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 306.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 306.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 306.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 303.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 303.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 303.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 301 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 301 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 301 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 298.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 298.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 298.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 295.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 295.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 295.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 292.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 292.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 292.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 289.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 289.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 289.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 287 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 287 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 287 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 284.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 284.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 284.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 281.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 281.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 281.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 278.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 278.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 278.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 275.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 275.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 275.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 273 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 273 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 273 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 270.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 270.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 270.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 267.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 267.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 267.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 264.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 264.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 264.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 261.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 261.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 261.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 259 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 259 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 259 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 256.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 256.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 256.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 253.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 253.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 253.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 250.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 250.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 250.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 247.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 247.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 247.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 245 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 245 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 245 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 242.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 242.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 242.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 239.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 239.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 239.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 236.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 236.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 236.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 233.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 233.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 233.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 231 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 231 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 231 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 228.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 228.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 228.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 225.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 225.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 225.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 222.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 222.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 222.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 219.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 219.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 219.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 217 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 217 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 217 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 214.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 214.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 214.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 211.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 211.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 211.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 208.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 208.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 208.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 205.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 205.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 205.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 203 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 203 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 203 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 200.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 200.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 200.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 197.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 197.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 197.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 194.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 194.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 194.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 191.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 191.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 191.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 189 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 189 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 189 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 186.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 186.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 186.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 183.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 183.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 183.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 180.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 180.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 180.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 177.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 177.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 177.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 175 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 175 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 175 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 172.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 172.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 172.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 169.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 169.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 169.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 166.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 166.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 166.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 163.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 163.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 163.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 161 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 161 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 161 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 158.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 158.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 158.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 155.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 155.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 155.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 152.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 152.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 152.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 149.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 149.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 149.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 147 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 147 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 147 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 144.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 144.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 144.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 141.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 141.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 141.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 138.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 138.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 138.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 339.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 339.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 339.14 1.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 337.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 337.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 337.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 334.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 334.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 334.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 331.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 331.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 331.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 329 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 329 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 329 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 326.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 326.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 326.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 323.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 323.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 323.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 320.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 320.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 320.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 317.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 317.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 317.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 315 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 315 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 315 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 312.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 312.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 312.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 309.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 309.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 309.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 306.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 306.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 306.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 303.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 303.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 303.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 301 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 301 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 301 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 298.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 298.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 298.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 295.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 295.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 295.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 292.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 292.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 292.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 289.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 289.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 289.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 287 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 287 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 287 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 284.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 284.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 284.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 281.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 281.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 281.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 278.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 278.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 278.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 275.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 275.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 275.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 273 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 273 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 273 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 270.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 270.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 270.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 267.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 267.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 267.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 264.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 264.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 264.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 261.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 261.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 261.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 259 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 259 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 259 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 256.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 256.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 256.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 253.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 253.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 253.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 250.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 250.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 250.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 247.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 247.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 247.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 245 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 245 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 245 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 242.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 242.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 242.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 239.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 239.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 239.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 236.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 236.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 236.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 233.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 233.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 233.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 231 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 231 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 231 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 228.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 228.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 228.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 225.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 225.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 225.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 222.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 222.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 222.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 219.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 219.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 219.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 217 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 217 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 217 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 214.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 214.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 214.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 211.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 211.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 211.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 208.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 208.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 208.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 205.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 205.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 205.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 203 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 203 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 203 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 200.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 200.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 200.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 197.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 197.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 197.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 194.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 194.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 194.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 191.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 191.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 191.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 189 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 189 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 189 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 186.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 186.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 186.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 183.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 183.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 183.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 180.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 180.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 180.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 177.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 177.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 177.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 175 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 175 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 175 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 172.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 172.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 172.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 169.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 169.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 169.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 166.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 166.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 166.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 163.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 163.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 163.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 161 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 161 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 161 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 158.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 158.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 158.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 155.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 155.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 155.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 152.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 152.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 152.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 149.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 149.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 149.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 147 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 147 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 147 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 144.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 144.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 144.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 141.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 141.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 141.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 138.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 138.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 138.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 1.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 337.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 337.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 337.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 334.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 334.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 334.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 331.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 331.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 331.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 329 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 329 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 329 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 326.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 326.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 326.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 323.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 323.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 323.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 320.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 320.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 320.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 317.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 317.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 317.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 315 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 315 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 315 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 312.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 312.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 312.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 309.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 309.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 309.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 306.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 306.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 306.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 303.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 303.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 303.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 301 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 301 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 301 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 298.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 298.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 298.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 295.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 295.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 295.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 292.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 292.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 292.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 289.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 289.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 289.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 287 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 287 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 287 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 284.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 284.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 284.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 281.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 281.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 281.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 278.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 278.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 278.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 275.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 275.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 275.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 273 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 273 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 273 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 270.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 270.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 270.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 267.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 267.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 267.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 264.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 264.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 264.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 261.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 261.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 261.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 259 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 259 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 259 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 256.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 256.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 256.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 253.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 253.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 253.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 250.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 250.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 250.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 247.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 247.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 247.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 245 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 245 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 245 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 242.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 242.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 242.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 239.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 239.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 239.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 236.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 236.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 236.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 233.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 233.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 233.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 231 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 231 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 231 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 228.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 228.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 228.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 225.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 225.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 225.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 222.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 222.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 222.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 219.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 219.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 219.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 217 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 217 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 217 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 214.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 214.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 214.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 211.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 211.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 211.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 208.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 208.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 208.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 205.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 205.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 205.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 203 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 203 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 203 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 200.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 200.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 200.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 197.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 197.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 197.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 194.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 194.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 194.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 191.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 191.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 191.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 189 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 189 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 189 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 186.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 186.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 186.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 183.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 183.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 183.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 180.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 180.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 180.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 177.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 177.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 177.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 175 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 175 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 175 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 172.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 172.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 172.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 169.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 169.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 169.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 166.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 166.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 166.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 163.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 163.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 163.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 161 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 161 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 161 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 158.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 158.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 158.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 155.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 155.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 155.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 152.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 152.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 152.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 149.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 149.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 149.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 147 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 147 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 147 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 144.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 144.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 144.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 141.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 141.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 141.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 138.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 138.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 138.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 1.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 337.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 337.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 337.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 334.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 334.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 334.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 331.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 331.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 331.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 329 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 329 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 329 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 326.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 326.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 326.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 323.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 323.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 323.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 320.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 320.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 320.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 317.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 317.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 317.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 315 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 315 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 315 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 312.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 312.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 312.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 309.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 309.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 309.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 306.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 306.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 306.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 303.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 303.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 303.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 301 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 301 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 301 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 298.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 298.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 298.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 295.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 295.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 295.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 292.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 292.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 292.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 289.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 289.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 289.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 287 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 287 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 287 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 284.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 284.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 284.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 281.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 281.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 281.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 278.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 278.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 278.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 275.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 275.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 275.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 273 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 273 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 273 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 270.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 270.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 270.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 267.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 267.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 267.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 264.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 264.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 264.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 261.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 261.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 261.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 259 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 259 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 259 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 256.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 256.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 256.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 253.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 253.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 253.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 250.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 250.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 250.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 247.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 247.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 247.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 245 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 245 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 245 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 242.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 242.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 242.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 239.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 239.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 239.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 236.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 236.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 236.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 233.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 233.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 233.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 231 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 231 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 231 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 228.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 228.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 228.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 225.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 225.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 225.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 222.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 222.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 222.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 219.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 219.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 219.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 217 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 217 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 217 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 214.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 214.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 214.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 211.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 211.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 211.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 208.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 208.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 208.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 205.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 205.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 205.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 203 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 203 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 203 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 200.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 200.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 200.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 197.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 197.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 197.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 194.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 194.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 194.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 191.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 191.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 191.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 189 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 189 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 189 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 186.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 186.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 186.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 183.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 183.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 183.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 180.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 180.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 180.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 177.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 177.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 177.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 175 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 175 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 175 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 172.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 172.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 172.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 169.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 169.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 169.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 166.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 166.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 166.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 163.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 163.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 163.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 161 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 161 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 161 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 158.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 158.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 158.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 155.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 155.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 155.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 152.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 152.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 152.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 149.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 149.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 149.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 147 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 147 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 147 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 144.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 144.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 144.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 141.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 141.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 141.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 138.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 138.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 138.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 1.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 337.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 337.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 337.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 334.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 334.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 334.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 331.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 331.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 331.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 329 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 329 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 329 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 326.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 326.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 326.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 323.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 323.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 323.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 320.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 320.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 320.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 317.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 317.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 317.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 315 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 315 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 315 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 312.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 312.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 312.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 309.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 309.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 309.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 306.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 306.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 306.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 303.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 303.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 303.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 301 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 301 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 301 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 298.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 298.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 298.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 295.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 295.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 295.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 292.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 292.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 292.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 289.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 289.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 289.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 287 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 287 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 287 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 284.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 284.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 284.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 281.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 281.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 281.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 278.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 278.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 278.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 275.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 275.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 275.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 273 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 273 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 273 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 270.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 270.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 270.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 267.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 267.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 267.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 264.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 264.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 264.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 261.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 261.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 261.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 259 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 259 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 259 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 256.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 256.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 256.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 253.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 253.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 253.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 250.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 250.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 250.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 247.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 247.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 247.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 245 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 245 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 245 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 242.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 242.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 242.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 239.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 239.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 239.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 236.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 236.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 236.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 233.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 233.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 233.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 231 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 231 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 231 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 228.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 228.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 228.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 225.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 225.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 225.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 222.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 222.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 222.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 219.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 219.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 219.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 217 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 217 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 217 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 214.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 214.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 214.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 211.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 211.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 211.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 208.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 208.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 208.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 205.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 205.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 205.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 203 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 203 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 203 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 200.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 200.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 200.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 197.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 197.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 197.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 194.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 194.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 194.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 191.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 191.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 191.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 189 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 189 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 189 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 186.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 186.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 186.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 183.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 183.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 183.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 180.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 180.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 180.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 177.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 177.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 177.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 175 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 175 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 175 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 172.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 172.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 172.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 169.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 169.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 169.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 166.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 166.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 166.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 163.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 163.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 163.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 161 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 161 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 161 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 158.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 158.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 158.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 155.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 155.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 155.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 152.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 152.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 152.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 149.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 149.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 149.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 147 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 147 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 147 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 144.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 144.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 144.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 141.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 141.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 141.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 138.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 138.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 138.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 1.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 337.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 337.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 337.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 334.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 334.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 334.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 331.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 331.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 331.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 329 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 329 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 329 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 326.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 326.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 326.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 323.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 323.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 323.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 320.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 320.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 320.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 317.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 317.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 317.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 315 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 315 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 315 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 312.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 312.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 312.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 309.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 309.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 309.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 306.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 306.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 306.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 303.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 303.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 303.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 301 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 301 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 301 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 298.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 298.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 298.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 295.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 295.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 295.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 292.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 292.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 292.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 289.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 289.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 289.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 287 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 287 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 287 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 284.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 284.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 284.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 281.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 281.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 281.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 278.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 278.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 278.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 275.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 275.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 275.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 273 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 273 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 273 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 270.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 270.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 270.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 267.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 267.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 267.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 264.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 264.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 264.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 261.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 261.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 261.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 259 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 259 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 259 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 256.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 256.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 256.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 253.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 253.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 253.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 250.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 250.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 250.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 247.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 247.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 247.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 245 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 245 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 245 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 242.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 242.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 242.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 239.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 239.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 239.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 236.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 236.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 236.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 233.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 233.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 233.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 231 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 231 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 231 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 228.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 228.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 228.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 225.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 225.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 225.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 222.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 222.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 222.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 219.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 219.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 219.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 217 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 217 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 217 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 214.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 214.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 214.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 211.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 211.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 211.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 208.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 208.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 208.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 205.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 205.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 205.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 203 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 203 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 203 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 200.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 200.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 200.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 197.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 197.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 197.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 194.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 194.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 194.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 191.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 191.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 191.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 189 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 189 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 189 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 186.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 186.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 186.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 183.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 183.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 183.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 180.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 180.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 180.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 177.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 177.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 177.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 175 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 175 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 175 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 172.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 172.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 172.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 169.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 169.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 169.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 166.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 166.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 166.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 163.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 163.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 163.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 161 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 161 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 161 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 158.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 158.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 158.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 155.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 155.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 155.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 152.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 152.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 152.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 149.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 149.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 149.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 147 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 147 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 147 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 144.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 144.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 144.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 141.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 141.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 141.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 138.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 138.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 138.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 1.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 337.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 337.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 337.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 334.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 334.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 334.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 331.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 331.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 331.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 329 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 329 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 329 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 326.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 326.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 326.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 323.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 323.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 323.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 320.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 320.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 320.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 317.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 317.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 317.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 315 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 315 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 315 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 312.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 312.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 312.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 309.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 309.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 309.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 306.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 306.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 306.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 303.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 303.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 303.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 301 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 301 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 301 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 298.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 298.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 298.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 295.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 295.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 295.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 292.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 292.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 292.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 289.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 289.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 289.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 287 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 287 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 287 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 284.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 284.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 284.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 281.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 281.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 281.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 278.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 278.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 278.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 275.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 275.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 275.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 273 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 273 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 273 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 270.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 270.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 270.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 267.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 267.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 267.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 264.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 264.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 264.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 261.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 261.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 261.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 259 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 259 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 259 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 256.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 256.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 256.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 253.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 253.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 253.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 250.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 250.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 250.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 247.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 247.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 247.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 245 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 245 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 245 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 242.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 242.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 242.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 239.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 239.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 239.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 236.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 236.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 236.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 233.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 233.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 233.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 231 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 231 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 231 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 228.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 228.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 228.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 225.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 225.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 225.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 222.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 222.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 222.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 219.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 219.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 219.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 217 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 217 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 217 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 214.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 214.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 214.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 211.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 211.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 211.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 208.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 208.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 208.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 205.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 205.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 205.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 203 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 203 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 203 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 200.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 200.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 200.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 197.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 197.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 197.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 194.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 194.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 194.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 191.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 191.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 191.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 189 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 189 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 189 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 186.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 186.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 186.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 183.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 183.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 183.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 180.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 180.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 180.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 177.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 177.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 177.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 175 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 175 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 175 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 172.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 172.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 172.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 169.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 169.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 169.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 166.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 166.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 166.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 163.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 163.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 163.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 161 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 161 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 161 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 158.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 158.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 158.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 155.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 155.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 155.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 152.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 152.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 152.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 149.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 149.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 149.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 147 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 147 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 147 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 144.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 144.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 144.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 141.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 141.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 141.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 138.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 138.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 138.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 1.4 via1_2_400_200_1_1_300_300 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal7 ;
        RECT  30.94 302.7 311.34 304.1 ;
        RECT  30.94 262.7 311.34 264.1 ;
        RECT  30.94 222.7 311.34 224.1 ;
        RECT  30.94 182.7 311.34 184.1 ;
        RECT  30.94 142.7 311.34 144.1 ;
        RECT  30.94 102.7 311.34 104.1 ;
        RECT  30.94 62.7 311.34 64.1 ;
        RECT  30.94 22.7 311.34 24.1 ;
      LAYER metal4 ;
        RECT  311.04 2.73 311.24 338.87 ;
        RECT  255.04 2.73 255.24 338.87 ;
        RECT  199.04 2.73 199.24 338.87 ;
        RECT  143.04 2.73 143.24 338.87 ;
        RECT  87.04 2.73 87.24 338.87 ;
        RECT  31.04 2.73 31.24 338.87 ;
      LAYER metal1 ;
        RECT  1.14 338.75 339.53 338.85 ;
        RECT  1.14 335.95 339.53 336.05 ;
        RECT  1.14 333.15 339.53 333.25 ;
        RECT  1.14 330.35 339.53 330.45 ;
        RECT  1.14 327.55 339.53 327.65 ;
        RECT  1.14 324.75 339.53 324.85 ;
        RECT  1.14 321.95 339.53 322.05 ;
        RECT  1.14 319.15 339.53 319.25 ;
        RECT  1.14 316.35 339.53 316.45 ;
        RECT  1.14 313.55 339.53 313.65 ;
        RECT  1.14 310.75 339.53 310.85 ;
        RECT  1.14 307.95 339.53 308.05 ;
        RECT  1.14 305.15 339.53 305.25 ;
        RECT  1.14 302.35 339.53 302.45 ;
        RECT  1.14 299.55 339.53 299.65 ;
        RECT  1.14 296.75 339.53 296.85 ;
        RECT  1.14 293.95 339.53 294.05 ;
        RECT  1.14 291.15 339.53 291.25 ;
        RECT  1.14 288.35 339.53 288.45 ;
        RECT  1.14 285.55 339.53 285.65 ;
        RECT  1.14 282.75 339.53 282.85 ;
        RECT  1.14 279.95 339.53 280.05 ;
        RECT  1.14 277.15 339.53 277.25 ;
        RECT  1.14 274.35 339.53 274.45 ;
        RECT  1.14 271.55 339.53 271.65 ;
        RECT  1.14 268.75 339.53 268.85 ;
        RECT  1.14 265.95 339.53 266.05 ;
        RECT  1.14 263.15 339.53 263.25 ;
        RECT  1.14 260.35 339.53 260.45 ;
        RECT  1.14 257.55 339.53 257.65 ;
        RECT  1.14 254.75 339.53 254.85 ;
        RECT  1.14 251.95 339.53 252.05 ;
        RECT  1.14 249.15 339.53 249.25 ;
        RECT  1.14 246.35 339.53 246.45 ;
        RECT  1.14 243.55 339.53 243.65 ;
        RECT  1.14 240.75 339.53 240.85 ;
        RECT  1.14 237.95 339.53 238.05 ;
        RECT  1.14 235.15 339.53 235.25 ;
        RECT  1.14 232.35 339.53 232.45 ;
        RECT  1.14 229.55 339.53 229.65 ;
        RECT  1.14 226.75 339.53 226.85 ;
        RECT  1.14 223.95 339.53 224.05 ;
        RECT  1.14 221.15 339.53 221.25 ;
        RECT  1.14 218.35 339.53 218.45 ;
        RECT  1.14 215.55 339.53 215.65 ;
        RECT  1.14 212.75 339.53 212.85 ;
        RECT  1.14 209.95 339.53 210.05 ;
        RECT  1.14 207.15 339.53 207.25 ;
        RECT  1.14 204.35 339.53 204.45 ;
        RECT  1.14 201.55 339.53 201.65 ;
        RECT  1.14 198.75 339.53 198.85 ;
        RECT  1.14 195.95 339.53 196.05 ;
        RECT  1.14 193.15 339.53 193.25 ;
        RECT  1.14 190.35 339.53 190.45 ;
        RECT  1.14 187.55 339.53 187.65 ;
        RECT  1.14 184.75 339.53 184.85 ;
        RECT  1.14 181.95 339.53 182.05 ;
        RECT  1.14 179.15 339.53 179.25 ;
        RECT  1.14 176.35 339.53 176.45 ;
        RECT  1.14 173.55 339.53 173.65 ;
        RECT  1.14 170.75 339.53 170.85 ;
        RECT  1.14 167.95 339.53 168.05 ;
        RECT  1.14 165.15 339.53 165.25 ;
        RECT  1.14 162.35 339.53 162.45 ;
        RECT  1.14 159.55 339.53 159.65 ;
        RECT  1.14 156.75 339.53 156.85 ;
        RECT  1.14 153.95 339.53 154.05 ;
        RECT  1.14 151.15 339.53 151.25 ;
        RECT  1.14 148.35 339.53 148.45 ;
        RECT  1.14 145.55 339.53 145.65 ;
        RECT  1.14 142.75 339.53 142.85 ;
        RECT  1.14 139.95 339.53 140.05 ;
        RECT  1.14 137.15 339.53 137.25 ;
        RECT  1.14 134.35 339.53 134.45 ;
        RECT  1.14 131.55 339.53 131.65 ;
        RECT  1.14 128.75 339.53 128.85 ;
        RECT  1.14 125.95 339.53 126.05 ;
        RECT  1.14 123.15 339.53 123.25 ;
        RECT  1.14 120.35 339.53 120.45 ;
        RECT  1.14 117.55 339.53 117.65 ;
        RECT  1.14 114.75 339.53 114.85 ;
        RECT  1.14 111.95 339.53 112.05 ;
        RECT  1.14 109.15 339.53 109.25 ;
        RECT  1.14 106.35 339.53 106.45 ;
        RECT  1.14 103.55 339.53 103.65 ;
        RECT  1.14 100.75 339.53 100.85 ;
        RECT  1.14 97.95 339.53 98.05 ;
        RECT  1.14 95.15 339.53 95.25 ;
        RECT  1.14 92.35 339.53 92.45 ;
        RECT  1.14 89.55 339.53 89.65 ;
        RECT  1.14 86.75 339.53 86.85 ;
        RECT  1.14 83.95 339.53 84.05 ;
        RECT  1.14 81.15 339.53 81.25 ;
        RECT  1.14 78.35 339.53 78.45 ;
        RECT  1.14 75.55 339.53 75.65 ;
        RECT  1.14 72.75 339.53 72.85 ;
        RECT  1.14 69.95 339.53 70.05 ;
        RECT  1.14 67.15 339.53 67.25 ;
        RECT  1.14 64.35 339.53 64.45 ;
        RECT  1.14 61.55 339.53 61.65 ;
        RECT  1.14 58.75 339.53 58.85 ;
        RECT  1.14 55.95 339.53 56.05 ;
        RECT  1.14 53.15 339.53 53.25 ;
        RECT  1.14 50.35 339.53 50.45 ;
        RECT  1.14 47.55 339.53 47.65 ;
        RECT  1.14 44.75 339.53 44.85 ;
        RECT  1.14 41.95 339.53 42.05 ;
        RECT  1.14 39.15 339.53 39.25 ;
        RECT  1.14 36.35 339.53 36.45 ;
        RECT  1.14 33.55 339.53 33.65 ;
        RECT  1.14 30.75 339.53 30.85 ;
        RECT  1.14 27.95 339.53 28.05 ;
        RECT  1.14 25.15 339.53 25.25 ;
        RECT  1.14 22.35 339.53 22.45 ;
        RECT  1.14 19.55 339.53 19.65 ;
        RECT  1.14 16.75 339.53 16.85 ;
        RECT  1.14 13.95 339.53 14.05 ;
        RECT  1.14 11.15 339.53 11.25 ;
        RECT  1.14 8.35 339.53 8.45 ;
        RECT  1.14 5.55 339.53 5.65 ;
        RECT  1.14 2.75 339.53 2.85 ;
      VIA 311.14 303.4 via6_7_400_2800_4_1_600_600 ;
      VIA 311.14 303.4 via5_6_400_2800_5_1_600_600 ;
      VIA 311.14 303.4 via4_5_400_2800_5_1_600_600 ;
      VIA 311.14 263.4 via6_7_400_2800_4_1_600_600 ;
      VIA 311.14 263.4 via5_6_400_2800_5_1_600_600 ;
      VIA 311.14 263.4 via4_5_400_2800_5_1_600_600 ;
      VIA 311.14 223.4 via6_7_400_2800_4_1_600_600 ;
      VIA 311.14 223.4 via5_6_400_2800_5_1_600_600 ;
      VIA 311.14 223.4 via4_5_400_2800_5_1_600_600 ;
      VIA 311.14 183.4 via6_7_400_2800_4_1_600_600 ;
      VIA 311.14 183.4 via5_6_400_2800_5_1_600_600 ;
      VIA 311.14 183.4 via4_5_400_2800_5_1_600_600 ;
      VIA 311.14 143.4 via6_7_400_2800_4_1_600_600 ;
      VIA 311.14 143.4 via5_6_400_2800_5_1_600_600 ;
      VIA 311.14 143.4 via4_5_400_2800_5_1_600_600 ;
      VIA 311.14 103.4 via6_7_400_2800_4_1_600_600 ;
      VIA 311.14 103.4 via5_6_400_2800_5_1_600_600 ;
      VIA 311.14 103.4 via4_5_400_2800_5_1_600_600 ;
      VIA 311.14 63.4 via6_7_400_2800_4_1_600_600 ;
      VIA 311.14 63.4 via5_6_400_2800_5_1_600_600 ;
      VIA 311.14 63.4 via4_5_400_2800_5_1_600_600 ;
      VIA 311.14 23.4 via6_7_400_2800_4_1_600_600 ;
      VIA 311.14 23.4 via5_6_400_2800_5_1_600_600 ;
      VIA 311.14 23.4 via4_5_400_2800_5_1_600_600 ;
      VIA 255.14 303.4 via6_7_400_2800_4_1_600_600 ;
      VIA 255.14 303.4 via5_6_400_2800_5_1_600_600 ;
      VIA 255.14 303.4 via4_5_400_2800_5_1_600_600 ;
      VIA 255.14 263.4 via6_7_400_2800_4_1_600_600 ;
      VIA 255.14 263.4 via5_6_400_2800_5_1_600_600 ;
      VIA 255.14 263.4 via4_5_400_2800_5_1_600_600 ;
      VIA 255.14 223.4 via6_7_400_2800_4_1_600_600 ;
      VIA 255.14 223.4 via5_6_400_2800_5_1_600_600 ;
      VIA 255.14 223.4 via4_5_400_2800_5_1_600_600 ;
      VIA 255.14 183.4 via6_7_400_2800_4_1_600_600 ;
      VIA 255.14 183.4 via5_6_400_2800_5_1_600_600 ;
      VIA 255.14 183.4 via4_5_400_2800_5_1_600_600 ;
      VIA 255.14 143.4 via6_7_400_2800_4_1_600_600 ;
      VIA 255.14 143.4 via5_6_400_2800_5_1_600_600 ;
      VIA 255.14 143.4 via4_5_400_2800_5_1_600_600 ;
      VIA 255.14 103.4 via6_7_400_2800_4_1_600_600 ;
      VIA 255.14 103.4 via5_6_400_2800_5_1_600_600 ;
      VIA 255.14 103.4 via4_5_400_2800_5_1_600_600 ;
      VIA 255.14 63.4 via6_7_400_2800_4_1_600_600 ;
      VIA 255.14 63.4 via5_6_400_2800_5_1_600_600 ;
      VIA 255.14 63.4 via4_5_400_2800_5_1_600_600 ;
      VIA 255.14 23.4 via6_7_400_2800_4_1_600_600 ;
      VIA 255.14 23.4 via5_6_400_2800_5_1_600_600 ;
      VIA 255.14 23.4 via4_5_400_2800_5_1_600_600 ;
      VIA 199.14 303.4 via6_7_400_2800_4_1_600_600 ;
      VIA 199.14 303.4 via5_6_400_2800_5_1_600_600 ;
      VIA 199.14 303.4 via4_5_400_2800_5_1_600_600 ;
      VIA 199.14 263.4 via6_7_400_2800_4_1_600_600 ;
      VIA 199.14 263.4 via5_6_400_2800_5_1_600_600 ;
      VIA 199.14 263.4 via4_5_400_2800_5_1_600_600 ;
      VIA 199.14 223.4 via6_7_400_2800_4_1_600_600 ;
      VIA 199.14 223.4 via5_6_400_2800_5_1_600_600 ;
      VIA 199.14 223.4 via4_5_400_2800_5_1_600_600 ;
      VIA 199.14 183.4 via6_7_400_2800_4_1_600_600 ;
      VIA 199.14 183.4 via5_6_400_2800_5_1_600_600 ;
      VIA 199.14 183.4 via4_5_400_2800_5_1_600_600 ;
      VIA 199.14 143.4 via6_7_400_2800_4_1_600_600 ;
      VIA 199.14 143.4 via5_6_400_2800_5_1_600_600 ;
      VIA 199.14 143.4 via4_5_400_2800_5_1_600_600 ;
      VIA 199.14 103.4 via6_7_400_2800_4_1_600_600 ;
      VIA 199.14 103.4 via5_6_400_2800_5_1_600_600 ;
      VIA 199.14 103.4 via4_5_400_2800_5_1_600_600 ;
      VIA 199.14 63.4 via6_7_400_2800_4_1_600_600 ;
      VIA 199.14 63.4 via5_6_400_2800_5_1_600_600 ;
      VIA 199.14 63.4 via4_5_400_2800_5_1_600_600 ;
      VIA 199.14 23.4 via6_7_400_2800_4_1_600_600 ;
      VIA 199.14 23.4 via5_6_400_2800_5_1_600_600 ;
      VIA 199.14 23.4 via4_5_400_2800_5_1_600_600 ;
      VIA 143.14 303.4 via6_7_400_2800_4_1_600_600 ;
      VIA 143.14 303.4 via5_6_400_2800_5_1_600_600 ;
      VIA 143.14 303.4 via4_5_400_2800_5_1_600_600 ;
      VIA 143.14 263.4 via6_7_400_2800_4_1_600_600 ;
      VIA 143.14 263.4 via5_6_400_2800_5_1_600_600 ;
      VIA 143.14 263.4 via4_5_400_2800_5_1_600_600 ;
      VIA 143.14 223.4 via6_7_400_2800_4_1_600_600 ;
      VIA 143.14 223.4 via5_6_400_2800_5_1_600_600 ;
      VIA 143.14 223.4 via4_5_400_2800_5_1_600_600 ;
      VIA 143.14 183.4 via6_7_400_2800_4_1_600_600 ;
      VIA 143.14 183.4 via5_6_400_2800_5_1_600_600 ;
      VIA 143.14 183.4 via4_5_400_2800_5_1_600_600 ;
      VIA 143.14 143.4 via6_7_400_2800_4_1_600_600 ;
      VIA 143.14 143.4 via5_6_400_2800_5_1_600_600 ;
      VIA 143.14 143.4 via4_5_400_2800_5_1_600_600 ;
      VIA 143.14 103.4 via6_7_400_2800_4_1_600_600 ;
      VIA 143.14 103.4 via5_6_400_2800_5_1_600_600 ;
      VIA 143.14 103.4 via4_5_400_2800_5_1_600_600 ;
      VIA 143.14 63.4 via6_7_400_2800_4_1_600_600 ;
      VIA 143.14 63.4 via5_6_400_2800_5_1_600_600 ;
      VIA 143.14 63.4 via4_5_400_2800_5_1_600_600 ;
      VIA 143.14 23.4 via6_7_400_2800_4_1_600_600 ;
      VIA 143.14 23.4 via5_6_400_2800_5_1_600_600 ;
      VIA 143.14 23.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 303.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 303.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 303.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 263.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 263.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 263.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 223.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 223.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 223.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 183.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 183.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 183.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 143.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 143.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 143.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 103.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 103.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 103.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 63.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 63.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 63.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 23.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 23.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 23.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 303.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 303.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 303.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 263.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 263.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 263.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 223.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 223.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 223.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 183.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 183.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 183.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 143.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 143.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 143.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 103.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 103.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 103.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 63.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 63.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 63.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 23.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 23.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 23.4 via4_5_400_2800_5_1_600_600 ;
      VIA 311.14 338.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 338.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 338.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 336 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 336 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 336 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 333.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 333.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 333.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 330.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 330.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 330.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 327.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 327.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 327.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 324.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 324.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 324.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 322 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 322 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 322 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 319.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 319.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 319.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 316.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 316.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 316.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 313.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 313.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 313.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 310.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 310.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 310.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 308 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 308 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 308 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 305.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 305.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 305.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 302.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 302.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 302.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 299.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 299.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 299.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 296.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 296.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 296.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 294 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 294 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 294 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 291.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 291.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 291.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 288.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 288.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 288.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 285.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 285.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 285.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 282.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 282.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 282.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 280 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 280 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 280 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 277.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 277.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 277.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 274.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 274.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 274.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 271.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 271.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 271.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 268.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 268.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 268.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 266 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 266 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 266 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 263.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 263.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 263.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 260.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 260.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 260.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 257.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 257.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 257.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 254.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 254.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 254.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 252 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 252 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 252 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 249.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 249.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 249.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 246.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 246.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 246.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 243.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 243.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 243.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 240.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 240.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 240.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 238 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 238 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 238 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 235.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 235.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 235.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 232.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 232.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 232.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 229.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 229.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 229.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 226.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 226.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 226.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 224 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 224 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 224 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 221.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 221.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 221.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 218.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 218.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 218.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 215.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 215.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 215.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 212.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 212.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 212.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 210 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 210 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 210 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 207.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 207.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 207.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 204.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 204.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 204.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 201.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 201.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 201.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 198.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 198.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 198.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 196 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 196 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 196 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 193.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 193.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 193.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 190.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 190.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 190.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 187.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 187.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 187.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 184.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 184.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 184.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 182 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 182 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 182 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 179.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 179.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 179.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 176.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 176.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 176.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 173.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 173.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 173.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 170.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 170.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 170.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 168 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 168 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 168 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 165.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 165.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 165.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 162.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 162.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 162.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 159.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 159.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 159.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 156.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 156.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 156.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 154 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 154 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 154 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 151.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 151.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 151.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 148.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 148.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 148.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 145.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 145.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 145.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 142.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 142.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 142.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 140 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 140 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 140 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 137.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 137.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 137.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 134.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 134.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 134.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 131.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 131.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 131.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 128.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 128.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 128.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 126 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 126 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 126 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 123.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 123.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 123.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 120.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 120.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 120.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 117.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 117.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 117.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 114.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 114.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 114.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 112 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 112 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 112 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 109.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 109.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 109.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 106.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 106.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 106.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 103.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 103.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 103.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 100.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 100.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 100.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 98 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 98 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 98 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 95.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 95.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 95.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 92.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 92.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 92.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 89.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 89.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 89.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 86.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 86.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 86.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 84 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 84 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 84 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 81.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 81.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 81.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 78.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 78.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 78.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 75.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 75.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 75.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 72.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 72.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 72.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 70 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 70 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 70 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 67.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 67.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 67.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 64.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 64.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 64.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 61.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 61.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 61.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 58.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 58.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 58.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 56 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 56 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 56 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 53.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 53.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 53.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 50.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 50.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 50.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 47.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 47.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 47.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 44.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 44.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 44.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 42 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 42 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 42 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 39.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 39.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 39.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 36.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 36.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 36.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 33.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 33.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 33.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 30.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 30.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 30.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 28 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 28 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 28 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 25.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 25.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 25.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 22.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 22.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 22.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 19.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 19.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 19.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 16.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 16.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 16.8 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 14 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 14 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 14 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 11.2 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 11.2 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 11.2 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 8.4 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 8.4 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 8.4 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 5.6 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 5.6 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 5.6 via1_2_400_200_1_1_300_300 ;
      VIA 311.14 2.8 via3_4_400_200_1_1_320_320 ;
      VIA 311.14 2.8 via2_3_400_200_1_1_320_320 ;
      VIA 311.14 2.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 338.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 338.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 338.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 336 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 336 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 336 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 333.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 333.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 333.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 330.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 330.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 330.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 327.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 327.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 327.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 324.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 324.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 324.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 322 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 322 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 322 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 319.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 319.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 319.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 316.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 316.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 316.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 313.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 313.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 313.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 310.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 310.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 310.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 308 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 308 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 308 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 305.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 305.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 305.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 302.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 302.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 302.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 299.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 299.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 299.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 296.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 296.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 296.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 294 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 294 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 294 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 291.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 291.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 291.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 288.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 288.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 288.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 285.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 285.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 285.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 282.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 282.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 282.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 280 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 280 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 280 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 277.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 277.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 277.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 274.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 274.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 274.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 271.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 271.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 271.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 268.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 268.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 268.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 266 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 266 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 266 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 263.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 263.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 263.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 260.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 260.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 260.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 257.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 257.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 257.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 254.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 254.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 254.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 252 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 252 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 252 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 249.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 249.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 249.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 246.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 246.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 246.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 243.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 243.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 243.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 240.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 240.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 240.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 238 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 238 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 238 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 235.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 235.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 235.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 232.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 232.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 232.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 229.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 229.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 229.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 226.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 226.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 226.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 224 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 224 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 224 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 221.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 221.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 221.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 218.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 218.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 218.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 215.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 215.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 215.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 212.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 212.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 212.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 210 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 210 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 210 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 207.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 207.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 207.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 204.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 204.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 204.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 201.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 201.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 201.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 198.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 198.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 198.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 196 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 196 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 196 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 193.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 193.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 193.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 190.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 190.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 190.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 187.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 187.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 187.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 184.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 184.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 184.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 182 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 182 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 182 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 179.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 179.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 179.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 176.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 176.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 176.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 173.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 173.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 173.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 170.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 170.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 170.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 168 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 168 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 168 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 165.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 165.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 165.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 162.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 162.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 162.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 159.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 159.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 159.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 156.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 156.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 156.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 154 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 154 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 154 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 151.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 151.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 151.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 148.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 148.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 148.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 145.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 145.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 145.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 142.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 142.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 142.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 140 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 140 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 140 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 137.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 137.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 137.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 134.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 134.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 134.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 131.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 131.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 131.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 128.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 128.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 128.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 126 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 126 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 126 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 123.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 123.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 123.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 120.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 120.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 120.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 117.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 117.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 117.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 114.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 114.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 114.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 112 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 112 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 112 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 109.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 109.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 109.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 106.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 106.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 106.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 103.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 103.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 103.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 100.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 100.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 100.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 98 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 98 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 98 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 95.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 95.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 95.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 92.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 92.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 92.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 89.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 89.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 89.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 86.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 86.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 86.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 84 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 84 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 84 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 81.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 81.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 81.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 78.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 78.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 78.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 75.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 75.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 75.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 72.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 72.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 72.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 70 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 70 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 70 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 67.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 67.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 67.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 64.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 64.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 64.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 61.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 61.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 61.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 58.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 58.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 58.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 56 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 56 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 56 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 53.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 53.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 53.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 50.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 50.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 50.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 47.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 47.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 47.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 44.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 44.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 44.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 42 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 42 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 42 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 39.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 39.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 39.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 36.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 36.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 36.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 33.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 33.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 33.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 30.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 30.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 30.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 28 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 28 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 28 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 25.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 25.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 25.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 22.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 22.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 22.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 19.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 19.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 19.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 16.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 16.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 16.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 14 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 14 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 14 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 11.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 11.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 11.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 8.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 8.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 8.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 5.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 5.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 5.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 2.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 2.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 2.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 338.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 338.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 338.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 336 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 336 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 336 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 333.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 333.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 333.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 330.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 330.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 330.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 327.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 327.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 327.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 324.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 324.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 324.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 322 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 322 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 322 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 319.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 319.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 319.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 316.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 316.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 316.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 313.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 313.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 313.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 310.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 310.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 310.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 308 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 308 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 308 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 305.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 305.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 305.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 302.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 302.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 302.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 299.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 299.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 299.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 296.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 296.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 296.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 294 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 294 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 294 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 291.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 291.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 291.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 288.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 288.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 288.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 285.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 285.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 285.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 282.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 282.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 282.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 280 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 280 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 280 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 277.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 277.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 277.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 274.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 274.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 274.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 271.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 271.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 271.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 268.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 268.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 268.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 266 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 266 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 266 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 263.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 263.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 263.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 260.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 260.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 260.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 257.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 257.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 257.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 254.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 254.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 254.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 252 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 252 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 252 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 249.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 249.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 249.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 246.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 246.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 246.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 243.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 243.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 243.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 240.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 240.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 240.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 238 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 238 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 238 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 235.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 235.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 235.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 232.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 232.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 232.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 229.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 229.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 229.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 226.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 226.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 226.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 224 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 224 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 224 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 221.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 221.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 221.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 218.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 218.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 218.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 215.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 215.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 215.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 212.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 212.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 212.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 210 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 210 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 210 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 207.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 207.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 207.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 204.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 204.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 204.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 201.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 201.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 201.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 198.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 198.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 198.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 196 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 196 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 196 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 193.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 193.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 193.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 190.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 190.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 190.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 187.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 187.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 187.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 184.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 184.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 184.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 182 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 182 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 182 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 179.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 179.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 179.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 176.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 176.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 176.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 173.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 173.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 173.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 170.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 170.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 170.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 168 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 168 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 168 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 165.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 165.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 165.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 162.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 162.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 162.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 159.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 159.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 159.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 156.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 156.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 156.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 154 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 154 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 154 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 151.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 151.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 151.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 148.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 148.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 148.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 145.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 145.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 145.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 142.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 142.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 142.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 140 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 140 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 140 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 137.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 137.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 137.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 134.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 134.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 134.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 131.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 131.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 131.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 128.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 128.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 128.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 126 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 126 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 126 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 123.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 123.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 123.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 120.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 120.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 120.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 117.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 117.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 117.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 114.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 114.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 114.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 112 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 112 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 112 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 109.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 109.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 109.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 106.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 106.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 106.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 103.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 103.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 103.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 100.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 100.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 100.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 98 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 98 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 98 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 95.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 95.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 95.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 92.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 92.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 92.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 89.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 89.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 89.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 86.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 86.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 86.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 84 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 84 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 84 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 81.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 81.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 81.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 78.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 78.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 78.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 75.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 75.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 75.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 72.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 72.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 72.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 70 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 70 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 70 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 67.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 67.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 67.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 64.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 64.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 64.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 61.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 61.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 61.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 58.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 58.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 58.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 56 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 56 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 56 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 53.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 53.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 53.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 50.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 50.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 50.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 47.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 47.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 47.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 44.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 44.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 44.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 42 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 42 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 42 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 39.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 39.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 39.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 36.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 36.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 36.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 33.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 33.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 33.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 30.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 30.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 30.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 28 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 28 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 28 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 25.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 25.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 25.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 22.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 22.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 22.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 19.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 19.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 19.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 16.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 16.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 16.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 14 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 14 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 14 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 11.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 11.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 11.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 8.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 8.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 8.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 5.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 5.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 5.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 2.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 2.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 2.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 338.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 338.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 338.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 336 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 336 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 336 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 333.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 333.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 333.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 330.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 330.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 330.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 327.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 327.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 327.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 324.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 324.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 324.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 322 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 322 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 322 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 319.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 319.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 319.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 316.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 316.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 316.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 313.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 313.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 313.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 310.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 310.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 310.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 308 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 308 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 308 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 305.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 305.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 305.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 302.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 302.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 302.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 299.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 299.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 299.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 296.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 296.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 296.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 294 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 294 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 294 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 291.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 291.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 291.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 288.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 288.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 288.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 285.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 285.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 285.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 282.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 282.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 282.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 280 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 280 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 280 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 277.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 277.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 277.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 274.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 274.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 274.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 271.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 271.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 271.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 268.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 268.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 268.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 266 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 266 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 266 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 263.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 263.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 263.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 260.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 260.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 260.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 257.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 257.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 257.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 254.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 254.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 254.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 252 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 252 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 252 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 249.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 249.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 249.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 246.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 246.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 246.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 243.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 243.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 243.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 240.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 240.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 240.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 238 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 238 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 238 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 235.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 235.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 235.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 232.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 232.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 232.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 229.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 229.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 229.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 226.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 226.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 226.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 224 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 224 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 224 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 221.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 221.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 221.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 218.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 218.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 218.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 215.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 215.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 215.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 212.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 212.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 212.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 210 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 210 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 210 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 207.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 207.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 207.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 204.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 204.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 204.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 201.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 201.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 201.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 198.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 198.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 198.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 196 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 196 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 196 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 193.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 193.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 193.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 190.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 190.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 190.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 187.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 187.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 187.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 184.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 184.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 184.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 182 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 182 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 182 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 179.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 179.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 179.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 176.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 176.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 176.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 173.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 173.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 173.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 170.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 170.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 170.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 168 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 168 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 168 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 165.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 165.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 165.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 162.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 162.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 162.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 159.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 159.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 159.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 156.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 156.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 156.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 154 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 154 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 154 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 151.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 151.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 151.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 148.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 148.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 148.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 145.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 145.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 145.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 142.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 142.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 142.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 140 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 140 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 140 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 137.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 137.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 137.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 134.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 134.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 134.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 131.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 131.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 131.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 128.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 128.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 128.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 126 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 126 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 126 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 123.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 123.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 123.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 120.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 120.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 120.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 117.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 117.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 117.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 114.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 114.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 114.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 112 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 112 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 112 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 109.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 109.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 109.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 106.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 106.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 106.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 103.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 103.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 103.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 100.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 100.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 100.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 98 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 98 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 98 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 95.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 95.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 95.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 92.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 92.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 92.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 89.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 89.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 89.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 86.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 86.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 86.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 84 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 84 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 84 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 81.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 81.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 81.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 78.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 78.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 78.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 75.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 75.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 75.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 72.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 72.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 72.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 70 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 70 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 70 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 67.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 67.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 67.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 64.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 64.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 64.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 61.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 61.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 61.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 58.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 58.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 58.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 56 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 56 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 56 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 53.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 53.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 53.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 50.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 50.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 50.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 47.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 47.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 47.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 44.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 44.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 44.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 42 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 42 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 42 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 39.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 39.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 39.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 36.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 36.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 36.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 33.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 33.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 33.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 30.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 30.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 30.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 28 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 28 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 28 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 25.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 25.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 25.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 22.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 22.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 22.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 19.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 19.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 19.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 16.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 16.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 16.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 14 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 14 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 14 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 11.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 11.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 11.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 8.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 8.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 8.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 5.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 5.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 5.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 2.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 2.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 2.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 338.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 338.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 338.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 336 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 336 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 336 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 333.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 333.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 333.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 330.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 330.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 330.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 327.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 327.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 327.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 324.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 324.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 324.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 322 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 322 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 322 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 319.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 319.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 319.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 316.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 316.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 316.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 313.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 313.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 313.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 310.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 310.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 310.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 308 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 308 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 308 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 305.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 305.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 305.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 302.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 302.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 302.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 299.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 299.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 299.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 296.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 296.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 296.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 294 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 294 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 294 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 291.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 291.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 291.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 288.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 288.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 288.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 285.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 285.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 285.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 282.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 282.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 282.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 280 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 280 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 280 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 277.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 277.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 277.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 274.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 274.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 274.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 271.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 271.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 271.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 268.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 268.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 268.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 266 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 266 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 266 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 263.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 263.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 263.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 260.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 260.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 260.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 257.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 257.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 257.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 254.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 254.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 254.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 252 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 252 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 252 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 249.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 249.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 249.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 246.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 246.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 246.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 243.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 243.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 243.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 240.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 240.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 240.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 238 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 238 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 238 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 235.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 235.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 235.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 232.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 232.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 232.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 229.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 229.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 229.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 226.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 226.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 226.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 224 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 224 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 224 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 221.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 221.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 221.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 218.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 218.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 218.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 215.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 215.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 215.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 212.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 212.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 212.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 210 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 210 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 210 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 207.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 207.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 207.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 204.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 204.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 204.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 201.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 201.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 201.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 198.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 198.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 198.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 196 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 196 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 196 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 193.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 193.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 193.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 190.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 190.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 190.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 187.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 187.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 187.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 184.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 184.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 184.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 182 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 182 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 182 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 179.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 179.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 179.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 176.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 176.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 176.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 173.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 173.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 173.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 170.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 170.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 170.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 168 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 168 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 168 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 165.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 165.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 165.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 162.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 162.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 162.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 159.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 159.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 159.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 156.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 156.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 156.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 154 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 154 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 154 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 151.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 151.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 151.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 148.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 148.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 148.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 145.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 145.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 145.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 142.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 142.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 142.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 140 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 140 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 140 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 137.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 137.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 137.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 134.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 134.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 134.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 131.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 131.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 131.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 128.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 128.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 128.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 126 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 126 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 126 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 123.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 123.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 123.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 120.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 120.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 120.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 117.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 117.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 117.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 114.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 114.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 114.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 112 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 112 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 112 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 109.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 109.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 109.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 106.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 106.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 106.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 103.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 103.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 103.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 100.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 100.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 100.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 98 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 98 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 98 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 95.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 95.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 95.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 92.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 92.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 92.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 89.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 89.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 89.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 86.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 86.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 86.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 84 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 84 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 84 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 81.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 81.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 81.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 78.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 78.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 78.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 75.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 75.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 75.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 72.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 72.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 72.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 70 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 70 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 70 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 67.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 67.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 67.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 64.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 64.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 64.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 61.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 61.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 61.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 58.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 58.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 58.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 56 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 56 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 56 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 53.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 53.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 53.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 50.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 50.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 50.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 47.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 47.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 47.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 44.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 44.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 44.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 42 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 42 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 42 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 39.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 39.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 39.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 36.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 36.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 36.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 33.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 33.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 33.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 30.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 30.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 30.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 28 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 28 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 28 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 25.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 25.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 25.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 22.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 22.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 22.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 19.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 19.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 19.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 16.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 16.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 16.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 14 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 14 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 14 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 11.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 11.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 11.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 8.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 8.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 8.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 5.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 5.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 5.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 2.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 2.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 2.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 338.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 338.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 338.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 336 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 336 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 336 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 333.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 333.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 333.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 330.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 330.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 330.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 327.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 327.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 327.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 324.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 324.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 324.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 322 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 322 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 322 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 319.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 319.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 319.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 316.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 316.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 316.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 313.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 313.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 313.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 310.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 310.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 310.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 308 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 308 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 308 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 305.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 305.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 305.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 302.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 302.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 302.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 299.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 299.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 299.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 296.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 296.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 296.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 294 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 294 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 294 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 291.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 291.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 291.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 288.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 288.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 288.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 285.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 285.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 285.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 282.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 282.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 282.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 280 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 280 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 280 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 277.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 277.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 277.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 274.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 274.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 274.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 271.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 271.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 271.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 268.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 268.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 268.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 266 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 266 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 266 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 263.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 263.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 263.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 260.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 260.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 260.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 257.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 257.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 257.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 254.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 254.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 254.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 252 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 252 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 252 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 249.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 249.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 249.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 246.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 246.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 246.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 243.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 243.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 243.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 240.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 240.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 240.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 238 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 238 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 238 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 235.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 235.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 235.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 232.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 232.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 232.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 229.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 229.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 229.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 226.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 226.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 226.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 224 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 224 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 224 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 221.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 221.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 221.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 218.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 218.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 218.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 215.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 215.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 215.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 212.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 212.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 212.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 210 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 210 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 210 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 207.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 207.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 207.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 204.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 204.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 204.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 201.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 201.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 201.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 198.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 198.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 198.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 196 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 196 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 196 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 193.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 193.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 193.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 190.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 190.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 190.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 187.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 187.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 187.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 184.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 184.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 184.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 182 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 182 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 182 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 179.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 179.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 179.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 176.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 176.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 176.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 173.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 173.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 173.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 170.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 170.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 170.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 168 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 168 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 168 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 165.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 165.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 165.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 162.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 162.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 162.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 159.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 159.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 159.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 156.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 156.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 156.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 154 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 154 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 154 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 151.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 151.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 151.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 148.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 148.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 148.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 145.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 145.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 145.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 142.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 142.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 142.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 140 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 140 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 140 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 137.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 137.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 137.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 134.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 134.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 134.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 131.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 131.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 131.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 128.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 128.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 128.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 126 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 126 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 126 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 123.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 123.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 123.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 120.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 120.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 120.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 117.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 117.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 117.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 114.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 114.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 114.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 112 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 112 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 112 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 109.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 109.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 109.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 106.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 106.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 106.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 103.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 103.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 103.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 100.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 100.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 100.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 98 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 98 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 98 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 95.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 95.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 95.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 92.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 92.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 92.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 89.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 89.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 89.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 86.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 86.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 86.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 84 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 84 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 84 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 81.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 81.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 81.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 78.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 78.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 78.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 75.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 75.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 75.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 72.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 72.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 72.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 70 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 70 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 70 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 67.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 67.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 67.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 64.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 64.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 64.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 61.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 61.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 61.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 58.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 58.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 58.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 56 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 56 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 56 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 53.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 53.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 53.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 50.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 50.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 50.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 47.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 47.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 47.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 44.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 44.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 44.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 42 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 42 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 42 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 39.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 39.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 39.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 36.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 36.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 36.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 33.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 33.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 33.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 30.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 30.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 30.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 28 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 28 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 28 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 25.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 25.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 25.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 22.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 22.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 22.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 19.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 19.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 19.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 16.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 16.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 16.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 14 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 14 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 14 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 11.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 11.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 11.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 8.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 8.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 8.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 5.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 5.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 5.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 2.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 2.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 2.8 via1_2_400_200_1_1_300_300 ;
    END
  END VDD
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 209.44 0.14 209.58 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  78.985 0 79.125 0.14 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 104.72 0.14 104.86 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  261.545 0 261.685 0.14 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  26.345 340.58 26.485 340.72 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  340.58 131.04 340.72 131.18 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  287.865 340.58 288.005 340.72 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 339.92 0.14 340.06 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  340.58 26.32 340.72 26.46 ;
    END
  END addr[8]
  PIN ce
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  235.785 340.58 235.925 340.72 ;
    END
  END ce
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  340.58 0.56 340.72 0.7 ;
    END
  END clk
  PIN di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  183.145 0 183.285 0.14 ;
    END
  END di[0]
  PIN di[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  340.58 52.64 340.72 52.78 ;
    END
  END di[10]
  PIN di[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  52.665 340.58 52.805 340.72 ;
    END
  END di[11]
  PIN di[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  340.58 78.96 340.72 79.1 ;
    END
  END di[12]
  PIN di[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 261.52 0.14 261.66 ;
    END
  END di[13]
  PIN di[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  157.385 340.58 157.525 340.72 ;
    END
  END di[14]
  PIN di[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  235.785 0 235.925 0.14 ;
    END
  END di[15]
  PIN di[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  287.865 0 288.005 0.14 ;
    END
  END di[16]
  PIN di[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 287.84 0.14 287.98 ;
    END
  END di[17]
  PIN di[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 157.36 0.14 157.5 ;
    END
  END di[18]
  PIN di[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 183.12 0.14 183.26 ;
    END
  END di[19]
  PIN di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  340.58 235.76 340.72 235.9 ;
    END
  END di[1]
  PIN di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 52.64 0.14 52.78 ;
    END
  END di[2]
  PIN di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  209.465 340.58 209.605 340.72 ;
    END
  END di[3]
  PIN di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  131.065 340.58 131.205 340.72 ;
    END
  END di[4]
  PIN di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  340.58 314.16 340.72 314.3 ;
    END
  END di[5]
  PIN di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  340.58 261.52 340.72 261.66 ;
    END
  END di[6]
  PIN di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  340.58 183.12 340.72 183.26 ;
    END
  END di[7]
  PIN di[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  261.545 340.58 261.685 340.72 ;
    END
  END di[8]
  PIN di[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  26.345 0 26.485 0.14 ;
    END
  END di[9]
  PIN doq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  0.585 0 0.725 0.14 ;
    END
  END doq[0]
  PIN doq[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 78.96 0.14 79.1 ;
    END
  END doq[10]
  PIN doq[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  340.58 287.84 340.72 287.98 ;
    END
  END doq[11]
  PIN doq[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  131.065 0 131.205 0.14 ;
    END
  END doq[12]
  PIN doq[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  340.58 209.44 340.72 209.58 ;
    END
  END doq[13]
  PIN doq[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  314.185 0 314.325 0.14 ;
    END
  END doq[14]
  PIN doq[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  183.145 340.58 183.285 340.72 ;
    END
  END doq[15]
  PIN doq[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  340.58 104.72 340.72 104.86 ;
    END
  END doq[16]
  PIN doq[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  52.665 0 52.805 0.14 ;
    END
  END doq[17]
  PIN doq[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  104.745 0 104.885 0.14 ;
    END
  END doq[18]
  PIN doq[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 235.76 0.14 235.9 ;
    END
  END doq[19]
  PIN doq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 26.32 0.14 26.46 ;
    END
  END doq[1]
  PIN doq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  157.385 0 157.525 0.14 ;
    END
  END doq[2]
  PIN doq[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  339.945 340.58 340.085 340.72 ;
    END
  END doq[3]
  PIN doq[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  314.185 340.58 314.325 340.72 ;
    END
  END doq[4]
  PIN doq[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  78.985 340.58 79.125 340.72 ;
    END
  END doq[5]
  PIN doq[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  104.745 340.58 104.885 340.72 ;
    END
  END doq[6]
  PIN doq[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  209.465 0 209.605 0.14 ;
    END
  END doq[7]
  PIN doq[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 131.04 0.14 131.18 ;
    END
  END doq[8]
  PIN doq[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 314.16 0.14 314.3 ;
    END
  END doq[9]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  340.58 157.36 340.72 157.5 ;
    END
  END we
  OBS
    LAYER metal1 ;
     RECT  0 0 340.72 340.72 ;
    LAYER metal2 ;
     RECT  0 0 340.72 340.72 ;
    LAYER metal3 ;
     RECT  0 0 340.72 340.72 ;
    LAYER metal4 ;
     RECT  0 0 340.72 340.72 ;
    LAYER metal5 ;
     RECT  0 0 340.72 340.72 ;
    LAYER metal6 ;
     RECT  0 0 340.72 340.72 ;
    LAYER metal7 ;
     RECT  0 0 340.72 340.72 ;
    LAYER metal8 ;
     RECT  0 0 340.72 340.72 ;
    LAYER metal9 ;
     RECT  0 0 340.72 340.72 ;
  END
END or1200_spram2
END LIBRARY
