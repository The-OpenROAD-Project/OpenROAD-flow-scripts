(* blackbox *) module A2O1A1Ixp33_ASAP7_75t_L (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module A2O1A1O1Ixp25_ASAP7_75t_L (Y, A1, A2, B, C, D);
	output Y;
	input A1, A2, B, C, D;
endmodule
(* blackbox *) module AO211x2_ASAP7_75t_L (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module AO21x1_ASAP7_75t_L (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AO21x2_ASAP7_75t_L (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AO221x1_ASAP7_75t_L (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module AO221x2_ASAP7_75t_L (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module AO222x2_ASAP7_75t_L (Y, A1, A2, B1, B2, C1, C2);
	output Y;
	input A1, A2, B1, B2, C1, C2;
endmodule
(* blackbox *) module AO22x1_ASAP7_75t_L (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AO22x2_ASAP7_75t_L (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AO31x2_ASAP7_75t_L (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module AO322x2_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, C1, C2;
endmodule
(* blackbox *) module AO32x1_ASAP7_75t_L (Y, A1, A2, A3, B1, B2);
	output Y;
	input A1, A2, A3, B1, B2;
endmodule
(* blackbox *) module AO32x2_ASAP7_75t_L (Y, A1, A2, A3, B1, B2);
	output Y;
	input A1, A2, A3, B1, B2;
endmodule
(* blackbox *) module AO331x1_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C);
	output Y;
	input A1, A2, A3, B1, B2, B3, C;
endmodule
(* blackbox *) module AO331x2_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C);
	output Y;
	input A1, A2, A3, B1, B2, B3, C;
endmodule
(* blackbox *) module AO332x1_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module AO332x2_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module AO333x1_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module AO333x2_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module AO33x2_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3);
	output Y;
	input A1, A2, A3, B1, B2, B3;
endmodule
(* blackbox *) module AOI211x1_ASAP7_75t_L (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module AOI211xp5_ASAP7_75t_L (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module AOI21x1_ASAP7_75t_L (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AOI21xp33_ASAP7_75t_L (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AOI21xp5_ASAP7_75t_L (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AOI221x1_ASAP7_75t_L (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module AOI221xp5_ASAP7_75t_L (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module AOI222xp33_ASAP7_75t_L (Y, A1, A2, B1, B2, C1, C2);
	output Y;
	input A1, A2, B1, B2, C1, C2;
endmodule
(* blackbox *) module AOI22x1_ASAP7_75t_L (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AOI22xp33_ASAP7_75t_L (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AOI22xp5_ASAP7_75t_L (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AOI311xp33_ASAP7_75t_L (Y, A1, A2, A3, B, C);
	output Y;
	input A1, A2, A3, B, C;
endmodule
(* blackbox *) module AOI31xp33_ASAP7_75t_L (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module AOI31xp67_ASAP7_75t_L (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module AOI321xp33_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, C);
	output Y;
	input A1, A2, A3, B1, B2, C;
endmodule
(* blackbox *) module AOI322xp5_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, C1, C2;
endmodule
(* blackbox *) module AOI32xp33_ASAP7_75t_L (Y, A1, A2, A3, B1, B2);
	output Y;
	input A1, A2, A3, B1, B2;
endmodule
(* blackbox *) module AOI331xp33_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C1);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1;
endmodule
(* blackbox *) module AOI332xp33_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module AOI333xp33_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module AOI33xp33_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3);
	output Y;
	input A1, A2, A3, B1, B2, B3;
endmodule
