module RegisterFile(
  input         clock,
  input  [6:0]  io_read_0_address,
                io_read_1_address,
                io_read_2_address,
                io_read_3_address,
                io_read_4_address,
                io_read_5_address,
                io_read_6_address,
                io_read_7_address,
  input         io_write_0_write,
  input  [6:0]  io_write_0_address,
  input  [63:0] io_write_0_value,
  input         io_write_0_byteMask_0,
                io_write_0_byteMask_1,
                io_write_0_byteMask_2,
                io_write_0_byteMask_3,
                io_write_0_byteMask_4,
                io_write_0_byteMask_5,
                io_write_0_byteMask_6,
                io_write_0_byteMask_7,
                io_write_1_write,
  input  [6:0]  io_write_1_address,
  input  [63:0] io_write_1_value,
  input         io_write_1_byteMask_0,
                io_write_1_byteMask_1,
                io_write_1_byteMask_2,
                io_write_1_byteMask_3,
                io_write_1_byteMask_4,
                io_write_1_byteMask_5,
                io_write_1_byteMask_6,
                io_write_1_byteMask_7,
                io_write_2_write,
  input  [6:0]  io_write_2_address,
  input  [63:0] io_write_2_value,
  input         io_write_2_byteMask_0,
                io_write_2_byteMask_1,
                io_write_2_byteMask_2,
                io_write_2_byteMask_3,
                io_write_2_byteMask_4,
                io_write_2_byteMask_5,
                io_write_2_byteMask_6,
                io_write_2_byteMask_7,
                io_write_3_write,
  input  [6:0]  io_write_3_address,
  input  [63:0] io_write_3_value,
  input         io_write_3_byteMask_0,
                io_write_3_byteMask_1,
                io_write_3_byteMask_2,
                io_write_3_byteMask_3,
                io_write_3_byteMask_4,
                io_write_3_byteMask_5,
                io_write_3_byteMask_6,
                io_write_3_byteMask_7,
  output [63:0] io_read_0_value,
                io_read_1_value,
                io_read_2_value,
                io_read_3_value,
                io_read_4_value,
                io_read_5_value,
                io_read_6_value,
                io_read_7_value
);

  wire [63:0] _registers_15_ext_R0_data;
  wire [63:0] _registers_15_ext_R1_data;
  wire [63:0] _registers_15_ext_R2_data;
  wire [63:0] _registers_15_ext_R3_data;
  wire [63:0] _registers_15_ext_R4_data;
  wire [63:0] _registers_15_ext_R5_data;
  wire [63:0] _registers_15_ext_R6_data;
  wire [63:0] _registers_15_ext_R7_data;
  wire [63:0] _registers_14_ext_R0_data;
  wire [63:0] _registers_14_ext_R1_data;
  wire [63:0] _registers_14_ext_R2_data;
  wire [63:0] _registers_14_ext_R3_data;
  wire [63:0] _registers_14_ext_R4_data;
  wire [63:0] _registers_14_ext_R5_data;
  wire [63:0] _registers_14_ext_R6_data;
  wire [63:0] _registers_14_ext_R7_data;
  wire [63:0] _registers_13_ext_R0_data;
  wire [63:0] _registers_13_ext_R1_data;
  wire [63:0] _registers_13_ext_R2_data;
  wire [63:0] _registers_13_ext_R3_data;
  wire [63:0] _registers_13_ext_R4_data;
  wire [63:0] _registers_13_ext_R5_data;
  wire [63:0] _registers_13_ext_R6_data;
  wire [63:0] _registers_13_ext_R7_data;
  wire [63:0] _registers_12_ext_R0_data;
  wire [63:0] _registers_12_ext_R1_data;
  wire [63:0] _registers_12_ext_R2_data;
  wire [63:0] _registers_12_ext_R3_data;
  wire [63:0] _registers_12_ext_R4_data;
  wire [63:0] _registers_12_ext_R5_data;
  wire [63:0] _registers_12_ext_R6_data;
  wire [63:0] _registers_12_ext_R7_data;
  wire [63:0] _registers_11_ext_R0_data;
  wire [63:0] _registers_11_ext_R1_data;
  wire [63:0] _registers_11_ext_R2_data;
  wire [63:0] _registers_11_ext_R3_data;
  wire [63:0] _registers_11_ext_R4_data;
  wire [63:0] _registers_11_ext_R5_data;
  wire [63:0] _registers_11_ext_R6_data;
  wire [63:0] _registers_11_ext_R7_data;
  wire [63:0] _registers_10_ext_R0_data;
  wire [63:0] _registers_10_ext_R1_data;
  wire [63:0] _registers_10_ext_R2_data;
  wire [63:0] _registers_10_ext_R3_data;
  wire [63:0] _registers_10_ext_R4_data;
  wire [63:0] _registers_10_ext_R5_data;
  wire [63:0] _registers_10_ext_R6_data;
  wire [63:0] _registers_10_ext_R7_data;
  wire [63:0] _registers_9_ext_R0_data;
  wire [63:0] _registers_9_ext_R1_data;
  wire [63:0] _registers_9_ext_R2_data;
  wire [63:0] _registers_9_ext_R3_data;
  wire [63:0] _registers_9_ext_R4_data;
  wire [63:0] _registers_9_ext_R5_data;
  wire [63:0] _registers_9_ext_R6_data;
  wire [63:0] _registers_9_ext_R7_data;
  wire [63:0] _registers_8_ext_R0_data;
  wire [63:0] _registers_8_ext_R1_data;
  wire [63:0] _registers_8_ext_R2_data;
  wire [63:0] _registers_8_ext_R3_data;
  wire [63:0] _registers_8_ext_R4_data;
  wire [63:0] _registers_8_ext_R5_data;
  wire [63:0] _registers_8_ext_R6_data;
  wire [63:0] _registers_8_ext_R7_data;
  wire [63:0] _registers_7_ext_R0_data;
  wire [63:0] _registers_7_ext_R1_data;
  wire [63:0] _registers_7_ext_R2_data;
  wire [63:0] _registers_7_ext_R3_data;
  wire [63:0] _registers_7_ext_R4_data;
  wire [63:0] _registers_7_ext_R5_data;
  wire [63:0] _registers_7_ext_R6_data;
  wire [63:0] _registers_7_ext_R7_data;
  wire [63:0] _registers_6_ext_R0_data;
  wire [63:0] _registers_6_ext_R1_data;
  wire [63:0] _registers_6_ext_R2_data;
  wire [63:0] _registers_6_ext_R3_data;
  wire [63:0] _registers_6_ext_R4_data;
  wire [63:0] _registers_6_ext_R5_data;
  wire [63:0] _registers_6_ext_R6_data;
  wire [63:0] _registers_6_ext_R7_data;
  wire [63:0] _registers_5_ext_R0_data;
  wire [63:0] _registers_5_ext_R1_data;
  wire [63:0] _registers_5_ext_R2_data;
  wire [63:0] _registers_5_ext_R3_data;
  wire [63:0] _registers_5_ext_R4_data;
  wire [63:0] _registers_5_ext_R5_data;
  wire [63:0] _registers_5_ext_R6_data;
  wire [63:0] _registers_5_ext_R7_data;
  wire [63:0] _registers_4_ext_R0_data;
  wire [63:0] _registers_4_ext_R1_data;
  wire [63:0] _registers_4_ext_R2_data;
  wire [63:0] _registers_4_ext_R3_data;
  wire [63:0] _registers_4_ext_R4_data;
  wire [63:0] _registers_4_ext_R5_data;
  wire [63:0] _registers_4_ext_R6_data;
  wire [63:0] _registers_4_ext_R7_data;
  wire [63:0] _registers_3_ext_R0_data;
  wire [63:0] _registers_3_ext_R1_data;
  wire [63:0] _registers_3_ext_R2_data;
  wire [63:0] _registers_3_ext_R3_data;
  wire [63:0] _registers_3_ext_R4_data;
  wire [63:0] _registers_3_ext_R5_data;
  wire [63:0] _registers_3_ext_R6_data;
  wire [63:0] _registers_3_ext_R7_data;
  wire [63:0] _registers_2_ext_R0_data;
  wire [63:0] _registers_2_ext_R1_data;
  wire [63:0] _registers_2_ext_R2_data;
  wire [63:0] _registers_2_ext_R3_data;
  wire [63:0] _registers_2_ext_R4_data;
  wire [63:0] _registers_2_ext_R5_data;
  wire [63:0] _registers_2_ext_R6_data;
  wire [63:0] _registers_2_ext_R7_data;
  wire [63:0] _registers_1_ext_R0_data;
  wire [63:0] _registers_1_ext_R1_data;
  wire [63:0] _registers_1_ext_R2_data;
  wire [63:0] _registers_1_ext_R3_data;
  wire [63:0] _registers_1_ext_R4_data;
  wire [63:0] _registers_1_ext_R5_data;
  wire [63:0] _registers_1_ext_R6_data;
  wire [63:0] _registers_1_ext_R7_data;
  wire [63:0] _registers_0_ext_R0_data;
  wire [63:0] _registers_0_ext_R1_data;
  wire [63:0] _registers_0_ext_R2_data;
  wire [63:0] _registers_0_ext_R3_data;
  wire [63:0] _registers_0_ext_R4_data;
  wire [63:0] _registers_0_ext_R5_data;
  wire [63:0] _registers_0_ext_R6_data;
  wire [63:0] _registers_0_ext_R7_data;
  reg  [7:0]  casez_tmp;
  reg  [7:0]  casez_tmp_0;
  reg  [7:0]  casez_tmp_1;
  reg  [7:0]  casez_tmp_2;
  reg  [7:0]  casez_tmp_3;
  reg  [7:0]  casez_tmp_4;
  reg  [7:0]  casez_tmp_5;
  reg  [7:0]  casez_tmp_6;
  reg  [7:0]  casez_tmp_7;
  reg  [7:0]  casez_tmp_8;
  reg  [7:0]  casez_tmp_9;
  reg  [7:0]  casez_tmp_10;
  reg  [7:0]  casez_tmp_11;
  reg  [7:0]  casez_tmp_12;
  reg  [7:0]  casez_tmp_13;
  reg  [7:0]  casez_tmp_14;
  reg  [7:0]  casez_tmp_15;
  reg  [7:0]  casez_tmp_16;
  reg  [7:0]  casez_tmp_17;
  reg  [7:0]  casez_tmp_18;
  reg  [7:0]  casez_tmp_19;
  reg  [7:0]  casez_tmp_20;
  reg  [7:0]  casez_tmp_21;
  reg  [7:0]  casez_tmp_22;
  reg  [7:0]  casez_tmp_23;
  reg  [7:0]  casez_tmp_24;
  reg  [7:0]  casez_tmp_25;
  reg  [7:0]  casez_tmp_26;
  reg  [7:0]  casez_tmp_27;
  reg  [7:0]  casez_tmp_28;
  reg  [7:0]  casez_tmp_29;
  reg  [7:0]  casez_tmp_30;
  reg  [7:0]  casez_tmp_31;
  reg  [7:0]  casez_tmp_32;
  reg  [7:0]  casez_tmp_33;
  reg  [7:0]  casez_tmp_34;
  reg  [7:0]  casez_tmp_35;
  reg  [7:0]  casez_tmp_36;
  reg  [7:0]  casez_tmp_37;
  reg  [7:0]  casez_tmp_38;
  reg  [7:0]  casez_tmp_39;
  reg  [7:0]  casez_tmp_40;
  reg  [7:0]  casez_tmp_41;
  reg  [7:0]  casez_tmp_42;
  reg  [7:0]  casez_tmp_43;
  reg  [7:0]  casez_tmp_44;
  reg  [7:0]  casez_tmp_45;
  reg  [7:0]  casez_tmp_46;
  reg  [7:0]  casez_tmp_47;
  reg  [7:0]  casez_tmp_48;
  reg  [7:0]  casez_tmp_49;
  reg  [7:0]  casez_tmp_50;
  reg  [7:0]  casez_tmp_51;
  reg  [7:0]  casez_tmp_52;
  reg  [7:0]  casez_tmp_53;
  reg  [7:0]  casez_tmp_54;
  reg  [7:0]  casez_tmp_55;
  reg  [7:0]  casez_tmp_56;
  reg  [7:0]  casez_tmp_57;
  reg  [7:0]  casez_tmp_58;
  reg  [7:0]  casez_tmp_59;
  reg  [7:0]  casez_tmp_60;
  reg  [7:0]  casez_tmp_61;
  reg  [7:0]  casez_tmp_62;
  wire [7:0]  _GEN =
    {io_write_0_byteMask_7,
     io_write_0_byteMask_6,
     io_write_0_byteMask_5,
     io_write_0_byteMask_4,
     io_write_0_byteMask_3,
     io_write_0_byteMask_2,
     io_write_0_byteMask_1,
     io_write_0_byteMask_0};
  wire [7:0]  _GEN_0 =
    {io_write_1_byteMask_7,
     io_write_1_byteMask_6,
     io_write_1_byteMask_5,
     io_write_1_byteMask_4,
     io_write_1_byteMask_3,
     io_write_1_byteMask_2,
     io_write_1_byteMask_1,
     io_write_1_byteMask_0};
  wire [7:0]  _GEN_1 =
    {io_write_2_byteMask_7,
     io_write_2_byteMask_6,
     io_write_2_byteMask_5,
     io_write_2_byteMask_4,
     io_write_2_byteMask_3,
     io_write_2_byteMask_2,
     io_write_2_byteMask_1,
     io_write_2_byteMask_0};
  wire [7:0]  _GEN_2 =
    {io_write_3_byteMask_7,
     io_write_3_byteMask_6,
     io_write_3_byteMask_5,
     io_write_3_byteMask_4,
     io_write_3_byteMask_3,
     io_write_3_byteMask_2,
     io_write_3_byteMask_1,
     io_write_3_byteMask_0};
  wire [6:0]  _GEN_3 = io_write_0_address / 7'h8;
  wire [6:0]  _GEN_4 = io_write_1_address / 7'h8;
  wire [6:0]  _GEN_5 = io_write_2_address / 7'h8;
  wire [6:0]  _GEN_6 = io_write_3_address / 7'h8;
  wire [6:0]  _io_read_0_value_T_16 = io_read_0_address / 7'h8;
  always @(*) begin
    casez (_io_read_0_value_T_16[3:0])
      4'b0000:
        casez_tmp = _registers_0_ext_R7_data[7:0];
      4'b0001:
        casez_tmp = _registers_1_ext_R7_data[7:0];
      4'b0010:
        casez_tmp = _registers_2_ext_R7_data[7:0];
      4'b0011:
        casez_tmp = _registers_3_ext_R7_data[7:0];
      4'b0100:
        casez_tmp = _registers_4_ext_R7_data[7:0];
      4'b0101:
        casez_tmp = _registers_5_ext_R7_data[7:0];
      4'b0110:
        casez_tmp = _registers_6_ext_R7_data[7:0];
      4'b0111:
        casez_tmp = _registers_7_ext_R7_data[7:0];
      4'b1000:
        casez_tmp = _registers_8_ext_R7_data[7:0];
      4'b1001:
        casez_tmp = _registers_9_ext_R7_data[7:0];
      4'b1010:
        casez_tmp = _registers_10_ext_R7_data[7:0];
      4'b1011:
        casez_tmp = _registers_11_ext_R7_data[7:0];
      4'b1100:
        casez_tmp = _registers_12_ext_R7_data[7:0];
      4'b1101:
        casez_tmp = _registers_13_ext_R7_data[7:0];
      4'b1110:
        casez_tmp = _registers_14_ext_R7_data[7:0];
      default:
        casez_tmp = _registers_15_ext_R7_data[7:0];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_0_value_T_16[3:0])
      4'b0000:
        casez_tmp_0 = _registers_0_ext_R7_data[15:8];
      4'b0001:
        casez_tmp_0 = _registers_1_ext_R7_data[15:8];
      4'b0010:
        casez_tmp_0 = _registers_2_ext_R7_data[15:8];
      4'b0011:
        casez_tmp_0 = _registers_3_ext_R7_data[15:8];
      4'b0100:
        casez_tmp_0 = _registers_4_ext_R7_data[15:8];
      4'b0101:
        casez_tmp_0 = _registers_5_ext_R7_data[15:8];
      4'b0110:
        casez_tmp_0 = _registers_6_ext_R7_data[15:8];
      4'b0111:
        casez_tmp_0 = _registers_7_ext_R7_data[15:8];
      4'b1000:
        casez_tmp_0 = _registers_8_ext_R7_data[15:8];
      4'b1001:
        casez_tmp_0 = _registers_9_ext_R7_data[15:8];
      4'b1010:
        casez_tmp_0 = _registers_10_ext_R7_data[15:8];
      4'b1011:
        casez_tmp_0 = _registers_11_ext_R7_data[15:8];
      4'b1100:
        casez_tmp_0 = _registers_12_ext_R7_data[15:8];
      4'b1101:
        casez_tmp_0 = _registers_13_ext_R7_data[15:8];
      4'b1110:
        casez_tmp_0 = _registers_14_ext_R7_data[15:8];
      default:
        casez_tmp_0 = _registers_15_ext_R7_data[15:8];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_0_value_T_16[3:0])
      4'b0000:
        casez_tmp_1 = _registers_0_ext_R7_data[23:16];
      4'b0001:
        casez_tmp_1 = _registers_1_ext_R7_data[23:16];
      4'b0010:
        casez_tmp_1 = _registers_2_ext_R7_data[23:16];
      4'b0011:
        casez_tmp_1 = _registers_3_ext_R7_data[23:16];
      4'b0100:
        casez_tmp_1 = _registers_4_ext_R7_data[23:16];
      4'b0101:
        casez_tmp_1 = _registers_5_ext_R7_data[23:16];
      4'b0110:
        casez_tmp_1 = _registers_6_ext_R7_data[23:16];
      4'b0111:
        casez_tmp_1 = _registers_7_ext_R7_data[23:16];
      4'b1000:
        casez_tmp_1 = _registers_8_ext_R7_data[23:16];
      4'b1001:
        casez_tmp_1 = _registers_9_ext_R7_data[23:16];
      4'b1010:
        casez_tmp_1 = _registers_10_ext_R7_data[23:16];
      4'b1011:
        casez_tmp_1 = _registers_11_ext_R7_data[23:16];
      4'b1100:
        casez_tmp_1 = _registers_12_ext_R7_data[23:16];
      4'b1101:
        casez_tmp_1 = _registers_13_ext_R7_data[23:16];
      4'b1110:
        casez_tmp_1 = _registers_14_ext_R7_data[23:16];
      default:
        casez_tmp_1 = _registers_15_ext_R7_data[23:16];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_0_value_T_16[3:0])
      4'b0000:
        casez_tmp_2 = _registers_0_ext_R7_data[31:24];
      4'b0001:
        casez_tmp_2 = _registers_1_ext_R7_data[31:24];
      4'b0010:
        casez_tmp_2 = _registers_2_ext_R7_data[31:24];
      4'b0011:
        casez_tmp_2 = _registers_3_ext_R7_data[31:24];
      4'b0100:
        casez_tmp_2 = _registers_4_ext_R7_data[31:24];
      4'b0101:
        casez_tmp_2 = _registers_5_ext_R7_data[31:24];
      4'b0110:
        casez_tmp_2 = _registers_6_ext_R7_data[31:24];
      4'b0111:
        casez_tmp_2 = _registers_7_ext_R7_data[31:24];
      4'b1000:
        casez_tmp_2 = _registers_8_ext_R7_data[31:24];
      4'b1001:
        casez_tmp_2 = _registers_9_ext_R7_data[31:24];
      4'b1010:
        casez_tmp_2 = _registers_10_ext_R7_data[31:24];
      4'b1011:
        casez_tmp_2 = _registers_11_ext_R7_data[31:24];
      4'b1100:
        casez_tmp_2 = _registers_12_ext_R7_data[31:24];
      4'b1101:
        casez_tmp_2 = _registers_13_ext_R7_data[31:24];
      4'b1110:
        casez_tmp_2 = _registers_14_ext_R7_data[31:24];
      default:
        casez_tmp_2 = _registers_15_ext_R7_data[31:24];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_0_value_T_16[3:0])
      4'b0000:
        casez_tmp_3 = _registers_0_ext_R7_data[39:32];
      4'b0001:
        casez_tmp_3 = _registers_1_ext_R7_data[39:32];
      4'b0010:
        casez_tmp_3 = _registers_2_ext_R7_data[39:32];
      4'b0011:
        casez_tmp_3 = _registers_3_ext_R7_data[39:32];
      4'b0100:
        casez_tmp_3 = _registers_4_ext_R7_data[39:32];
      4'b0101:
        casez_tmp_3 = _registers_5_ext_R7_data[39:32];
      4'b0110:
        casez_tmp_3 = _registers_6_ext_R7_data[39:32];
      4'b0111:
        casez_tmp_3 = _registers_7_ext_R7_data[39:32];
      4'b1000:
        casez_tmp_3 = _registers_8_ext_R7_data[39:32];
      4'b1001:
        casez_tmp_3 = _registers_9_ext_R7_data[39:32];
      4'b1010:
        casez_tmp_3 = _registers_10_ext_R7_data[39:32];
      4'b1011:
        casez_tmp_3 = _registers_11_ext_R7_data[39:32];
      4'b1100:
        casez_tmp_3 = _registers_12_ext_R7_data[39:32];
      4'b1101:
        casez_tmp_3 = _registers_13_ext_R7_data[39:32];
      4'b1110:
        casez_tmp_3 = _registers_14_ext_R7_data[39:32];
      default:
        casez_tmp_3 = _registers_15_ext_R7_data[39:32];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_0_value_T_16[3:0])
      4'b0000:
        casez_tmp_4 = _registers_0_ext_R7_data[47:40];
      4'b0001:
        casez_tmp_4 = _registers_1_ext_R7_data[47:40];
      4'b0010:
        casez_tmp_4 = _registers_2_ext_R7_data[47:40];
      4'b0011:
        casez_tmp_4 = _registers_3_ext_R7_data[47:40];
      4'b0100:
        casez_tmp_4 = _registers_4_ext_R7_data[47:40];
      4'b0101:
        casez_tmp_4 = _registers_5_ext_R7_data[47:40];
      4'b0110:
        casez_tmp_4 = _registers_6_ext_R7_data[47:40];
      4'b0111:
        casez_tmp_4 = _registers_7_ext_R7_data[47:40];
      4'b1000:
        casez_tmp_4 = _registers_8_ext_R7_data[47:40];
      4'b1001:
        casez_tmp_4 = _registers_9_ext_R7_data[47:40];
      4'b1010:
        casez_tmp_4 = _registers_10_ext_R7_data[47:40];
      4'b1011:
        casez_tmp_4 = _registers_11_ext_R7_data[47:40];
      4'b1100:
        casez_tmp_4 = _registers_12_ext_R7_data[47:40];
      4'b1101:
        casez_tmp_4 = _registers_13_ext_R7_data[47:40];
      4'b1110:
        casez_tmp_4 = _registers_14_ext_R7_data[47:40];
      default:
        casez_tmp_4 = _registers_15_ext_R7_data[47:40];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_0_value_T_16[3:0])
      4'b0000:
        casez_tmp_5 = _registers_0_ext_R7_data[55:48];
      4'b0001:
        casez_tmp_5 = _registers_1_ext_R7_data[55:48];
      4'b0010:
        casez_tmp_5 = _registers_2_ext_R7_data[55:48];
      4'b0011:
        casez_tmp_5 = _registers_3_ext_R7_data[55:48];
      4'b0100:
        casez_tmp_5 = _registers_4_ext_R7_data[55:48];
      4'b0101:
        casez_tmp_5 = _registers_5_ext_R7_data[55:48];
      4'b0110:
        casez_tmp_5 = _registers_6_ext_R7_data[55:48];
      4'b0111:
        casez_tmp_5 = _registers_7_ext_R7_data[55:48];
      4'b1000:
        casez_tmp_5 = _registers_8_ext_R7_data[55:48];
      4'b1001:
        casez_tmp_5 = _registers_9_ext_R7_data[55:48];
      4'b1010:
        casez_tmp_5 = _registers_10_ext_R7_data[55:48];
      4'b1011:
        casez_tmp_5 = _registers_11_ext_R7_data[55:48];
      4'b1100:
        casez_tmp_5 = _registers_12_ext_R7_data[55:48];
      4'b1101:
        casez_tmp_5 = _registers_13_ext_R7_data[55:48];
      4'b1110:
        casez_tmp_5 = _registers_14_ext_R7_data[55:48];
      default:
        casez_tmp_5 = _registers_15_ext_R7_data[55:48];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_0_value_T_16[3:0])
      4'b0000:
        casez_tmp_6 = _registers_0_ext_R7_data[63:56];
      4'b0001:
        casez_tmp_6 = _registers_1_ext_R7_data[63:56];
      4'b0010:
        casez_tmp_6 = _registers_2_ext_R7_data[63:56];
      4'b0011:
        casez_tmp_6 = _registers_3_ext_R7_data[63:56];
      4'b0100:
        casez_tmp_6 = _registers_4_ext_R7_data[63:56];
      4'b0101:
        casez_tmp_6 = _registers_5_ext_R7_data[63:56];
      4'b0110:
        casez_tmp_6 = _registers_6_ext_R7_data[63:56];
      4'b0111:
        casez_tmp_6 = _registers_7_ext_R7_data[63:56];
      4'b1000:
        casez_tmp_6 = _registers_8_ext_R7_data[63:56];
      4'b1001:
        casez_tmp_6 = _registers_9_ext_R7_data[63:56];
      4'b1010:
        casez_tmp_6 = _registers_10_ext_R7_data[63:56];
      4'b1011:
        casez_tmp_6 = _registers_11_ext_R7_data[63:56];
      4'b1100:
        casez_tmp_6 = _registers_12_ext_R7_data[63:56];
      4'b1101:
        casez_tmp_6 = _registers_13_ext_R7_data[63:56];
      4'b1110:
        casez_tmp_6 = _registers_14_ext_R7_data[63:56];
      default:
        casez_tmp_6 = _registers_15_ext_R7_data[63:56];
    endcase
  end // always @(*)
  wire [6:0]  _io_read_1_value_T_16 = io_read_1_address / 7'h8;
  always @(*) begin
    casez (_io_read_1_value_T_16[3:0])
      4'b0000:
        casez_tmp_7 = _registers_0_ext_R6_data[7:0];
      4'b0001:
        casez_tmp_7 = _registers_1_ext_R6_data[7:0];
      4'b0010:
        casez_tmp_7 = _registers_2_ext_R6_data[7:0];
      4'b0011:
        casez_tmp_7 = _registers_3_ext_R6_data[7:0];
      4'b0100:
        casez_tmp_7 = _registers_4_ext_R6_data[7:0];
      4'b0101:
        casez_tmp_7 = _registers_5_ext_R6_data[7:0];
      4'b0110:
        casez_tmp_7 = _registers_6_ext_R6_data[7:0];
      4'b0111:
        casez_tmp_7 = _registers_7_ext_R6_data[7:0];
      4'b1000:
        casez_tmp_7 = _registers_8_ext_R6_data[7:0];
      4'b1001:
        casez_tmp_7 = _registers_9_ext_R6_data[7:0];
      4'b1010:
        casez_tmp_7 = _registers_10_ext_R6_data[7:0];
      4'b1011:
        casez_tmp_7 = _registers_11_ext_R6_data[7:0];
      4'b1100:
        casez_tmp_7 = _registers_12_ext_R6_data[7:0];
      4'b1101:
        casez_tmp_7 = _registers_13_ext_R6_data[7:0];
      4'b1110:
        casez_tmp_7 = _registers_14_ext_R6_data[7:0];
      default:
        casez_tmp_7 = _registers_15_ext_R6_data[7:0];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_1_value_T_16[3:0])
      4'b0000:
        casez_tmp_8 = _registers_0_ext_R6_data[15:8];
      4'b0001:
        casez_tmp_8 = _registers_1_ext_R6_data[15:8];
      4'b0010:
        casez_tmp_8 = _registers_2_ext_R6_data[15:8];
      4'b0011:
        casez_tmp_8 = _registers_3_ext_R6_data[15:8];
      4'b0100:
        casez_tmp_8 = _registers_4_ext_R6_data[15:8];
      4'b0101:
        casez_tmp_8 = _registers_5_ext_R6_data[15:8];
      4'b0110:
        casez_tmp_8 = _registers_6_ext_R6_data[15:8];
      4'b0111:
        casez_tmp_8 = _registers_7_ext_R6_data[15:8];
      4'b1000:
        casez_tmp_8 = _registers_8_ext_R6_data[15:8];
      4'b1001:
        casez_tmp_8 = _registers_9_ext_R6_data[15:8];
      4'b1010:
        casez_tmp_8 = _registers_10_ext_R6_data[15:8];
      4'b1011:
        casez_tmp_8 = _registers_11_ext_R6_data[15:8];
      4'b1100:
        casez_tmp_8 = _registers_12_ext_R6_data[15:8];
      4'b1101:
        casez_tmp_8 = _registers_13_ext_R6_data[15:8];
      4'b1110:
        casez_tmp_8 = _registers_14_ext_R6_data[15:8];
      default:
        casez_tmp_8 = _registers_15_ext_R6_data[15:8];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_1_value_T_16[3:0])
      4'b0000:
        casez_tmp_9 = _registers_0_ext_R6_data[23:16];
      4'b0001:
        casez_tmp_9 = _registers_1_ext_R6_data[23:16];
      4'b0010:
        casez_tmp_9 = _registers_2_ext_R6_data[23:16];
      4'b0011:
        casez_tmp_9 = _registers_3_ext_R6_data[23:16];
      4'b0100:
        casez_tmp_9 = _registers_4_ext_R6_data[23:16];
      4'b0101:
        casez_tmp_9 = _registers_5_ext_R6_data[23:16];
      4'b0110:
        casez_tmp_9 = _registers_6_ext_R6_data[23:16];
      4'b0111:
        casez_tmp_9 = _registers_7_ext_R6_data[23:16];
      4'b1000:
        casez_tmp_9 = _registers_8_ext_R6_data[23:16];
      4'b1001:
        casez_tmp_9 = _registers_9_ext_R6_data[23:16];
      4'b1010:
        casez_tmp_9 = _registers_10_ext_R6_data[23:16];
      4'b1011:
        casez_tmp_9 = _registers_11_ext_R6_data[23:16];
      4'b1100:
        casez_tmp_9 = _registers_12_ext_R6_data[23:16];
      4'b1101:
        casez_tmp_9 = _registers_13_ext_R6_data[23:16];
      4'b1110:
        casez_tmp_9 = _registers_14_ext_R6_data[23:16];
      default:
        casez_tmp_9 = _registers_15_ext_R6_data[23:16];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_1_value_T_16[3:0])
      4'b0000:
        casez_tmp_10 = _registers_0_ext_R6_data[31:24];
      4'b0001:
        casez_tmp_10 = _registers_1_ext_R6_data[31:24];
      4'b0010:
        casez_tmp_10 = _registers_2_ext_R6_data[31:24];
      4'b0011:
        casez_tmp_10 = _registers_3_ext_R6_data[31:24];
      4'b0100:
        casez_tmp_10 = _registers_4_ext_R6_data[31:24];
      4'b0101:
        casez_tmp_10 = _registers_5_ext_R6_data[31:24];
      4'b0110:
        casez_tmp_10 = _registers_6_ext_R6_data[31:24];
      4'b0111:
        casez_tmp_10 = _registers_7_ext_R6_data[31:24];
      4'b1000:
        casez_tmp_10 = _registers_8_ext_R6_data[31:24];
      4'b1001:
        casez_tmp_10 = _registers_9_ext_R6_data[31:24];
      4'b1010:
        casez_tmp_10 = _registers_10_ext_R6_data[31:24];
      4'b1011:
        casez_tmp_10 = _registers_11_ext_R6_data[31:24];
      4'b1100:
        casez_tmp_10 = _registers_12_ext_R6_data[31:24];
      4'b1101:
        casez_tmp_10 = _registers_13_ext_R6_data[31:24];
      4'b1110:
        casez_tmp_10 = _registers_14_ext_R6_data[31:24];
      default:
        casez_tmp_10 = _registers_15_ext_R6_data[31:24];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_1_value_T_16[3:0])
      4'b0000:
        casez_tmp_11 = _registers_0_ext_R6_data[39:32];
      4'b0001:
        casez_tmp_11 = _registers_1_ext_R6_data[39:32];
      4'b0010:
        casez_tmp_11 = _registers_2_ext_R6_data[39:32];
      4'b0011:
        casez_tmp_11 = _registers_3_ext_R6_data[39:32];
      4'b0100:
        casez_tmp_11 = _registers_4_ext_R6_data[39:32];
      4'b0101:
        casez_tmp_11 = _registers_5_ext_R6_data[39:32];
      4'b0110:
        casez_tmp_11 = _registers_6_ext_R6_data[39:32];
      4'b0111:
        casez_tmp_11 = _registers_7_ext_R6_data[39:32];
      4'b1000:
        casez_tmp_11 = _registers_8_ext_R6_data[39:32];
      4'b1001:
        casez_tmp_11 = _registers_9_ext_R6_data[39:32];
      4'b1010:
        casez_tmp_11 = _registers_10_ext_R6_data[39:32];
      4'b1011:
        casez_tmp_11 = _registers_11_ext_R6_data[39:32];
      4'b1100:
        casez_tmp_11 = _registers_12_ext_R6_data[39:32];
      4'b1101:
        casez_tmp_11 = _registers_13_ext_R6_data[39:32];
      4'b1110:
        casez_tmp_11 = _registers_14_ext_R6_data[39:32];
      default:
        casez_tmp_11 = _registers_15_ext_R6_data[39:32];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_1_value_T_16[3:0])
      4'b0000:
        casez_tmp_12 = _registers_0_ext_R6_data[47:40];
      4'b0001:
        casez_tmp_12 = _registers_1_ext_R6_data[47:40];
      4'b0010:
        casez_tmp_12 = _registers_2_ext_R6_data[47:40];
      4'b0011:
        casez_tmp_12 = _registers_3_ext_R6_data[47:40];
      4'b0100:
        casez_tmp_12 = _registers_4_ext_R6_data[47:40];
      4'b0101:
        casez_tmp_12 = _registers_5_ext_R6_data[47:40];
      4'b0110:
        casez_tmp_12 = _registers_6_ext_R6_data[47:40];
      4'b0111:
        casez_tmp_12 = _registers_7_ext_R6_data[47:40];
      4'b1000:
        casez_tmp_12 = _registers_8_ext_R6_data[47:40];
      4'b1001:
        casez_tmp_12 = _registers_9_ext_R6_data[47:40];
      4'b1010:
        casez_tmp_12 = _registers_10_ext_R6_data[47:40];
      4'b1011:
        casez_tmp_12 = _registers_11_ext_R6_data[47:40];
      4'b1100:
        casez_tmp_12 = _registers_12_ext_R6_data[47:40];
      4'b1101:
        casez_tmp_12 = _registers_13_ext_R6_data[47:40];
      4'b1110:
        casez_tmp_12 = _registers_14_ext_R6_data[47:40];
      default:
        casez_tmp_12 = _registers_15_ext_R6_data[47:40];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_1_value_T_16[3:0])
      4'b0000:
        casez_tmp_13 = _registers_0_ext_R6_data[55:48];
      4'b0001:
        casez_tmp_13 = _registers_1_ext_R6_data[55:48];
      4'b0010:
        casez_tmp_13 = _registers_2_ext_R6_data[55:48];
      4'b0011:
        casez_tmp_13 = _registers_3_ext_R6_data[55:48];
      4'b0100:
        casez_tmp_13 = _registers_4_ext_R6_data[55:48];
      4'b0101:
        casez_tmp_13 = _registers_5_ext_R6_data[55:48];
      4'b0110:
        casez_tmp_13 = _registers_6_ext_R6_data[55:48];
      4'b0111:
        casez_tmp_13 = _registers_7_ext_R6_data[55:48];
      4'b1000:
        casez_tmp_13 = _registers_8_ext_R6_data[55:48];
      4'b1001:
        casez_tmp_13 = _registers_9_ext_R6_data[55:48];
      4'b1010:
        casez_tmp_13 = _registers_10_ext_R6_data[55:48];
      4'b1011:
        casez_tmp_13 = _registers_11_ext_R6_data[55:48];
      4'b1100:
        casez_tmp_13 = _registers_12_ext_R6_data[55:48];
      4'b1101:
        casez_tmp_13 = _registers_13_ext_R6_data[55:48];
      4'b1110:
        casez_tmp_13 = _registers_14_ext_R6_data[55:48];
      default:
        casez_tmp_13 = _registers_15_ext_R6_data[55:48];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_1_value_T_16[3:0])
      4'b0000:
        casez_tmp_14 = _registers_0_ext_R6_data[63:56];
      4'b0001:
        casez_tmp_14 = _registers_1_ext_R6_data[63:56];
      4'b0010:
        casez_tmp_14 = _registers_2_ext_R6_data[63:56];
      4'b0011:
        casez_tmp_14 = _registers_3_ext_R6_data[63:56];
      4'b0100:
        casez_tmp_14 = _registers_4_ext_R6_data[63:56];
      4'b0101:
        casez_tmp_14 = _registers_5_ext_R6_data[63:56];
      4'b0110:
        casez_tmp_14 = _registers_6_ext_R6_data[63:56];
      4'b0111:
        casez_tmp_14 = _registers_7_ext_R6_data[63:56];
      4'b1000:
        casez_tmp_14 = _registers_8_ext_R6_data[63:56];
      4'b1001:
        casez_tmp_14 = _registers_9_ext_R6_data[63:56];
      4'b1010:
        casez_tmp_14 = _registers_10_ext_R6_data[63:56];
      4'b1011:
        casez_tmp_14 = _registers_11_ext_R6_data[63:56];
      4'b1100:
        casez_tmp_14 = _registers_12_ext_R6_data[63:56];
      4'b1101:
        casez_tmp_14 = _registers_13_ext_R6_data[63:56];
      4'b1110:
        casez_tmp_14 = _registers_14_ext_R6_data[63:56];
      default:
        casez_tmp_14 = _registers_15_ext_R6_data[63:56];
    endcase
  end // always @(*)
  wire [6:0]  _io_read_2_value_T_16 = io_read_2_address / 7'h8;
  always @(*) begin
    casez (_io_read_2_value_T_16[3:0])
      4'b0000:
        casez_tmp_15 = _registers_0_ext_R5_data[7:0];
      4'b0001:
        casez_tmp_15 = _registers_1_ext_R5_data[7:0];
      4'b0010:
        casez_tmp_15 = _registers_2_ext_R5_data[7:0];
      4'b0011:
        casez_tmp_15 = _registers_3_ext_R5_data[7:0];
      4'b0100:
        casez_tmp_15 = _registers_4_ext_R5_data[7:0];
      4'b0101:
        casez_tmp_15 = _registers_5_ext_R5_data[7:0];
      4'b0110:
        casez_tmp_15 = _registers_6_ext_R5_data[7:0];
      4'b0111:
        casez_tmp_15 = _registers_7_ext_R5_data[7:0];
      4'b1000:
        casez_tmp_15 = _registers_8_ext_R5_data[7:0];
      4'b1001:
        casez_tmp_15 = _registers_9_ext_R5_data[7:0];
      4'b1010:
        casez_tmp_15 = _registers_10_ext_R5_data[7:0];
      4'b1011:
        casez_tmp_15 = _registers_11_ext_R5_data[7:0];
      4'b1100:
        casez_tmp_15 = _registers_12_ext_R5_data[7:0];
      4'b1101:
        casez_tmp_15 = _registers_13_ext_R5_data[7:0];
      4'b1110:
        casez_tmp_15 = _registers_14_ext_R5_data[7:0];
      default:
        casez_tmp_15 = _registers_15_ext_R5_data[7:0];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_2_value_T_16[3:0])
      4'b0000:
        casez_tmp_16 = _registers_0_ext_R5_data[15:8];
      4'b0001:
        casez_tmp_16 = _registers_1_ext_R5_data[15:8];
      4'b0010:
        casez_tmp_16 = _registers_2_ext_R5_data[15:8];
      4'b0011:
        casez_tmp_16 = _registers_3_ext_R5_data[15:8];
      4'b0100:
        casez_tmp_16 = _registers_4_ext_R5_data[15:8];
      4'b0101:
        casez_tmp_16 = _registers_5_ext_R5_data[15:8];
      4'b0110:
        casez_tmp_16 = _registers_6_ext_R5_data[15:8];
      4'b0111:
        casez_tmp_16 = _registers_7_ext_R5_data[15:8];
      4'b1000:
        casez_tmp_16 = _registers_8_ext_R5_data[15:8];
      4'b1001:
        casez_tmp_16 = _registers_9_ext_R5_data[15:8];
      4'b1010:
        casez_tmp_16 = _registers_10_ext_R5_data[15:8];
      4'b1011:
        casez_tmp_16 = _registers_11_ext_R5_data[15:8];
      4'b1100:
        casez_tmp_16 = _registers_12_ext_R5_data[15:8];
      4'b1101:
        casez_tmp_16 = _registers_13_ext_R5_data[15:8];
      4'b1110:
        casez_tmp_16 = _registers_14_ext_R5_data[15:8];
      default:
        casez_tmp_16 = _registers_15_ext_R5_data[15:8];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_2_value_T_16[3:0])
      4'b0000:
        casez_tmp_17 = _registers_0_ext_R5_data[23:16];
      4'b0001:
        casez_tmp_17 = _registers_1_ext_R5_data[23:16];
      4'b0010:
        casez_tmp_17 = _registers_2_ext_R5_data[23:16];
      4'b0011:
        casez_tmp_17 = _registers_3_ext_R5_data[23:16];
      4'b0100:
        casez_tmp_17 = _registers_4_ext_R5_data[23:16];
      4'b0101:
        casez_tmp_17 = _registers_5_ext_R5_data[23:16];
      4'b0110:
        casez_tmp_17 = _registers_6_ext_R5_data[23:16];
      4'b0111:
        casez_tmp_17 = _registers_7_ext_R5_data[23:16];
      4'b1000:
        casez_tmp_17 = _registers_8_ext_R5_data[23:16];
      4'b1001:
        casez_tmp_17 = _registers_9_ext_R5_data[23:16];
      4'b1010:
        casez_tmp_17 = _registers_10_ext_R5_data[23:16];
      4'b1011:
        casez_tmp_17 = _registers_11_ext_R5_data[23:16];
      4'b1100:
        casez_tmp_17 = _registers_12_ext_R5_data[23:16];
      4'b1101:
        casez_tmp_17 = _registers_13_ext_R5_data[23:16];
      4'b1110:
        casez_tmp_17 = _registers_14_ext_R5_data[23:16];
      default:
        casez_tmp_17 = _registers_15_ext_R5_data[23:16];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_2_value_T_16[3:0])
      4'b0000:
        casez_tmp_18 = _registers_0_ext_R5_data[31:24];
      4'b0001:
        casez_tmp_18 = _registers_1_ext_R5_data[31:24];
      4'b0010:
        casez_tmp_18 = _registers_2_ext_R5_data[31:24];
      4'b0011:
        casez_tmp_18 = _registers_3_ext_R5_data[31:24];
      4'b0100:
        casez_tmp_18 = _registers_4_ext_R5_data[31:24];
      4'b0101:
        casez_tmp_18 = _registers_5_ext_R5_data[31:24];
      4'b0110:
        casez_tmp_18 = _registers_6_ext_R5_data[31:24];
      4'b0111:
        casez_tmp_18 = _registers_7_ext_R5_data[31:24];
      4'b1000:
        casez_tmp_18 = _registers_8_ext_R5_data[31:24];
      4'b1001:
        casez_tmp_18 = _registers_9_ext_R5_data[31:24];
      4'b1010:
        casez_tmp_18 = _registers_10_ext_R5_data[31:24];
      4'b1011:
        casez_tmp_18 = _registers_11_ext_R5_data[31:24];
      4'b1100:
        casez_tmp_18 = _registers_12_ext_R5_data[31:24];
      4'b1101:
        casez_tmp_18 = _registers_13_ext_R5_data[31:24];
      4'b1110:
        casez_tmp_18 = _registers_14_ext_R5_data[31:24];
      default:
        casez_tmp_18 = _registers_15_ext_R5_data[31:24];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_2_value_T_16[3:0])
      4'b0000:
        casez_tmp_19 = _registers_0_ext_R5_data[39:32];
      4'b0001:
        casez_tmp_19 = _registers_1_ext_R5_data[39:32];
      4'b0010:
        casez_tmp_19 = _registers_2_ext_R5_data[39:32];
      4'b0011:
        casez_tmp_19 = _registers_3_ext_R5_data[39:32];
      4'b0100:
        casez_tmp_19 = _registers_4_ext_R5_data[39:32];
      4'b0101:
        casez_tmp_19 = _registers_5_ext_R5_data[39:32];
      4'b0110:
        casez_tmp_19 = _registers_6_ext_R5_data[39:32];
      4'b0111:
        casez_tmp_19 = _registers_7_ext_R5_data[39:32];
      4'b1000:
        casez_tmp_19 = _registers_8_ext_R5_data[39:32];
      4'b1001:
        casez_tmp_19 = _registers_9_ext_R5_data[39:32];
      4'b1010:
        casez_tmp_19 = _registers_10_ext_R5_data[39:32];
      4'b1011:
        casez_tmp_19 = _registers_11_ext_R5_data[39:32];
      4'b1100:
        casez_tmp_19 = _registers_12_ext_R5_data[39:32];
      4'b1101:
        casez_tmp_19 = _registers_13_ext_R5_data[39:32];
      4'b1110:
        casez_tmp_19 = _registers_14_ext_R5_data[39:32];
      default:
        casez_tmp_19 = _registers_15_ext_R5_data[39:32];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_2_value_T_16[3:0])
      4'b0000:
        casez_tmp_20 = _registers_0_ext_R5_data[47:40];
      4'b0001:
        casez_tmp_20 = _registers_1_ext_R5_data[47:40];
      4'b0010:
        casez_tmp_20 = _registers_2_ext_R5_data[47:40];
      4'b0011:
        casez_tmp_20 = _registers_3_ext_R5_data[47:40];
      4'b0100:
        casez_tmp_20 = _registers_4_ext_R5_data[47:40];
      4'b0101:
        casez_tmp_20 = _registers_5_ext_R5_data[47:40];
      4'b0110:
        casez_tmp_20 = _registers_6_ext_R5_data[47:40];
      4'b0111:
        casez_tmp_20 = _registers_7_ext_R5_data[47:40];
      4'b1000:
        casez_tmp_20 = _registers_8_ext_R5_data[47:40];
      4'b1001:
        casez_tmp_20 = _registers_9_ext_R5_data[47:40];
      4'b1010:
        casez_tmp_20 = _registers_10_ext_R5_data[47:40];
      4'b1011:
        casez_tmp_20 = _registers_11_ext_R5_data[47:40];
      4'b1100:
        casez_tmp_20 = _registers_12_ext_R5_data[47:40];
      4'b1101:
        casez_tmp_20 = _registers_13_ext_R5_data[47:40];
      4'b1110:
        casez_tmp_20 = _registers_14_ext_R5_data[47:40];
      default:
        casez_tmp_20 = _registers_15_ext_R5_data[47:40];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_2_value_T_16[3:0])
      4'b0000:
        casez_tmp_21 = _registers_0_ext_R5_data[55:48];
      4'b0001:
        casez_tmp_21 = _registers_1_ext_R5_data[55:48];
      4'b0010:
        casez_tmp_21 = _registers_2_ext_R5_data[55:48];
      4'b0011:
        casez_tmp_21 = _registers_3_ext_R5_data[55:48];
      4'b0100:
        casez_tmp_21 = _registers_4_ext_R5_data[55:48];
      4'b0101:
        casez_tmp_21 = _registers_5_ext_R5_data[55:48];
      4'b0110:
        casez_tmp_21 = _registers_6_ext_R5_data[55:48];
      4'b0111:
        casez_tmp_21 = _registers_7_ext_R5_data[55:48];
      4'b1000:
        casez_tmp_21 = _registers_8_ext_R5_data[55:48];
      4'b1001:
        casez_tmp_21 = _registers_9_ext_R5_data[55:48];
      4'b1010:
        casez_tmp_21 = _registers_10_ext_R5_data[55:48];
      4'b1011:
        casez_tmp_21 = _registers_11_ext_R5_data[55:48];
      4'b1100:
        casez_tmp_21 = _registers_12_ext_R5_data[55:48];
      4'b1101:
        casez_tmp_21 = _registers_13_ext_R5_data[55:48];
      4'b1110:
        casez_tmp_21 = _registers_14_ext_R5_data[55:48];
      default:
        casez_tmp_21 = _registers_15_ext_R5_data[55:48];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_2_value_T_16[3:0])
      4'b0000:
        casez_tmp_22 = _registers_0_ext_R5_data[63:56];
      4'b0001:
        casez_tmp_22 = _registers_1_ext_R5_data[63:56];
      4'b0010:
        casez_tmp_22 = _registers_2_ext_R5_data[63:56];
      4'b0011:
        casez_tmp_22 = _registers_3_ext_R5_data[63:56];
      4'b0100:
        casez_tmp_22 = _registers_4_ext_R5_data[63:56];
      4'b0101:
        casez_tmp_22 = _registers_5_ext_R5_data[63:56];
      4'b0110:
        casez_tmp_22 = _registers_6_ext_R5_data[63:56];
      4'b0111:
        casez_tmp_22 = _registers_7_ext_R5_data[63:56];
      4'b1000:
        casez_tmp_22 = _registers_8_ext_R5_data[63:56];
      4'b1001:
        casez_tmp_22 = _registers_9_ext_R5_data[63:56];
      4'b1010:
        casez_tmp_22 = _registers_10_ext_R5_data[63:56];
      4'b1011:
        casez_tmp_22 = _registers_11_ext_R5_data[63:56];
      4'b1100:
        casez_tmp_22 = _registers_12_ext_R5_data[63:56];
      4'b1101:
        casez_tmp_22 = _registers_13_ext_R5_data[63:56];
      4'b1110:
        casez_tmp_22 = _registers_14_ext_R5_data[63:56];
      default:
        casez_tmp_22 = _registers_15_ext_R5_data[63:56];
    endcase
  end // always @(*)
  wire [6:0]  _io_read_3_value_T_16 = io_read_3_address / 7'h8;
  always @(*) begin
    casez (_io_read_3_value_T_16[3:0])
      4'b0000:
        casez_tmp_23 = _registers_0_ext_R4_data[7:0];
      4'b0001:
        casez_tmp_23 = _registers_1_ext_R4_data[7:0];
      4'b0010:
        casez_tmp_23 = _registers_2_ext_R4_data[7:0];
      4'b0011:
        casez_tmp_23 = _registers_3_ext_R4_data[7:0];
      4'b0100:
        casez_tmp_23 = _registers_4_ext_R4_data[7:0];
      4'b0101:
        casez_tmp_23 = _registers_5_ext_R4_data[7:0];
      4'b0110:
        casez_tmp_23 = _registers_6_ext_R4_data[7:0];
      4'b0111:
        casez_tmp_23 = _registers_7_ext_R4_data[7:0];
      4'b1000:
        casez_tmp_23 = _registers_8_ext_R4_data[7:0];
      4'b1001:
        casez_tmp_23 = _registers_9_ext_R4_data[7:0];
      4'b1010:
        casez_tmp_23 = _registers_10_ext_R4_data[7:0];
      4'b1011:
        casez_tmp_23 = _registers_11_ext_R4_data[7:0];
      4'b1100:
        casez_tmp_23 = _registers_12_ext_R4_data[7:0];
      4'b1101:
        casez_tmp_23 = _registers_13_ext_R4_data[7:0];
      4'b1110:
        casez_tmp_23 = _registers_14_ext_R4_data[7:0];
      default:
        casez_tmp_23 = _registers_15_ext_R4_data[7:0];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_3_value_T_16[3:0])
      4'b0000:
        casez_tmp_24 = _registers_0_ext_R4_data[15:8];
      4'b0001:
        casez_tmp_24 = _registers_1_ext_R4_data[15:8];
      4'b0010:
        casez_tmp_24 = _registers_2_ext_R4_data[15:8];
      4'b0011:
        casez_tmp_24 = _registers_3_ext_R4_data[15:8];
      4'b0100:
        casez_tmp_24 = _registers_4_ext_R4_data[15:8];
      4'b0101:
        casez_tmp_24 = _registers_5_ext_R4_data[15:8];
      4'b0110:
        casez_tmp_24 = _registers_6_ext_R4_data[15:8];
      4'b0111:
        casez_tmp_24 = _registers_7_ext_R4_data[15:8];
      4'b1000:
        casez_tmp_24 = _registers_8_ext_R4_data[15:8];
      4'b1001:
        casez_tmp_24 = _registers_9_ext_R4_data[15:8];
      4'b1010:
        casez_tmp_24 = _registers_10_ext_R4_data[15:8];
      4'b1011:
        casez_tmp_24 = _registers_11_ext_R4_data[15:8];
      4'b1100:
        casez_tmp_24 = _registers_12_ext_R4_data[15:8];
      4'b1101:
        casez_tmp_24 = _registers_13_ext_R4_data[15:8];
      4'b1110:
        casez_tmp_24 = _registers_14_ext_R4_data[15:8];
      default:
        casez_tmp_24 = _registers_15_ext_R4_data[15:8];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_3_value_T_16[3:0])
      4'b0000:
        casez_tmp_25 = _registers_0_ext_R4_data[23:16];
      4'b0001:
        casez_tmp_25 = _registers_1_ext_R4_data[23:16];
      4'b0010:
        casez_tmp_25 = _registers_2_ext_R4_data[23:16];
      4'b0011:
        casez_tmp_25 = _registers_3_ext_R4_data[23:16];
      4'b0100:
        casez_tmp_25 = _registers_4_ext_R4_data[23:16];
      4'b0101:
        casez_tmp_25 = _registers_5_ext_R4_data[23:16];
      4'b0110:
        casez_tmp_25 = _registers_6_ext_R4_data[23:16];
      4'b0111:
        casez_tmp_25 = _registers_7_ext_R4_data[23:16];
      4'b1000:
        casez_tmp_25 = _registers_8_ext_R4_data[23:16];
      4'b1001:
        casez_tmp_25 = _registers_9_ext_R4_data[23:16];
      4'b1010:
        casez_tmp_25 = _registers_10_ext_R4_data[23:16];
      4'b1011:
        casez_tmp_25 = _registers_11_ext_R4_data[23:16];
      4'b1100:
        casez_tmp_25 = _registers_12_ext_R4_data[23:16];
      4'b1101:
        casez_tmp_25 = _registers_13_ext_R4_data[23:16];
      4'b1110:
        casez_tmp_25 = _registers_14_ext_R4_data[23:16];
      default:
        casez_tmp_25 = _registers_15_ext_R4_data[23:16];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_3_value_T_16[3:0])
      4'b0000:
        casez_tmp_26 = _registers_0_ext_R4_data[31:24];
      4'b0001:
        casez_tmp_26 = _registers_1_ext_R4_data[31:24];
      4'b0010:
        casez_tmp_26 = _registers_2_ext_R4_data[31:24];
      4'b0011:
        casez_tmp_26 = _registers_3_ext_R4_data[31:24];
      4'b0100:
        casez_tmp_26 = _registers_4_ext_R4_data[31:24];
      4'b0101:
        casez_tmp_26 = _registers_5_ext_R4_data[31:24];
      4'b0110:
        casez_tmp_26 = _registers_6_ext_R4_data[31:24];
      4'b0111:
        casez_tmp_26 = _registers_7_ext_R4_data[31:24];
      4'b1000:
        casez_tmp_26 = _registers_8_ext_R4_data[31:24];
      4'b1001:
        casez_tmp_26 = _registers_9_ext_R4_data[31:24];
      4'b1010:
        casez_tmp_26 = _registers_10_ext_R4_data[31:24];
      4'b1011:
        casez_tmp_26 = _registers_11_ext_R4_data[31:24];
      4'b1100:
        casez_tmp_26 = _registers_12_ext_R4_data[31:24];
      4'b1101:
        casez_tmp_26 = _registers_13_ext_R4_data[31:24];
      4'b1110:
        casez_tmp_26 = _registers_14_ext_R4_data[31:24];
      default:
        casez_tmp_26 = _registers_15_ext_R4_data[31:24];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_3_value_T_16[3:0])
      4'b0000:
        casez_tmp_27 = _registers_0_ext_R4_data[39:32];
      4'b0001:
        casez_tmp_27 = _registers_1_ext_R4_data[39:32];
      4'b0010:
        casez_tmp_27 = _registers_2_ext_R4_data[39:32];
      4'b0011:
        casez_tmp_27 = _registers_3_ext_R4_data[39:32];
      4'b0100:
        casez_tmp_27 = _registers_4_ext_R4_data[39:32];
      4'b0101:
        casez_tmp_27 = _registers_5_ext_R4_data[39:32];
      4'b0110:
        casez_tmp_27 = _registers_6_ext_R4_data[39:32];
      4'b0111:
        casez_tmp_27 = _registers_7_ext_R4_data[39:32];
      4'b1000:
        casez_tmp_27 = _registers_8_ext_R4_data[39:32];
      4'b1001:
        casez_tmp_27 = _registers_9_ext_R4_data[39:32];
      4'b1010:
        casez_tmp_27 = _registers_10_ext_R4_data[39:32];
      4'b1011:
        casez_tmp_27 = _registers_11_ext_R4_data[39:32];
      4'b1100:
        casez_tmp_27 = _registers_12_ext_R4_data[39:32];
      4'b1101:
        casez_tmp_27 = _registers_13_ext_R4_data[39:32];
      4'b1110:
        casez_tmp_27 = _registers_14_ext_R4_data[39:32];
      default:
        casez_tmp_27 = _registers_15_ext_R4_data[39:32];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_3_value_T_16[3:0])
      4'b0000:
        casez_tmp_28 = _registers_0_ext_R4_data[47:40];
      4'b0001:
        casez_tmp_28 = _registers_1_ext_R4_data[47:40];
      4'b0010:
        casez_tmp_28 = _registers_2_ext_R4_data[47:40];
      4'b0011:
        casez_tmp_28 = _registers_3_ext_R4_data[47:40];
      4'b0100:
        casez_tmp_28 = _registers_4_ext_R4_data[47:40];
      4'b0101:
        casez_tmp_28 = _registers_5_ext_R4_data[47:40];
      4'b0110:
        casez_tmp_28 = _registers_6_ext_R4_data[47:40];
      4'b0111:
        casez_tmp_28 = _registers_7_ext_R4_data[47:40];
      4'b1000:
        casez_tmp_28 = _registers_8_ext_R4_data[47:40];
      4'b1001:
        casez_tmp_28 = _registers_9_ext_R4_data[47:40];
      4'b1010:
        casez_tmp_28 = _registers_10_ext_R4_data[47:40];
      4'b1011:
        casez_tmp_28 = _registers_11_ext_R4_data[47:40];
      4'b1100:
        casez_tmp_28 = _registers_12_ext_R4_data[47:40];
      4'b1101:
        casez_tmp_28 = _registers_13_ext_R4_data[47:40];
      4'b1110:
        casez_tmp_28 = _registers_14_ext_R4_data[47:40];
      default:
        casez_tmp_28 = _registers_15_ext_R4_data[47:40];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_3_value_T_16[3:0])
      4'b0000:
        casez_tmp_29 = _registers_0_ext_R4_data[55:48];
      4'b0001:
        casez_tmp_29 = _registers_1_ext_R4_data[55:48];
      4'b0010:
        casez_tmp_29 = _registers_2_ext_R4_data[55:48];
      4'b0011:
        casez_tmp_29 = _registers_3_ext_R4_data[55:48];
      4'b0100:
        casez_tmp_29 = _registers_4_ext_R4_data[55:48];
      4'b0101:
        casez_tmp_29 = _registers_5_ext_R4_data[55:48];
      4'b0110:
        casez_tmp_29 = _registers_6_ext_R4_data[55:48];
      4'b0111:
        casez_tmp_29 = _registers_7_ext_R4_data[55:48];
      4'b1000:
        casez_tmp_29 = _registers_8_ext_R4_data[55:48];
      4'b1001:
        casez_tmp_29 = _registers_9_ext_R4_data[55:48];
      4'b1010:
        casez_tmp_29 = _registers_10_ext_R4_data[55:48];
      4'b1011:
        casez_tmp_29 = _registers_11_ext_R4_data[55:48];
      4'b1100:
        casez_tmp_29 = _registers_12_ext_R4_data[55:48];
      4'b1101:
        casez_tmp_29 = _registers_13_ext_R4_data[55:48];
      4'b1110:
        casez_tmp_29 = _registers_14_ext_R4_data[55:48];
      default:
        casez_tmp_29 = _registers_15_ext_R4_data[55:48];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_3_value_T_16[3:0])
      4'b0000:
        casez_tmp_30 = _registers_0_ext_R4_data[63:56];
      4'b0001:
        casez_tmp_30 = _registers_1_ext_R4_data[63:56];
      4'b0010:
        casez_tmp_30 = _registers_2_ext_R4_data[63:56];
      4'b0011:
        casez_tmp_30 = _registers_3_ext_R4_data[63:56];
      4'b0100:
        casez_tmp_30 = _registers_4_ext_R4_data[63:56];
      4'b0101:
        casez_tmp_30 = _registers_5_ext_R4_data[63:56];
      4'b0110:
        casez_tmp_30 = _registers_6_ext_R4_data[63:56];
      4'b0111:
        casez_tmp_30 = _registers_7_ext_R4_data[63:56];
      4'b1000:
        casez_tmp_30 = _registers_8_ext_R4_data[63:56];
      4'b1001:
        casez_tmp_30 = _registers_9_ext_R4_data[63:56];
      4'b1010:
        casez_tmp_30 = _registers_10_ext_R4_data[63:56];
      4'b1011:
        casez_tmp_30 = _registers_11_ext_R4_data[63:56];
      4'b1100:
        casez_tmp_30 = _registers_12_ext_R4_data[63:56];
      4'b1101:
        casez_tmp_30 = _registers_13_ext_R4_data[63:56];
      4'b1110:
        casez_tmp_30 = _registers_14_ext_R4_data[63:56];
      default:
        casez_tmp_30 = _registers_15_ext_R4_data[63:56];
    endcase
  end // always @(*)
  wire [6:0]  _io_read_4_value_T_16 = io_read_4_address / 7'h8;
  always @(*) begin
    casez (_io_read_4_value_T_16[3:0])
      4'b0000:
        casez_tmp_31 = _registers_0_ext_R3_data[7:0];
      4'b0001:
        casez_tmp_31 = _registers_1_ext_R3_data[7:0];
      4'b0010:
        casez_tmp_31 = _registers_2_ext_R3_data[7:0];
      4'b0011:
        casez_tmp_31 = _registers_3_ext_R3_data[7:0];
      4'b0100:
        casez_tmp_31 = _registers_4_ext_R3_data[7:0];
      4'b0101:
        casez_tmp_31 = _registers_5_ext_R3_data[7:0];
      4'b0110:
        casez_tmp_31 = _registers_6_ext_R3_data[7:0];
      4'b0111:
        casez_tmp_31 = _registers_7_ext_R3_data[7:0];
      4'b1000:
        casez_tmp_31 = _registers_8_ext_R3_data[7:0];
      4'b1001:
        casez_tmp_31 = _registers_9_ext_R3_data[7:0];
      4'b1010:
        casez_tmp_31 = _registers_10_ext_R3_data[7:0];
      4'b1011:
        casez_tmp_31 = _registers_11_ext_R3_data[7:0];
      4'b1100:
        casez_tmp_31 = _registers_12_ext_R3_data[7:0];
      4'b1101:
        casez_tmp_31 = _registers_13_ext_R3_data[7:0];
      4'b1110:
        casez_tmp_31 = _registers_14_ext_R3_data[7:0];
      default:
        casez_tmp_31 = _registers_15_ext_R3_data[7:0];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_4_value_T_16[3:0])
      4'b0000:
        casez_tmp_32 = _registers_0_ext_R3_data[15:8];
      4'b0001:
        casez_tmp_32 = _registers_1_ext_R3_data[15:8];
      4'b0010:
        casez_tmp_32 = _registers_2_ext_R3_data[15:8];
      4'b0011:
        casez_tmp_32 = _registers_3_ext_R3_data[15:8];
      4'b0100:
        casez_tmp_32 = _registers_4_ext_R3_data[15:8];
      4'b0101:
        casez_tmp_32 = _registers_5_ext_R3_data[15:8];
      4'b0110:
        casez_tmp_32 = _registers_6_ext_R3_data[15:8];
      4'b0111:
        casez_tmp_32 = _registers_7_ext_R3_data[15:8];
      4'b1000:
        casez_tmp_32 = _registers_8_ext_R3_data[15:8];
      4'b1001:
        casez_tmp_32 = _registers_9_ext_R3_data[15:8];
      4'b1010:
        casez_tmp_32 = _registers_10_ext_R3_data[15:8];
      4'b1011:
        casez_tmp_32 = _registers_11_ext_R3_data[15:8];
      4'b1100:
        casez_tmp_32 = _registers_12_ext_R3_data[15:8];
      4'b1101:
        casez_tmp_32 = _registers_13_ext_R3_data[15:8];
      4'b1110:
        casez_tmp_32 = _registers_14_ext_R3_data[15:8];
      default:
        casez_tmp_32 = _registers_15_ext_R3_data[15:8];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_4_value_T_16[3:0])
      4'b0000:
        casez_tmp_33 = _registers_0_ext_R3_data[23:16];
      4'b0001:
        casez_tmp_33 = _registers_1_ext_R3_data[23:16];
      4'b0010:
        casez_tmp_33 = _registers_2_ext_R3_data[23:16];
      4'b0011:
        casez_tmp_33 = _registers_3_ext_R3_data[23:16];
      4'b0100:
        casez_tmp_33 = _registers_4_ext_R3_data[23:16];
      4'b0101:
        casez_tmp_33 = _registers_5_ext_R3_data[23:16];
      4'b0110:
        casez_tmp_33 = _registers_6_ext_R3_data[23:16];
      4'b0111:
        casez_tmp_33 = _registers_7_ext_R3_data[23:16];
      4'b1000:
        casez_tmp_33 = _registers_8_ext_R3_data[23:16];
      4'b1001:
        casez_tmp_33 = _registers_9_ext_R3_data[23:16];
      4'b1010:
        casez_tmp_33 = _registers_10_ext_R3_data[23:16];
      4'b1011:
        casez_tmp_33 = _registers_11_ext_R3_data[23:16];
      4'b1100:
        casez_tmp_33 = _registers_12_ext_R3_data[23:16];
      4'b1101:
        casez_tmp_33 = _registers_13_ext_R3_data[23:16];
      4'b1110:
        casez_tmp_33 = _registers_14_ext_R3_data[23:16];
      default:
        casez_tmp_33 = _registers_15_ext_R3_data[23:16];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_4_value_T_16[3:0])
      4'b0000:
        casez_tmp_34 = _registers_0_ext_R3_data[31:24];
      4'b0001:
        casez_tmp_34 = _registers_1_ext_R3_data[31:24];
      4'b0010:
        casez_tmp_34 = _registers_2_ext_R3_data[31:24];
      4'b0011:
        casez_tmp_34 = _registers_3_ext_R3_data[31:24];
      4'b0100:
        casez_tmp_34 = _registers_4_ext_R3_data[31:24];
      4'b0101:
        casez_tmp_34 = _registers_5_ext_R3_data[31:24];
      4'b0110:
        casez_tmp_34 = _registers_6_ext_R3_data[31:24];
      4'b0111:
        casez_tmp_34 = _registers_7_ext_R3_data[31:24];
      4'b1000:
        casez_tmp_34 = _registers_8_ext_R3_data[31:24];
      4'b1001:
        casez_tmp_34 = _registers_9_ext_R3_data[31:24];
      4'b1010:
        casez_tmp_34 = _registers_10_ext_R3_data[31:24];
      4'b1011:
        casez_tmp_34 = _registers_11_ext_R3_data[31:24];
      4'b1100:
        casez_tmp_34 = _registers_12_ext_R3_data[31:24];
      4'b1101:
        casez_tmp_34 = _registers_13_ext_R3_data[31:24];
      4'b1110:
        casez_tmp_34 = _registers_14_ext_R3_data[31:24];
      default:
        casez_tmp_34 = _registers_15_ext_R3_data[31:24];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_4_value_T_16[3:0])
      4'b0000:
        casez_tmp_35 = _registers_0_ext_R3_data[39:32];
      4'b0001:
        casez_tmp_35 = _registers_1_ext_R3_data[39:32];
      4'b0010:
        casez_tmp_35 = _registers_2_ext_R3_data[39:32];
      4'b0011:
        casez_tmp_35 = _registers_3_ext_R3_data[39:32];
      4'b0100:
        casez_tmp_35 = _registers_4_ext_R3_data[39:32];
      4'b0101:
        casez_tmp_35 = _registers_5_ext_R3_data[39:32];
      4'b0110:
        casez_tmp_35 = _registers_6_ext_R3_data[39:32];
      4'b0111:
        casez_tmp_35 = _registers_7_ext_R3_data[39:32];
      4'b1000:
        casez_tmp_35 = _registers_8_ext_R3_data[39:32];
      4'b1001:
        casez_tmp_35 = _registers_9_ext_R3_data[39:32];
      4'b1010:
        casez_tmp_35 = _registers_10_ext_R3_data[39:32];
      4'b1011:
        casez_tmp_35 = _registers_11_ext_R3_data[39:32];
      4'b1100:
        casez_tmp_35 = _registers_12_ext_R3_data[39:32];
      4'b1101:
        casez_tmp_35 = _registers_13_ext_R3_data[39:32];
      4'b1110:
        casez_tmp_35 = _registers_14_ext_R3_data[39:32];
      default:
        casez_tmp_35 = _registers_15_ext_R3_data[39:32];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_4_value_T_16[3:0])
      4'b0000:
        casez_tmp_36 = _registers_0_ext_R3_data[47:40];
      4'b0001:
        casez_tmp_36 = _registers_1_ext_R3_data[47:40];
      4'b0010:
        casez_tmp_36 = _registers_2_ext_R3_data[47:40];
      4'b0011:
        casez_tmp_36 = _registers_3_ext_R3_data[47:40];
      4'b0100:
        casez_tmp_36 = _registers_4_ext_R3_data[47:40];
      4'b0101:
        casez_tmp_36 = _registers_5_ext_R3_data[47:40];
      4'b0110:
        casez_tmp_36 = _registers_6_ext_R3_data[47:40];
      4'b0111:
        casez_tmp_36 = _registers_7_ext_R3_data[47:40];
      4'b1000:
        casez_tmp_36 = _registers_8_ext_R3_data[47:40];
      4'b1001:
        casez_tmp_36 = _registers_9_ext_R3_data[47:40];
      4'b1010:
        casez_tmp_36 = _registers_10_ext_R3_data[47:40];
      4'b1011:
        casez_tmp_36 = _registers_11_ext_R3_data[47:40];
      4'b1100:
        casez_tmp_36 = _registers_12_ext_R3_data[47:40];
      4'b1101:
        casez_tmp_36 = _registers_13_ext_R3_data[47:40];
      4'b1110:
        casez_tmp_36 = _registers_14_ext_R3_data[47:40];
      default:
        casez_tmp_36 = _registers_15_ext_R3_data[47:40];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_4_value_T_16[3:0])
      4'b0000:
        casez_tmp_37 = _registers_0_ext_R3_data[55:48];
      4'b0001:
        casez_tmp_37 = _registers_1_ext_R3_data[55:48];
      4'b0010:
        casez_tmp_37 = _registers_2_ext_R3_data[55:48];
      4'b0011:
        casez_tmp_37 = _registers_3_ext_R3_data[55:48];
      4'b0100:
        casez_tmp_37 = _registers_4_ext_R3_data[55:48];
      4'b0101:
        casez_tmp_37 = _registers_5_ext_R3_data[55:48];
      4'b0110:
        casez_tmp_37 = _registers_6_ext_R3_data[55:48];
      4'b0111:
        casez_tmp_37 = _registers_7_ext_R3_data[55:48];
      4'b1000:
        casez_tmp_37 = _registers_8_ext_R3_data[55:48];
      4'b1001:
        casez_tmp_37 = _registers_9_ext_R3_data[55:48];
      4'b1010:
        casez_tmp_37 = _registers_10_ext_R3_data[55:48];
      4'b1011:
        casez_tmp_37 = _registers_11_ext_R3_data[55:48];
      4'b1100:
        casez_tmp_37 = _registers_12_ext_R3_data[55:48];
      4'b1101:
        casez_tmp_37 = _registers_13_ext_R3_data[55:48];
      4'b1110:
        casez_tmp_37 = _registers_14_ext_R3_data[55:48];
      default:
        casez_tmp_37 = _registers_15_ext_R3_data[55:48];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_4_value_T_16[3:0])
      4'b0000:
        casez_tmp_38 = _registers_0_ext_R3_data[63:56];
      4'b0001:
        casez_tmp_38 = _registers_1_ext_R3_data[63:56];
      4'b0010:
        casez_tmp_38 = _registers_2_ext_R3_data[63:56];
      4'b0011:
        casez_tmp_38 = _registers_3_ext_R3_data[63:56];
      4'b0100:
        casez_tmp_38 = _registers_4_ext_R3_data[63:56];
      4'b0101:
        casez_tmp_38 = _registers_5_ext_R3_data[63:56];
      4'b0110:
        casez_tmp_38 = _registers_6_ext_R3_data[63:56];
      4'b0111:
        casez_tmp_38 = _registers_7_ext_R3_data[63:56];
      4'b1000:
        casez_tmp_38 = _registers_8_ext_R3_data[63:56];
      4'b1001:
        casez_tmp_38 = _registers_9_ext_R3_data[63:56];
      4'b1010:
        casez_tmp_38 = _registers_10_ext_R3_data[63:56];
      4'b1011:
        casez_tmp_38 = _registers_11_ext_R3_data[63:56];
      4'b1100:
        casez_tmp_38 = _registers_12_ext_R3_data[63:56];
      4'b1101:
        casez_tmp_38 = _registers_13_ext_R3_data[63:56];
      4'b1110:
        casez_tmp_38 = _registers_14_ext_R3_data[63:56];
      default:
        casez_tmp_38 = _registers_15_ext_R3_data[63:56];
    endcase
  end // always @(*)
  wire [6:0]  _io_read_5_value_T_16 = io_read_5_address / 7'h8;
  always @(*) begin
    casez (_io_read_5_value_T_16[3:0])
      4'b0000:
        casez_tmp_39 = _registers_0_ext_R2_data[7:0];
      4'b0001:
        casez_tmp_39 = _registers_1_ext_R2_data[7:0];
      4'b0010:
        casez_tmp_39 = _registers_2_ext_R2_data[7:0];
      4'b0011:
        casez_tmp_39 = _registers_3_ext_R2_data[7:0];
      4'b0100:
        casez_tmp_39 = _registers_4_ext_R2_data[7:0];
      4'b0101:
        casez_tmp_39 = _registers_5_ext_R2_data[7:0];
      4'b0110:
        casez_tmp_39 = _registers_6_ext_R2_data[7:0];
      4'b0111:
        casez_tmp_39 = _registers_7_ext_R2_data[7:0];
      4'b1000:
        casez_tmp_39 = _registers_8_ext_R2_data[7:0];
      4'b1001:
        casez_tmp_39 = _registers_9_ext_R2_data[7:0];
      4'b1010:
        casez_tmp_39 = _registers_10_ext_R2_data[7:0];
      4'b1011:
        casez_tmp_39 = _registers_11_ext_R2_data[7:0];
      4'b1100:
        casez_tmp_39 = _registers_12_ext_R2_data[7:0];
      4'b1101:
        casez_tmp_39 = _registers_13_ext_R2_data[7:0];
      4'b1110:
        casez_tmp_39 = _registers_14_ext_R2_data[7:0];
      default:
        casez_tmp_39 = _registers_15_ext_R2_data[7:0];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_5_value_T_16[3:0])
      4'b0000:
        casez_tmp_40 = _registers_0_ext_R2_data[15:8];
      4'b0001:
        casez_tmp_40 = _registers_1_ext_R2_data[15:8];
      4'b0010:
        casez_tmp_40 = _registers_2_ext_R2_data[15:8];
      4'b0011:
        casez_tmp_40 = _registers_3_ext_R2_data[15:8];
      4'b0100:
        casez_tmp_40 = _registers_4_ext_R2_data[15:8];
      4'b0101:
        casez_tmp_40 = _registers_5_ext_R2_data[15:8];
      4'b0110:
        casez_tmp_40 = _registers_6_ext_R2_data[15:8];
      4'b0111:
        casez_tmp_40 = _registers_7_ext_R2_data[15:8];
      4'b1000:
        casez_tmp_40 = _registers_8_ext_R2_data[15:8];
      4'b1001:
        casez_tmp_40 = _registers_9_ext_R2_data[15:8];
      4'b1010:
        casez_tmp_40 = _registers_10_ext_R2_data[15:8];
      4'b1011:
        casez_tmp_40 = _registers_11_ext_R2_data[15:8];
      4'b1100:
        casez_tmp_40 = _registers_12_ext_R2_data[15:8];
      4'b1101:
        casez_tmp_40 = _registers_13_ext_R2_data[15:8];
      4'b1110:
        casez_tmp_40 = _registers_14_ext_R2_data[15:8];
      default:
        casez_tmp_40 = _registers_15_ext_R2_data[15:8];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_5_value_T_16[3:0])
      4'b0000:
        casez_tmp_41 = _registers_0_ext_R2_data[23:16];
      4'b0001:
        casez_tmp_41 = _registers_1_ext_R2_data[23:16];
      4'b0010:
        casez_tmp_41 = _registers_2_ext_R2_data[23:16];
      4'b0011:
        casez_tmp_41 = _registers_3_ext_R2_data[23:16];
      4'b0100:
        casez_tmp_41 = _registers_4_ext_R2_data[23:16];
      4'b0101:
        casez_tmp_41 = _registers_5_ext_R2_data[23:16];
      4'b0110:
        casez_tmp_41 = _registers_6_ext_R2_data[23:16];
      4'b0111:
        casez_tmp_41 = _registers_7_ext_R2_data[23:16];
      4'b1000:
        casez_tmp_41 = _registers_8_ext_R2_data[23:16];
      4'b1001:
        casez_tmp_41 = _registers_9_ext_R2_data[23:16];
      4'b1010:
        casez_tmp_41 = _registers_10_ext_R2_data[23:16];
      4'b1011:
        casez_tmp_41 = _registers_11_ext_R2_data[23:16];
      4'b1100:
        casez_tmp_41 = _registers_12_ext_R2_data[23:16];
      4'b1101:
        casez_tmp_41 = _registers_13_ext_R2_data[23:16];
      4'b1110:
        casez_tmp_41 = _registers_14_ext_R2_data[23:16];
      default:
        casez_tmp_41 = _registers_15_ext_R2_data[23:16];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_5_value_T_16[3:0])
      4'b0000:
        casez_tmp_42 = _registers_0_ext_R2_data[31:24];
      4'b0001:
        casez_tmp_42 = _registers_1_ext_R2_data[31:24];
      4'b0010:
        casez_tmp_42 = _registers_2_ext_R2_data[31:24];
      4'b0011:
        casez_tmp_42 = _registers_3_ext_R2_data[31:24];
      4'b0100:
        casez_tmp_42 = _registers_4_ext_R2_data[31:24];
      4'b0101:
        casez_tmp_42 = _registers_5_ext_R2_data[31:24];
      4'b0110:
        casez_tmp_42 = _registers_6_ext_R2_data[31:24];
      4'b0111:
        casez_tmp_42 = _registers_7_ext_R2_data[31:24];
      4'b1000:
        casez_tmp_42 = _registers_8_ext_R2_data[31:24];
      4'b1001:
        casez_tmp_42 = _registers_9_ext_R2_data[31:24];
      4'b1010:
        casez_tmp_42 = _registers_10_ext_R2_data[31:24];
      4'b1011:
        casez_tmp_42 = _registers_11_ext_R2_data[31:24];
      4'b1100:
        casez_tmp_42 = _registers_12_ext_R2_data[31:24];
      4'b1101:
        casez_tmp_42 = _registers_13_ext_R2_data[31:24];
      4'b1110:
        casez_tmp_42 = _registers_14_ext_R2_data[31:24];
      default:
        casez_tmp_42 = _registers_15_ext_R2_data[31:24];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_5_value_T_16[3:0])
      4'b0000:
        casez_tmp_43 = _registers_0_ext_R2_data[39:32];
      4'b0001:
        casez_tmp_43 = _registers_1_ext_R2_data[39:32];
      4'b0010:
        casez_tmp_43 = _registers_2_ext_R2_data[39:32];
      4'b0011:
        casez_tmp_43 = _registers_3_ext_R2_data[39:32];
      4'b0100:
        casez_tmp_43 = _registers_4_ext_R2_data[39:32];
      4'b0101:
        casez_tmp_43 = _registers_5_ext_R2_data[39:32];
      4'b0110:
        casez_tmp_43 = _registers_6_ext_R2_data[39:32];
      4'b0111:
        casez_tmp_43 = _registers_7_ext_R2_data[39:32];
      4'b1000:
        casez_tmp_43 = _registers_8_ext_R2_data[39:32];
      4'b1001:
        casez_tmp_43 = _registers_9_ext_R2_data[39:32];
      4'b1010:
        casez_tmp_43 = _registers_10_ext_R2_data[39:32];
      4'b1011:
        casez_tmp_43 = _registers_11_ext_R2_data[39:32];
      4'b1100:
        casez_tmp_43 = _registers_12_ext_R2_data[39:32];
      4'b1101:
        casez_tmp_43 = _registers_13_ext_R2_data[39:32];
      4'b1110:
        casez_tmp_43 = _registers_14_ext_R2_data[39:32];
      default:
        casez_tmp_43 = _registers_15_ext_R2_data[39:32];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_5_value_T_16[3:0])
      4'b0000:
        casez_tmp_44 = _registers_0_ext_R2_data[47:40];
      4'b0001:
        casez_tmp_44 = _registers_1_ext_R2_data[47:40];
      4'b0010:
        casez_tmp_44 = _registers_2_ext_R2_data[47:40];
      4'b0011:
        casez_tmp_44 = _registers_3_ext_R2_data[47:40];
      4'b0100:
        casez_tmp_44 = _registers_4_ext_R2_data[47:40];
      4'b0101:
        casez_tmp_44 = _registers_5_ext_R2_data[47:40];
      4'b0110:
        casez_tmp_44 = _registers_6_ext_R2_data[47:40];
      4'b0111:
        casez_tmp_44 = _registers_7_ext_R2_data[47:40];
      4'b1000:
        casez_tmp_44 = _registers_8_ext_R2_data[47:40];
      4'b1001:
        casez_tmp_44 = _registers_9_ext_R2_data[47:40];
      4'b1010:
        casez_tmp_44 = _registers_10_ext_R2_data[47:40];
      4'b1011:
        casez_tmp_44 = _registers_11_ext_R2_data[47:40];
      4'b1100:
        casez_tmp_44 = _registers_12_ext_R2_data[47:40];
      4'b1101:
        casez_tmp_44 = _registers_13_ext_R2_data[47:40];
      4'b1110:
        casez_tmp_44 = _registers_14_ext_R2_data[47:40];
      default:
        casez_tmp_44 = _registers_15_ext_R2_data[47:40];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_5_value_T_16[3:0])
      4'b0000:
        casez_tmp_45 = _registers_0_ext_R2_data[55:48];
      4'b0001:
        casez_tmp_45 = _registers_1_ext_R2_data[55:48];
      4'b0010:
        casez_tmp_45 = _registers_2_ext_R2_data[55:48];
      4'b0011:
        casez_tmp_45 = _registers_3_ext_R2_data[55:48];
      4'b0100:
        casez_tmp_45 = _registers_4_ext_R2_data[55:48];
      4'b0101:
        casez_tmp_45 = _registers_5_ext_R2_data[55:48];
      4'b0110:
        casez_tmp_45 = _registers_6_ext_R2_data[55:48];
      4'b0111:
        casez_tmp_45 = _registers_7_ext_R2_data[55:48];
      4'b1000:
        casez_tmp_45 = _registers_8_ext_R2_data[55:48];
      4'b1001:
        casez_tmp_45 = _registers_9_ext_R2_data[55:48];
      4'b1010:
        casez_tmp_45 = _registers_10_ext_R2_data[55:48];
      4'b1011:
        casez_tmp_45 = _registers_11_ext_R2_data[55:48];
      4'b1100:
        casez_tmp_45 = _registers_12_ext_R2_data[55:48];
      4'b1101:
        casez_tmp_45 = _registers_13_ext_R2_data[55:48];
      4'b1110:
        casez_tmp_45 = _registers_14_ext_R2_data[55:48];
      default:
        casez_tmp_45 = _registers_15_ext_R2_data[55:48];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_5_value_T_16[3:0])
      4'b0000:
        casez_tmp_46 = _registers_0_ext_R2_data[63:56];
      4'b0001:
        casez_tmp_46 = _registers_1_ext_R2_data[63:56];
      4'b0010:
        casez_tmp_46 = _registers_2_ext_R2_data[63:56];
      4'b0011:
        casez_tmp_46 = _registers_3_ext_R2_data[63:56];
      4'b0100:
        casez_tmp_46 = _registers_4_ext_R2_data[63:56];
      4'b0101:
        casez_tmp_46 = _registers_5_ext_R2_data[63:56];
      4'b0110:
        casez_tmp_46 = _registers_6_ext_R2_data[63:56];
      4'b0111:
        casez_tmp_46 = _registers_7_ext_R2_data[63:56];
      4'b1000:
        casez_tmp_46 = _registers_8_ext_R2_data[63:56];
      4'b1001:
        casez_tmp_46 = _registers_9_ext_R2_data[63:56];
      4'b1010:
        casez_tmp_46 = _registers_10_ext_R2_data[63:56];
      4'b1011:
        casez_tmp_46 = _registers_11_ext_R2_data[63:56];
      4'b1100:
        casez_tmp_46 = _registers_12_ext_R2_data[63:56];
      4'b1101:
        casez_tmp_46 = _registers_13_ext_R2_data[63:56];
      4'b1110:
        casez_tmp_46 = _registers_14_ext_R2_data[63:56];
      default:
        casez_tmp_46 = _registers_15_ext_R2_data[63:56];
    endcase
  end // always @(*)
  wire [6:0]  _io_read_6_value_T_16 = io_read_6_address / 7'h8;
  always @(*) begin
    casez (_io_read_6_value_T_16[3:0])
      4'b0000:
        casez_tmp_47 = _registers_0_ext_R1_data[7:0];
      4'b0001:
        casez_tmp_47 = _registers_1_ext_R1_data[7:0];
      4'b0010:
        casez_tmp_47 = _registers_2_ext_R1_data[7:0];
      4'b0011:
        casez_tmp_47 = _registers_3_ext_R1_data[7:0];
      4'b0100:
        casez_tmp_47 = _registers_4_ext_R1_data[7:0];
      4'b0101:
        casez_tmp_47 = _registers_5_ext_R1_data[7:0];
      4'b0110:
        casez_tmp_47 = _registers_6_ext_R1_data[7:0];
      4'b0111:
        casez_tmp_47 = _registers_7_ext_R1_data[7:0];
      4'b1000:
        casez_tmp_47 = _registers_8_ext_R1_data[7:0];
      4'b1001:
        casez_tmp_47 = _registers_9_ext_R1_data[7:0];
      4'b1010:
        casez_tmp_47 = _registers_10_ext_R1_data[7:0];
      4'b1011:
        casez_tmp_47 = _registers_11_ext_R1_data[7:0];
      4'b1100:
        casez_tmp_47 = _registers_12_ext_R1_data[7:0];
      4'b1101:
        casez_tmp_47 = _registers_13_ext_R1_data[7:0];
      4'b1110:
        casez_tmp_47 = _registers_14_ext_R1_data[7:0];
      default:
        casez_tmp_47 = _registers_15_ext_R1_data[7:0];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_6_value_T_16[3:0])
      4'b0000:
        casez_tmp_48 = _registers_0_ext_R1_data[15:8];
      4'b0001:
        casez_tmp_48 = _registers_1_ext_R1_data[15:8];
      4'b0010:
        casez_tmp_48 = _registers_2_ext_R1_data[15:8];
      4'b0011:
        casez_tmp_48 = _registers_3_ext_R1_data[15:8];
      4'b0100:
        casez_tmp_48 = _registers_4_ext_R1_data[15:8];
      4'b0101:
        casez_tmp_48 = _registers_5_ext_R1_data[15:8];
      4'b0110:
        casez_tmp_48 = _registers_6_ext_R1_data[15:8];
      4'b0111:
        casez_tmp_48 = _registers_7_ext_R1_data[15:8];
      4'b1000:
        casez_tmp_48 = _registers_8_ext_R1_data[15:8];
      4'b1001:
        casez_tmp_48 = _registers_9_ext_R1_data[15:8];
      4'b1010:
        casez_tmp_48 = _registers_10_ext_R1_data[15:8];
      4'b1011:
        casez_tmp_48 = _registers_11_ext_R1_data[15:8];
      4'b1100:
        casez_tmp_48 = _registers_12_ext_R1_data[15:8];
      4'b1101:
        casez_tmp_48 = _registers_13_ext_R1_data[15:8];
      4'b1110:
        casez_tmp_48 = _registers_14_ext_R1_data[15:8];
      default:
        casez_tmp_48 = _registers_15_ext_R1_data[15:8];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_6_value_T_16[3:0])
      4'b0000:
        casez_tmp_49 = _registers_0_ext_R1_data[23:16];
      4'b0001:
        casez_tmp_49 = _registers_1_ext_R1_data[23:16];
      4'b0010:
        casez_tmp_49 = _registers_2_ext_R1_data[23:16];
      4'b0011:
        casez_tmp_49 = _registers_3_ext_R1_data[23:16];
      4'b0100:
        casez_tmp_49 = _registers_4_ext_R1_data[23:16];
      4'b0101:
        casez_tmp_49 = _registers_5_ext_R1_data[23:16];
      4'b0110:
        casez_tmp_49 = _registers_6_ext_R1_data[23:16];
      4'b0111:
        casez_tmp_49 = _registers_7_ext_R1_data[23:16];
      4'b1000:
        casez_tmp_49 = _registers_8_ext_R1_data[23:16];
      4'b1001:
        casez_tmp_49 = _registers_9_ext_R1_data[23:16];
      4'b1010:
        casez_tmp_49 = _registers_10_ext_R1_data[23:16];
      4'b1011:
        casez_tmp_49 = _registers_11_ext_R1_data[23:16];
      4'b1100:
        casez_tmp_49 = _registers_12_ext_R1_data[23:16];
      4'b1101:
        casez_tmp_49 = _registers_13_ext_R1_data[23:16];
      4'b1110:
        casez_tmp_49 = _registers_14_ext_R1_data[23:16];
      default:
        casez_tmp_49 = _registers_15_ext_R1_data[23:16];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_6_value_T_16[3:0])
      4'b0000:
        casez_tmp_50 = _registers_0_ext_R1_data[31:24];
      4'b0001:
        casez_tmp_50 = _registers_1_ext_R1_data[31:24];
      4'b0010:
        casez_tmp_50 = _registers_2_ext_R1_data[31:24];
      4'b0011:
        casez_tmp_50 = _registers_3_ext_R1_data[31:24];
      4'b0100:
        casez_tmp_50 = _registers_4_ext_R1_data[31:24];
      4'b0101:
        casez_tmp_50 = _registers_5_ext_R1_data[31:24];
      4'b0110:
        casez_tmp_50 = _registers_6_ext_R1_data[31:24];
      4'b0111:
        casez_tmp_50 = _registers_7_ext_R1_data[31:24];
      4'b1000:
        casez_tmp_50 = _registers_8_ext_R1_data[31:24];
      4'b1001:
        casez_tmp_50 = _registers_9_ext_R1_data[31:24];
      4'b1010:
        casez_tmp_50 = _registers_10_ext_R1_data[31:24];
      4'b1011:
        casez_tmp_50 = _registers_11_ext_R1_data[31:24];
      4'b1100:
        casez_tmp_50 = _registers_12_ext_R1_data[31:24];
      4'b1101:
        casez_tmp_50 = _registers_13_ext_R1_data[31:24];
      4'b1110:
        casez_tmp_50 = _registers_14_ext_R1_data[31:24];
      default:
        casez_tmp_50 = _registers_15_ext_R1_data[31:24];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_6_value_T_16[3:0])
      4'b0000:
        casez_tmp_51 = _registers_0_ext_R1_data[39:32];
      4'b0001:
        casez_tmp_51 = _registers_1_ext_R1_data[39:32];
      4'b0010:
        casez_tmp_51 = _registers_2_ext_R1_data[39:32];
      4'b0011:
        casez_tmp_51 = _registers_3_ext_R1_data[39:32];
      4'b0100:
        casez_tmp_51 = _registers_4_ext_R1_data[39:32];
      4'b0101:
        casez_tmp_51 = _registers_5_ext_R1_data[39:32];
      4'b0110:
        casez_tmp_51 = _registers_6_ext_R1_data[39:32];
      4'b0111:
        casez_tmp_51 = _registers_7_ext_R1_data[39:32];
      4'b1000:
        casez_tmp_51 = _registers_8_ext_R1_data[39:32];
      4'b1001:
        casez_tmp_51 = _registers_9_ext_R1_data[39:32];
      4'b1010:
        casez_tmp_51 = _registers_10_ext_R1_data[39:32];
      4'b1011:
        casez_tmp_51 = _registers_11_ext_R1_data[39:32];
      4'b1100:
        casez_tmp_51 = _registers_12_ext_R1_data[39:32];
      4'b1101:
        casez_tmp_51 = _registers_13_ext_R1_data[39:32];
      4'b1110:
        casez_tmp_51 = _registers_14_ext_R1_data[39:32];
      default:
        casez_tmp_51 = _registers_15_ext_R1_data[39:32];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_6_value_T_16[3:0])
      4'b0000:
        casez_tmp_52 = _registers_0_ext_R1_data[47:40];
      4'b0001:
        casez_tmp_52 = _registers_1_ext_R1_data[47:40];
      4'b0010:
        casez_tmp_52 = _registers_2_ext_R1_data[47:40];
      4'b0011:
        casez_tmp_52 = _registers_3_ext_R1_data[47:40];
      4'b0100:
        casez_tmp_52 = _registers_4_ext_R1_data[47:40];
      4'b0101:
        casez_tmp_52 = _registers_5_ext_R1_data[47:40];
      4'b0110:
        casez_tmp_52 = _registers_6_ext_R1_data[47:40];
      4'b0111:
        casez_tmp_52 = _registers_7_ext_R1_data[47:40];
      4'b1000:
        casez_tmp_52 = _registers_8_ext_R1_data[47:40];
      4'b1001:
        casez_tmp_52 = _registers_9_ext_R1_data[47:40];
      4'b1010:
        casez_tmp_52 = _registers_10_ext_R1_data[47:40];
      4'b1011:
        casez_tmp_52 = _registers_11_ext_R1_data[47:40];
      4'b1100:
        casez_tmp_52 = _registers_12_ext_R1_data[47:40];
      4'b1101:
        casez_tmp_52 = _registers_13_ext_R1_data[47:40];
      4'b1110:
        casez_tmp_52 = _registers_14_ext_R1_data[47:40];
      default:
        casez_tmp_52 = _registers_15_ext_R1_data[47:40];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_6_value_T_16[3:0])
      4'b0000:
        casez_tmp_53 = _registers_0_ext_R1_data[55:48];
      4'b0001:
        casez_tmp_53 = _registers_1_ext_R1_data[55:48];
      4'b0010:
        casez_tmp_53 = _registers_2_ext_R1_data[55:48];
      4'b0011:
        casez_tmp_53 = _registers_3_ext_R1_data[55:48];
      4'b0100:
        casez_tmp_53 = _registers_4_ext_R1_data[55:48];
      4'b0101:
        casez_tmp_53 = _registers_5_ext_R1_data[55:48];
      4'b0110:
        casez_tmp_53 = _registers_6_ext_R1_data[55:48];
      4'b0111:
        casez_tmp_53 = _registers_7_ext_R1_data[55:48];
      4'b1000:
        casez_tmp_53 = _registers_8_ext_R1_data[55:48];
      4'b1001:
        casez_tmp_53 = _registers_9_ext_R1_data[55:48];
      4'b1010:
        casez_tmp_53 = _registers_10_ext_R1_data[55:48];
      4'b1011:
        casez_tmp_53 = _registers_11_ext_R1_data[55:48];
      4'b1100:
        casez_tmp_53 = _registers_12_ext_R1_data[55:48];
      4'b1101:
        casez_tmp_53 = _registers_13_ext_R1_data[55:48];
      4'b1110:
        casez_tmp_53 = _registers_14_ext_R1_data[55:48];
      default:
        casez_tmp_53 = _registers_15_ext_R1_data[55:48];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_6_value_T_16[3:0])
      4'b0000:
        casez_tmp_54 = _registers_0_ext_R1_data[63:56];
      4'b0001:
        casez_tmp_54 = _registers_1_ext_R1_data[63:56];
      4'b0010:
        casez_tmp_54 = _registers_2_ext_R1_data[63:56];
      4'b0011:
        casez_tmp_54 = _registers_3_ext_R1_data[63:56];
      4'b0100:
        casez_tmp_54 = _registers_4_ext_R1_data[63:56];
      4'b0101:
        casez_tmp_54 = _registers_5_ext_R1_data[63:56];
      4'b0110:
        casez_tmp_54 = _registers_6_ext_R1_data[63:56];
      4'b0111:
        casez_tmp_54 = _registers_7_ext_R1_data[63:56];
      4'b1000:
        casez_tmp_54 = _registers_8_ext_R1_data[63:56];
      4'b1001:
        casez_tmp_54 = _registers_9_ext_R1_data[63:56];
      4'b1010:
        casez_tmp_54 = _registers_10_ext_R1_data[63:56];
      4'b1011:
        casez_tmp_54 = _registers_11_ext_R1_data[63:56];
      4'b1100:
        casez_tmp_54 = _registers_12_ext_R1_data[63:56];
      4'b1101:
        casez_tmp_54 = _registers_13_ext_R1_data[63:56];
      4'b1110:
        casez_tmp_54 = _registers_14_ext_R1_data[63:56];
      default:
        casez_tmp_54 = _registers_15_ext_R1_data[63:56];
    endcase
  end // always @(*)
  wire [6:0]  _io_read_7_value_T_16 = io_read_7_address / 7'h8;
  always @(*) begin
    casez (_io_read_7_value_T_16[3:0])
      4'b0000:
        casez_tmp_55 = _registers_0_ext_R0_data[7:0];
      4'b0001:
        casez_tmp_55 = _registers_1_ext_R0_data[7:0];
      4'b0010:
        casez_tmp_55 = _registers_2_ext_R0_data[7:0];
      4'b0011:
        casez_tmp_55 = _registers_3_ext_R0_data[7:0];
      4'b0100:
        casez_tmp_55 = _registers_4_ext_R0_data[7:0];
      4'b0101:
        casez_tmp_55 = _registers_5_ext_R0_data[7:0];
      4'b0110:
        casez_tmp_55 = _registers_6_ext_R0_data[7:0];
      4'b0111:
        casez_tmp_55 = _registers_7_ext_R0_data[7:0];
      4'b1000:
        casez_tmp_55 = _registers_8_ext_R0_data[7:0];
      4'b1001:
        casez_tmp_55 = _registers_9_ext_R0_data[7:0];
      4'b1010:
        casez_tmp_55 = _registers_10_ext_R0_data[7:0];
      4'b1011:
        casez_tmp_55 = _registers_11_ext_R0_data[7:0];
      4'b1100:
        casez_tmp_55 = _registers_12_ext_R0_data[7:0];
      4'b1101:
        casez_tmp_55 = _registers_13_ext_R0_data[7:0];
      4'b1110:
        casez_tmp_55 = _registers_14_ext_R0_data[7:0];
      default:
        casez_tmp_55 = _registers_15_ext_R0_data[7:0];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_7_value_T_16[3:0])
      4'b0000:
        casez_tmp_56 = _registers_0_ext_R0_data[15:8];
      4'b0001:
        casez_tmp_56 = _registers_1_ext_R0_data[15:8];
      4'b0010:
        casez_tmp_56 = _registers_2_ext_R0_data[15:8];
      4'b0011:
        casez_tmp_56 = _registers_3_ext_R0_data[15:8];
      4'b0100:
        casez_tmp_56 = _registers_4_ext_R0_data[15:8];
      4'b0101:
        casez_tmp_56 = _registers_5_ext_R0_data[15:8];
      4'b0110:
        casez_tmp_56 = _registers_6_ext_R0_data[15:8];
      4'b0111:
        casez_tmp_56 = _registers_7_ext_R0_data[15:8];
      4'b1000:
        casez_tmp_56 = _registers_8_ext_R0_data[15:8];
      4'b1001:
        casez_tmp_56 = _registers_9_ext_R0_data[15:8];
      4'b1010:
        casez_tmp_56 = _registers_10_ext_R0_data[15:8];
      4'b1011:
        casez_tmp_56 = _registers_11_ext_R0_data[15:8];
      4'b1100:
        casez_tmp_56 = _registers_12_ext_R0_data[15:8];
      4'b1101:
        casez_tmp_56 = _registers_13_ext_R0_data[15:8];
      4'b1110:
        casez_tmp_56 = _registers_14_ext_R0_data[15:8];
      default:
        casez_tmp_56 = _registers_15_ext_R0_data[15:8];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_7_value_T_16[3:0])
      4'b0000:
        casez_tmp_57 = _registers_0_ext_R0_data[23:16];
      4'b0001:
        casez_tmp_57 = _registers_1_ext_R0_data[23:16];
      4'b0010:
        casez_tmp_57 = _registers_2_ext_R0_data[23:16];
      4'b0011:
        casez_tmp_57 = _registers_3_ext_R0_data[23:16];
      4'b0100:
        casez_tmp_57 = _registers_4_ext_R0_data[23:16];
      4'b0101:
        casez_tmp_57 = _registers_5_ext_R0_data[23:16];
      4'b0110:
        casez_tmp_57 = _registers_6_ext_R0_data[23:16];
      4'b0111:
        casez_tmp_57 = _registers_7_ext_R0_data[23:16];
      4'b1000:
        casez_tmp_57 = _registers_8_ext_R0_data[23:16];
      4'b1001:
        casez_tmp_57 = _registers_9_ext_R0_data[23:16];
      4'b1010:
        casez_tmp_57 = _registers_10_ext_R0_data[23:16];
      4'b1011:
        casez_tmp_57 = _registers_11_ext_R0_data[23:16];
      4'b1100:
        casez_tmp_57 = _registers_12_ext_R0_data[23:16];
      4'b1101:
        casez_tmp_57 = _registers_13_ext_R0_data[23:16];
      4'b1110:
        casez_tmp_57 = _registers_14_ext_R0_data[23:16];
      default:
        casez_tmp_57 = _registers_15_ext_R0_data[23:16];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_7_value_T_16[3:0])
      4'b0000:
        casez_tmp_58 = _registers_0_ext_R0_data[31:24];
      4'b0001:
        casez_tmp_58 = _registers_1_ext_R0_data[31:24];
      4'b0010:
        casez_tmp_58 = _registers_2_ext_R0_data[31:24];
      4'b0011:
        casez_tmp_58 = _registers_3_ext_R0_data[31:24];
      4'b0100:
        casez_tmp_58 = _registers_4_ext_R0_data[31:24];
      4'b0101:
        casez_tmp_58 = _registers_5_ext_R0_data[31:24];
      4'b0110:
        casez_tmp_58 = _registers_6_ext_R0_data[31:24];
      4'b0111:
        casez_tmp_58 = _registers_7_ext_R0_data[31:24];
      4'b1000:
        casez_tmp_58 = _registers_8_ext_R0_data[31:24];
      4'b1001:
        casez_tmp_58 = _registers_9_ext_R0_data[31:24];
      4'b1010:
        casez_tmp_58 = _registers_10_ext_R0_data[31:24];
      4'b1011:
        casez_tmp_58 = _registers_11_ext_R0_data[31:24];
      4'b1100:
        casez_tmp_58 = _registers_12_ext_R0_data[31:24];
      4'b1101:
        casez_tmp_58 = _registers_13_ext_R0_data[31:24];
      4'b1110:
        casez_tmp_58 = _registers_14_ext_R0_data[31:24];
      default:
        casez_tmp_58 = _registers_15_ext_R0_data[31:24];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_7_value_T_16[3:0])
      4'b0000:
        casez_tmp_59 = _registers_0_ext_R0_data[39:32];
      4'b0001:
        casez_tmp_59 = _registers_1_ext_R0_data[39:32];
      4'b0010:
        casez_tmp_59 = _registers_2_ext_R0_data[39:32];
      4'b0011:
        casez_tmp_59 = _registers_3_ext_R0_data[39:32];
      4'b0100:
        casez_tmp_59 = _registers_4_ext_R0_data[39:32];
      4'b0101:
        casez_tmp_59 = _registers_5_ext_R0_data[39:32];
      4'b0110:
        casez_tmp_59 = _registers_6_ext_R0_data[39:32];
      4'b0111:
        casez_tmp_59 = _registers_7_ext_R0_data[39:32];
      4'b1000:
        casez_tmp_59 = _registers_8_ext_R0_data[39:32];
      4'b1001:
        casez_tmp_59 = _registers_9_ext_R0_data[39:32];
      4'b1010:
        casez_tmp_59 = _registers_10_ext_R0_data[39:32];
      4'b1011:
        casez_tmp_59 = _registers_11_ext_R0_data[39:32];
      4'b1100:
        casez_tmp_59 = _registers_12_ext_R0_data[39:32];
      4'b1101:
        casez_tmp_59 = _registers_13_ext_R0_data[39:32];
      4'b1110:
        casez_tmp_59 = _registers_14_ext_R0_data[39:32];
      default:
        casez_tmp_59 = _registers_15_ext_R0_data[39:32];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_7_value_T_16[3:0])
      4'b0000:
        casez_tmp_60 = _registers_0_ext_R0_data[47:40];
      4'b0001:
        casez_tmp_60 = _registers_1_ext_R0_data[47:40];
      4'b0010:
        casez_tmp_60 = _registers_2_ext_R0_data[47:40];
      4'b0011:
        casez_tmp_60 = _registers_3_ext_R0_data[47:40];
      4'b0100:
        casez_tmp_60 = _registers_4_ext_R0_data[47:40];
      4'b0101:
        casez_tmp_60 = _registers_5_ext_R0_data[47:40];
      4'b0110:
        casez_tmp_60 = _registers_6_ext_R0_data[47:40];
      4'b0111:
        casez_tmp_60 = _registers_7_ext_R0_data[47:40];
      4'b1000:
        casez_tmp_60 = _registers_8_ext_R0_data[47:40];
      4'b1001:
        casez_tmp_60 = _registers_9_ext_R0_data[47:40];
      4'b1010:
        casez_tmp_60 = _registers_10_ext_R0_data[47:40];
      4'b1011:
        casez_tmp_60 = _registers_11_ext_R0_data[47:40];
      4'b1100:
        casez_tmp_60 = _registers_12_ext_R0_data[47:40];
      4'b1101:
        casez_tmp_60 = _registers_13_ext_R0_data[47:40];
      4'b1110:
        casez_tmp_60 = _registers_14_ext_R0_data[47:40];
      default:
        casez_tmp_60 = _registers_15_ext_R0_data[47:40];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_7_value_T_16[3:0])
      4'b0000:
        casez_tmp_61 = _registers_0_ext_R0_data[55:48];
      4'b0001:
        casez_tmp_61 = _registers_1_ext_R0_data[55:48];
      4'b0010:
        casez_tmp_61 = _registers_2_ext_R0_data[55:48];
      4'b0011:
        casez_tmp_61 = _registers_3_ext_R0_data[55:48];
      4'b0100:
        casez_tmp_61 = _registers_4_ext_R0_data[55:48];
      4'b0101:
        casez_tmp_61 = _registers_5_ext_R0_data[55:48];
      4'b0110:
        casez_tmp_61 = _registers_6_ext_R0_data[55:48];
      4'b0111:
        casez_tmp_61 = _registers_7_ext_R0_data[55:48];
      4'b1000:
        casez_tmp_61 = _registers_8_ext_R0_data[55:48];
      4'b1001:
        casez_tmp_61 = _registers_9_ext_R0_data[55:48];
      4'b1010:
        casez_tmp_61 = _registers_10_ext_R0_data[55:48];
      4'b1011:
        casez_tmp_61 = _registers_11_ext_R0_data[55:48];
      4'b1100:
        casez_tmp_61 = _registers_12_ext_R0_data[55:48];
      4'b1101:
        casez_tmp_61 = _registers_13_ext_R0_data[55:48];
      4'b1110:
        casez_tmp_61 = _registers_14_ext_R0_data[55:48];
      default:
        casez_tmp_61 = _registers_15_ext_R0_data[55:48];
    endcase
  end // always @(*)
  always @(*) begin
    casez (_io_read_7_value_T_16[3:0])
      4'b0000:
        casez_tmp_62 = _registers_0_ext_R0_data[63:56];
      4'b0001:
        casez_tmp_62 = _registers_1_ext_R0_data[63:56];
      4'b0010:
        casez_tmp_62 = _registers_2_ext_R0_data[63:56];
      4'b0011:
        casez_tmp_62 = _registers_3_ext_R0_data[63:56];
      4'b0100:
        casez_tmp_62 = _registers_4_ext_R0_data[63:56];
      4'b0101:
        casez_tmp_62 = _registers_5_ext_R0_data[63:56];
      4'b0110:
        casez_tmp_62 = _registers_6_ext_R0_data[63:56];
      4'b0111:
        casez_tmp_62 = _registers_7_ext_R0_data[63:56];
      4'b1000:
        casez_tmp_62 = _registers_8_ext_R0_data[63:56];
      4'b1001:
        casez_tmp_62 = _registers_9_ext_R0_data[63:56];
      4'b1010:
        casez_tmp_62 = _registers_10_ext_R0_data[63:56];
      4'b1011:
        casez_tmp_62 = _registers_11_ext_R0_data[63:56];
      4'b1100:
        casez_tmp_62 = _registers_12_ext_R0_data[63:56];
      4'b1101:
        casez_tmp_62 = _registers_13_ext_R0_data[63:56];
      4'b1110:
        casez_tmp_62 = _registers_14_ext_R0_data[63:56];
      default:
        casez_tmp_62 = _registers_15_ext_R0_data[63:56];
    endcase
  end // always @(*)
  registers_8x64 registers_0_ext (
    .R0_addr (io_read_7_address[2:0]),
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .R1_addr (io_read_6_address[2:0]),
    .R1_en   (1'h1),
    .R1_clk  (clock),
    .R2_addr (io_read_5_address[2:0]),
    .R2_en   (1'h1),
    .R2_clk  (clock),
    .R3_addr (io_read_4_address[2:0]),
    .R3_en   (1'h1),
    .R3_clk  (clock),
    .R4_addr (io_read_3_address[2:0]),
    .R4_en   (1'h1),
    .R4_clk  (clock),
    .R5_addr (io_read_2_address[2:0]),
    .R5_en   (1'h1),
    .R5_clk  (clock),
    .R6_addr (io_read_1_address[2:0]),
    .R6_en   (1'h1),
    .R6_clk  (clock),
    .R7_addr (io_read_0_address[2:0]),
    .R7_en   (1'h1),
    .R7_clk  (clock),
    .W0_addr (io_write_3_address[2:0]),
    .W0_en   (io_write_3_write & _GEN_6 == 7'h0),
    .W0_clk  (clock),
    .W0_data (io_write_3_value),
    .W0_mask (_GEN_2),
    .W1_addr (io_write_2_address[2:0]),
    .W1_en   (io_write_2_write & _GEN_5 == 7'h0),
    .W1_clk  (clock),
    .W1_data (io_write_2_value),
    .W1_mask (_GEN_1),
    .W2_addr (io_write_1_address[2:0]),
    .W2_en   (io_write_1_write & _GEN_4 == 7'h0),
    .W2_clk  (clock),
    .W2_data (io_write_1_value),
    .W2_mask (_GEN_0),
    .W3_addr (io_write_0_address[2:0]),
    .W3_en   (io_write_0_write & _GEN_3 == 7'h0),
    .W3_clk  (clock),
    .W3_data (io_write_0_value),
    .W3_mask (_GEN),
    .R0_data (_registers_0_ext_R0_data),
    .R1_data (_registers_0_ext_R1_data),
    .R2_data (_registers_0_ext_R2_data),
    .R3_data (_registers_0_ext_R3_data),
    .R4_data (_registers_0_ext_R4_data),
    .R5_data (_registers_0_ext_R5_data),
    .R6_data (_registers_0_ext_R6_data),
    .R7_data (_registers_0_ext_R7_data)
  );
  registers_8x64 registers_1_ext (
    .R0_addr (io_read_7_address[2:0]),
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .R1_addr (io_read_6_address[2:0]),
    .R1_en   (1'h1),
    .R1_clk  (clock),
    .R2_addr (io_read_5_address[2:0]),
    .R2_en   (1'h1),
    .R2_clk  (clock),
    .R3_addr (io_read_4_address[2:0]),
    .R3_en   (1'h1),
    .R3_clk  (clock),
    .R4_addr (io_read_3_address[2:0]),
    .R4_en   (1'h1),
    .R4_clk  (clock),
    .R5_addr (io_read_2_address[2:0]),
    .R5_en   (1'h1),
    .R5_clk  (clock),
    .R6_addr (io_read_1_address[2:0]),
    .R6_en   (1'h1),
    .R6_clk  (clock),
    .R7_addr (io_read_0_address[2:0]),
    .R7_en   (1'h1),
    .R7_clk  (clock),
    .W0_addr (io_write_3_address[2:0]),
    .W0_en   (io_write_3_write & _GEN_6 == 7'h1),
    .W0_clk  (clock),
    .W0_data (io_write_3_value),
    .W0_mask (_GEN_2),
    .W1_addr (io_write_2_address[2:0]),
    .W1_en   (io_write_2_write & _GEN_5 == 7'h1),
    .W1_clk  (clock),
    .W1_data (io_write_2_value),
    .W1_mask (_GEN_1),
    .W2_addr (io_write_1_address[2:0]),
    .W2_en   (io_write_1_write & _GEN_4 == 7'h1),
    .W2_clk  (clock),
    .W2_data (io_write_1_value),
    .W2_mask (_GEN_0),
    .W3_addr (io_write_0_address[2:0]),
    .W3_en   (io_write_0_write & _GEN_3 == 7'h1),
    .W3_clk  (clock),
    .W3_data (io_write_0_value),
    .W3_mask (_GEN),
    .R0_data (_registers_1_ext_R0_data),
    .R1_data (_registers_1_ext_R1_data),
    .R2_data (_registers_1_ext_R2_data),
    .R3_data (_registers_1_ext_R3_data),
    .R4_data (_registers_1_ext_R4_data),
    .R5_data (_registers_1_ext_R5_data),
    .R6_data (_registers_1_ext_R6_data),
    .R7_data (_registers_1_ext_R7_data)
  );
  registers_8x64 registers_2_ext (
    .R0_addr (io_read_7_address[2:0]),
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .R1_addr (io_read_6_address[2:0]),
    .R1_en   (1'h1),
    .R1_clk  (clock),
    .R2_addr (io_read_5_address[2:0]),
    .R2_en   (1'h1),
    .R2_clk  (clock),
    .R3_addr (io_read_4_address[2:0]),
    .R3_en   (1'h1),
    .R3_clk  (clock),
    .R4_addr (io_read_3_address[2:0]),
    .R4_en   (1'h1),
    .R4_clk  (clock),
    .R5_addr (io_read_2_address[2:0]),
    .R5_en   (1'h1),
    .R5_clk  (clock),
    .R6_addr (io_read_1_address[2:0]),
    .R6_en   (1'h1),
    .R6_clk  (clock),
    .R7_addr (io_read_0_address[2:0]),
    .R7_en   (1'h1),
    .R7_clk  (clock),
    .W0_addr (io_write_2_address[2:0]),
    .W0_en   (io_write_2_write & _GEN_5 == 7'h2),
    .W0_clk  (clock),
    .W0_data (io_write_2_value),
    .W0_mask (_GEN_1),
    .W1_addr (io_write_0_address[2:0]),
    .W1_en   (io_write_0_write & _GEN_3 == 7'h2),
    .W1_clk  (clock),
    .W1_data (io_write_0_value),
    .W1_mask (_GEN),
    .W2_addr (io_write_1_address[2:0]),
    .W2_en   (io_write_1_write & _GEN_4 == 7'h2),
    .W2_clk  (clock),
    .W2_data (io_write_1_value),
    .W2_mask (_GEN_0),
    .W3_addr (io_write_3_address[2:0]),
    .W3_en   (io_write_3_write & _GEN_6 == 7'h2),
    .W3_clk  (clock),
    .W3_data (io_write_3_value),
    .W3_mask (_GEN_2),
    .R0_data (_registers_2_ext_R0_data),
    .R1_data (_registers_2_ext_R1_data),
    .R2_data (_registers_2_ext_R2_data),
    .R3_data (_registers_2_ext_R3_data),
    .R4_data (_registers_2_ext_R4_data),
    .R5_data (_registers_2_ext_R5_data),
    .R6_data (_registers_2_ext_R6_data),
    .R7_data (_registers_2_ext_R7_data)
  );
  registers_8x64 registers_3_ext (
    .R0_addr (io_read_7_address[2:0]),
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .R1_addr (io_read_6_address[2:0]),
    .R1_en   (1'h1),
    .R1_clk  (clock),
    .R2_addr (io_read_5_address[2:0]),
    .R2_en   (1'h1),
    .R2_clk  (clock),
    .R3_addr (io_read_4_address[2:0]),
    .R3_en   (1'h1),
    .R3_clk  (clock),
    .R4_addr (io_read_3_address[2:0]),
    .R4_en   (1'h1),
    .R4_clk  (clock),
    .R5_addr (io_read_2_address[2:0]),
    .R5_en   (1'h1),
    .R5_clk  (clock),
    .R6_addr (io_read_1_address[2:0]),
    .R6_en   (1'h1),
    .R6_clk  (clock),
    .R7_addr (io_read_0_address[2:0]),
    .R7_en   (1'h1),
    .R7_clk  (clock),
    .W0_addr (io_write_2_address[2:0]),
    .W0_en   (io_write_2_write & _GEN_5 == 7'h3),
    .W0_clk  (clock),
    .W0_data (io_write_2_value),
    .W0_mask (_GEN_1),
    .W1_addr (io_write_0_address[2:0]),
    .W1_en   (io_write_0_write & _GEN_3 == 7'h3),
    .W1_clk  (clock),
    .W1_data (io_write_0_value),
    .W1_mask (_GEN),
    .W2_addr (io_write_1_address[2:0]),
    .W2_en   (io_write_1_write & _GEN_4 == 7'h3),
    .W2_clk  (clock),
    .W2_data (io_write_1_value),
    .W2_mask (_GEN_0),
    .W3_addr (io_write_3_address[2:0]),
    .W3_en   (io_write_3_write & _GEN_6 == 7'h3),
    .W3_clk  (clock),
    .W3_data (io_write_3_value),
    .W3_mask (_GEN_2),
    .R0_data (_registers_3_ext_R0_data),
    .R1_data (_registers_3_ext_R1_data),
    .R2_data (_registers_3_ext_R2_data),
    .R3_data (_registers_3_ext_R3_data),
    .R4_data (_registers_3_ext_R4_data),
    .R5_data (_registers_3_ext_R5_data),
    .R6_data (_registers_3_ext_R6_data),
    .R7_data (_registers_3_ext_R7_data)
  );
  registers_8x64 registers_4_ext (
    .R0_addr (io_read_7_address[2:0]),
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .R1_addr (io_read_6_address[2:0]),
    .R1_en   (1'h1),
    .R1_clk  (clock),
    .R2_addr (io_read_5_address[2:0]),
    .R2_en   (1'h1),
    .R2_clk  (clock),
    .R3_addr (io_read_4_address[2:0]),
    .R3_en   (1'h1),
    .R3_clk  (clock),
    .R4_addr (io_read_3_address[2:0]),
    .R4_en   (1'h1),
    .R4_clk  (clock),
    .R5_addr (io_read_2_address[2:0]),
    .R5_en   (1'h1),
    .R5_clk  (clock),
    .R6_addr (io_read_1_address[2:0]),
    .R6_en   (1'h1),
    .R6_clk  (clock),
    .R7_addr (io_read_0_address[2:0]),
    .R7_en   (1'h1),
    .R7_clk  (clock),
    .W0_addr (io_write_0_address[2:0]),
    .W0_en   (io_write_0_write & _GEN_3 == 7'h4),
    .W0_clk  (clock),
    .W0_data (io_write_0_value),
    .W0_mask (_GEN),
    .W1_addr (io_write_2_address[2:0]),
    .W1_en   (io_write_2_write & _GEN_5 == 7'h4),
    .W1_clk  (clock),
    .W1_data (io_write_2_value),
    .W1_mask (_GEN_1),
    .W2_addr (io_write_1_address[2:0]),
    .W2_en   (io_write_1_write & _GEN_4 == 7'h4),
    .W2_clk  (clock),
    .W2_data (io_write_1_value),
    .W2_mask (_GEN_0),
    .W3_addr (io_write_3_address[2:0]),
    .W3_en   (io_write_3_write & _GEN_6 == 7'h4),
    .W3_clk  (clock),
    .W3_data (io_write_3_value),
    .W3_mask (_GEN_2),
    .R0_data (_registers_4_ext_R0_data),
    .R1_data (_registers_4_ext_R1_data),
    .R2_data (_registers_4_ext_R2_data),
    .R3_data (_registers_4_ext_R3_data),
    .R4_data (_registers_4_ext_R4_data),
    .R5_data (_registers_4_ext_R5_data),
    .R6_data (_registers_4_ext_R6_data),
    .R7_data (_registers_4_ext_R7_data)
  );
  registers_8x64 registers_5_ext (
    .R0_addr (io_read_7_address[2:0]),
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .R1_addr (io_read_6_address[2:0]),
    .R1_en   (1'h1),
    .R1_clk  (clock),
    .R2_addr (io_read_5_address[2:0]),
    .R2_en   (1'h1),
    .R2_clk  (clock),
    .R3_addr (io_read_4_address[2:0]),
    .R3_en   (1'h1),
    .R3_clk  (clock),
    .R4_addr (io_read_3_address[2:0]),
    .R4_en   (1'h1),
    .R4_clk  (clock),
    .R5_addr (io_read_2_address[2:0]),
    .R5_en   (1'h1),
    .R5_clk  (clock),
    .R6_addr (io_read_1_address[2:0]),
    .R6_en   (1'h1),
    .R6_clk  (clock),
    .R7_addr (io_read_0_address[2:0]),
    .R7_en   (1'h1),
    .R7_clk  (clock),
    .W0_addr (io_write_2_address[2:0]),
    .W0_en   (io_write_2_write & _GEN_5 == 7'h5),
    .W0_clk  (clock),
    .W0_data (io_write_2_value),
    .W0_mask (_GEN_1),
    .W1_addr (io_write_1_address[2:0]),
    .W1_en   (io_write_1_write & _GEN_4 == 7'h5),
    .W1_clk  (clock),
    .W1_data (io_write_1_value),
    .W1_mask (_GEN_0),
    .W2_addr (io_write_0_address[2:0]),
    .W2_en   (io_write_0_write & _GEN_3 == 7'h5),
    .W2_clk  (clock),
    .W2_data (io_write_0_value),
    .W2_mask (_GEN),
    .W3_addr (io_write_3_address[2:0]),
    .W3_en   (io_write_3_write & _GEN_6 == 7'h5),
    .W3_clk  (clock),
    .W3_data (io_write_3_value),
    .W3_mask (_GEN_2),
    .R0_data (_registers_5_ext_R0_data),
    .R1_data (_registers_5_ext_R1_data),
    .R2_data (_registers_5_ext_R2_data),
    .R3_data (_registers_5_ext_R3_data),
    .R4_data (_registers_5_ext_R4_data),
    .R5_data (_registers_5_ext_R5_data),
    .R6_data (_registers_5_ext_R6_data),
    .R7_data (_registers_5_ext_R7_data)
  );
  registers_8x64 registers_6_ext (
    .R0_addr (io_read_7_address[2:0]),
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .R1_addr (io_read_6_address[2:0]),
    .R1_en   (1'h1),
    .R1_clk  (clock),
    .R2_addr (io_read_5_address[2:0]),
    .R2_en   (1'h1),
    .R2_clk  (clock),
    .R3_addr (io_read_4_address[2:0]),
    .R3_en   (1'h1),
    .R3_clk  (clock),
    .R4_addr (io_read_3_address[2:0]),
    .R4_en   (1'h1),
    .R4_clk  (clock),
    .R5_addr (io_read_2_address[2:0]),
    .R5_en   (1'h1),
    .R5_clk  (clock),
    .R6_addr (io_read_1_address[2:0]),
    .R6_en   (1'h1),
    .R6_clk  (clock),
    .R7_addr (io_read_0_address[2:0]),
    .R7_en   (1'h1),
    .R7_clk  (clock),
    .W0_addr (io_write_2_address[2:0]),
    .W0_en   (io_write_2_write & _GEN_5 == 7'h6),
    .W0_clk  (clock),
    .W0_data (io_write_2_value),
    .W0_mask (_GEN_1),
    .W1_addr (io_write_1_address[2:0]),
    .W1_en   (io_write_1_write & _GEN_4 == 7'h6),
    .W1_clk  (clock),
    .W1_data (io_write_1_value),
    .W1_mask (_GEN_0),
    .W2_addr (io_write_0_address[2:0]),
    .W2_en   (io_write_0_write & _GEN_3 == 7'h6),
    .W2_clk  (clock),
    .W2_data (io_write_0_value),
    .W2_mask (_GEN),
    .W3_addr (io_write_3_address[2:0]),
    .W3_en   (io_write_3_write & _GEN_6 == 7'h6),
    .W3_clk  (clock),
    .W3_data (io_write_3_value),
    .W3_mask (_GEN_2),
    .R0_data (_registers_6_ext_R0_data),
    .R1_data (_registers_6_ext_R1_data),
    .R2_data (_registers_6_ext_R2_data),
    .R3_data (_registers_6_ext_R3_data),
    .R4_data (_registers_6_ext_R4_data),
    .R5_data (_registers_6_ext_R5_data),
    .R6_data (_registers_6_ext_R6_data),
    .R7_data (_registers_6_ext_R7_data)
  );
  registers_8x64 registers_7_ext (
    .R0_addr (io_read_7_address[2:0]),
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .R1_addr (io_read_6_address[2:0]),
    .R1_en   (1'h1),
    .R1_clk  (clock),
    .R2_addr (io_read_5_address[2:0]),
    .R2_en   (1'h1),
    .R2_clk  (clock),
    .R3_addr (io_read_4_address[2:0]),
    .R3_en   (1'h1),
    .R3_clk  (clock),
    .R4_addr (io_read_3_address[2:0]),
    .R4_en   (1'h1),
    .R4_clk  (clock),
    .R5_addr (io_read_2_address[2:0]),
    .R5_en   (1'h1),
    .R5_clk  (clock),
    .R6_addr (io_read_1_address[2:0]),
    .R6_en   (1'h1),
    .R6_clk  (clock),
    .R7_addr (io_read_0_address[2:0]),
    .R7_en   (1'h1),
    .R7_clk  (clock),
    .W0_addr (io_write_2_address[2:0]),
    .W0_en   (io_write_2_write & _GEN_5 == 7'h7),
    .W0_clk  (clock),
    .W0_data (io_write_2_value),
    .W0_mask (_GEN_1),
    .W1_addr (io_write_1_address[2:0]),
    .W1_en   (io_write_1_write & _GEN_4 == 7'h7),
    .W1_clk  (clock),
    .W1_data (io_write_1_value),
    .W1_mask (_GEN_0),
    .W2_addr (io_write_0_address[2:0]),
    .W2_en   (io_write_0_write & _GEN_3 == 7'h7),
    .W2_clk  (clock),
    .W2_data (io_write_0_value),
    .W2_mask (_GEN),
    .W3_addr (io_write_3_address[2:0]),
    .W3_en   (io_write_3_write & _GEN_6 == 7'h7),
    .W3_clk  (clock),
    .W3_data (io_write_3_value),
    .W3_mask (_GEN_2),
    .R0_data (_registers_7_ext_R0_data),
    .R1_data (_registers_7_ext_R1_data),
    .R2_data (_registers_7_ext_R2_data),
    .R3_data (_registers_7_ext_R3_data),
    .R4_data (_registers_7_ext_R4_data),
    .R5_data (_registers_7_ext_R5_data),
    .R6_data (_registers_7_ext_R6_data),
    .R7_data (_registers_7_ext_R7_data)
  );
  registers_8x64 registers_8_ext (
    .R0_addr (io_read_7_address[2:0]),
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .R1_addr (io_read_6_address[2:0]),
    .R1_en   (1'h1),
    .R1_clk  (clock),
    .R2_addr (io_read_5_address[2:0]),
    .R2_en   (1'h1),
    .R2_clk  (clock),
    .R3_addr (io_read_4_address[2:0]),
    .R3_en   (1'h1),
    .R3_clk  (clock),
    .R4_addr (io_read_3_address[2:0]),
    .R4_en   (1'h1),
    .R4_clk  (clock),
    .R5_addr (io_read_2_address[2:0]),
    .R5_en   (1'h1),
    .R5_clk  (clock),
    .R6_addr (io_read_1_address[2:0]),
    .R6_en   (1'h1),
    .R6_clk  (clock),
    .R7_addr (io_read_0_address[2:0]),
    .R7_en   (1'h1),
    .R7_clk  (clock),
    .W0_addr (io_write_2_address[2:0]),
    .W0_en   (io_write_2_write & _GEN_5 == 7'h8),
    .W0_clk  (clock),
    .W0_data (io_write_2_value),
    .W0_mask (_GEN_1),
    .W1_addr (io_write_1_address[2:0]),
    .W1_en   (io_write_1_write & _GEN_4 == 7'h8),
    .W1_clk  (clock),
    .W1_data (io_write_1_value),
    .W1_mask (_GEN_0),
    .W2_addr (io_write_0_address[2:0]),
    .W2_en   (io_write_0_write & _GEN_3 == 7'h8),
    .W2_clk  (clock),
    .W2_data (io_write_0_value),
    .W2_mask (_GEN),
    .W3_addr (io_write_3_address[2:0]),
    .W3_en   (io_write_3_write & _GEN_6 == 7'h8),
    .W3_clk  (clock),
    .W3_data (io_write_3_value),
    .W3_mask (_GEN_2),
    .R0_data (_registers_8_ext_R0_data),
    .R1_data (_registers_8_ext_R1_data),
    .R2_data (_registers_8_ext_R2_data),
    .R3_data (_registers_8_ext_R3_data),
    .R4_data (_registers_8_ext_R4_data),
    .R5_data (_registers_8_ext_R5_data),
    .R6_data (_registers_8_ext_R6_data),
    .R7_data (_registers_8_ext_R7_data)
  );
  registers_8x64 registers_9_ext (
    .R0_addr (io_read_7_address[2:0]),
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .R1_addr (io_read_6_address[2:0]),
    .R1_en   (1'h1),
    .R1_clk  (clock),
    .R2_addr (io_read_5_address[2:0]),
    .R2_en   (1'h1),
    .R2_clk  (clock),
    .R3_addr (io_read_4_address[2:0]),
    .R3_en   (1'h1),
    .R3_clk  (clock),
    .R4_addr (io_read_3_address[2:0]),
    .R4_en   (1'h1),
    .R4_clk  (clock),
    .R5_addr (io_read_2_address[2:0]),
    .R5_en   (1'h1),
    .R5_clk  (clock),
    .R6_addr (io_read_1_address[2:0]),
    .R6_en   (1'h1),
    .R6_clk  (clock),
    .R7_addr (io_read_0_address[2:0]),
    .R7_en   (1'h1),
    .R7_clk  (clock),
    .W0_addr (io_write_2_address[2:0]),
    .W0_en   (io_write_2_write & _GEN_5 == 7'h9),
    .W0_clk  (clock),
    .W0_data (io_write_2_value),
    .W0_mask (_GEN_1),
    .W1_addr (io_write_1_address[2:0]),
    .W1_en   (io_write_1_write & _GEN_4 == 7'h9),
    .W1_clk  (clock),
    .W1_data (io_write_1_value),
    .W1_mask (_GEN_0),
    .W2_addr (io_write_0_address[2:0]),
    .W2_en   (io_write_0_write & _GEN_3 == 7'h9),
    .W2_clk  (clock),
    .W2_data (io_write_0_value),
    .W2_mask (_GEN),
    .W3_addr (io_write_3_address[2:0]),
    .W3_en   (io_write_3_write & _GEN_6 == 7'h9),
    .W3_clk  (clock),
    .W3_data (io_write_3_value),
    .W3_mask (_GEN_2),
    .R0_data (_registers_9_ext_R0_data),
    .R1_data (_registers_9_ext_R1_data),
    .R2_data (_registers_9_ext_R2_data),
    .R3_data (_registers_9_ext_R3_data),
    .R4_data (_registers_9_ext_R4_data),
    .R5_data (_registers_9_ext_R5_data),
    .R6_data (_registers_9_ext_R6_data),
    .R7_data (_registers_9_ext_R7_data)
  );
  registers_8x64 registers_10_ext (
    .R0_addr (io_read_7_address[2:0]),
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .R1_addr (io_read_6_address[2:0]),
    .R1_en   (1'h1),
    .R1_clk  (clock),
    .R2_addr (io_read_5_address[2:0]),
    .R2_en   (1'h1),
    .R2_clk  (clock),
    .R3_addr (io_read_4_address[2:0]),
    .R3_en   (1'h1),
    .R3_clk  (clock),
    .R4_addr (io_read_3_address[2:0]),
    .R4_en   (1'h1),
    .R4_clk  (clock),
    .R5_addr (io_read_2_address[2:0]),
    .R5_en   (1'h1),
    .R5_clk  (clock),
    .R6_addr (io_read_1_address[2:0]),
    .R6_en   (1'h1),
    .R6_clk  (clock),
    .R7_addr (io_read_0_address[2:0]),
    .R7_en   (1'h1),
    .R7_clk  (clock),
    .W0_addr (io_write_2_address[2:0]),
    .W0_en   (io_write_2_write & _GEN_5 == 7'hA),
    .W0_clk  (clock),
    .W0_data (io_write_2_value),
    .W0_mask (_GEN_1),
    .W1_addr (io_write_1_address[2:0]),
    .W1_en   (io_write_1_write & _GEN_4 == 7'hA),
    .W1_clk  (clock),
    .W1_data (io_write_1_value),
    .W1_mask (_GEN_0),
    .W2_addr (io_write_0_address[2:0]),
    .W2_en   (io_write_0_write & _GEN_3 == 7'hA),
    .W2_clk  (clock),
    .W2_data (io_write_0_value),
    .W2_mask (_GEN),
    .W3_addr (io_write_3_address[2:0]),
    .W3_en   (io_write_3_write & _GEN_6 == 7'hA),
    .W3_clk  (clock),
    .W3_data (io_write_3_value),
    .W3_mask (_GEN_2),
    .R0_data (_registers_10_ext_R0_data),
    .R1_data (_registers_10_ext_R1_data),
    .R2_data (_registers_10_ext_R2_data),
    .R3_data (_registers_10_ext_R3_data),
    .R4_data (_registers_10_ext_R4_data),
    .R5_data (_registers_10_ext_R5_data),
    .R6_data (_registers_10_ext_R6_data),
    .R7_data (_registers_10_ext_R7_data)
  );
  registers_8x64 registers_11_ext (
    .R0_addr (io_read_7_address[2:0]),
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .R1_addr (io_read_6_address[2:0]),
    .R1_en   (1'h1),
    .R1_clk  (clock),
    .R2_addr (io_read_5_address[2:0]),
    .R2_en   (1'h1),
    .R2_clk  (clock),
    .R3_addr (io_read_4_address[2:0]),
    .R3_en   (1'h1),
    .R3_clk  (clock),
    .R4_addr (io_read_3_address[2:0]),
    .R4_en   (1'h1),
    .R4_clk  (clock),
    .R5_addr (io_read_2_address[2:0]),
    .R5_en   (1'h1),
    .R5_clk  (clock),
    .R6_addr (io_read_1_address[2:0]),
    .R6_en   (1'h1),
    .R6_clk  (clock),
    .R7_addr (io_read_0_address[2:0]),
    .R7_en   (1'h1),
    .R7_clk  (clock),
    .W0_addr (io_write_2_address[2:0]),
    .W0_en   (io_write_2_write & _GEN_5 == 7'hB),
    .W0_clk  (clock),
    .W0_data (io_write_2_value),
    .W0_mask (_GEN_1),
    .W1_addr (io_write_1_address[2:0]),
    .W1_en   (io_write_1_write & _GEN_4 == 7'hB),
    .W1_clk  (clock),
    .W1_data (io_write_1_value),
    .W1_mask (_GEN_0),
    .W2_addr (io_write_0_address[2:0]),
    .W2_en   (io_write_0_write & _GEN_3 == 7'hB),
    .W2_clk  (clock),
    .W2_data (io_write_0_value),
    .W2_mask (_GEN),
    .W3_addr (io_write_3_address[2:0]),
    .W3_en   (io_write_3_write & _GEN_6 == 7'hB),
    .W3_clk  (clock),
    .W3_data (io_write_3_value),
    .W3_mask (_GEN_2),
    .R0_data (_registers_11_ext_R0_data),
    .R1_data (_registers_11_ext_R1_data),
    .R2_data (_registers_11_ext_R2_data),
    .R3_data (_registers_11_ext_R3_data),
    .R4_data (_registers_11_ext_R4_data),
    .R5_data (_registers_11_ext_R5_data),
    .R6_data (_registers_11_ext_R6_data),
    .R7_data (_registers_11_ext_R7_data)
  );
  registers_8x64 registers_12_ext (
    .R0_addr (io_read_7_address[2:0]),
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .R1_addr (io_read_6_address[2:0]),
    .R1_en   (1'h1),
    .R1_clk  (clock),
    .R2_addr (io_read_5_address[2:0]),
    .R2_en   (1'h1),
    .R2_clk  (clock),
    .R3_addr (io_read_4_address[2:0]),
    .R3_en   (1'h1),
    .R3_clk  (clock),
    .R4_addr (io_read_3_address[2:0]),
    .R4_en   (1'h1),
    .R4_clk  (clock),
    .R5_addr (io_read_2_address[2:0]),
    .R5_en   (1'h1),
    .R5_clk  (clock),
    .R6_addr (io_read_1_address[2:0]),
    .R6_en   (1'h1),
    .R6_clk  (clock),
    .R7_addr (io_read_0_address[2:0]),
    .R7_en   (1'h1),
    .R7_clk  (clock),
    .W0_addr (io_write_2_address[2:0]),
    .W0_en   (io_write_2_write & _GEN_5 == 7'hC),
    .W0_clk  (clock),
    .W0_data (io_write_2_value),
    .W0_mask (_GEN_1),
    .W1_addr (io_write_1_address[2:0]),
    .W1_en   (io_write_1_write & _GEN_4 == 7'hC),
    .W1_clk  (clock),
    .W1_data (io_write_1_value),
    .W1_mask (_GEN_0),
    .W2_addr (io_write_0_address[2:0]),
    .W2_en   (io_write_0_write & _GEN_3 == 7'hC),
    .W2_clk  (clock),
    .W2_data (io_write_0_value),
    .W2_mask (_GEN),
    .W3_addr (io_write_3_address[2:0]),
    .W3_en   (io_write_3_write & _GEN_6 == 7'hC),
    .W3_clk  (clock),
    .W3_data (io_write_3_value),
    .W3_mask (_GEN_2),
    .R0_data (_registers_12_ext_R0_data),
    .R1_data (_registers_12_ext_R1_data),
    .R2_data (_registers_12_ext_R2_data),
    .R3_data (_registers_12_ext_R3_data),
    .R4_data (_registers_12_ext_R4_data),
    .R5_data (_registers_12_ext_R5_data),
    .R6_data (_registers_12_ext_R6_data),
    .R7_data (_registers_12_ext_R7_data)
  );
  registers_8x64 registers_13_ext (
    .R0_addr (io_read_7_address[2:0]),
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .R1_addr (io_read_6_address[2:0]),
    .R1_en   (1'h1),
    .R1_clk  (clock),
    .R2_addr (io_read_5_address[2:0]),
    .R2_en   (1'h1),
    .R2_clk  (clock),
    .R3_addr (io_read_4_address[2:0]),
    .R3_en   (1'h1),
    .R3_clk  (clock),
    .R4_addr (io_read_3_address[2:0]),
    .R4_en   (1'h1),
    .R4_clk  (clock),
    .R5_addr (io_read_2_address[2:0]),
    .R5_en   (1'h1),
    .R5_clk  (clock),
    .R6_addr (io_read_1_address[2:0]),
    .R6_en   (1'h1),
    .R6_clk  (clock),
    .R7_addr (io_read_0_address[2:0]),
    .R7_en   (1'h1),
    .R7_clk  (clock),
    .W0_addr (io_write_2_address[2:0]),
    .W0_en   (io_write_2_write & _GEN_5 == 7'hD),
    .W0_clk  (clock),
    .W0_data (io_write_2_value),
    .W0_mask (_GEN_1),
    .W1_addr (io_write_1_address[2:0]),
    .W1_en   (io_write_1_write & _GEN_4 == 7'hD),
    .W1_clk  (clock),
    .W1_data (io_write_1_value),
    .W1_mask (_GEN_0),
    .W2_addr (io_write_0_address[2:0]),
    .W2_en   (io_write_0_write & _GEN_3 == 7'hD),
    .W2_clk  (clock),
    .W2_data (io_write_0_value),
    .W2_mask (_GEN),
    .W3_addr (io_write_3_address[2:0]),
    .W3_en   (io_write_3_write & _GEN_6 == 7'hD),
    .W3_clk  (clock),
    .W3_data (io_write_3_value),
    .W3_mask (_GEN_2),
    .R0_data (_registers_13_ext_R0_data),
    .R1_data (_registers_13_ext_R1_data),
    .R2_data (_registers_13_ext_R2_data),
    .R3_data (_registers_13_ext_R3_data),
    .R4_data (_registers_13_ext_R4_data),
    .R5_data (_registers_13_ext_R5_data),
    .R6_data (_registers_13_ext_R6_data),
    .R7_data (_registers_13_ext_R7_data)
  );
  registers_8x64 registers_14_ext (
    .R0_addr (io_read_7_address[2:0]),
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .R1_addr (io_read_6_address[2:0]),
    .R1_en   (1'h1),
    .R1_clk  (clock),
    .R2_addr (io_read_5_address[2:0]),
    .R2_en   (1'h1),
    .R2_clk  (clock),
    .R3_addr (io_read_4_address[2:0]),
    .R3_en   (1'h1),
    .R3_clk  (clock),
    .R4_addr (io_read_3_address[2:0]),
    .R4_en   (1'h1),
    .R4_clk  (clock),
    .R5_addr (io_read_2_address[2:0]),
    .R5_en   (1'h1),
    .R5_clk  (clock),
    .R6_addr (io_read_1_address[2:0]),
    .R6_en   (1'h1),
    .R6_clk  (clock),
    .R7_addr (io_read_0_address[2:0]),
    .R7_en   (1'h1),
    .R7_clk  (clock),
    .W0_addr (io_write_2_address[2:0]),
    .W0_en   (io_write_2_write & _GEN_5 == 7'hE),
    .W0_clk  (clock),
    .W0_data (io_write_2_value),
    .W0_mask (_GEN_1),
    .W1_addr (io_write_1_address[2:0]),
    .W1_en   (io_write_1_write & _GEN_4 == 7'hE),
    .W1_clk  (clock),
    .W1_data (io_write_1_value),
    .W1_mask (_GEN_0),
    .W2_addr (io_write_0_address[2:0]),
    .W2_en   (io_write_0_write & _GEN_3 == 7'hE),
    .W2_clk  (clock),
    .W2_data (io_write_0_value),
    .W2_mask (_GEN),
    .W3_addr (io_write_3_address[2:0]),
    .W3_en   (io_write_3_write & _GEN_6 == 7'hE),
    .W3_clk  (clock),
    .W3_data (io_write_3_value),
    .W3_mask (_GEN_2),
    .R0_data (_registers_14_ext_R0_data),
    .R1_data (_registers_14_ext_R1_data),
    .R2_data (_registers_14_ext_R2_data),
    .R3_data (_registers_14_ext_R3_data),
    .R4_data (_registers_14_ext_R4_data),
    .R5_data (_registers_14_ext_R5_data),
    .R6_data (_registers_14_ext_R6_data),
    .R7_data (_registers_14_ext_R7_data)
  );
  registers_8x64 registers_15_ext (
    .R0_addr (io_read_7_address[2:0]),
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .R1_addr (io_read_6_address[2:0]),
    .R1_en   (1'h1),
    .R1_clk  (clock),
    .R2_addr (io_read_5_address[2:0]),
    .R2_en   (1'h1),
    .R2_clk  (clock),
    .R3_addr (io_read_4_address[2:0]),
    .R3_en   (1'h1),
    .R3_clk  (clock),
    .R4_addr (io_read_3_address[2:0]),
    .R4_en   (1'h1),
    .R4_clk  (clock),
    .R5_addr (io_read_2_address[2:0]),
    .R5_en   (1'h1),
    .R5_clk  (clock),
    .R6_addr (io_read_1_address[2:0]),
    .R6_en   (1'h1),
    .R6_clk  (clock),
    .R7_addr (io_read_0_address[2:0]),
    .R7_en   (1'h1),
    .R7_clk  (clock),
    .W0_addr (io_write_2_address[2:0]),
    .W0_en   (io_write_2_write & _GEN_5 == 7'hF),
    .W0_clk  (clock),
    .W0_data (io_write_2_value),
    .W0_mask (_GEN_1),
    .W1_addr (io_write_1_address[2:0]),
    .W1_en   (io_write_1_write & _GEN_4 == 7'hF),
    .W1_clk  (clock),
    .W1_data (io_write_1_value),
    .W1_mask (_GEN_0),
    .W2_addr (io_write_0_address[2:0]),
    .W2_en   (io_write_0_write & _GEN_3 == 7'hF),
    .W2_clk  (clock),
    .W2_data (io_write_0_value),
    .W2_mask (_GEN),
    .W3_addr (io_write_3_address[2:0]),
    .W3_en   (io_write_3_write & _GEN_6 == 7'hF),
    .W3_clk  (clock),
    .W3_data (io_write_3_value),
    .W3_mask (_GEN_2),
    .R0_data (_registers_15_ext_R0_data),
    .R1_data (_registers_15_ext_R1_data),
    .R2_data (_registers_15_ext_R2_data),
    .R3_data (_registers_15_ext_R3_data),
    .R4_data (_registers_15_ext_R4_data),
    .R5_data (_registers_15_ext_R5_data),
    .R6_data (_registers_15_ext_R6_data),
    .R7_data (_registers_15_ext_R7_data)
  );
  assign io_read_0_value =
    {casez_tmp_6,
     casez_tmp_5,
     casez_tmp_4,
     casez_tmp_3,
     casez_tmp_2,
     casez_tmp_1,
     casez_tmp_0,
     casez_tmp};
  assign io_read_1_value =
    {casez_tmp_14,
     casez_tmp_13,
     casez_tmp_12,
     casez_tmp_11,
     casez_tmp_10,
     casez_tmp_9,
     casez_tmp_8,
     casez_tmp_7};
  assign io_read_2_value =
    {casez_tmp_22,
     casez_tmp_21,
     casez_tmp_20,
     casez_tmp_19,
     casez_tmp_18,
     casez_tmp_17,
     casez_tmp_16,
     casez_tmp_15};
  assign io_read_3_value =
    {casez_tmp_30,
     casez_tmp_29,
     casez_tmp_28,
     casez_tmp_27,
     casez_tmp_26,
     casez_tmp_25,
     casez_tmp_24,
     casez_tmp_23};
  assign io_read_4_value =
    {casez_tmp_38,
     casez_tmp_37,
     casez_tmp_36,
     casez_tmp_35,
     casez_tmp_34,
     casez_tmp_33,
     casez_tmp_32,
     casez_tmp_31};
  assign io_read_5_value =
    {casez_tmp_46,
     casez_tmp_45,
     casez_tmp_44,
     casez_tmp_43,
     casez_tmp_42,
     casez_tmp_41,
     casez_tmp_40,
     casez_tmp_39};
  assign io_read_6_value =
    {casez_tmp_54,
     casez_tmp_53,
     casez_tmp_52,
     casez_tmp_51,
     casez_tmp_50,
     casez_tmp_49,
     casez_tmp_48,
     casez_tmp_47};
  assign io_read_7_value =
    {casez_tmp_62,
     casez_tmp_61,
     casez_tmp_60,
     casez_tmp_59,
     casez_tmp_58,
     casez_tmp_57,
     casez_tmp_56,
     casez_tmp_55};
endmodule

