VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_2048x39
  FOREIGN fakeram45_2048x39 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 206.910 BY 219.800 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.400 0.070 1.470 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.940 0.070 3.010 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.480 0.070 4.550 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.020 0.070 6.090 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.560 0.070 7.630 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.100 0.070 9.170 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.640 0.070 10.710 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.180 0.070 12.250 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.720 0.070 13.790 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.260 0.070 15.330 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.800 0.070 16.870 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.340 0.070 18.410 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.880 0.070 19.950 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.420 0.070 21.490 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.960 0.070 23.030 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.500 0.070 24.570 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.040 0.070 26.110 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.580 0.070 27.650 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.120 0.070 29.190 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.660 0.070 30.730 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.200 0.070 32.270 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.740 0.070 33.810 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.280 0.070 35.350 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.820 0.070 36.890 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.360 0.070 38.430 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.900 0.070 39.970 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.440 0.070 41.510 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.980 0.070 43.050 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.520 0.070 44.590 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.060 0.070 46.130 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.600 0.070 47.670 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.140 0.070 49.210 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.680 0.070 50.750 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.220 0.070 52.290 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.760 0.070 53.830 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.300 0.070 55.370 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.840 0.070 56.910 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.380 0.070 58.450 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.920 0.070 59.990 ;
    END
  END w_mask_in[38]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.700 0.070 63.770 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.240 0.070 65.310 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.780 0.070 66.850 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.320 0.070 68.390 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.860 0.070 69.930 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.400 0.070 71.470 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.940 0.070 73.010 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.480 0.070 74.550 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.020 0.070 76.090 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.560 0.070 77.630 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.100 0.070 79.170 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.640 0.070 80.710 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.180 0.070 82.250 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.720 0.070 83.790 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.260 0.070 85.330 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.800 0.070 86.870 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.340 0.070 88.410 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.880 0.070 89.950 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.420 0.070 91.490 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.960 0.070 93.030 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.500 0.070 94.570 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.040 0.070 96.110 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.580 0.070 97.650 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.120 0.070 99.190 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.660 0.070 100.730 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.200 0.070 102.270 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.740 0.070 103.810 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.280 0.070 105.350 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.820 0.070 106.890 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.360 0.070 108.430 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.900 0.070 109.970 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.440 0.070 111.510 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.980 0.070 113.050 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.520 0.070 114.590 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.060 0.070 116.130 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.600 0.070 117.670 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.140 0.070 119.210 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.680 0.070 120.750 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.220 0.070 122.290 ;
    END
  END rd_out[38]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.000 0.070 126.070 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.540 0.070 127.610 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.080 0.070 129.150 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 130.620 0.070 130.690 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.160 0.070 132.230 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 133.700 0.070 133.770 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 135.240 0.070 135.310 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.780 0.070 136.850 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.320 0.070 138.390 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.860 0.070 139.930 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 141.400 0.070 141.470 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.940 0.070 143.010 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.480 0.070 144.550 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.020 0.070 146.090 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.560 0.070 147.630 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 149.100 0.070 149.170 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.640 0.070 150.710 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.180 0.070 152.250 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.720 0.070 153.790 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.260 0.070 155.330 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.800 0.070 156.870 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.340 0.070 158.410 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.880 0.070 159.950 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.420 0.070 161.490 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.960 0.070 163.030 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.500 0.070 164.570 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.040 0.070 166.110 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.580 0.070 167.650 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.120 0.070 169.190 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.660 0.070 170.730 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.200 0.070 172.270 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.740 0.070 173.810 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.280 0.070 175.350 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.820 0.070 176.890 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.360 0.070 178.430 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.900 0.070 179.970 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.440 0.070 181.510 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 182.980 0.070 183.050 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.520 0.070 184.590 ;
    END
  END wd_in[38]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.300 0.070 188.370 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.840 0.070 189.910 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.380 0.070 191.450 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.920 0.070 192.990 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.460 0.070 194.530 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.000 0.070 196.070 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.540 0.070 197.610 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 199.080 0.070 199.150 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 200.620 0.070 200.690 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 202.160 0.070 202.230 ;
    END
  END addr_in[9]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 203.700 0.070 203.770 ;
    END
  END addr_in[10]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 207.480 0.070 207.550 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.020 0.070 209.090 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 210.560 0.070 210.630 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 218.400 ;
      RECT 3.500 1.400 3.780 218.400 ;
      RECT 5.740 1.400 6.020 218.400 ;
      RECT 7.980 1.400 8.260 218.400 ;
      RECT 10.220 1.400 10.500 218.400 ;
      RECT 12.460 1.400 12.740 218.400 ;
      RECT 14.700 1.400 14.980 218.400 ;
      RECT 16.940 1.400 17.220 218.400 ;
      RECT 19.180 1.400 19.460 218.400 ;
      RECT 21.420 1.400 21.700 218.400 ;
      RECT 23.660 1.400 23.940 218.400 ;
      RECT 25.900 1.400 26.180 218.400 ;
      RECT 28.140 1.400 28.420 218.400 ;
      RECT 30.380 1.400 30.660 218.400 ;
      RECT 32.620 1.400 32.900 218.400 ;
      RECT 34.860 1.400 35.140 218.400 ;
      RECT 37.100 1.400 37.380 218.400 ;
      RECT 39.340 1.400 39.620 218.400 ;
      RECT 41.580 1.400 41.860 218.400 ;
      RECT 43.820 1.400 44.100 218.400 ;
      RECT 46.060 1.400 46.340 218.400 ;
      RECT 48.300 1.400 48.580 218.400 ;
      RECT 50.540 1.400 50.820 218.400 ;
      RECT 52.780 1.400 53.060 218.400 ;
      RECT 55.020 1.400 55.300 218.400 ;
      RECT 57.260 1.400 57.540 218.400 ;
      RECT 59.500 1.400 59.780 218.400 ;
      RECT 61.740 1.400 62.020 218.400 ;
      RECT 63.980 1.400 64.260 218.400 ;
      RECT 66.220 1.400 66.500 218.400 ;
      RECT 68.460 1.400 68.740 218.400 ;
      RECT 70.700 1.400 70.980 218.400 ;
      RECT 72.940 1.400 73.220 218.400 ;
      RECT 75.180 1.400 75.460 218.400 ;
      RECT 77.420 1.400 77.700 218.400 ;
      RECT 79.660 1.400 79.940 218.400 ;
      RECT 81.900 1.400 82.180 218.400 ;
      RECT 84.140 1.400 84.420 218.400 ;
      RECT 86.380 1.400 86.660 218.400 ;
      RECT 88.620 1.400 88.900 218.400 ;
      RECT 90.860 1.400 91.140 218.400 ;
      RECT 93.100 1.400 93.380 218.400 ;
      RECT 95.340 1.400 95.620 218.400 ;
      RECT 97.580 1.400 97.860 218.400 ;
      RECT 99.820 1.400 100.100 218.400 ;
      RECT 102.060 1.400 102.340 218.400 ;
      RECT 104.300 1.400 104.580 218.400 ;
      RECT 106.540 1.400 106.820 218.400 ;
      RECT 108.780 1.400 109.060 218.400 ;
      RECT 111.020 1.400 111.300 218.400 ;
      RECT 113.260 1.400 113.540 218.400 ;
      RECT 115.500 1.400 115.780 218.400 ;
      RECT 117.740 1.400 118.020 218.400 ;
      RECT 119.980 1.400 120.260 218.400 ;
      RECT 122.220 1.400 122.500 218.400 ;
      RECT 124.460 1.400 124.740 218.400 ;
      RECT 126.700 1.400 126.980 218.400 ;
      RECT 128.940 1.400 129.220 218.400 ;
      RECT 131.180 1.400 131.460 218.400 ;
      RECT 133.420 1.400 133.700 218.400 ;
      RECT 135.660 1.400 135.940 218.400 ;
      RECT 137.900 1.400 138.180 218.400 ;
      RECT 140.140 1.400 140.420 218.400 ;
      RECT 142.380 1.400 142.660 218.400 ;
      RECT 144.620 1.400 144.900 218.400 ;
      RECT 146.860 1.400 147.140 218.400 ;
      RECT 149.100 1.400 149.380 218.400 ;
      RECT 151.340 1.400 151.620 218.400 ;
      RECT 153.580 1.400 153.860 218.400 ;
      RECT 155.820 1.400 156.100 218.400 ;
      RECT 158.060 1.400 158.340 218.400 ;
      RECT 160.300 1.400 160.580 218.400 ;
      RECT 162.540 1.400 162.820 218.400 ;
      RECT 164.780 1.400 165.060 218.400 ;
      RECT 167.020 1.400 167.300 218.400 ;
      RECT 169.260 1.400 169.540 218.400 ;
      RECT 171.500 1.400 171.780 218.400 ;
      RECT 173.740 1.400 174.020 218.400 ;
      RECT 175.980 1.400 176.260 218.400 ;
      RECT 178.220 1.400 178.500 218.400 ;
      RECT 180.460 1.400 180.740 218.400 ;
      RECT 182.700 1.400 182.980 218.400 ;
      RECT 184.940 1.400 185.220 218.400 ;
      RECT 187.180 1.400 187.460 218.400 ;
      RECT 189.420 1.400 189.700 218.400 ;
      RECT 191.660 1.400 191.940 218.400 ;
      RECT 193.900 1.400 194.180 218.400 ;
      RECT 196.140 1.400 196.420 218.400 ;
      RECT 198.380 1.400 198.660 218.400 ;
      RECT 200.620 1.400 200.900 218.400 ;
      RECT 202.860 1.400 203.140 218.400 ;
      RECT 205.100 1.400 205.380 218.400 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 218.400 ;
      RECT 4.620 1.400 4.900 218.400 ;
      RECT 6.860 1.400 7.140 218.400 ;
      RECT 9.100 1.400 9.380 218.400 ;
      RECT 11.340 1.400 11.620 218.400 ;
      RECT 13.580 1.400 13.860 218.400 ;
      RECT 15.820 1.400 16.100 218.400 ;
      RECT 18.060 1.400 18.340 218.400 ;
      RECT 20.300 1.400 20.580 218.400 ;
      RECT 22.540 1.400 22.820 218.400 ;
      RECT 24.780 1.400 25.060 218.400 ;
      RECT 27.020 1.400 27.300 218.400 ;
      RECT 29.260 1.400 29.540 218.400 ;
      RECT 31.500 1.400 31.780 218.400 ;
      RECT 33.740 1.400 34.020 218.400 ;
      RECT 35.980 1.400 36.260 218.400 ;
      RECT 38.220 1.400 38.500 218.400 ;
      RECT 40.460 1.400 40.740 218.400 ;
      RECT 42.700 1.400 42.980 218.400 ;
      RECT 44.940 1.400 45.220 218.400 ;
      RECT 47.180 1.400 47.460 218.400 ;
      RECT 49.420 1.400 49.700 218.400 ;
      RECT 51.660 1.400 51.940 218.400 ;
      RECT 53.900 1.400 54.180 218.400 ;
      RECT 56.140 1.400 56.420 218.400 ;
      RECT 58.380 1.400 58.660 218.400 ;
      RECT 60.620 1.400 60.900 218.400 ;
      RECT 62.860 1.400 63.140 218.400 ;
      RECT 65.100 1.400 65.380 218.400 ;
      RECT 67.340 1.400 67.620 218.400 ;
      RECT 69.580 1.400 69.860 218.400 ;
      RECT 71.820 1.400 72.100 218.400 ;
      RECT 74.060 1.400 74.340 218.400 ;
      RECT 76.300 1.400 76.580 218.400 ;
      RECT 78.540 1.400 78.820 218.400 ;
      RECT 80.780 1.400 81.060 218.400 ;
      RECT 83.020 1.400 83.300 218.400 ;
      RECT 85.260 1.400 85.540 218.400 ;
      RECT 87.500 1.400 87.780 218.400 ;
      RECT 89.740 1.400 90.020 218.400 ;
      RECT 91.980 1.400 92.260 218.400 ;
      RECT 94.220 1.400 94.500 218.400 ;
      RECT 96.460 1.400 96.740 218.400 ;
      RECT 98.700 1.400 98.980 218.400 ;
      RECT 100.940 1.400 101.220 218.400 ;
      RECT 103.180 1.400 103.460 218.400 ;
      RECT 105.420 1.400 105.700 218.400 ;
      RECT 107.660 1.400 107.940 218.400 ;
      RECT 109.900 1.400 110.180 218.400 ;
      RECT 112.140 1.400 112.420 218.400 ;
      RECT 114.380 1.400 114.660 218.400 ;
      RECT 116.620 1.400 116.900 218.400 ;
      RECT 118.860 1.400 119.140 218.400 ;
      RECT 121.100 1.400 121.380 218.400 ;
      RECT 123.340 1.400 123.620 218.400 ;
      RECT 125.580 1.400 125.860 218.400 ;
      RECT 127.820 1.400 128.100 218.400 ;
      RECT 130.060 1.400 130.340 218.400 ;
      RECT 132.300 1.400 132.580 218.400 ;
      RECT 134.540 1.400 134.820 218.400 ;
      RECT 136.780 1.400 137.060 218.400 ;
      RECT 139.020 1.400 139.300 218.400 ;
      RECT 141.260 1.400 141.540 218.400 ;
      RECT 143.500 1.400 143.780 218.400 ;
      RECT 145.740 1.400 146.020 218.400 ;
      RECT 147.980 1.400 148.260 218.400 ;
      RECT 150.220 1.400 150.500 218.400 ;
      RECT 152.460 1.400 152.740 218.400 ;
      RECT 154.700 1.400 154.980 218.400 ;
      RECT 156.940 1.400 157.220 218.400 ;
      RECT 159.180 1.400 159.460 218.400 ;
      RECT 161.420 1.400 161.700 218.400 ;
      RECT 163.660 1.400 163.940 218.400 ;
      RECT 165.900 1.400 166.180 218.400 ;
      RECT 168.140 1.400 168.420 218.400 ;
      RECT 170.380 1.400 170.660 218.400 ;
      RECT 172.620 1.400 172.900 218.400 ;
      RECT 174.860 1.400 175.140 218.400 ;
      RECT 177.100 1.400 177.380 218.400 ;
      RECT 179.340 1.400 179.620 218.400 ;
      RECT 181.580 1.400 181.860 218.400 ;
      RECT 183.820 1.400 184.100 218.400 ;
      RECT 186.060 1.400 186.340 218.400 ;
      RECT 188.300 1.400 188.580 218.400 ;
      RECT 190.540 1.400 190.820 218.400 ;
      RECT 192.780 1.400 193.060 218.400 ;
      RECT 195.020 1.400 195.300 218.400 ;
      RECT 197.260 1.400 197.540 218.400 ;
      RECT 199.500 1.400 199.780 218.400 ;
      RECT 201.740 1.400 202.020 218.400 ;
      RECT 203.980 1.400 204.260 218.400 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 206.910 219.800 ;
    LAYER metal2 ;
    RECT 0 0 206.910 219.800 ;
    LAYER metal3 ;
    RECT 0.070 0 206.910 219.800 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 2.905 ;
    RECT 0 2.975 0.070 4.445 ;
    RECT 0 4.515 0.070 5.985 ;
    RECT 0 6.055 0.070 7.525 ;
    RECT 0 7.595 0.070 9.065 ;
    RECT 0 9.135 0.070 10.605 ;
    RECT 0 10.675 0.070 12.145 ;
    RECT 0 12.215 0.070 13.685 ;
    RECT 0 13.755 0.070 15.225 ;
    RECT 0 15.295 0.070 16.765 ;
    RECT 0 16.835 0.070 18.305 ;
    RECT 0 18.375 0.070 19.845 ;
    RECT 0 19.915 0.070 21.385 ;
    RECT 0 21.455 0.070 22.925 ;
    RECT 0 22.995 0.070 24.465 ;
    RECT 0 24.535 0.070 26.005 ;
    RECT 0 26.075 0.070 27.545 ;
    RECT 0 27.615 0.070 29.085 ;
    RECT 0 29.155 0.070 30.625 ;
    RECT 0 30.695 0.070 32.165 ;
    RECT 0 32.235 0.070 33.705 ;
    RECT 0 33.775 0.070 35.245 ;
    RECT 0 35.315 0.070 36.785 ;
    RECT 0 36.855 0.070 38.325 ;
    RECT 0 38.395 0.070 39.865 ;
    RECT 0 39.935 0.070 41.405 ;
    RECT 0 41.475 0.070 42.945 ;
    RECT 0 43.015 0.070 44.485 ;
    RECT 0 44.555 0.070 46.025 ;
    RECT 0 46.095 0.070 47.565 ;
    RECT 0 47.635 0.070 49.105 ;
    RECT 0 49.175 0.070 50.645 ;
    RECT 0 50.715 0.070 52.185 ;
    RECT 0 52.255 0.070 53.725 ;
    RECT 0 53.795 0.070 55.265 ;
    RECT 0 55.335 0.070 56.805 ;
    RECT 0 56.875 0.070 58.345 ;
    RECT 0 58.415 0.070 59.885 ;
    RECT 0 59.955 0.070 63.665 ;
    RECT 0 63.735 0.070 65.205 ;
    RECT 0 65.275 0.070 66.745 ;
    RECT 0 66.815 0.070 68.285 ;
    RECT 0 68.355 0.070 69.825 ;
    RECT 0 69.895 0.070 71.365 ;
    RECT 0 71.435 0.070 72.905 ;
    RECT 0 72.975 0.070 74.445 ;
    RECT 0 74.515 0.070 75.985 ;
    RECT 0 76.055 0.070 77.525 ;
    RECT 0 77.595 0.070 79.065 ;
    RECT 0 79.135 0.070 80.605 ;
    RECT 0 80.675 0.070 82.145 ;
    RECT 0 82.215 0.070 83.685 ;
    RECT 0 83.755 0.070 85.225 ;
    RECT 0 85.295 0.070 86.765 ;
    RECT 0 86.835 0.070 88.305 ;
    RECT 0 88.375 0.070 89.845 ;
    RECT 0 89.915 0.070 91.385 ;
    RECT 0 91.455 0.070 92.925 ;
    RECT 0 92.995 0.070 94.465 ;
    RECT 0 94.535 0.070 96.005 ;
    RECT 0 96.075 0.070 97.545 ;
    RECT 0 97.615 0.070 99.085 ;
    RECT 0 99.155 0.070 100.625 ;
    RECT 0 100.695 0.070 102.165 ;
    RECT 0 102.235 0.070 103.705 ;
    RECT 0 103.775 0.070 105.245 ;
    RECT 0 105.315 0.070 106.785 ;
    RECT 0 106.855 0.070 108.325 ;
    RECT 0 108.395 0.070 109.865 ;
    RECT 0 109.935 0.070 111.405 ;
    RECT 0 111.475 0.070 112.945 ;
    RECT 0 113.015 0.070 114.485 ;
    RECT 0 114.555 0.070 116.025 ;
    RECT 0 116.095 0.070 117.565 ;
    RECT 0 117.635 0.070 119.105 ;
    RECT 0 119.175 0.070 120.645 ;
    RECT 0 120.715 0.070 122.185 ;
    RECT 0 122.255 0.070 125.965 ;
    RECT 0 126.035 0.070 127.505 ;
    RECT 0 127.575 0.070 129.045 ;
    RECT 0 129.115 0.070 130.585 ;
    RECT 0 130.655 0.070 132.125 ;
    RECT 0 132.195 0.070 133.665 ;
    RECT 0 133.735 0.070 135.205 ;
    RECT 0 135.275 0.070 136.745 ;
    RECT 0 136.815 0.070 138.285 ;
    RECT 0 138.355 0.070 139.825 ;
    RECT 0 139.895 0.070 141.365 ;
    RECT 0 141.435 0.070 142.905 ;
    RECT 0 142.975 0.070 144.445 ;
    RECT 0 144.515 0.070 145.985 ;
    RECT 0 146.055 0.070 147.525 ;
    RECT 0 147.595 0.070 149.065 ;
    RECT 0 149.135 0.070 150.605 ;
    RECT 0 150.675 0.070 152.145 ;
    RECT 0 152.215 0.070 153.685 ;
    RECT 0 153.755 0.070 155.225 ;
    RECT 0 155.295 0.070 156.765 ;
    RECT 0 156.835 0.070 158.305 ;
    RECT 0 158.375 0.070 159.845 ;
    RECT 0 159.915 0.070 161.385 ;
    RECT 0 161.455 0.070 162.925 ;
    RECT 0 162.995 0.070 164.465 ;
    RECT 0 164.535 0.070 166.005 ;
    RECT 0 166.075 0.070 167.545 ;
    RECT 0 167.615 0.070 169.085 ;
    RECT 0 169.155 0.070 170.625 ;
    RECT 0 170.695 0.070 172.165 ;
    RECT 0 172.235 0.070 173.705 ;
    RECT 0 173.775 0.070 175.245 ;
    RECT 0 175.315 0.070 176.785 ;
    RECT 0 176.855 0.070 178.325 ;
    RECT 0 178.395 0.070 179.865 ;
    RECT 0 179.935 0.070 181.405 ;
    RECT 0 181.475 0.070 182.945 ;
    RECT 0 183.015 0.070 184.485 ;
    RECT 0 184.555 0.070 188.265 ;
    RECT 0 188.335 0.070 189.805 ;
    RECT 0 189.875 0.070 191.345 ;
    RECT 0 191.415 0.070 192.885 ;
    RECT 0 192.955 0.070 194.425 ;
    RECT 0 194.495 0.070 195.965 ;
    RECT 0 196.035 0.070 197.505 ;
    RECT 0 197.575 0.070 199.045 ;
    RECT 0 199.115 0.070 200.585 ;
    RECT 0 200.655 0.070 202.125 ;
    RECT 0 202.195 0.070 203.665 ;
    RECT 0 203.735 0.070 207.445 ;
    RECT 0 207.515 0.070 208.985 ;
    RECT 0 209.055 0.070 210.525 ;
    RECT 0 210.595 0.070 219.800 ;
    LAYER metal4 ;
    RECT 0 0 206.910 1.400 ;
    RECT 0 218.400 206.910 219.800 ;
    RECT 0.000 1.400 1.260 218.400 ;
    RECT 1.540 1.400 2.380 218.400 ;
    RECT 2.660 1.400 3.500 218.400 ;
    RECT 3.780 1.400 4.620 218.400 ;
    RECT 4.900 1.400 5.740 218.400 ;
    RECT 6.020 1.400 6.860 218.400 ;
    RECT 7.140 1.400 7.980 218.400 ;
    RECT 8.260 1.400 9.100 218.400 ;
    RECT 9.380 1.400 10.220 218.400 ;
    RECT 10.500 1.400 11.340 218.400 ;
    RECT 11.620 1.400 12.460 218.400 ;
    RECT 12.740 1.400 13.580 218.400 ;
    RECT 13.860 1.400 14.700 218.400 ;
    RECT 14.980 1.400 15.820 218.400 ;
    RECT 16.100 1.400 16.940 218.400 ;
    RECT 17.220 1.400 18.060 218.400 ;
    RECT 18.340 1.400 19.180 218.400 ;
    RECT 19.460 1.400 20.300 218.400 ;
    RECT 20.580 1.400 21.420 218.400 ;
    RECT 21.700 1.400 22.540 218.400 ;
    RECT 22.820 1.400 23.660 218.400 ;
    RECT 23.940 1.400 24.780 218.400 ;
    RECT 25.060 1.400 25.900 218.400 ;
    RECT 26.180 1.400 27.020 218.400 ;
    RECT 27.300 1.400 28.140 218.400 ;
    RECT 28.420 1.400 29.260 218.400 ;
    RECT 29.540 1.400 30.380 218.400 ;
    RECT 30.660 1.400 31.500 218.400 ;
    RECT 31.780 1.400 32.620 218.400 ;
    RECT 32.900 1.400 33.740 218.400 ;
    RECT 34.020 1.400 34.860 218.400 ;
    RECT 35.140 1.400 35.980 218.400 ;
    RECT 36.260 1.400 37.100 218.400 ;
    RECT 37.380 1.400 38.220 218.400 ;
    RECT 38.500 1.400 39.340 218.400 ;
    RECT 39.620 1.400 40.460 218.400 ;
    RECT 40.740 1.400 41.580 218.400 ;
    RECT 41.860 1.400 42.700 218.400 ;
    RECT 42.980 1.400 43.820 218.400 ;
    RECT 44.100 1.400 44.940 218.400 ;
    RECT 45.220 1.400 46.060 218.400 ;
    RECT 46.340 1.400 47.180 218.400 ;
    RECT 47.460 1.400 48.300 218.400 ;
    RECT 48.580 1.400 49.420 218.400 ;
    RECT 49.700 1.400 50.540 218.400 ;
    RECT 50.820 1.400 51.660 218.400 ;
    RECT 51.940 1.400 52.780 218.400 ;
    RECT 53.060 1.400 53.900 218.400 ;
    RECT 54.180 1.400 55.020 218.400 ;
    RECT 55.300 1.400 56.140 218.400 ;
    RECT 56.420 1.400 57.260 218.400 ;
    RECT 57.540 1.400 58.380 218.400 ;
    RECT 58.660 1.400 59.500 218.400 ;
    RECT 59.780 1.400 60.620 218.400 ;
    RECT 60.900 1.400 61.740 218.400 ;
    RECT 62.020 1.400 62.860 218.400 ;
    RECT 63.140 1.400 63.980 218.400 ;
    RECT 64.260 1.400 65.100 218.400 ;
    RECT 65.380 1.400 66.220 218.400 ;
    RECT 66.500 1.400 67.340 218.400 ;
    RECT 67.620 1.400 68.460 218.400 ;
    RECT 68.740 1.400 69.580 218.400 ;
    RECT 69.860 1.400 70.700 218.400 ;
    RECT 70.980 1.400 71.820 218.400 ;
    RECT 72.100 1.400 72.940 218.400 ;
    RECT 73.220 1.400 74.060 218.400 ;
    RECT 74.340 1.400 75.180 218.400 ;
    RECT 75.460 1.400 76.300 218.400 ;
    RECT 76.580 1.400 77.420 218.400 ;
    RECT 77.700 1.400 78.540 218.400 ;
    RECT 78.820 1.400 79.660 218.400 ;
    RECT 79.940 1.400 80.780 218.400 ;
    RECT 81.060 1.400 81.900 218.400 ;
    RECT 82.180 1.400 83.020 218.400 ;
    RECT 83.300 1.400 84.140 218.400 ;
    RECT 84.420 1.400 85.260 218.400 ;
    RECT 85.540 1.400 86.380 218.400 ;
    RECT 86.660 1.400 87.500 218.400 ;
    RECT 87.780 1.400 88.620 218.400 ;
    RECT 88.900 1.400 89.740 218.400 ;
    RECT 90.020 1.400 90.860 218.400 ;
    RECT 91.140 1.400 91.980 218.400 ;
    RECT 92.260 1.400 93.100 218.400 ;
    RECT 93.380 1.400 94.220 218.400 ;
    RECT 94.500 1.400 95.340 218.400 ;
    RECT 95.620 1.400 96.460 218.400 ;
    RECT 96.740 1.400 97.580 218.400 ;
    RECT 97.860 1.400 98.700 218.400 ;
    RECT 98.980 1.400 99.820 218.400 ;
    RECT 100.100 1.400 100.940 218.400 ;
    RECT 101.220 1.400 102.060 218.400 ;
    RECT 102.340 1.400 103.180 218.400 ;
    RECT 103.460 1.400 104.300 218.400 ;
    RECT 104.580 1.400 105.420 218.400 ;
    RECT 105.700 1.400 106.540 218.400 ;
    RECT 106.820 1.400 107.660 218.400 ;
    RECT 107.940 1.400 108.780 218.400 ;
    RECT 109.060 1.400 109.900 218.400 ;
    RECT 110.180 1.400 111.020 218.400 ;
    RECT 111.300 1.400 112.140 218.400 ;
    RECT 112.420 1.400 113.260 218.400 ;
    RECT 113.540 1.400 114.380 218.400 ;
    RECT 114.660 1.400 115.500 218.400 ;
    RECT 115.780 1.400 116.620 218.400 ;
    RECT 116.900 1.400 117.740 218.400 ;
    RECT 118.020 1.400 118.860 218.400 ;
    RECT 119.140 1.400 119.980 218.400 ;
    RECT 120.260 1.400 121.100 218.400 ;
    RECT 121.380 1.400 122.220 218.400 ;
    RECT 122.500 1.400 123.340 218.400 ;
    RECT 123.620 1.400 124.460 218.400 ;
    RECT 124.740 1.400 125.580 218.400 ;
    RECT 125.860 1.400 126.700 218.400 ;
    RECT 126.980 1.400 127.820 218.400 ;
    RECT 128.100 1.400 128.940 218.400 ;
    RECT 129.220 1.400 130.060 218.400 ;
    RECT 130.340 1.400 131.180 218.400 ;
    RECT 131.460 1.400 132.300 218.400 ;
    RECT 132.580 1.400 133.420 218.400 ;
    RECT 133.700 1.400 134.540 218.400 ;
    RECT 134.820 1.400 135.660 218.400 ;
    RECT 135.940 1.400 136.780 218.400 ;
    RECT 137.060 1.400 137.900 218.400 ;
    RECT 138.180 1.400 139.020 218.400 ;
    RECT 139.300 1.400 140.140 218.400 ;
    RECT 140.420 1.400 141.260 218.400 ;
    RECT 141.540 1.400 142.380 218.400 ;
    RECT 142.660 1.400 143.500 218.400 ;
    RECT 143.780 1.400 144.620 218.400 ;
    RECT 144.900 1.400 145.740 218.400 ;
    RECT 146.020 1.400 146.860 218.400 ;
    RECT 147.140 1.400 147.980 218.400 ;
    RECT 148.260 1.400 149.100 218.400 ;
    RECT 149.380 1.400 150.220 218.400 ;
    RECT 150.500 1.400 151.340 218.400 ;
    RECT 151.620 1.400 152.460 218.400 ;
    RECT 152.740 1.400 153.580 218.400 ;
    RECT 153.860 1.400 154.700 218.400 ;
    RECT 154.980 1.400 155.820 218.400 ;
    RECT 156.100 1.400 156.940 218.400 ;
    RECT 157.220 1.400 158.060 218.400 ;
    RECT 158.340 1.400 159.180 218.400 ;
    RECT 159.460 1.400 160.300 218.400 ;
    RECT 160.580 1.400 161.420 218.400 ;
    RECT 161.700 1.400 162.540 218.400 ;
    RECT 162.820 1.400 163.660 218.400 ;
    RECT 163.940 1.400 164.780 218.400 ;
    RECT 165.060 1.400 165.900 218.400 ;
    RECT 166.180 1.400 167.020 218.400 ;
    RECT 167.300 1.400 168.140 218.400 ;
    RECT 168.420 1.400 169.260 218.400 ;
    RECT 169.540 1.400 170.380 218.400 ;
    RECT 170.660 1.400 171.500 218.400 ;
    RECT 171.780 1.400 172.620 218.400 ;
    RECT 172.900 1.400 173.740 218.400 ;
    RECT 174.020 1.400 174.860 218.400 ;
    RECT 175.140 1.400 175.980 218.400 ;
    RECT 176.260 1.400 177.100 218.400 ;
    RECT 177.380 1.400 178.220 218.400 ;
    RECT 178.500 1.400 179.340 218.400 ;
    RECT 179.620 1.400 180.460 218.400 ;
    RECT 180.740 1.400 181.580 218.400 ;
    RECT 181.860 1.400 182.700 218.400 ;
    RECT 182.980 1.400 183.820 218.400 ;
    RECT 184.100 1.400 184.940 218.400 ;
    RECT 185.220 1.400 186.060 218.400 ;
    RECT 186.340 1.400 187.180 218.400 ;
    RECT 187.460 1.400 188.300 218.400 ;
    RECT 188.580 1.400 189.420 218.400 ;
    RECT 189.700 1.400 190.540 218.400 ;
    RECT 190.820 1.400 191.660 218.400 ;
    RECT 191.940 1.400 192.780 218.400 ;
    RECT 193.060 1.400 193.900 218.400 ;
    RECT 194.180 1.400 195.020 218.400 ;
    RECT 195.300 1.400 196.140 218.400 ;
    RECT 196.420 1.400 197.260 218.400 ;
    RECT 197.540 1.400 198.380 218.400 ;
    RECT 198.660 1.400 199.500 218.400 ;
    RECT 199.780 1.400 200.620 218.400 ;
    RECT 200.900 1.400 201.740 218.400 ;
    RECT 202.020 1.400 202.860 218.400 ;
    RECT 203.140 1.400 203.980 218.400 ;
    RECT 204.260 1.400 205.100 218.400 ;
    RECT 205.380 1.400 206.910 218.400 ;
    LAYER OVERLAP ;
    RECT 0 0 206.910 219.800 ;
  END
END fakeram45_2048x39

END LIBRARY
