// Standard header to adapt well known macros for prints and assertions.

// Users can define 'ASSERT_VERBOSE_COND' to add an extra gate to assert error printing.
`ifndef ASSERT_VERBOSE_COND_
  `ifdef ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ (`ASSERT_VERBOSE_COND)
  `else  // ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ 1
  `endif // ASSERT_VERBOSE_COND
`endif // not def ASSERT_VERBOSE_COND_

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifndef STOP_COND_
  `ifdef STOP_COND
    `define STOP_COND_ (`STOP_COND)
  `else  // STOP_COND
    `define STOP_COND_ 1
  `endif // STOP_COND
`endif // not def STOP_COND_

module Rob(
  input         clock,
                reset,
                io_enq_valids_0,
                io_enq_valids_1,
                io_enq_valids_2,
                io_enq_valids_3,
  input  [6:0]  io_enq_uops_0_uopc,
  input         io_enq_uops_0_is_rvc,
                io_enq_uops_0_is_br,
                io_enq_uops_0_is_jalr,
                io_enq_uops_0_is_jal,
  input  [19:0] io_enq_uops_0_br_mask,
  input  [5:0]  io_enq_uops_0_ftq_idx,
  input         io_enq_uops_0_edge_inst,
  input  [5:0]  io_enq_uops_0_pc_lob,
  input  [6:0]  io_enq_uops_0_rob_idx,
                io_enq_uops_0_pdst,
                io_enq_uops_0_stale_pdst,
  input         io_enq_uops_0_exception,
  input  [63:0] io_enq_uops_0_exc_cause,
  input         io_enq_uops_0_is_fence,
                io_enq_uops_0_is_fencei,
                io_enq_uops_0_uses_ldq,
                io_enq_uops_0_uses_stq,
                io_enq_uops_0_is_sys_pc2epc,
                io_enq_uops_0_is_unique,
                io_enq_uops_0_flush_on_commit,
  input  [5:0]  io_enq_uops_0_ldst,
  input         io_enq_uops_0_ldst_val,
  input  [1:0]  io_enq_uops_0_dst_rtype,
  input         io_enq_uops_0_fp_val,
  input  [1:0]  io_enq_uops_0_debug_fsrc,
  input  [6:0]  io_enq_uops_1_uopc,
  input         io_enq_uops_1_is_rvc,
                io_enq_uops_1_is_br,
                io_enq_uops_1_is_jalr,
                io_enq_uops_1_is_jal,
  input  [19:0] io_enq_uops_1_br_mask,
  input  [5:0]  io_enq_uops_1_ftq_idx,
  input         io_enq_uops_1_edge_inst,
  input  [5:0]  io_enq_uops_1_pc_lob,
  input  [6:0]  io_enq_uops_1_rob_idx,
                io_enq_uops_1_pdst,
                io_enq_uops_1_stale_pdst,
  input         io_enq_uops_1_exception,
  input  [63:0] io_enq_uops_1_exc_cause,
  input         io_enq_uops_1_is_fence,
                io_enq_uops_1_is_fencei,
                io_enq_uops_1_uses_ldq,
                io_enq_uops_1_uses_stq,
                io_enq_uops_1_is_sys_pc2epc,
                io_enq_uops_1_is_unique,
                io_enq_uops_1_flush_on_commit,
  input  [5:0]  io_enq_uops_1_ldst,
  input         io_enq_uops_1_ldst_val,
  input  [1:0]  io_enq_uops_1_dst_rtype,
  input         io_enq_uops_1_fp_val,
  input  [1:0]  io_enq_uops_1_debug_fsrc,
  input  [6:0]  io_enq_uops_2_uopc,
  input         io_enq_uops_2_is_rvc,
                io_enq_uops_2_is_br,
                io_enq_uops_2_is_jalr,
                io_enq_uops_2_is_jal,
  input  [19:0] io_enq_uops_2_br_mask,
  input  [5:0]  io_enq_uops_2_ftq_idx,
  input         io_enq_uops_2_edge_inst,
  input  [5:0]  io_enq_uops_2_pc_lob,
  input  [6:0]  io_enq_uops_2_rob_idx,
                io_enq_uops_2_pdst,
                io_enq_uops_2_stale_pdst,
  input         io_enq_uops_2_exception,
  input  [63:0] io_enq_uops_2_exc_cause,
  input         io_enq_uops_2_is_fence,
                io_enq_uops_2_is_fencei,
                io_enq_uops_2_uses_ldq,
                io_enq_uops_2_uses_stq,
                io_enq_uops_2_is_sys_pc2epc,
                io_enq_uops_2_is_unique,
                io_enq_uops_2_flush_on_commit,
  input  [5:0]  io_enq_uops_2_ldst,
  input         io_enq_uops_2_ldst_val,
  input  [1:0]  io_enq_uops_2_dst_rtype,
  input         io_enq_uops_2_fp_val,
  input  [1:0]  io_enq_uops_2_debug_fsrc,
  input  [6:0]  io_enq_uops_3_uopc,
  input         io_enq_uops_3_is_rvc,
                io_enq_uops_3_is_br,
                io_enq_uops_3_is_jalr,
                io_enq_uops_3_is_jal,
  input  [19:0] io_enq_uops_3_br_mask,
  input  [5:0]  io_enq_uops_3_ftq_idx,
  input         io_enq_uops_3_edge_inst,
  input  [5:0]  io_enq_uops_3_pc_lob,
  input  [6:0]  io_enq_uops_3_rob_idx,
                io_enq_uops_3_pdst,
                io_enq_uops_3_stale_pdst,
  input         io_enq_uops_3_exception,
  input  [63:0] io_enq_uops_3_exc_cause,
  input         io_enq_uops_3_is_fence,
                io_enq_uops_3_is_fencei,
                io_enq_uops_3_uses_ldq,
                io_enq_uops_3_uses_stq,
                io_enq_uops_3_is_sys_pc2epc,
                io_enq_uops_3_is_unique,
                io_enq_uops_3_flush_on_commit,
  input  [5:0]  io_enq_uops_3_ldst,
  input         io_enq_uops_3_ldst_val,
  input  [1:0]  io_enq_uops_3_dst_rtype,
  input         io_enq_uops_3_fp_val,
  input  [1:0]  io_enq_uops_3_debug_fsrc,
  input         io_enq_partial_stall,
  input  [39:0] io_xcpt_fetch_pc,
  output [6:0]  io_rob_tail_idx,
                io_rob_head_idx,
  input  [19:0] io_brupdate_b1_resolve_mask,
                io_brupdate_b1_mispredict_mask,
  input  [6:0]  io_brupdate_b2_uop_rob_idx,
  input         io_brupdate_b2_mispredict,
                io_wb_resps_0_valid,
  input  [6:0]  io_wb_resps_0_bits_uop_rob_idx,
                io_wb_resps_0_bits_uop_pdst,
  input         io_wb_resps_0_bits_predicated,
                io_wb_resps_1_valid,
  input  [6:0]  io_wb_resps_1_bits_uop_rob_idx,
                io_wb_resps_1_bits_uop_pdst,
  input         io_wb_resps_2_valid,
  input  [6:0]  io_wb_resps_2_bits_uop_rob_idx,
                io_wb_resps_2_bits_uop_pdst,
  input         io_wb_resps_3_valid,
  input  [6:0]  io_wb_resps_3_bits_uop_rob_idx,
                io_wb_resps_3_bits_uop_pdst,
  input         io_wb_resps_4_valid,
  input  [6:0]  io_wb_resps_4_bits_uop_rob_idx,
                io_wb_resps_4_bits_uop_pdst,
  input         io_wb_resps_5_valid,
  input  [6:0]  io_wb_resps_5_bits_uop_rob_idx,
                io_wb_resps_5_bits_uop_pdst,
  input         io_wb_resps_6_valid,
  input  [6:0]  io_wb_resps_6_bits_uop_rob_idx,
                io_wb_resps_6_bits_uop_pdst,
  input         io_wb_resps_6_bits_predicated,
                io_wb_resps_7_valid,
  input  [6:0]  io_wb_resps_7_bits_uop_rob_idx,
                io_wb_resps_7_bits_uop_pdst,
  input         io_wb_resps_8_valid,
  input  [6:0]  io_wb_resps_8_bits_uop_rob_idx,
                io_wb_resps_8_bits_uop_pdst,
  input         io_wb_resps_9_valid,
  input  [6:0]  io_wb_resps_9_bits_uop_rob_idx,
                io_wb_resps_9_bits_uop_pdst,
  input         io_lsu_clr_bsy_0_valid,
  input  [6:0]  io_lsu_clr_bsy_0_bits,
  input         io_lsu_clr_bsy_1_valid,
  input  [6:0]  io_lsu_clr_bsy_1_bits,
  input         io_lsu_clr_bsy_2_valid,
  input  [6:0]  io_lsu_clr_bsy_2_bits,
  input         io_fflags_0_valid,
  input  [6:0]  io_fflags_0_bits_uop_rob_idx,
  input  [4:0]  io_fflags_0_bits_flags,
  input         io_fflags_2_valid,
  input  [6:0]  io_fflags_2_bits_uop_rob_idx,
  input  [4:0]  io_fflags_2_bits_flags,
  input         io_fflags_3_valid,
  input  [6:0]  io_fflags_3_bits_uop_rob_idx,
  input  [4:0]  io_fflags_3_bits_flags,
  input         io_lxcpt_valid,
  input  [19:0] io_lxcpt_bits_uop_br_mask,
  input  [6:0]  io_lxcpt_bits_uop_rob_idx,
  input  [4:0]  io_lxcpt_bits_cause,
  input  [39:0] io_lxcpt_bits_badvaddr,
  output        io_commit_valids_0,
                io_commit_valids_1,
                io_commit_valids_2,
                io_commit_valids_3,
                io_commit_arch_valids_0,
                io_commit_arch_valids_1,
                io_commit_arch_valids_2,
                io_commit_arch_valids_3,
                io_commit_uops_0_is_br,
                io_commit_uops_0_is_jalr,
                io_commit_uops_0_is_jal,
  output [5:0]  io_commit_uops_0_ftq_idx,
  output [6:0]  io_commit_uops_0_pdst,
                io_commit_uops_0_stale_pdst,
  output        io_commit_uops_0_is_fencei,
                io_commit_uops_0_uses_ldq,
                io_commit_uops_0_uses_stq,
  output [5:0]  io_commit_uops_0_ldst,
  output        io_commit_uops_0_ldst_val,
  output [1:0]  io_commit_uops_0_dst_rtype,
                io_commit_uops_0_debug_fsrc,
  output        io_commit_uops_1_is_br,
                io_commit_uops_1_is_jalr,
                io_commit_uops_1_is_jal,
  output [5:0]  io_commit_uops_1_ftq_idx,
  output [6:0]  io_commit_uops_1_pdst,
                io_commit_uops_1_stale_pdst,
  output        io_commit_uops_1_is_fencei,
                io_commit_uops_1_uses_ldq,
                io_commit_uops_1_uses_stq,
  output [5:0]  io_commit_uops_1_ldst,
  output        io_commit_uops_1_ldst_val,
  output [1:0]  io_commit_uops_1_dst_rtype,
                io_commit_uops_1_debug_fsrc,
  output        io_commit_uops_2_is_br,
                io_commit_uops_2_is_jalr,
                io_commit_uops_2_is_jal,
  output [5:0]  io_commit_uops_2_ftq_idx,
  output [6:0]  io_commit_uops_2_pdst,
                io_commit_uops_2_stale_pdst,
  output        io_commit_uops_2_is_fencei,
                io_commit_uops_2_uses_ldq,
                io_commit_uops_2_uses_stq,
  output [5:0]  io_commit_uops_2_ldst,
  output        io_commit_uops_2_ldst_val,
  output [1:0]  io_commit_uops_2_dst_rtype,
                io_commit_uops_2_debug_fsrc,
  output        io_commit_uops_3_is_br,
                io_commit_uops_3_is_jalr,
                io_commit_uops_3_is_jal,
  output [5:0]  io_commit_uops_3_ftq_idx,
  output [6:0]  io_commit_uops_3_pdst,
                io_commit_uops_3_stale_pdst,
  output        io_commit_uops_3_is_fencei,
                io_commit_uops_3_uses_ldq,
                io_commit_uops_3_uses_stq,
  output [5:0]  io_commit_uops_3_ldst,
  output        io_commit_uops_3_ldst_val,
  output [1:0]  io_commit_uops_3_dst_rtype,
                io_commit_uops_3_debug_fsrc,
  output        io_commit_fflags_valid,
  output [4:0]  io_commit_fflags_bits,
  output        io_commit_rbk_valids_0,
                io_commit_rbk_valids_1,
                io_commit_rbk_valids_2,
                io_commit_rbk_valids_3,
                io_commit_rollback,
                io_com_load_is_at_rob_head,
                io_com_xcpt_valid,
  output [5:0]  io_com_xcpt_bits_ftq_idx,
  output        io_com_xcpt_bits_edge_inst,
  output [5:0]  io_com_xcpt_bits_pc_lob,
  output [63:0] io_com_xcpt_bits_cause,
                io_com_xcpt_bits_badvaddr,
  input         io_csr_stall,
  output        io_flush_valid,
  output [5:0]  io_flush_bits_ftq_idx,
  output        io_flush_bits_edge_inst,
                io_flush_bits_is_rvc,
  output [5:0]  io_flush_bits_pc_lob,
  output [2:0]  io_flush_bits_flush_typ,
  output        io_empty,
                io_ready,
                io_flush_frontend
);

  wire        empty;
  wire        full;
  wire        will_commit_3;
  wire        will_commit_2;
  wire        will_commit_1;
  wire        will_commit_0;
  reg  [1:0]  rob_state;
  reg  [4:0]  rob_head;
  reg  [1:0]  rob_head_lsb;
  wire [6:0]  rob_head_idx = {rob_head, rob_head_lsb};
  reg  [4:0]  rob_tail;
  reg  [1:0]  rob_tail_lsb;
  wire [6:0]  rob_tail_idx = {rob_tail, rob_tail_lsb};
  reg  [4:0]  rob_pnr;
  reg  [1:0]  rob_pnr_lsb;
  wire        _io_commit_rollback_T_3 = rob_state == 2'h2;
  wire [4:0]  com_idx = _io_commit_rollback_T_3 ? rob_tail : rob_head;
  reg         maybe_full;
  reg         r_xcpt_val;
  reg  [19:0] r_xcpt_uop_br_mask;
  reg  [6:0]  r_xcpt_uop_rob_idx;
  reg  [63:0] r_xcpt_uop_exc_cause;
  reg  [39:0] r_xcpt_badvaddr;
  reg  [4:0]  rob_fflags_0_0;
  reg  [4:0]  rob_fflags_0_1;
  reg  [4:0]  rob_fflags_0_2;
  reg  [4:0]  rob_fflags_0_3;
  reg  [4:0]  rob_fflags_0_4;
  reg  [4:0]  rob_fflags_0_5;
  reg  [4:0]  rob_fflags_0_6;
  reg  [4:0]  rob_fflags_0_7;
  reg  [4:0]  rob_fflags_0_8;
  reg  [4:0]  rob_fflags_0_9;
  reg  [4:0]  rob_fflags_0_10;
  reg  [4:0]  rob_fflags_0_11;
  reg  [4:0]  rob_fflags_0_12;
  reg  [4:0]  rob_fflags_0_13;
  reg  [4:0]  rob_fflags_0_14;
  reg  [4:0]  rob_fflags_0_15;
  reg  [4:0]  rob_fflags_0_16;
  reg  [4:0]  rob_fflags_0_17;
  reg  [4:0]  rob_fflags_0_18;
  reg  [4:0]  rob_fflags_0_19;
  reg  [4:0]  rob_fflags_0_20;
  reg  [4:0]  rob_fflags_0_21;
  reg  [4:0]  rob_fflags_0_22;
  reg  [4:0]  rob_fflags_0_23;
  reg  [4:0]  rob_fflags_0_24;
  reg  [4:0]  rob_fflags_0_25;
  reg  [4:0]  rob_fflags_0_26;
  reg  [4:0]  rob_fflags_0_27;
  reg  [4:0]  rob_fflags_0_28;
  reg  [4:0]  rob_fflags_0_29;
  reg  [4:0]  rob_fflags_0_30;
  reg  [4:0]  rob_fflags_0_31;
  reg  [4:0]  rob_fflags_1_0;
  reg  [4:0]  rob_fflags_1_1;
  reg  [4:0]  rob_fflags_1_2;
  reg  [4:0]  rob_fflags_1_3;
  reg  [4:0]  rob_fflags_1_4;
  reg  [4:0]  rob_fflags_1_5;
  reg  [4:0]  rob_fflags_1_6;
  reg  [4:0]  rob_fflags_1_7;
  reg  [4:0]  rob_fflags_1_8;
  reg  [4:0]  rob_fflags_1_9;
  reg  [4:0]  rob_fflags_1_10;
  reg  [4:0]  rob_fflags_1_11;
  reg  [4:0]  rob_fflags_1_12;
  reg  [4:0]  rob_fflags_1_13;
  reg  [4:0]  rob_fflags_1_14;
  reg  [4:0]  rob_fflags_1_15;
  reg  [4:0]  rob_fflags_1_16;
  reg  [4:0]  rob_fflags_1_17;
  reg  [4:0]  rob_fflags_1_18;
  reg  [4:0]  rob_fflags_1_19;
  reg  [4:0]  rob_fflags_1_20;
  reg  [4:0]  rob_fflags_1_21;
  reg  [4:0]  rob_fflags_1_22;
  reg  [4:0]  rob_fflags_1_23;
  reg  [4:0]  rob_fflags_1_24;
  reg  [4:0]  rob_fflags_1_25;
  reg  [4:0]  rob_fflags_1_26;
  reg  [4:0]  rob_fflags_1_27;
  reg  [4:0]  rob_fflags_1_28;
  reg  [4:0]  rob_fflags_1_29;
  reg  [4:0]  rob_fflags_1_30;
  reg  [4:0]  rob_fflags_1_31;
  reg  [4:0]  rob_fflags_2_0;
  reg  [4:0]  rob_fflags_2_1;
  reg  [4:0]  rob_fflags_2_2;
  reg  [4:0]  rob_fflags_2_3;
  reg  [4:0]  rob_fflags_2_4;
  reg  [4:0]  rob_fflags_2_5;
  reg  [4:0]  rob_fflags_2_6;
  reg  [4:0]  rob_fflags_2_7;
  reg  [4:0]  rob_fflags_2_8;
  reg  [4:0]  rob_fflags_2_9;
  reg  [4:0]  rob_fflags_2_10;
  reg  [4:0]  rob_fflags_2_11;
  reg  [4:0]  rob_fflags_2_12;
  reg  [4:0]  rob_fflags_2_13;
  reg  [4:0]  rob_fflags_2_14;
  reg  [4:0]  rob_fflags_2_15;
  reg  [4:0]  rob_fflags_2_16;
  reg  [4:0]  rob_fflags_2_17;
  reg  [4:0]  rob_fflags_2_18;
  reg  [4:0]  rob_fflags_2_19;
  reg  [4:0]  rob_fflags_2_20;
  reg  [4:0]  rob_fflags_2_21;
  reg  [4:0]  rob_fflags_2_22;
  reg  [4:0]  rob_fflags_2_23;
  reg  [4:0]  rob_fflags_2_24;
  reg  [4:0]  rob_fflags_2_25;
  reg  [4:0]  rob_fflags_2_26;
  reg  [4:0]  rob_fflags_2_27;
  reg  [4:0]  rob_fflags_2_28;
  reg  [4:0]  rob_fflags_2_29;
  reg  [4:0]  rob_fflags_2_30;
  reg  [4:0]  rob_fflags_2_31;
  reg  [4:0]  rob_fflags_3_0;
  reg  [4:0]  rob_fflags_3_1;
  reg  [4:0]  rob_fflags_3_2;
  reg  [4:0]  rob_fflags_3_3;
  reg  [4:0]  rob_fflags_3_4;
  reg  [4:0]  rob_fflags_3_5;
  reg  [4:0]  rob_fflags_3_6;
  reg  [4:0]  rob_fflags_3_7;
  reg  [4:0]  rob_fflags_3_8;
  reg  [4:0]  rob_fflags_3_9;
  reg  [4:0]  rob_fflags_3_10;
  reg  [4:0]  rob_fflags_3_11;
  reg  [4:0]  rob_fflags_3_12;
  reg  [4:0]  rob_fflags_3_13;
  reg  [4:0]  rob_fflags_3_14;
  reg  [4:0]  rob_fflags_3_15;
  reg  [4:0]  rob_fflags_3_16;
  reg  [4:0]  rob_fflags_3_17;
  reg  [4:0]  rob_fflags_3_18;
  reg  [4:0]  rob_fflags_3_19;
  reg  [4:0]  rob_fflags_3_20;
  reg  [4:0]  rob_fflags_3_21;
  reg  [4:0]  rob_fflags_3_22;
  reg  [4:0]  rob_fflags_3_23;
  reg  [4:0]  rob_fflags_3_24;
  reg  [4:0]  rob_fflags_3_25;
  reg  [4:0]  rob_fflags_3_26;
  reg  [4:0]  rob_fflags_3_27;
  reg  [4:0]  rob_fflags_3_28;
  reg  [4:0]  rob_fflags_3_29;
  reg  [4:0]  rob_fflags_3_30;
  reg  [4:0]  rob_fflags_3_31;
  reg         rob_val_0;
  reg         rob_val_1;
  reg         rob_val_2;
  reg         rob_val_3;
  reg         rob_val_4;
  reg         rob_val_5;
  reg         rob_val_6;
  reg         rob_val_7;
  reg         rob_val_8;
  reg         rob_val_9;
  reg         rob_val_10;
  reg         rob_val_11;
  reg         rob_val_12;
  reg         rob_val_13;
  reg         rob_val_14;
  reg         rob_val_15;
  reg         rob_val_16;
  reg         rob_val_17;
  reg         rob_val_18;
  reg         rob_val_19;
  reg         rob_val_20;
  reg         rob_val_21;
  reg         rob_val_22;
  reg         rob_val_23;
  reg         rob_val_24;
  reg         rob_val_25;
  reg         rob_val_26;
  reg         rob_val_27;
  reg         rob_val_28;
  reg         rob_val_29;
  reg         rob_val_30;
  reg         rob_val_31;
  reg         rob_bsy_0;
  reg         rob_bsy_1;
  reg         rob_bsy_2;
  reg         rob_bsy_3;
  reg         rob_bsy_4;
  reg         rob_bsy_5;
  reg         rob_bsy_6;
  reg         rob_bsy_7;
  reg         rob_bsy_8;
  reg         rob_bsy_9;
  reg         rob_bsy_10;
  reg         rob_bsy_11;
  reg         rob_bsy_12;
  reg         rob_bsy_13;
  reg         rob_bsy_14;
  reg         rob_bsy_15;
  reg         rob_bsy_16;
  reg         rob_bsy_17;
  reg         rob_bsy_18;
  reg         rob_bsy_19;
  reg         rob_bsy_20;
  reg         rob_bsy_21;
  reg         rob_bsy_22;
  reg         rob_bsy_23;
  reg         rob_bsy_24;
  reg         rob_bsy_25;
  reg         rob_bsy_26;
  reg         rob_bsy_27;
  reg         rob_bsy_28;
  reg         rob_bsy_29;
  reg         rob_bsy_30;
  reg         rob_bsy_31;
  reg         rob_unsafe_0;
  reg         rob_unsafe_1;
  reg         rob_unsafe_2;
  reg         rob_unsafe_3;
  reg         rob_unsafe_4;
  reg         rob_unsafe_5;
  reg         rob_unsafe_6;
  reg         rob_unsafe_7;
  reg         rob_unsafe_8;
  reg         rob_unsafe_9;
  reg         rob_unsafe_10;
  reg         rob_unsafe_11;
  reg         rob_unsafe_12;
  reg         rob_unsafe_13;
  reg         rob_unsafe_14;
  reg         rob_unsafe_15;
  reg         rob_unsafe_16;
  reg         rob_unsafe_17;
  reg         rob_unsafe_18;
  reg         rob_unsafe_19;
  reg         rob_unsafe_20;
  reg         rob_unsafe_21;
  reg         rob_unsafe_22;
  reg         rob_unsafe_23;
  reg         rob_unsafe_24;
  reg         rob_unsafe_25;
  reg         rob_unsafe_26;
  reg         rob_unsafe_27;
  reg         rob_unsafe_28;
  reg         rob_unsafe_29;
  reg         rob_unsafe_30;
  reg         rob_unsafe_31;
  reg  [6:0]  rob_uop_0_uopc;
  reg         rob_uop_0_is_rvc;
  reg         rob_uop_0_is_br;
  reg         rob_uop_0_is_jalr;
  reg         rob_uop_0_is_jal;
  reg  [19:0] rob_uop_0_br_mask;
  reg  [5:0]  rob_uop_0_ftq_idx;
  reg         rob_uop_0_edge_inst;
  reg  [5:0]  rob_uop_0_pc_lob;
  reg  [6:0]  rob_uop_0_pdst;
  reg  [6:0]  rob_uop_0_stale_pdst;
  reg         rob_uop_0_is_fencei;
  reg         rob_uop_0_uses_ldq;
  reg         rob_uop_0_uses_stq;
  reg         rob_uop_0_is_sys_pc2epc;
  reg         rob_uop_0_flush_on_commit;
  reg  [5:0]  rob_uop_0_ldst;
  reg         rob_uop_0_ldst_val;
  reg  [1:0]  rob_uop_0_dst_rtype;
  reg         rob_uop_0_fp_val;
  reg  [1:0]  rob_uop_0_debug_fsrc;
  reg  [6:0]  rob_uop_1_uopc;
  reg         rob_uop_1_is_rvc;
  reg         rob_uop_1_is_br;
  reg         rob_uop_1_is_jalr;
  reg         rob_uop_1_is_jal;
  reg  [19:0] rob_uop_1_br_mask;
  reg  [5:0]  rob_uop_1_ftq_idx;
  reg         rob_uop_1_edge_inst;
  reg  [5:0]  rob_uop_1_pc_lob;
  reg  [6:0]  rob_uop_1_pdst;
  reg  [6:0]  rob_uop_1_stale_pdst;
  reg         rob_uop_1_is_fencei;
  reg         rob_uop_1_uses_ldq;
  reg         rob_uop_1_uses_stq;
  reg         rob_uop_1_is_sys_pc2epc;
  reg         rob_uop_1_flush_on_commit;
  reg  [5:0]  rob_uop_1_ldst;
  reg         rob_uop_1_ldst_val;
  reg  [1:0]  rob_uop_1_dst_rtype;
  reg         rob_uop_1_fp_val;
  reg  [1:0]  rob_uop_1_debug_fsrc;
  reg  [6:0]  rob_uop_2_uopc;
  reg         rob_uop_2_is_rvc;
  reg         rob_uop_2_is_br;
  reg         rob_uop_2_is_jalr;
  reg         rob_uop_2_is_jal;
  reg  [19:0] rob_uop_2_br_mask;
  reg  [5:0]  rob_uop_2_ftq_idx;
  reg         rob_uop_2_edge_inst;
  reg  [5:0]  rob_uop_2_pc_lob;
  reg  [6:0]  rob_uop_2_pdst;
  reg  [6:0]  rob_uop_2_stale_pdst;
  reg         rob_uop_2_is_fencei;
  reg         rob_uop_2_uses_ldq;
  reg         rob_uop_2_uses_stq;
  reg         rob_uop_2_is_sys_pc2epc;
  reg         rob_uop_2_flush_on_commit;
  reg  [5:0]  rob_uop_2_ldst;
  reg         rob_uop_2_ldst_val;
  reg  [1:0]  rob_uop_2_dst_rtype;
  reg         rob_uop_2_fp_val;
  reg  [1:0]  rob_uop_2_debug_fsrc;
  reg  [6:0]  rob_uop_3_uopc;
  reg         rob_uop_3_is_rvc;
  reg         rob_uop_3_is_br;
  reg         rob_uop_3_is_jalr;
  reg         rob_uop_3_is_jal;
  reg  [19:0] rob_uop_3_br_mask;
  reg  [5:0]  rob_uop_3_ftq_idx;
  reg         rob_uop_3_edge_inst;
  reg  [5:0]  rob_uop_3_pc_lob;
  reg  [6:0]  rob_uop_3_pdst;
  reg  [6:0]  rob_uop_3_stale_pdst;
  reg         rob_uop_3_is_fencei;
  reg         rob_uop_3_uses_ldq;
  reg         rob_uop_3_uses_stq;
  reg         rob_uop_3_is_sys_pc2epc;
  reg         rob_uop_3_flush_on_commit;
  reg  [5:0]  rob_uop_3_ldst;
  reg         rob_uop_3_ldst_val;
  reg  [1:0]  rob_uop_3_dst_rtype;
  reg         rob_uop_3_fp_val;
  reg  [1:0]  rob_uop_3_debug_fsrc;
  reg  [6:0]  rob_uop_4_uopc;
  reg         rob_uop_4_is_rvc;
  reg         rob_uop_4_is_br;
  reg         rob_uop_4_is_jalr;
  reg         rob_uop_4_is_jal;
  reg  [19:0] rob_uop_4_br_mask;
  reg  [5:0]  rob_uop_4_ftq_idx;
  reg         rob_uop_4_edge_inst;
  reg  [5:0]  rob_uop_4_pc_lob;
  reg  [6:0]  rob_uop_4_pdst;
  reg  [6:0]  rob_uop_4_stale_pdst;
  reg         rob_uop_4_is_fencei;
  reg         rob_uop_4_uses_ldq;
  reg         rob_uop_4_uses_stq;
  reg         rob_uop_4_is_sys_pc2epc;
  reg         rob_uop_4_flush_on_commit;
  reg  [5:0]  rob_uop_4_ldst;
  reg         rob_uop_4_ldst_val;
  reg  [1:0]  rob_uop_4_dst_rtype;
  reg         rob_uop_4_fp_val;
  reg  [1:0]  rob_uop_4_debug_fsrc;
  reg  [6:0]  rob_uop_5_uopc;
  reg         rob_uop_5_is_rvc;
  reg         rob_uop_5_is_br;
  reg         rob_uop_5_is_jalr;
  reg         rob_uop_5_is_jal;
  reg  [19:0] rob_uop_5_br_mask;
  reg  [5:0]  rob_uop_5_ftq_idx;
  reg         rob_uop_5_edge_inst;
  reg  [5:0]  rob_uop_5_pc_lob;
  reg  [6:0]  rob_uop_5_pdst;
  reg  [6:0]  rob_uop_5_stale_pdst;
  reg         rob_uop_5_is_fencei;
  reg         rob_uop_5_uses_ldq;
  reg         rob_uop_5_uses_stq;
  reg         rob_uop_5_is_sys_pc2epc;
  reg         rob_uop_5_flush_on_commit;
  reg  [5:0]  rob_uop_5_ldst;
  reg         rob_uop_5_ldst_val;
  reg  [1:0]  rob_uop_5_dst_rtype;
  reg         rob_uop_5_fp_val;
  reg  [1:0]  rob_uop_5_debug_fsrc;
  reg  [6:0]  rob_uop_6_uopc;
  reg         rob_uop_6_is_rvc;
  reg         rob_uop_6_is_br;
  reg         rob_uop_6_is_jalr;
  reg         rob_uop_6_is_jal;
  reg  [19:0] rob_uop_6_br_mask;
  reg  [5:0]  rob_uop_6_ftq_idx;
  reg         rob_uop_6_edge_inst;
  reg  [5:0]  rob_uop_6_pc_lob;
  reg  [6:0]  rob_uop_6_pdst;
  reg  [6:0]  rob_uop_6_stale_pdst;
  reg         rob_uop_6_is_fencei;
  reg         rob_uop_6_uses_ldq;
  reg         rob_uop_6_uses_stq;
  reg         rob_uop_6_is_sys_pc2epc;
  reg         rob_uop_6_flush_on_commit;
  reg  [5:0]  rob_uop_6_ldst;
  reg         rob_uop_6_ldst_val;
  reg  [1:0]  rob_uop_6_dst_rtype;
  reg         rob_uop_6_fp_val;
  reg  [1:0]  rob_uop_6_debug_fsrc;
  reg  [6:0]  rob_uop_7_uopc;
  reg         rob_uop_7_is_rvc;
  reg         rob_uop_7_is_br;
  reg         rob_uop_7_is_jalr;
  reg         rob_uop_7_is_jal;
  reg  [19:0] rob_uop_7_br_mask;
  reg  [5:0]  rob_uop_7_ftq_idx;
  reg         rob_uop_7_edge_inst;
  reg  [5:0]  rob_uop_7_pc_lob;
  reg  [6:0]  rob_uop_7_pdst;
  reg  [6:0]  rob_uop_7_stale_pdst;
  reg         rob_uop_7_is_fencei;
  reg         rob_uop_7_uses_ldq;
  reg         rob_uop_7_uses_stq;
  reg         rob_uop_7_is_sys_pc2epc;
  reg         rob_uop_7_flush_on_commit;
  reg  [5:0]  rob_uop_7_ldst;
  reg         rob_uop_7_ldst_val;
  reg  [1:0]  rob_uop_7_dst_rtype;
  reg         rob_uop_7_fp_val;
  reg  [1:0]  rob_uop_7_debug_fsrc;
  reg  [6:0]  rob_uop_8_uopc;
  reg         rob_uop_8_is_rvc;
  reg         rob_uop_8_is_br;
  reg         rob_uop_8_is_jalr;
  reg         rob_uop_8_is_jal;
  reg  [19:0] rob_uop_8_br_mask;
  reg  [5:0]  rob_uop_8_ftq_idx;
  reg         rob_uop_8_edge_inst;
  reg  [5:0]  rob_uop_8_pc_lob;
  reg  [6:0]  rob_uop_8_pdst;
  reg  [6:0]  rob_uop_8_stale_pdst;
  reg         rob_uop_8_is_fencei;
  reg         rob_uop_8_uses_ldq;
  reg         rob_uop_8_uses_stq;
  reg         rob_uop_8_is_sys_pc2epc;
  reg         rob_uop_8_flush_on_commit;
  reg  [5:0]  rob_uop_8_ldst;
  reg         rob_uop_8_ldst_val;
  reg  [1:0]  rob_uop_8_dst_rtype;
  reg         rob_uop_8_fp_val;
  reg  [1:0]  rob_uop_8_debug_fsrc;
  reg  [6:0]  rob_uop_9_uopc;
  reg         rob_uop_9_is_rvc;
  reg         rob_uop_9_is_br;
  reg         rob_uop_9_is_jalr;
  reg         rob_uop_9_is_jal;
  reg  [19:0] rob_uop_9_br_mask;
  reg  [5:0]  rob_uop_9_ftq_idx;
  reg         rob_uop_9_edge_inst;
  reg  [5:0]  rob_uop_9_pc_lob;
  reg  [6:0]  rob_uop_9_pdst;
  reg  [6:0]  rob_uop_9_stale_pdst;
  reg         rob_uop_9_is_fencei;
  reg         rob_uop_9_uses_ldq;
  reg         rob_uop_9_uses_stq;
  reg         rob_uop_9_is_sys_pc2epc;
  reg         rob_uop_9_flush_on_commit;
  reg  [5:0]  rob_uop_9_ldst;
  reg         rob_uop_9_ldst_val;
  reg  [1:0]  rob_uop_9_dst_rtype;
  reg         rob_uop_9_fp_val;
  reg  [1:0]  rob_uop_9_debug_fsrc;
  reg  [6:0]  rob_uop_10_uopc;
  reg         rob_uop_10_is_rvc;
  reg         rob_uop_10_is_br;
  reg         rob_uop_10_is_jalr;
  reg         rob_uop_10_is_jal;
  reg  [19:0] rob_uop_10_br_mask;
  reg  [5:0]  rob_uop_10_ftq_idx;
  reg         rob_uop_10_edge_inst;
  reg  [5:0]  rob_uop_10_pc_lob;
  reg  [6:0]  rob_uop_10_pdst;
  reg  [6:0]  rob_uop_10_stale_pdst;
  reg         rob_uop_10_is_fencei;
  reg         rob_uop_10_uses_ldq;
  reg         rob_uop_10_uses_stq;
  reg         rob_uop_10_is_sys_pc2epc;
  reg         rob_uop_10_flush_on_commit;
  reg  [5:0]  rob_uop_10_ldst;
  reg         rob_uop_10_ldst_val;
  reg  [1:0]  rob_uop_10_dst_rtype;
  reg         rob_uop_10_fp_val;
  reg  [1:0]  rob_uop_10_debug_fsrc;
  reg  [6:0]  rob_uop_11_uopc;
  reg         rob_uop_11_is_rvc;
  reg         rob_uop_11_is_br;
  reg         rob_uop_11_is_jalr;
  reg         rob_uop_11_is_jal;
  reg  [19:0] rob_uop_11_br_mask;
  reg  [5:0]  rob_uop_11_ftq_idx;
  reg         rob_uop_11_edge_inst;
  reg  [5:0]  rob_uop_11_pc_lob;
  reg  [6:0]  rob_uop_11_pdst;
  reg  [6:0]  rob_uop_11_stale_pdst;
  reg         rob_uop_11_is_fencei;
  reg         rob_uop_11_uses_ldq;
  reg         rob_uop_11_uses_stq;
  reg         rob_uop_11_is_sys_pc2epc;
  reg         rob_uop_11_flush_on_commit;
  reg  [5:0]  rob_uop_11_ldst;
  reg         rob_uop_11_ldst_val;
  reg  [1:0]  rob_uop_11_dst_rtype;
  reg         rob_uop_11_fp_val;
  reg  [1:0]  rob_uop_11_debug_fsrc;
  reg  [6:0]  rob_uop_12_uopc;
  reg         rob_uop_12_is_rvc;
  reg         rob_uop_12_is_br;
  reg         rob_uop_12_is_jalr;
  reg         rob_uop_12_is_jal;
  reg  [19:0] rob_uop_12_br_mask;
  reg  [5:0]  rob_uop_12_ftq_idx;
  reg         rob_uop_12_edge_inst;
  reg  [5:0]  rob_uop_12_pc_lob;
  reg  [6:0]  rob_uop_12_pdst;
  reg  [6:0]  rob_uop_12_stale_pdst;
  reg         rob_uop_12_is_fencei;
  reg         rob_uop_12_uses_ldq;
  reg         rob_uop_12_uses_stq;
  reg         rob_uop_12_is_sys_pc2epc;
  reg         rob_uop_12_flush_on_commit;
  reg  [5:0]  rob_uop_12_ldst;
  reg         rob_uop_12_ldst_val;
  reg  [1:0]  rob_uop_12_dst_rtype;
  reg         rob_uop_12_fp_val;
  reg  [1:0]  rob_uop_12_debug_fsrc;
  reg  [6:0]  rob_uop_13_uopc;
  reg         rob_uop_13_is_rvc;
  reg         rob_uop_13_is_br;
  reg         rob_uop_13_is_jalr;
  reg         rob_uop_13_is_jal;
  reg  [19:0] rob_uop_13_br_mask;
  reg  [5:0]  rob_uop_13_ftq_idx;
  reg         rob_uop_13_edge_inst;
  reg  [5:0]  rob_uop_13_pc_lob;
  reg  [6:0]  rob_uop_13_pdst;
  reg  [6:0]  rob_uop_13_stale_pdst;
  reg         rob_uop_13_is_fencei;
  reg         rob_uop_13_uses_ldq;
  reg         rob_uop_13_uses_stq;
  reg         rob_uop_13_is_sys_pc2epc;
  reg         rob_uop_13_flush_on_commit;
  reg  [5:0]  rob_uop_13_ldst;
  reg         rob_uop_13_ldst_val;
  reg  [1:0]  rob_uop_13_dst_rtype;
  reg         rob_uop_13_fp_val;
  reg  [1:0]  rob_uop_13_debug_fsrc;
  reg  [6:0]  rob_uop_14_uopc;
  reg         rob_uop_14_is_rvc;
  reg         rob_uop_14_is_br;
  reg         rob_uop_14_is_jalr;
  reg         rob_uop_14_is_jal;
  reg  [19:0] rob_uop_14_br_mask;
  reg  [5:0]  rob_uop_14_ftq_idx;
  reg         rob_uop_14_edge_inst;
  reg  [5:0]  rob_uop_14_pc_lob;
  reg  [6:0]  rob_uop_14_pdst;
  reg  [6:0]  rob_uop_14_stale_pdst;
  reg         rob_uop_14_is_fencei;
  reg         rob_uop_14_uses_ldq;
  reg         rob_uop_14_uses_stq;
  reg         rob_uop_14_is_sys_pc2epc;
  reg         rob_uop_14_flush_on_commit;
  reg  [5:0]  rob_uop_14_ldst;
  reg         rob_uop_14_ldst_val;
  reg  [1:0]  rob_uop_14_dst_rtype;
  reg         rob_uop_14_fp_val;
  reg  [1:0]  rob_uop_14_debug_fsrc;
  reg  [6:0]  rob_uop_15_uopc;
  reg         rob_uop_15_is_rvc;
  reg         rob_uop_15_is_br;
  reg         rob_uop_15_is_jalr;
  reg         rob_uop_15_is_jal;
  reg  [19:0] rob_uop_15_br_mask;
  reg  [5:0]  rob_uop_15_ftq_idx;
  reg         rob_uop_15_edge_inst;
  reg  [5:0]  rob_uop_15_pc_lob;
  reg  [6:0]  rob_uop_15_pdst;
  reg  [6:0]  rob_uop_15_stale_pdst;
  reg         rob_uop_15_is_fencei;
  reg         rob_uop_15_uses_ldq;
  reg         rob_uop_15_uses_stq;
  reg         rob_uop_15_is_sys_pc2epc;
  reg         rob_uop_15_flush_on_commit;
  reg  [5:0]  rob_uop_15_ldst;
  reg         rob_uop_15_ldst_val;
  reg  [1:0]  rob_uop_15_dst_rtype;
  reg         rob_uop_15_fp_val;
  reg  [1:0]  rob_uop_15_debug_fsrc;
  reg  [6:0]  rob_uop_16_uopc;
  reg         rob_uop_16_is_rvc;
  reg         rob_uop_16_is_br;
  reg         rob_uop_16_is_jalr;
  reg         rob_uop_16_is_jal;
  reg  [19:0] rob_uop_16_br_mask;
  reg  [5:0]  rob_uop_16_ftq_idx;
  reg         rob_uop_16_edge_inst;
  reg  [5:0]  rob_uop_16_pc_lob;
  reg  [6:0]  rob_uop_16_pdst;
  reg  [6:0]  rob_uop_16_stale_pdst;
  reg         rob_uop_16_is_fencei;
  reg         rob_uop_16_uses_ldq;
  reg         rob_uop_16_uses_stq;
  reg         rob_uop_16_is_sys_pc2epc;
  reg         rob_uop_16_flush_on_commit;
  reg  [5:0]  rob_uop_16_ldst;
  reg         rob_uop_16_ldst_val;
  reg  [1:0]  rob_uop_16_dst_rtype;
  reg         rob_uop_16_fp_val;
  reg  [1:0]  rob_uop_16_debug_fsrc;
  reg  [6:0]  rob_uop_17_uopc;
  reg         rob_uop_17_is_rvc;
  reg         rob_uop_17_is_br;
  reg         rob_uop_17_is_jalr;
  reg         rob_uop_17_is_jal;
  reg  [19:0] rob_uop_17_br_mask;
  reg  [5:0]  rob_uop_17_ftq_idx;
  reg         rob_uop_17_edge_inst;
  reg  [5:0]  rob_uop_17_pc_lob;
  reg  [6:0]  rob_uop_17_pdst;
  reg  [6:0]  rob_uop_17_stale_pdst;
  reg         rob_uop_17_is_fencei;
  reg         rob_uop_17_uses_ldq;
  reg         rob_uop_17_uses_stq;
  reg         rob_uop_17_is_sys_pc2epc;
  reg         rob_uop_17_flush_on_commit;
  reg  [5:0]  rob_uop_17_ldst;
  reg         rob_uop_17_ldst_val;
  reg  [1:0]  rob_uop_17_dst_rtype;
  reg         rob_uop_17_fp_val;
  reg  [1:0]  rob_uop_17_debug_fsrc;
  reg  [6:0]  rob_uop_18_uopc;
  reg         rob_uop_18_is_rvc;
  reg         rob_uop_18_is_br;
  reg         rob_uop_18_is_jalr;
  reg         rob_uop_18_is_jal;
  reg  [19:0] rob_uop_18_br_mask;
  reg  [5:0]  rob_uop_18_ftq_idx;
  reg         rob_uop_18_edge_inst;
  reg  [5:0]  rob_uop_18_pc_lob;
  reg  [6:0]  rob_uop_18_pdst;
  reg  [6:0]  rob_uop_18_stale_pdst;
  reg         rob_uop_18_is_fencei;
  reg         rob_uop_18_uses_ldq;
  reg         rob_uop_18_uses_stq;
  reg         rob_uop_18_is_sys_pc2epc;
  reg         rob_uop_18_flush_on_commit;
  reg  [5:0]  rob_uop_18_ldst;
  reg         rob_uop_18_ldst_val;
  reg  [1:0]  rob_uop_18_dst_rtype;
  reg         rob_uop_18_fp_val;
  reg  [1:0]  rob_uop_18_debug_fsrc;
  reg  [6:0]  rob_uop_19_uopc;
  reg         rob_uop_19_is_rvc;
  reg         rob_uop_19_is_br;
  reg         rob_uop_19_is_jalr;
  reg         rob_uop_19_is_jal;
  reg  [19:0] rob_uop_19_br_mask;
  reg  [5:0]  rob_uop_19_ftq_idx;
  reg         rob_uop_19_edge_inst;
  reg  [5:0]  rob_uop_19_pc_lob;
  reg  [6:0]  rob_uop_19_pdst;
  reg  [6:0]  rob_uop_19_stale_pdst;
  reg         rob_uop_19_is_fencei;
  reg         rob_uop_19_uses_ldq;
  reg         rob_uop_19_uses_stq;
  reg         rob_uop_19_is_sys_pc2epc;
  reg         rob_uop_19_flush_on_commit;
  reg  [5:0]  rob_uop_19_ldst;
  reg         rob_uop_19_ldst_val;
  reg  [1:0]  rob_uop_19_dst_rtype;
  reg         rob_uop_19_fp_val;
  reg  [1:0]  rob_uop_19_debug_fsrc;
  reg  [6:0]  rob_uop_20_uopc;
  reg         rob_uop_20_is_rvc;
  reg         rob_uop_20_is_br;
  reg         rob_uop_20_is_jalr;
  reg         rob_uop_20_is_jal;
  reg  [19:0] rob_uop_20_br_mask;
  reg  [5:0]  rob_uop_20_ftq_idx;
  reg         rob_uop_20_edge_inst;
  reg  [5:0]  rob_uop_20_pc_lob;
  reg  [6:0]  rob_uop_20_pdst;
  reg  [6:0]  rob_uop_20_stale_pdst;
  reg         rob_uop_20_is_fencei;
  reg         rob_uop_20_uses_ldq;
  reg         rob_uop_20_uses_stq;
  reg         rob_uop_20_is_sys_pc2epc;
  reg         rob_uop_20_flush_on_commit;
  reg  [5:0]  rob_uop_20_ldst;
  reg         rob_uop_20_ldst_val;
  reg  [1:0]  rob_uop_20_dst_rtype;
  reg         rob_uop_20_fp_val;
  reg  [1:0]  rob_uop_20_debug_fsrc;
  reg  [6:0]  rob_uop_21_uopc;
  reg         rob_uop_21_is_rvc;
  reg         rob_uop_21_is_br;
  reg         rob_uop_21_is_jalr;
  reg         rob_uop_21_is_jal;
  reg  [19:0] rob_uop_21_br_mask;
  reg  [5:0]  rob_uop_21_ftq_idx;
  reg         rob_uop_21_edge_inst;
  reg  [5:0]  rob_uop_21_pc_lob;
  reg  [6:0]  rob_uop_21_pdst;
  reg  [6:0]  rob_uop_21_stale_pdst;
  reg         rob_uop_21_is_fencei;
  reg         rob_uop_21_uses_ldq;
  reg         rob_uop_21_uses_stq;
  reg         rob_uop_21_is_sys_pc2epc;
  reg         rob_uop_21_flush_on_commit;
  reg  [5:0]  rob_uop_21_ldst;
  reg         rob_uop_21_ldst_val;
  reg  [1:0]  rob_uop_21_dst_rtype;
  reg         rob_uop_21_fp_val;
  reg  [1:0]  rob_uop_21_debug_fsrc;
  reg  [6:0]  rob_uop_22_uopc;
  reg         rob_uop_22_is_rvc;
  reg         rob_uop_22_is_br;
  reg         rob_uop_22_is_jalr;
  reg         rob_uop_22_is_jal;
  reg  [19:0] rob_uop_22_br_mask;
  reg  [5:0]  rob_uop_22_ftq_idx;
  reg         rob_uop_22_edge_inst;
  reg  [5:0]  rob_uop_22_pc_lob;
  reg  [6:0]  rob_uop_22_pdst;
  reg  [6:0]  rob_uop_22_stale_pdst;
  reg         rob_uop_22_is_fencei;
  reg         rob_uop_22_uses_ldq;
  reg         rob_uop_22_uses_stq;
  reg         rob_uop_22_is_sys_pc2epc;
  reg         rob_uop_22_flush_on_commit;
  reg  [5:0]  rob_uop_22_ldst;
  reg         rob_uop_22_ldst_val;
  reg  [1:0]  rob_uop_22_dst_rtype;
  reg         rob_uop_22_fp_val;
  reg  [1:0]  rob_uop_22_debug_fsrc;
  reg  [6:0]  rob_uop_23_uopc;
  reg         rob_uop_23_is_rvc;
  reg         rob_uop_23_is_br;
  reg         rob_uop_23_is_jalr;
  reg         rob_uop_23_is_jal;
  reg  [19:0] rob_uop_23_br_mask;
  reg  [5:0]  rob_uop_23_ftq_idx;
  reg         rob_uop_23_edge_inst;
  reg  [5:0]  rob_uop_23_pc_lob;
  reg  [6:0]  rob_uop_23_pdst;
  reg  [6:0]  rob_uop_23_stale_pdst;
  reg         rob_uop_23_is_fencei;
  reg         rob_uop_23_uses_ldq;
  reg         rob_uop_23_uses_stq;
  reg         rob_uop_23_is_sys_pc2epc;
  reg         rob_uop_23_flush_on_commit;
  reg  [5:0]  rob_uop_23_ldst;
  reg         rob_uop_23_ldst_val;
  reg  [1:0]  rob_uop_23_dst_rtype;
  reg         rob_uop_23_fp_val;
  reg  [1:0]  rob_uop_23_debug_fsrc;
  reg  [6:0]  rob_uop_24_uopc;
  reg         rob_uop_24_is_rvc;
  reg         rob_uop_24_is_br;
  reg         rob_uop_24_is_jalr;
  reg         rob_uop_24_is_jal;
  reg  [19:0] rob_uop_24_br_mask;
  reg  [5:0]  rob_uop_24_ftq_idx;
  reg         rob_uop_24_edge_inst;
  reg  [5:0]  rob_uop_24_pc_lob;
  reg  [6:0]  rob_uop_24_pdst;
  reg  [6:0]  rob_uop_24_stale_pdst;
  reg         rob_uop_24_is_fencei;
  reg         rob_uop_24_uses_ldq;
  reg         rob_uop_24_uses_stq;
  reg         rob_uop_24_is_sys_pc2epc;
  reg         rob_uop_24_flush_on_commit;
  reg  [5:0]  rob_uop_24_ldst;
  reg         rob_uop_24_ldst_val;
  reg  [1:0]  rob_uop_24_dst_rtype;
  reg         rob_uop_24_fp_val;
  reg  [1:0]  rob_uop_24_debug_fsrc;
  reg  [6:0]  rob_uop_25_uopc;
  reg         rob_uop_25_is_rvc;
  reg         rob_uop_25_is_br;
  reg         rob_uop_25_is_jalr;
  reg         rob_uop_25_is_jal;
  reg  [19:0] rob_uop_25_br_mask;
  reg  [5:0]  rob_uop_25_ftq_idx;
  reg         rob_uop_25_edge_inst;
  reg  [5:0]  rob_uop_25_pc_lob;
  reg  [6:0]  rob_uop_25_pdst;
  reg  [6:0]  rob_uop_25_stale_pdst;
  reg         rob_uop_25_is_fencei;
  reg         rob_uop_25_uses_ldq;
  reg         rob_uop_25_uses_stq;
  reg         rob_uop_25_is_sys_pc2epc;
  reg         rob_uop_25_flush_on_commit;
  reg  [5:0]  rob_uop_25_ldst;
  reg         rob_uop_25_ldst_val;
  reg  [1:0]  rob_uop_25_dst_rtype;
  reg         rob_uop_25_fp_val;
  reg  [1:0]  rob_uop_25_debug_fsrc;
  reg  [6:0]  rob_uop_26_uopc;
  reg         rob_uop_26_is_rvc;
  reg         rob_uop_26_is_br;
  reg         rob_uop_26_is_jalr;
  reg         rob_uop_26_is_jal;
  reg  [19:0] rob_uop_26_br_mask;
  reg  [5:0]  rob_uop_26_ftq_idx;
  reg         rob_uop_26_edge_inst;
  reg  [5:0]  rob_uop_26_pc_lob;
  reg  [6:0]  rob_uop_26_pdst;
  reg  [6:0]  rob_uop_26_stale_pdst;
  reg         rob_uop_26_is_fencei;
  reg         rob_uop_26_uses_ldq;
  reg         rob_uop_26_uses_stq;
  reg         rob_uop_26_is_sys_pc2epc;
  reg         rob_uop_26_flush_on_commit;
  reg  [5:0]  rob_uop_26_ldst;
  reg         rob_uop_26_ldst_val;
  reg  [1:0]  rob_uop_26_dst_rtype;
  reg         rob_uop_26_fp_val;
  reg  [1:0]  rob_uop_26_debug_fsrc;
  reg  [6:0]  rob_uop_27_uopc;
  reg         rob_uop_27_is_rvc;
  reg         rob_uop_27_is_br;
  reg         rob_uop_27_is_jalr;
  reg         rob_uop_27_is_jal;
  reg  [19:0] rob_uop_27_br_mask;
  reg  [5:0]  rob_uop_27_ftq_idx;
  reg         rob_uop_27_edge_inst;
  reg  [5:0]  rob_uop_27_pc_lob;
  reg  [6:0]  rob_uop_27_pdst;
  reg  [6:0]  rob_uop_27_stale_pdst;
  reg         rob_uop_27_is_fencei;
  reg         rob_uop_27_uses_ldq;
  reg         rob_uop_27_uses_stq;
  reg         rob_uop_27_is_sys_pc2epc;
  reg         rob_uop_27_flush_on_commit;
  reg  [5:0]  rob_uop_27_ldst;
  reg         rob_uop_27_ldst_val;
  reg  [1:0]  rob_uop_27_dst_rtype;
  reg         rob_uop_27_fp_val;
  reg  [1:0]  rob_uop_27_debug_fsrc;
  reg  [6:0]  rob_uop_28_uopc;
  reg         rob_uop_28_is_rvc;
  reg         rob_uop_28_is_br;
  reg         rob_uop_28_is_jalr;
  reg         rob_uop_28_is_jal;
  reg  [19:0] rob_uop_28_br_mask;
  reg  [5:0]  rob_uop_28_ftq_idx;
  reg         rob_uop_28_edge_inst;
  reg  [5:0]  rob_uop_28_pc_lob;
  reg  [6:0]  rob_uop_28_pdst;
  reg  [6:0]  rob_uop_28_stale_pdst;
  reg         rob_uop_28_is_fencei;
  reg         rob_uop_28_uses_ldq;
  reg         rob_uop_28_uses_stq;
  reg         rob_uop_28_is_sys_pc2epc;
  reg         rob_uop_28_flush_on_commit;
  reg  [5:0]  rob_uop_28_ldst;
  reg         rob_uop_28_ldst_val;
  reg  [1:0]  rob_uop_28_dst_rtype;
  reg         rob_uop_28_fp_val;
  reg  [1:0]  rob_uop_28_debug_fsrc;
  reg  [6:0]  rob_uop_29_uopc;
  reg         rob_uop_29_is_rvc;
  reg         rob_uop_29_is_br;
  reg         rob_uop_29_is_jalr;
  reg         rob_uop_29_is_jal;
  reg  [19:0] rob_uop_29_br_mask;
  reg  [5:0]  rob_uop_29_ftq_idx;
  reg         rob_uop_29_edge_inst;
  reg  [5:0]  rob_uop_29_pc_lob;
  reg  [6:0]  rob_uop_29_pdst;
  reg  [6:0]  rob_uop_29_stale_pdst;
  reg         rob_uop_29_is_fencei;
  reg         rob_uop_29_uses_ldq;
  reg         rob_uop_29_uses_stq;
  reg         rob_uop_29_is_sys_pc2epc;
  reg         rob_uop_29_flush_on_commit;
  reg  [5:0]  rob_uop_29_ldst;
  reg         rob_uop_29_ldst_val;
  reg  [1:0]  rob_uop_29_dst_rtype;
  reg         rob_uop_29_fp_val;
  reg  [1:0]  rob_uop_29_debug_fsrc;
  reg  [6:0]  rob_uop_30_uopc;
  reg         rob_uop_30_is_rvc;
  reg         rob_uop_30_is_br;
  reg         rob_uop_30_is_jalr;
  reg         rob_uop_30_is_jal;
  reg  [19:0] rob_uop_30_br_mask;
  reg  [5:0]  rob_uop_30_ftq_idx;
  reg         rob_uop_30_edge_inst;
  reg  [5:0]  rob_uop_30_pc_lob;
  reg  [6:0]  rob_uop_30_pdst;
  reg  [6:0]  rob_uop_30_stale_pdst;
  reg         rob_uop_30_is_fencei;
  reg         rob_uop_30_uses_ldq;
  reg         rob_uop_30_uses_stq;
  reg         rob_uop_30_is_sys_pc2epc;
  reg         rob_uop_30_flush_on_commit;
  reg  [5:0]  rob_uop_30_ldst;
  reg         rob_uop_30_ldst_val;
  reg  [1:0]  rob_uop_30_dst_rtype;
  reg         rob_uop_30_fp_val;
  reg  [1:0]  rob_uop_30_debug_fsrc;
  reg  [6:0]  rob_uop_31_uopc;
  reg         rob_uop_31_is_rvc;
  reg         rob_uop_31_is_br;
  reg         rob_uop_31_is_jalr;
  reg         rob_uop_31_is_jal;
  reg  [19:0] rob_uop_31_br_mask;
  reg  [5:0]  rob_uop_31_ftq_idx;
  reg         rob_uop_31_edge_inst;
  reg  [5:0]  rob_uop_31_pc_lob;
  reg  [6:0]  rob_uop_31_pdst;
  reg  [6:0]  rob_uop_31_stale_pdst;
  reg         rob_uop_31_is_fencei;
  reg         rob_uop_31_uses_ldq;
  reg         rob_uop_31_uses_stq;
  reg         rob_uop_31_is_sys_pc2epc;
  reg         rob_uop_31_flush_on_commit;
  reg  [5:0]  rob_uop_31_ldst;
  reg         rob_uop_31_ldst_val;
  reg  [1:0]  rob_uop_31_dst_rtype;
  reg         rob_uop_31_fp_val;
  reg  [1:0]  rob_uop_31_debug_fsrc;
  reg         rob_exception_0;
  reg         rob_exception_1;
  reg         rob_exception_2;
  reg         rob_exception_3;
  reg         rob_exception_4;
  reg         rob_exception_5;
  reg         rob_exception_6;
  reg         rob_exception_7;
  reg         rob_exception_8;
  reg         rob_exception_9;
  reg         rob_exception_10;
  reg         rob_exception_11;
  reg         rob_exception_12;
  reg         rob_exception_13;
  reg         rob_exception_14;
  reg         rob_exception_15;
  reg         rob_exception_16;
  reg         rob_exception_17;
  reg         rob_exception_18;
  reg         rob_exception_19;
  reg         rob_exception_20;
  reg         rob_exception_21;
  reg         rob_exception_22;
  reg         rob_exception_23;
  reg         rob_exception_24;
  reg         rob_exception_25;
  reg         rob_exception_26;
  reg         rob_exception_27;
  reg         rob_exception_28;
  reg         rob_exception_29;
  reg         rob_exception_30;
  reg         rob_exception_31;
  reg         rob_predicated_0;
  reg         rob_predicated_1;
  reg         rob_predicated_2;
  reg         rob_predicated_3;
  reg         rob_predicated_4;
  reg         rob_predicated_5;
  reg         rob_predicated_6;
  reg         rob_predicated_7;
  reg         rob_predicated_8;
  reg         rob_predicated_9;
  reg         rob_predicated_10;
  reg         rob_predicated_11;
  reg         rob_predicated_12;
  reg         rob_predicated_13;
  reg         rob_predicated_14;
  reg         rob_predicated_15;
  reg         rob_predicated_16;
  reg         rob_predicated_17;
  reg         rob_predicated_18;
  reg         rob_predicated_19;
  reg         rob_predicated_20;
  reg         rob_predicated_21;
  reg         rob_predicated_22;
  reg         rob_predicated_23;
  reg         rob_predicated_24;
  reg         rob_predicated_25;
  reg         rob_predicated_26;
  reg         rob_predicated_27;
  reg         rob_predicated_28;
  reg         rob_predicated_29;
  reg         rob_predicated_30;
  reg         rob_predicated_31;
  reg         casez_tmp;
  always @(*) begin
    casez (rob_tail)
      5'b00000:
        casez_tmp = rob_val_0;
      5'b00001:
        casez_tmp = rob_val_1;
      5'b00010:
        casez_tmp = rob_val_2;
      5'b00011:
        casez_tmp = rob_val_3;
      5'b00100:
        casez_tmp = rob_val_4;
      5'b00101:
        casez_tmp = rob_val_5;
      5'b00110:
        casez_tmp = rob_val_6;
      5'b00111:
        casez_tmp = rob_val_7;
      5'b01000:
        casez_tmp = rob_val_8;
      5'b01001:
        casez_tmp = rob_val_9;
      5'b01010:
        casez_tmp = rob_val_10;
      5'b01011:
        casez_tmp = rob_val_11;
      5'b01100:
        casez_tmp = rob_val_12;
      5'b01101:
        casez_tmp = rob_val_13;
      5'b01110:
        casez_tmp = rob_val_14;
      5'b01111:
        casez_tmp = rob_val_15;
      5'b10000:
        casez_tmp = rob_val_16;
      5'b10001:
        casez_tmp = rob_val_17;
      5'b10010:
        casez_tmp = rob_val_18;
      5'b10011:
        casez_tmp = rob_val_19;
      5'b10100:
        casez_tmp = rob_val_20;
      5'b10101:
        casez_tmp = rob_val_21;
      5'b10110:
        casez_tmp = rob_val_22;
      5'b10111:
        casez_tmp = rob_val_23;
      5'b11000:
        casez_tmp = rob_val_24;
      5'b11001:
        casez_tmp = rob_val_25;
      5'b11010:
        casez_tmp = rob_val_26;
      5'b11011:
        casez_tmp = rob_val_27;
      5'b11100:
        casez_tmp = rob_val_28;
      5'b11101:
        casez_tmp = rob_val_29;
      5'b11110:
        casez_tmp = rob_val_30;
      default:
        casez_tmp = rob_val_31;
    endcase
  end // always @(*)
  wire        _GEN = io_wb_resps_0_valid & io_wb_resps_0_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_0 = io_wb_resps_1_valid & io_wb_resps_1_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_1 = io_wb_resps_2_valid & io_wb_resps_2_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_2 = io_wb_resps_3_valid & io_wb_resps_3_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_3 = io_wb_resps_4_valid & io_wb_resps_4_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_4 = io_wb_resps_5_valid & io_wb_resps_5_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_5 = io_wb_resps_6_valid & io_wb_resps_6_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_6 = io_wb_resps_7_valid & io_wb_resps_7_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_7 = io_wb_resps_8_valid & io_wb_resps_8_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_8 = io_wb_resps_9_valid & io_wb_resps_9_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_9 = io_lsu_clr_bsy_0_valid & io_lsu_clr_bsy_0_bits[1:0] == 2'h0;
  reg         casez_tmp_0;
  always @(*) begin
    casez (io_lsu_clr_bsy_0_bits[6:2])
      5'b00000:
        casez_tmp_0 = rob_val_0;
      5'b00001:
        casez_tmp_0 = rob_val_1;
      5'b00010:
        casez_tmp_0 = rob_val_2;
      5'b00011:
        casez_tmp_0 = rob_val_3;
      5'b00100:
        casez_tmp_0 = rob_val_4;
      5'b00101:
        casez_tmp_0 = rob_val_5;
      5'b00110:
        casez_tmp_0 = rob_val_6;
      5'b00111:
        casez_tmp_0 = rob_val_7;
      5'b01000:
        casez_tmp_0 = rob_val_8;
      5'b01001:
        casez_tmp_0 = rob_val_9;
      5'b01010:
        casez_tmp_0 = rob_val_10;
      5'b01011:
        casez_tmp_0 = rob_val_11;
      5'b01100:
        casez_tmp_0 = rob_val_12;
      5'b01101:
        casez_tmp_0 = rob_val_13;
      5'b01110:
        casez_tmp_0 = rob_val_14;
      5'b01111:
        casez_tmp_0 = rob_val_15;
      5'b10000:
        casez_tmp_0 = rob_val_16;
      5'b10001:
        casez_tmp_0 = rob_val_17;
      5'b10010:
        casez_tmp_0 = rob_val_18;
      5'b10011:
        casez_tmp_0 = rob_val_19;
      5'b10100:
        casez_tmp_0 = rob_val_20;
      5'b10101:
        casez_tmp_0 = rob_val_21;
      5'b10110:
        casez_tmp_0 = rob_val_22;
      5'b10111:
        casez_tmp_0 = rob_val_23;
      5'b11000:
        casez_tmp_0 = rob_val_24;
      5'b11001:
        casez_tmp_0 = rob_val_25;
      5'b11010:
        casez_tmp_0 = rob_val_26;
      5'b11011:
        casez_tmp_0 = rob_val_27;
      5'b11100:
        casez_tmp_0 = rob_val_28;
      5'b11101:
        casez_tmp_0 = rob_val_29;
      5'b11110:
        casez_tmp_0 = rob_val_30;
      default:
        casez_tmp_0 = rob_val_31;
    endcase
  end // always @(*)
  reg         casez_tmp_1;
  always @(*) begin
    casez (io_lsu_clr_bsy_0_bits[6:2])
      5'b00000:
        casez_tmp_1 = rob_bsy_0;
      5'b00001:
        casez_tmp_1 = rob_bsy_1;
      5'b00010:
        casez_tmp_1 = rob_bsy_2;
      5'b00011:
        casez_tmp_1 = rob_bsy_3;
      5'b00100:
        casez_tmp_1 = rob_bsy_4;
      5'b00101:
        casez_tmp_1 = rob_bsy_5;
      5'b00110:
        casez_tmp_1 = rob_bsy_6;
      5'b00111:
        casez_tmp_1 = rob_bsy_7;
      5'b01000:
        casez_tmp_1 = rob_bsy_8;
      5'b01001:
        casez_tmp_1 = rob_bsy_9;
      5'b01010:
        casez_tmp_1 = rob_bsy_10;
      5'b01011:
        casez_tmp_1 = rob_bsy_11;
      5'b01100:
        casez_tmp_1 = rob_bsy_12;
      5'b01101:
        casez_tmp_1 = rob_bsy_13;
      5'b01110:
        casez_tmp_1 = rob_bsy_14;
      5'b01111:
        casez_tmp_1 = rob_bsy_15;
      5'b10000:
        casez_tmp_1 = rob_bsy_16;
      5'b10001:
        casez_tmp_1 = rob_bsy_17;
      5'b10010:
        casez_tmp_1 = rob_bsy_18;
      5'b10011:
        casez_tmp_1 = rob_bsy_19;
      5'b10100:
        casez_tmp_1 = rob_bsy_20;
      5'b10101:
        casez_tmp_1 = rob_bsy_21;
      5'b10110:
        casez_tmp_1 = rob_bsy_22;
      5'b10111:
        casez_tmp_1 = rob_bsy_23;
      5'b11000:
        casez_tmp_1 = rob_bsy_24;
      5'b11001:
        casez_tmp_1 = rob_bsy_25;
      5'b11010:
        casez_tmp_1 = rob_bsy_26;
      5'b11011:
        casez_tmp_1 = rob_bsy_27;
      5'b11100:
        casez_tmp_1 = rob_bsy_28;
      5'b11101:
        casez_tmp_1 = rob_bsy_29;
      5'b11110:
        casez_tmp_1 = rob_bsy_30;
      default:
        casez_tmp_1 = rob_bsy_31;
    endcase
  end // always @(*)
  wire        _GEN_10 = io_lsu_clr_bsy_1_valid & io_lsu_clr_bsy_1_bits[1:0] == 2'h0;
  reg         casez_tmp_2;
  always @(*) begin
    casez (io_lsu_clr_bsy_1_bits[6:2])
      5'b00000:
        casez_tmp_2 = rob_val_0;
      5'b00001:
        casez_tmp_2 = rob_val_1;
      5'b00010:
        casez_tmp_2 = rob_val_2;
      5'b00011:
        casez_tmp_2 = rob_val_3;
      5'b00100:
        casez_tmp_2 = rob_val_4;
      5'b00101:
        casez_tmp_2 = rob_val_5;
      5'b00110:
        casez_tmp_2 = rob_val_6;
      5'b00111:
        casez_tmp_2 = rob_val_7;
      5'b01000:
        casez_tmp_2 = rob_val_8;
      5'b01001:
        casez_tmp_2 = rob_val_9;
      5'b01010:
        casez_tmp_2 = rob_val_10;
      5'b01011:
        casez_tmp_2 = rob_val_11;
      5'b01100:
        casez_tmp_2 = rob_val_12;
      5'b01101:
        casez_tmp_2 = rob_val_13;
      5'b01110:
        casez_tmp_2 = rob_val_14;
      5'b01111:
        casez_tmp_2 = rob_val_15;
      5'b10000:
        casez_tmp_2 = rob_val_16;
      5'b10001:
        casez_tmp_2 = rob_val_17;
      5'b10010:
        casez_tmp_2 = rob_val_18;
      5'b10011:
        casez_tmp_2 = rob_val_19;
      5'b10100:
        casez_tmp_2 = rob_val_20;
      5'b10101:
        casez_tmp_2 = rob_val_21;
      5'b10110:
        casez_tmp_2 = rob_val_22;
      5'b10111:
        casez_tmp_2 = rob_val_23;
      5'b11000:
        casez_tmp_2 = rob_val_24;
      5'b11001:
        casez_tmp_2 = rob_val_25;
      5'b11010:
        casez_tmp_2 = rob_val_26;
      5'b11011:
        casez_tmp_2 = rob_val_27;
      5'b11100:
        casez_tmp_2 = rob_val_28;
      5'b11101:
        casez_tmp_2 = rob_val_29;
      5'b11110:
        casez_tmp_2 = rob_val_30;
      default:
        casez_tmp_2 = rob_val_31;
    endcase
  end // always @(*)
  reg         casez_tmp_3;
  always @(*) begin
    casez (io_lsu_clr_bsy_1_bits[6:2])
      5'b00000:
        casez_tmp_3 = rob_bsy_0;
      5'b00001:
        casez_tmp_3 = rob_bsy_1;
      5'b00010:
        casez_tmp_3 = rob_bsy_2;
      5'b00011:
        casez_tmp_3 = rob_bsy_3;
      5'b00100:
        casez_tmp_3 = rob_bsy_4;
      5'b00101:
        casez_tmp_3 = rob_bsy_5;
      5'b00110:
        casez_tmp_3 = rob_bsy_6;
      5'b00111:
        casez_tmp_3 = rob_bsy_7;
      5'b01000:
        casez_tmp_3 = rob_bsy_8;
      5'b01001:
        casez_tmp_3 = rob_bsy_9;
      5'b01010:
        casez_tmp_3 = rob_bsy_10;
      5'b01011:
        casez_tmp_3 = rob_bsy_11;
      5'b01100:
        casez_tmp_3 = rob_bsy_12;
      5'b01101:
        casez_tmp_3 = rob_bsy_13;
      5'b01110:
        casez_tmp_3 = rob_bsy_14;
      5'b01111:
        casez_tmp_3 = rob_bsy_15;
      5'b10000:
        casez_tmp_3 = rob_bsy_16;
      5'b10001:
        casez_tmp_3 = rob_bsy_17;
      5'b10010:
        casez_tmp_3 = rob_bsy_18;
      5'b10011:
        casez_tmp_3 = rob_bsy_19;
      5'b10100:
        casez_tmp_3 = rob_bsy_20;
      5'b10101:
        casez_tmp_3 = rob_bsy_21;
      5'b10110:
        casez_tmp_3 = rob_bsy_22;
      5'b10111:
        casez_tmp_3 = rob_bsy_23;
      5'b11000:
        casez_tmp_3 = rob_bsy_24;
      5'b11001:
        casez_tmp_3 = rob_bsy_25;
      5'b11010:
        casez_tmp_3 = rob_bsy_26;
      5'b11011:
        casez_tmp_3 = rob_bsy_27;
      5'b11100:
        casez_tmp_3 = rob_bsy_28;
      5'b11101:
        casez_tmp_3 = rob_bsy_29;
      5'b11110:
        casez_tmp_3 = rob_bsy_30;
      default:
        casez_tmp_3 = rob_bsy_31;
    endcase
  end // always @(*)
  wire        _GEN_11 = io_lsu_clr_bsy_2_valid & io_lsu_clr_bsy_2_bits[1:0] == 2'h0;
  reg         casez_tmp_4;
  always @(*) begin
    casez (io_lsu_clr_bsy_2_bits[6:2])
      5'b00000:
        casez_tmp_4 = rob_val_0;
      5'b00001:
        casez_tmp_4 = rob_val_1;
      5'b00010:
        casez_tmp_4 = rob_val_2;
      5'b00011:
        casez_tmp_4 = rob_val_3;
      5'b00100:
        casez_tmp_4 = rob_val_4;
      5'b00101:
        casez_tmp_4 = rob_val_5;
      5'b00110:
        casez_tmp_4 = rob_val_6;
      5'b00111:
        casez_tmp_4 = rob_val_7;
      5'b01000:
        casez_tmp_4 = rob_val_8;
      5'b01001:
        casez_tmp_4 = rob_val_9;
      5'b01010:
        casez_tmp_4 = rob_val_10;
      5'b01011:
        casez_tmp_4 = rob_val_11;
      5'b01100:
        casez_tmp_4 = rob_val_12;
      5'b01101:
        casez_tmp_4 = rob_val_13;
      5'b01110:
        casez_tmp_4 = rob_val_14;
      5'b01111:
        casez_tmp_4 = rob_val_15;
      5'b10000:
        casez_tmp_4 = rob_val_16;
      5'b10001:
        casez_tmp_4 = rob_val_17;
      5'b10010:
        casez_tmp_4 = rob_val_18;
      5'b10011:
        casez_tmp_4 = rob_val_19;
      5'b10100:
        casez_tmp_4 = rob_val_20;
      5'b10101:
        casez_tmp_4 = rob_val_21;
      5'b10110:
        casez_tmp_4 = rob_val_22;
      5'b10111:
        casez_tmp_4 = rob_val_23;
      5'b11000:
        casez_tmp_4 = rob_val_24;
      5'b11001:
        casez_tmp_4 = rob_val_25;
      5'b11010:
        casez_tmp_4 = rob_val_26;
      5'b11011:
        casez_tmp_4 = rob_val_27;
      5'b11100:
        casez_tmp_4 = rob_val_28;
      5'b11101:
        casez_tmp_4 = rob_val_29;
      5'b11110:
        casez_tmp_4 = rob_val_30;
      default:
        casez_tmp_4 = rob_val_31;
    endcase
  end // always @(*)
  reg         casez_tmp_5;
  always @(*) begin
    casez (io_lsu_clr_bsy_2_bits[6:2])
      5'b00000:
        casez_tmp_5 = rob_bsy_0;
      5'b00001:
        casez_tmp_5 = rob_bsy_1;
      5'b00010:
        casez_tmp_5 = rob_bsy_2;
      5'b00011:
        casez_tmp_5 = rob_bsy_3;
      5'b00100:
        casez_tmp_5 = rob_bsy_4;
      5'b00101:
        casez_tmp_5 = rob_bsy_5;
      5'b00110:
        casez_tmp_5 = rob_bsy_6;
      5'b00111:
        casez_tmp_5 = rob_bsy_7;
      5'b01000:
        casez_tmp_5 = rob_bsy_8;
      5'b01001:
        casez_tmp_5 = rob_bsy_9;
      5'b01010:
        casez_tmp_5 = rob_bsy_10;
      5'b01011:
        casez_tmp_5 = rob_bsy_11;
      5'b01100:
        casez_tmp_5 = rob_bsy_12;
      5'b01101:
        casez_tmp_5 = rob_bsy_13;
      5'b01110:
        casez_tmp_5 = rob_bsy_14;
      5'b01111:
        casez_tmp_5 = rob_bsy_15;
      5'b10000:
        casez_tmp_5 = rob_bsy_16;
      5'b10001:
        casez_tmp_5 = rob_bsy_17;
      5'b10010:
        casez_tmp_5 = rob_bsy_18;
      5'b10011:
        casez_tmp_5 = rob_bsy_19;
      5'b10100:
        casez_tmp_5 = rob_bsy_20;
      5'b10101:
        casez_tmp_5 = rob_bsy_21;
      5'b10110:
        casez_tmp_5 = rob_bsy_22;
      5'b10111:
        casez_tmp_5 = rob_bsy_23;
      5'b11000:
        casez_tmp_5 = rob_bsy_24;
      5'b11001:
        casez_tmp_5 = rob_bsy_25;
      5'b11010:
        casez_tmp_5 = rob_bsy_26;
      5'b11011:
        casez_tmp_5 = rob_bsy_27;
      5'b11100:
        casez_tmp_5 = rob_bsy_28;
      5'b11101:
        casez_tmp_5 = rob_bsy_29;
      5'b11110:
        casez_tmp_5 = rob_bsy_30;
      default:
        casez_tmp_5 = rob_bsy_31;
    endcase
  end // always @(*)
  wire        _GEN_12 = io_lxcpt_valid & io_lxcpt_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_13 = io_lxcpt_bits_cause != 5'h10;
  wire        _GEN_14 = _GEN_12 & _GEN_13 & ~reset;
  reg         casez_tmp_6;
  always @(*) begin
    casez (io_lxcpt_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_6 = rob_unsafe_0;
      5'b00001:
        casez_tmp_6 = rob_unsafe_1;
      5'b00010:
        casez_tmp_6 = rob_unsafe_2;
      5'b00011:
        casez_tmp_6 = rob_unsafe_3;
      5'b00100:
        casez_tmp_6 = rob_unsafe_4;
      5'b00101:
        casez_tmp_6 = rob_unsafe_5;
      5'b00110:
        casez_tmp_6 = rob_unsafe_6;
      5'b00111:
        casez_tmp_6 = rob_unsafe_7;
      5'b01000:
        casez_tmp_6 = rob_unsafe_8;
      5'b01001:
        casez_tmp_6 = rob_unsafe_9;
      5'b01010:
        casez_tmp_6 = rob_unsafe_10;
      5'b01011:
        casez_tmp_6 = rob_unsafe_11;
      5'b01100:
        casez_tmp_6 = rob_unsafe_12;
      5'b01101:
        casez_tmp_6 = rob_unsafe_13;
      5'b01110:
        casez_tmp_6 = rob_unsafe_14;
      5'b01111:
        casez_tmp_6 = rob_unsafe_15;
      5'b10000:
        casez_tmp_6 = rob_unsafe_16;
      5'b10001:
        casez_tmp_6 = rob_unsafe_17;
      5'b10010:
        casez_tmp_6 = rob_unsafe_18;
      5'b10011:
        casez_tmp_6 = rob_unsafe_19;
      5'b10100:
        casez_tmp_6 = rob_unsafe_20;
      5'b10101:
        casez_tmp_6 = rob_unsafe_21;
      5'b10110:
        casez_tmp_6 = rob_unsafe_22;
      5'b10111:
        casez_tmp_6 = rob_unsafe_23;
      5'b11000:
        casez_tmp_6 = rob_unsafe_24;
      5'b11001:
        casez_tmp_6 = rob_unsafe_25;
      5'b11010:
        casez_tmp_6 = rob_unsafe_26;
      5'b11011:
        casez_tmp_6 = rob_unsafe_27;
      5'b11100:
        casez_tmp_6 = rob_unsafe_28;
      5'b11101:
        casez_tmp_6 = rob_unsafe_29;
      5'b11110:
        casez_tmp_6 = rob_unsafe_30;
      default:
        casez_tmp_6 = rob_unsafe_31;
    endcase
  end // always @(*)
  reg         casez_tmp_7;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_7 = rob_val_0;
      5'b00001:
        casez_tmp_7 = rob_val_1;
      5'b00010:
        casez_tmp_7 = rob_val_2;
      5'b00011:
        casez_tmp_7 = rob_val_3;
      5'b00100:
        casez_tmp_7 = rob_val_4;
      5'b00101:
        casez_tmp_7 = rob_val_5;
      5'b00110:
        casez_tmp_7 = rob_val_6;
      5'b00111:
        casez_tmp_7 = rob_val_7;
      5'b01000:
        casez_tmp_7 = rob_val_8;
      5'b01001:
        casez_tmp_7 = rob_val_9;
      5'b01010:
        casez_tmp_7 = rob_val_10;
      5'b01011:
        casez_tmp_7 = rob_val_11;
      5'b01100:
        casez_tmp_7 = rob_val_12;
      5'b01101:
        casez_tmp_7 = rob_val_13;
      5'b01110:
        casez_tmp_7 = rob_val_14;
      5'b01111:
        casez_tmp_7 = rob_val_15;
      5'b10000:
        casez_tmp_7 = rob_val_16;
      5'b10001:
        casez_tmp_7 = rob_val_17;
      5'b10010:
        casez_tmp_7 = rob_val_18;
      5'b10011:
        casez_tmp_7 = rob_val_19;
      5'b10100:
        casez_tmp_7 = rob_val_20;
      5'b10101:
        casez_tmp_7 = rob_val_21;
      5'b10110:
        casez_tmp_7 = rob_val_22;
      5'b10111:
        casez_tmp_7 = rob_val_23;
      5'b11000:
        casez_tmp_7 = rob_val_24;
      5'b11001:
        casez_tmp_7 = rob_val_25;
      5'b11010:
        casez_tmp_7 = rob_val_26;
      5'b11011:
        casez_tmp_7 = rob_val_27;
      5'b11100:
        casez_tmp_7 = rob_val_28;
      5'b11101:
        casez_tmp_7 = rob_val_29;
      5'b11110:
        casez_tmp_7 = rob_val_30;
      default:
        casez_tmp_7 = rob_val_31;
    endcase
  end // always @(*)
  reg         casez_tmp_8;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_8 = rob_exception_0;
      5'b00001:
        casez_tmp_8 = rob_exception_1;
      5'b00010:
        casez_tmp_8 = rob_exception_2;
      5'b00011:
        casez_tmp_8 = rob_exception_3;
      5'b00100:
        casez_tmp_8 = rob_exception_4;
      5'b00101:
        casez_tmp_8 = rob_exception_5;
      5'b00110:
        casez_tmp_8 = rob_exception_6;
      5'b00111:
        casez_tmp_8 = rob_exception_7;
      5'b01000:
        casez_tmp_8 = rob_exception_8;
      5'b01001:
        casez_tmp_8 = rob_exception_9;
      5'b01010:
        casez_tmp_8 = rob_exception_10;
      5'b01011:
        casez_tmp_8 = rob_exception_11;
      5'b01100:
        casez_tmp_8 = rob_exception_12;
      5'b01101:
        casez_tmp_8 = rob_exception_13;
      5'b01110:
        casez_tmp_8 = rob_exception_14;
      5'b01111:
        casez_tmp_8 = rob_exception_15;
      5'b10000:
        casez_tmp_8 = rob_exception_16;
      5'b10001:
        casez_tmp_8 = rob_exception_17;
      5'b10010:
        casez_tmp_8 = rob_exception_18;
      5'b10011:
        casez_tmp_8 = rob_exception_19;
      5'b10100:
        casez_tmp_8 = rob_exception_20;
      5'b10101:
        casez_tmp_8 = rob_exception_21;
      5'b10110:
        casez_tmp_8 = rob_exception_22;
      5'b10111:
        casez_tmp_8 = rob_exception_23;
      5'b11000:
        casez_tmp_8 = rob_exception_24;
      5'b11001:
        casez_tmp_8 = rob_exception_25;
      5'b11010:
        casez_tmp_8 = rob_exception_26;
      5'b11011:
        casez_tmp_8 = rob_exception_27;
      5'b11100:
        casez_tmp_8 = rob_exception_28;
      5'b11101:
        casez_tmp_8 = rob_exception_29;
      5'b11110:
        casez_tmp_8 = rob_exception_30;
      default:
        casez_tmp_8 = rob_exception_31;
    endcase
  end // always @(*)
  wire        can_throw_exception_0 = casez_tmp_7 & casez_tmp_8;
  reg         casez_tmp_9;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_9 = rob_bsy_0;
      5'b00001:
        casez_tmp_9 = rob_bsy_1;
      5'b00010:
        casez_tmp_9 = rob_bsy_2;
      5'b00011:
        casez_tmp_9 = rob_bsy_3;
      5'b00100:
        casez_tmp_9 = rob_bsy_4;
      5'b00101:
        casez_tmp_9 = rob_bsy_5;
      5'b00110:
        casez_tmp_9 = rob_bsy_6;
      5'b00111:
        casez_tmp_9 = rob_bsy_7;
      5'b01000:
        casez_tmp_9 = rob_bsy_8;
      5'b01001:
        casez_tmp_9 = rob_bsy_9;
      5'b01010:
        casez_tmp_9 = rob_bsy_10;
      5'b01011:
        casez_tmp_9 = rob_bsy_11;
      5'b01100:
        casez_tmp_9 = rob_bsy_12;
      5'b01101:
        casez_tmp_9 = rob_bsy_13;
      5'b01110:
        casez_tmp_9 = rob_bsy_14;
      5'b01111:
        casez_tmp_9 = rob_bsy_15;
      5'b10000:
        casez_tmp_9 = rob_bsy_16;
      5'b10001:
        casez_tmp_9 = rob_bsy_17;
      5'b10010:
        casez_tmp_9 = rob_bsy_18;
      5'b10011:
        casez_tmp_9 = rob_bsy_19;
      5'b10100:
        casez_tmp_9 = rob_bsy_20;
      5'b10101:
        casez_tmp_9 = rob_bsy_21;
      5'b10110:
        casez_tmp_9 = rob_bsy_22;
      5'b10111:
        casez_tmp_9 = rob_bsy_23;
      5'b11000:
        casez_tmp_9 = rob_bsy_24;
      5'b11001:
        casez_tmp_9 = rob_bsy_25;
      5'b11010:
        casez_tmp_9 = rob_bsy_26;
      5'b11011:
        casez_tmp_9 = rob_bsy_27;
      5'b11100:
        casez_tmp_9 = rob_bsy_28;
      5'b11101:
        casez_tmp_9 = rob_bsy_29;
      5'b11110:
        casez_tmp_9 = rob_bsy_30;
      default:
        casez_tmp_9 = rob_bsy_31;
    endcase
  end // always @(*)
  wire        can_commit_0 = casez_tmp_7 & ~casez_tmp_9 & ~io_csr_stall;
  reg         casez_tmp_10;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_10 = rob_predicated_0;
      5'b00001:
        casez_tmp_10 = rob_predicated_1;
      5'b00010:
        casez_tmp_10 = rob_predicated_2;
      5'b00011:
        casez_tmp_10 = rob_predicated_3;
      5'b00100:
        casez_tmp_10 = rob_predicated_4;
      5'b00101:
        casez_tmp_10 = rob_predicated_5;
      5'b00110:
        casez_tmp_10 = rob_predicated_6;
      5'b00111:
        casez_tmp_10 = rob_predicated_7;
      5'b01000:
        casez_tmp_10 = rob_predicated_8;
      5'b01001:
        casez_tmp_10 = rob_predicated_9;
      5'b01010:
        casez_tmp_10 = rob_predicated_10;
      5'b01011:
        casez_tmp_10 = rob_predicated_11;
      5'b01100:
        casez_tmp_10 = rob_predicated_12;
      5'b01101:
        casez_tmp_10 = rob_predicated_13;
      5'b01110:
        casez_tmp_10 = rob_predicated_14;
      5'b01111:
        casez_tmp_10 = rob_predicated_15;
      5'b10000:
        casez_tmp_10 = rob_predicated_16;
      5'b10001:
        casez_tmp_10 = rob_predicated_17;
      5'b10010:
        casez_tmp_10 = rob_predicated_18;
      5'b10011:
        casez_tmp_10 = rob_predicated_19;
      5'b10100:
        casez_tmp_10 = rob_predicated_20;
      5'b10101:
        casez_tmp_10 = rob_predicated_21;
      5'b10110:
        casez_tmp_10 = rob_predicated_22;
      5'b10111:
        casez_tmp_10 = rob_predicated_23;
      5'b11000:
        casez_tmp_10 = rob_predicated_24;
      5'b11001:
        casez_tmp_10 = rob_predicated_25;
      5'b11010:
        casez_tmp_10 = rob_predicated_26;
      5'b11011:
        casez_tmp_10 = rob_predicated_27;
      5'b11100:
        casez_tmp_10 = rob_predicated_28;
      5'b11101:
        casez_tmp_10 = rob_predicated_29;
      5'b11110:
        casez_tmp_10 = rob_predicated_30;
      default:
        casez_tmp_10 = rob_predicated_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_11;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_11 = rob_uop_0_uopc;
      5'b00001:
        casez_tmp_11 = rob_uop_1_uopc;
      5'b00010:
        casez_tmp_11 = rob_uop_2_uopc;
      5'b00011:
        casez_tmp_11 = rob_uop_3_uopc;
      5'b00100:
        casez_tmp_11 = rob_uop_4_uopc;
      5'b00101:
        casez_tmp_11 = rob_uop_5_uopc;
      5'b00110:
        casez_tmp_11 = rob_uop_6_uopc;
      5'b00111:
        casez_tmp_11 = rob_uop_7_uopc;
      5'b01000:
        casez_tmp_11 = rob_uop_8_uopc;
      5'b01001:
        casez_tmp_11 = rob_uop_9_uopc;
      5'b01010:
        casez_tmp_11 = rob_uop_10_uopc;
      5'b01011:
        casez_tmp_11 = rob_uop_11_uopc;
      5'b01100:
        casez_tmp_11 = rob_uop_12_uopc;
      5'b01101:
        casez_tmp_11 = rob_uop_13_uopc;
      5'b01110:
        casez_tmp_11 = rob_uop_14_uopc;
      5'b01111:
        casez_tmp_11 = rob_uop_15_uopc;
      5'b10000:
        casez_tmp_11 = rob_uop_16_uopc;
      5'b10001:
        casez_tmp_11 = rob_uop_17_uopc;
      5'b10010:
        casez_tmp_11 = rob_uop_18_uopc;
      5'b10011:
        casez_tmp_11 = rob_uop_19_uopc;
      5'b10100:
        casez_tmp_11 = rob_uop_20_uopc;
      5'b10101:
        casez_tmp_11 = rob_uop_21_uopc;
      5'b10110:
        casez_tmp_11 = rob_uop_22_uopc;
      5'b10111:
        casez_tmp_11 = rob_uop_23_uopc;
      5'b11000:
        casez_tmp_11 = rob_uop_24_uopc;
      5'b11001:
        casez_tmp_11 = rob_uop_25_uopc;
      5'b11010:
        casez_tmp_11 = rob_uop_26_uopc;
      5'b11011:
        casez_tmp_11 = rob_uop_27_uopc;
      5'b11100:
        casez_tmp_11 = rob_uop_28_uopc;
      5'b11101:
        casez_tmp_11 = rob_uop_29_uopc;
      5'b11110:
        casez_tmp_11 = rob_uop_30_uopc;
      default:
        casez_tmp_11 = rob_uop_31_uopc;
    endcase
  end // always @(*)
  reg         casez_tmp_12;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_12 = rob_uop_0_is_rvc;
      5'b00001:
        casez_tmp_12 = rob_uop_1_is_rvc;
      5'b00010:
        casez_tmp_12 = rob_uop_2_is_rvc;
      5'b00011:
        casez_tmp_12 = rob_uop_3_is_rvc;
      5'b00100:
        casez_tmp_12 = rob_uop_4_is_rvc;
      5'b00101:
        casez_tmp_12 = rob_uop_5_is_rvc;
      5'b00110:
        casez_tmp_12 = rob_uop_6_is_rvc;
      5'b00111:
        casez_tmp_12 = rob_uop_7_is_rvc;
      5'b01000:
        casez_tmp_12 = rob_uop_8_is_rvc;
      5'b01001:
        casez_tmp_12 = rob_uop_9_is_rvc;
      5'b01010:
        casez_tmp_12 = rob_uop_10_is_rvc;
      5'b01011:
        casez_tmp_12 = rob_uop_11_is_rvc;
      5'b01100:
        casez_tmp_12 = rob_uop_12_is_rvc;
      5'b01101:
        casez_tmp_12 = rob_uop_13_is_rvc;
      5'b01110:
        casez_tmp_12 = rob_uop_14_is_rvc;
      5'b01111:
        casez_tmp_12 = rob_uop_15_is_rvc;
      5'b10000:
        casez_tmp_12 = rob_uop_16_is_rvc;
      5'b10001:
        casez_tmp_12 = rob_uop_17_is_rvc;
      5'b10010:
        casez_tmp_12 = rob_uop_18_is_rvc;
      5'b10011:
        casez_tmp_12 = rob_uop_19_is_rvc;
      5'b10100:
        casez_tmp_12 = rob_uop_20_is_rvc;
      5'b10101:
        casez_tmp_12 = rob_uop_21_is_rvc;
      5'b10110:
        casez_tmp_12 = rob_uop_22_is_rvc;
      5'b10111:
        casez_tmp_12 = rob_uop_23_is_rvc;
      5'b11000:
        casez_tmp_12 = rob_uop_24_is_rvc;
      5'b11001:
        casez_tmp_12 = rob_uop_25_is_rvc;
      5'b11010:
        casez_tmp_12 = rob_uop_26_is_rvc;
      5'b11011:
        casez_tmp_12 = rob_uop_27_is_rvc;
      5'b11100:
        casez_tmp_12 = rob_uop_28_is_rvc;
      5'b11101:
        casez_tmp_12 = rob_uop_29_is_rvc;
      5'b11110:
        casez_tmp_12 = rob_uop_30_is_rvc;
      default:
        casez_tmp_12 = rob_uop_31_is_rvc;
    endcase
  end // always @(*)
  reg         casez_tmp_13;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_13 = rob_uop_0_is_br;
      5'b00001:
        casez_tmp_13 = rob_uop_1_is_br;
      5'b00010:
        casez_tmp_13 = rob_uop_2_is_br;
      5'b00011:
        casez_tmp_13 = rob_uop_3_is_br;
      5'b00100:
        casez_tmp_13 = rob_uop_4_is_br;
      5'b00101:
        casez_tmp_13 = rob_uop_5_is_br;
      5'b00110:
        casez_tmp_13 = rob_uop_6_is_br;
      5'b00111:
        casez_tmp_13 = rob_uop_7_is_br;
      5'b01000:
        casez_tmp_13 = rob_uop_8_is_br;
      5'b01001:
        casez_tmp_13 = rob_uop_9_is_br;
      5'b01010:
        casez_tmp_13 = rob_uop_10_is_br;
      5'b01011:
        casez_tmp_13 = rob_uop_11_is_br;
      5'b01100:
        casez_tmp_13 = rob_uop_12_is_br;
      5'b01101:
        casez_tmp_13 = rob_uop_13_is_br;
      5'b01110:
        casez_tmp_13 = rob_uop_14_is_br;
      5'b01111:
        casez_tmp_13 = rob_uop_15_is_br;
      5'b10000:
        casez_tmp_13 = rob_uop_16_is_br;
      5'b10001:
        casez_tmp_13 = rob_uop_17_is_br;
      5'b10010:
        casez_tmp_13 = rob_uop_18_is_br;
      5'b10011:
        casez_tmp_13 = rob_uop_19_is_br;
      5'b10100:
        casez_tmp_13 = rob_uop_20_is_br;
      5'b10101:
        casez_tmp_13 = rob_uop_21_is_br;
      5'b10110:
        casez_tmp_13 = rob_uop_22_is_br;
      5'b10111:
        casez_tmp_13 = rob_uop_23_is_br;
      5'b11000:
        casez_tmp_13 = rob_uop_24_is_br;
      5'b11001:
        casez_tmp_13 = rob_uop_25_is_br;
      5'b11010:
        casez_tmp_13 = rob_uop_26_is_br;
      5'b11011:
        casez_tmp_13 = rob_uop_27_is_br;
      5'b11100:
        casez_tmp_13 = rob_uop_28_is_br;
      5'b11101:
        casez_tmp_13 = rob_uop_29_is_br;
      5'b11110:
        casez_tmp_13 = rob_uop_30_is_br;
      default:
        casez_tmp_13 = rob_uop_31_is_br;
    endcase
  end // always @(*)
  reg         casez_tmp_14;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_14 = rob_uop_0_is_jalr;
      5'b00001:
        casez_tmp_14 = rob_uop_1_is_jalr;
      5'b00010:
        casez_tmp_14 = rob_uop_2_is_jalr;
      5'b00011:
        casez_tmp_14 = rob_uop_3_is_jalr;
      5'b00100:
        casez_tmp_14 = rob_uop_4_is_jalr;
      5'b00101:
        casez_tmp_14 = rob_uop_5_is_jalr;
      5'b00110:
        casez_tmp_14 = rob_uop_6_is_jalr;
      5'b00111:
        casez_tmp_14 = rob_uop_7_is_jalr;
      5'b01000:
        casez_tmp_14 = rob_uop_8_is_jalr;
      5'b01001:
        casez_tmp_14 = rob_uop_9_is_jalr;
      5'b01010:
        casez_tmp_14 = rob_uop_10_is_jalr;
      5'b01011:
        casez_tmp_14 = rob_uop_11_is_jalr;
      5'b01100:
        casez_tmp_14 = rob_uop_12_is_jalr;
      5'b01101:
        casez_tmp_14 = rob_uop_13_is_jalr;
      5'b01110:
        casez_tmp_14 = rob_uop_14_is_jalr;
      5'b01111:
        casez_tmp_14 = rob_uop_15_is_jalr;
      5'b10000:
        casez_tmp_14 = rob_uop_16_is_jalr;
      5'b10001:
        casez_tmp_14 = rob_uop_17_is_jalr;
      5'b10010:
        casez_tmp_14 = rob_uop_18_is_jalr;
      5'b10011:
        casez_tmp_14 = rob_uop_19_is_jalr;
      5'b10100:
        casez_tmp_14 = rob_uop_20_is_jalr;
      5'b10101:
        casez_tmp_14 = rob_uop_21_is_jalr;
      5'b10110:
        casez_tmp_14 = rob_uop_22_is_jalr;
      5'b10111:
        casez_tmp_14 = rob_uop_23_is_jalr;
      5'b11000:
        casez_tmp_14 = rob_uop_24_is_jalr;
      5'b11001:
        casez_tmp_14 = rob_uop_25_is_jalr;
      5'b11010:
        casez_tmp_14 = rob_uop_26_is_jalr;
      5'b11011:
        casez_tmp_14 = rob_uop_27_is_jalr;
      5'b11100:
        casez_tmp_14 = rob_uop_28_is_jalr;
      5'b11101:
        casez_tmp_14 = rob_uop_29_is_jalr;
      5'b11110:
        casez_tmp_14 = rob_uop_30_is_jalr;
      default:
        casez_tmp_14 = rob_uop_31_is_jalr;
    endcase
  end // always @(*)
  reg         casez_tmp_15;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_15 = rob_uop_0_is_jal;
      5'b00001:
        casez_tmp_15 = rob_uop_1_is_jal;
      5'b00010:
        casez_tmp_15 = rob_uop_2_is_jal;
      5'b00011:
        casez_tmp_15 = rob_uop_3_is_jal;
      5'b00100:
        casez_tmp_15 = rob_uop_4_is_jal;
      5'b00101:
        casez_tmp_15 = rob_uop_5_is_jal;
      5'b00110:
        casez_tmp_15 = rob_uop_6_is_jal;
      5'b00111:
        casez_tmp_15 = rob_uop_7_is_jal;
      5'b01000:
        casez_tmp_15 = rob_uop_8_is_jal;
      5'b01001:
        casez_tmp_15 = rob_uop_9_is_jal;
      5'b01010:
        casez_tmp_15 = rob_uop_10_is_jal;
      5'b01011:
        casez_tmp_15 = rob_uop_11_is_jal;
      5'b01100:
        casez_tmp_15 = rob_uop_12_is_jal;
      5'b01101:
        casez_tmp_15 = rob_uop_13_is_jal;
      5'b01110:
        casez_tmp_15 = rob_uop_14_is_jal;
      5'b01111:
        casez_tmp_15 = rob_uop_15_is_jal;
      5'b10000:
        casez_tmp_15 = rob_uop_16_is_jal;
      5'b10001:
        casez_tmp_15 = rob_uop_17_is_jal;
      5'b10010:
        casez_tmp_15 = rob_uop_18_is_jal;
      5'b10011:
        casez_tmp_15 = rob_uop_19_is_jal;
      5'b10100:
        casez_tmp_15 = rob_uop_20_is_jal;
      5'b10101:
        casez_tmp_15 = rob_uop_21_is_jal;
      5'b10110:
        casez_tmp_15 = rob_uop_22_is_jal;
      5'b10111:
        casez_tmp_15 = rob_uop_23_is_jal;
      5'b11000:
        casez_tmp_15 = rob_uop_24_is_jal;
      5'b11001:
        casez_tmp_15 = rob_uop_25_is_jal;
      5'b11010:
        casez_tmp_15 = rob_uop_26_is_jal;
      5'b11011:
        casez_tmp_15 = rob_uop_27_is_jal;
      5'b11100:
        casez_tmp_15 = rob_uop_28_is_jal;
      5'b11101:
        casez_tmp_15 = rob_uop_29_is_jal;
      5'b11110:
        casez_tmp_15 = rob_uop_30_is_jal;
      default:
        casez_tmp_15 = rob_uop_31_is_jal;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_16;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_16 = rob_uop_0_ftq_idx;
      5'b00001:
        casez_tmp_16 = rob_uop_1_ftq_idx;
      5'b00010:
        casez_tmp_16 = rob_uop_2_ftq_idx;
      5'b00011:
        casez_tmp_16 = rob_uop_3_ftq_idx;
      5'b00100:
        casez_tmp_16 = rob_uop_4_ftq_idx;
      5'b00101:
        casez_tmp_16 = rob_uop_5_ftq_idx;
      5'b00110:
        casez_tmp_16 = rob_uop_6_ftq_idx;
      5'b00111:
        casez_tmp_16 = rob_uop_7_ftq_idx;
      5'b01000:
        casez_tmp_16 = rob_uop_8_ftq_idx;
      5'b01001:
        casez_tmp_16 = rob_uop_9_ftq_idx;
      5'b01010:
        casez_tmp_16 = rob_uop_10_ftq_idx;
      5'b01011:
        casez_tmp_16 = rob_uop_11_ftq_idx;
      5'b01100:
        casez_tmp_16 = rob_uop_12_ftq_idx;
      5'b01101:
        casez_tmp_16 = rob_uop_13_ftq_idx;
      5'b01110:
        casez_tmp_16 = rob_uop_14_ftq_idx;
      5'b01111:
        casez_tmp_16 = rob_uop_15_ftq_idx;
      5'b10000:
        casez_tmp_16 = rob_uop_16_ftq_idx;
      5'b10001:
        casez_tmp_16 = rob_uop_17_ftq_idx;
      5'b10010:
        casez_tmp_16 = rob_uop_18_ftq_idx;
      5'b10011:
        casez_tmp_16 = rob_uop_19_ftq_idx;
      5'b10100:
        casez_tmp_16 = rob_uop_20_ftq_idx;
      5'b10101:
        casez_tmp_16 = rob_uop_21_ftq_idx;
      5'b10110:
        casez_tmp_16 = rob_uop_22_ftq_idx;
      5'b10111:
        casez_tmp_16 = rob_uop_23_ftq_idx;
      5'b11000:
        casez_tmp_16 = rob_uop_24_ftq_idx;
      5'b11001:
        casez_tmp_16 = rob_uop_25_ftq_idx;
      5'b11010:
        casez_tmp_16 = rob_uop_26_ftq_idx;
      5'b11011:
        casez_tmp_16 = rob_uop_27_ftq_idx;
      5'b11100:
        casez_tmp_16 = rob_uop_28_ftq_idx;
      5'b11101:
        casez_tmp_16 = rob_uop_29_ftq_idx;
      5'b11110:
        casez_tmp_16 = rob_uop_30_ftq_idx;
      default:
        casez_tmp_16 = rob_uop_31_ftq_idx;
    endcase
  end // always @(*)
  reg         casez_tmp_17;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_17 = rob_uop_0_edge_inst;
      5'b00001:
        casez_tmp_17 = rob_uop_1_edge_inst;
      5'b00010:
        casez_tmp_17 = rob_uop_2_edge_inst;
      5'b00011:
        casez_tmp_17 = rob_uop_3_edge_inst;
      5'b00100:
        casez_tmp_17 = rob_uop_4_edge_inst;
      5'b00101:
        casez_tmp_17 = rob_uop_5_edge_inst;
      5'b00110:
        casez_tmp_17 = rob_uop_6_edge_inst;
      5'b00111:
        casez_tmp_17 = rob_uop_7_edge_inst;
      5'b01000:
        casez_tmp_17 = rob_uop_8_edge_inst;
      5'b01001:
        casez_tmp_17 = rob_uop_9_edge_inst;
      5'b01010:
        casez_tmp_17 = rob_uop_10_edge_inst;
      5'b01011:
        casez_tmp_17 = rob_uop_11_edge_inst;
      5'b01100:
        casez_tmp_17 = rob_uop_12_edge_inst;
      5'b01101:
        casez_tmp_17 = rob_uop_13_edge_inst;
      5'b01110:
        casez_tmp_17 = rob_uop_14_edge_inst;
      5'b01111:
        casez_tmp_17 = rob_uop_15_edge_inst;
      5'b10000:
        casez_tmp_17 = rob_uop_16_edge_inst;
      5'b10001:
        casez_tmp_17 = rob_uop_17_edge_inst;
      5'b10010:
        casez_tmp_17 = rob_uop_18_edge_inst;
      5'b10011:
        casez_tmp_17 = rob_uop_19_edge_inst;
      5'b10100:
        casez_tmp_17 = rob_uop_20_edge_inst;
      5'b10101:
        casez_tmp_17 = rob_uop_21_edge_inst;
      5'b10110:
        casez_tmp_17 = rob_uop_22_edge_inst;
      5'b10111:
        casez_tmp_17 = rob_uop_23_edge_inst;
      5'b11000:
        casez_tmp_17 = rob_uop_24_edge_inst;
      5'b11001:
        casez_tmp_17 = rob_uop_25_edge_inst;
      5'b11010:
        casez_tmp_17 = rob_uop_26_edge_inst;
      5'b11011:
        casez_tmp_17 = rob_uop_27_edge_inst;
      5'b11100:
        casez_tmp_17 = rob_uop_28_edge_inst;
      5'b11101:
        casez_tmp_17 = rob_uop_29_edge_inst;
      5'b11110:
        casez_tmp_17 = rob_uop_30_edge_inst;
      default:
        casez_tmp_17 = rob_uop_31_edge_inst;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_18;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_18 = rob_uop_0_pc_lob;
      5'b00001:
        casez_tmp_18 = rob_uop_1_pc_lob;
      5'b00010:
        casez_tmp_18 = rob_uop_2_pc_lob;
      5'b00011:
        casez_tmp_18 = rob_uop_3_pc_lob;
      5'b00100:
        casez_tmp_18 = rob_uop_4_pc_lob;
      5'b00101:
        casez_tmp_18 = rob_uop_5_pc_lob;
      5'b00110:
        casez_tmp_18 = rob_uop_6_pc_lob;
      5'b00111:
        casez_tmp_18 = rob_uop_7_pc_lob;
      5'b01000:
        casez_tmp_18 = rob_uop_8_pc_lob;
      5'b01001:
        casez_tmp_18 = rob_uop_9_pc_lob;
      5'b01010:
        casez_tmp_18 = rob_uop_10_pc_lob;
      5'b01011:
        casez_tmp_18 = rob_uop_11_pc_lob;
      5'b01100:
        casez_tmp_18 = rob_uop_12_pc_lob;
      5'b01101:
        casez_tmp_18 = rob_uop_13_pc_lob;
      5'b01110:
        casez_tmp_18 = rob_uop_14_pc_lob;
      5'b01111:
        casez_tmp_18 = rob_uop_15_pc_lob;
      5'b10000:
        casez_tmp_18 = rob_uop_16_pc_lob;
      5'b10001:
        casez_tmp_18 = rob_uop_17_pc_lob;
      5'b10010:
        casez_tmp_18 = rob_uop_18_pc_lob;
      5'b10011:
        casez_tmp_18 = rob_uop_19_pc_lob;
      5'b10100:
        casez_tmp_18 = rob_uop_20_pc_lob;
      5'b10101:
        casez_tmp_18 = rob_uop_21_pc_lob;
      5'b10110:
        casez_tmp_18 = rob_uop_22_pc_lob;
      5'b10111:
        casez_tmp_18 = rob_uop_23_pc_lob;
      5'b11000:
        casez_tmp_18 = rob_uop_24_pc_lob;
      5'b11001:
        casez_tmp_18 = rob_uop_25_pc_lob;
      5'b11010:
        casez_tmp_18 = rob_uop_26_pc_lob;
      5'b11011:
        casez_tmp_18 = rob_uop_27_pc_lob;
      5'b11100:
        casez_tmp_18 = rob_uop_28_pc_lob;
      5'b11101:
        casez_tmp_18 = rob_uop_29_pc_lob;
      5'b11110:
        casez_tmp_18 = rob_uop_30_pc_lob;
      default:
        casez_tmp_18 = rob_uop_31_pc_lob;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_19;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_19 = rob_uop_0_pdst;
      5'b00001:
        casez_tmp_19 = rob_uop_1_pdst;
      5'b00010:
        casez_tmp_19 = rob_uop_2_pdst;
      5'b00011:
        casez_tmp_19 = rob_uop_3_pdst;
      5'b00100:
        casez_tmp_19 = rob_uop_4_pdst;
      5'b00101:
        casez_tmp_19 = rob_uop_5_pdst;
      5'b00110:
        casez_tmp_19 = rob_uop_6_pdst;
      5'b00111:
        casez_tmp_19 = rob_uop_7_pdst;
      5'b01000:
        casez_tmp_19 = rob_uop_8_pdst;
      5'b01001:
        casez_tmp_19 = rob_uop_9_pdst;
      5'b01010:
        casez_tmp_19 = rob_uop_10_pdst;
      5'b01011:
        casez_tmp_19 = rob_uop_11_pdst;
      5'b01100:
        casez_tmp_19 = rob_uop_12_pdst;
      5'b01101:
        casez_tmp_19 = rob_uop_13_pdst;
      5'b01110:
        casez_tmp_19 = rob_uop_14_pdst;
      5'b01111:
        casez_tmp_19 = rob_uop_15_pdst;
      5'b10000:
        casez_tmp_19 = rob_uop_16_pdst;
      5'b10001:
        casez_tmp_19 = rob_uop_17_pdst;
      5'b10010:
        casez_tmp_19 = rob_uop_18_pdst;
      5'b10011:
        casez_tmp_19 = rob_uop_19_pdst;
      5'b10100:
        casez_tmp_19 = rob_uop_20_pdst;
      5'b10101:
        casez_tmp_19 = rob_uop_21_pdst;
      5'b10110:
        casez_tmp_19 = rob_uop_22_pdst;
      5'b10111:
        casez_tmp_19 = rob_uop_23_pdst;
      5'b11000:
        casez_tmp_19 = rob_uop_24_pdst;
      5'b11001:
        casez_tmp_19 = rob_uop_25_pdst;
      5'b11010:
        casez_tmp_19 = rob_uop_26_pdst;
      5'b11011:
        casez_tmp_19 = rob_uop_27_pdst;
      5'b11100:
        casez_tmp_19 = rob_uop_28_pdst;
      5'b11101:
        casez_tmp_19 = rob_uop_29_pdst;
      5'b11110:
        casez_tmp_19 = rob_uop_30_pdst;
      default:
        casez_tmp_19 = rob_uop_31_pdst;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_20;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_20 = rob_uop_0_stale_pdst;
      5'b00001:
        casez_tmp_20 = rob_uop_1_stale_pdst;
      5'b00010:
        casez_tmp_20 = rob_uop_2_stale_pdst;
      5'b00011:
        casez_tmp_20 = rob_uop_3_stale_pdst;
      5'b00100:
        casez_tmp_20 = rob_uop_4_stale_pdst;
      5'b00101:
        casez_tmp_20 = rob_uop_5_stale_pdst;
      5'b00110:
        casez_tmp_20 = rob_uop_6_stale_pdst;
      5'b00111:
        casez_tmp_20 = rob_uop_7_stale_pdst;
      5'b01000:
        casez_tmp_20 = rob_uop_8_stale_pdst;
      5'b01001:
        casez_tmp_20 = rob_uop_9_stale_pdst;
      5'b01010:
        casez_tmp_20 = rob_uop_10_stale_pdst;
      5'b01011:
        casez_tmp_20 = rob_uop_11_stale_pdst;
      5'b01100:
        casez_tmp_20 = rob_uop_12_stale_pdst;
      5'b01101:
        casez_tmp_20 = rob_uop_13_stale_pdst;
      5'b01110:
        casez_tmp_20 = rob_uop_14_stale_pdst;
      5'b01111:
        casez_tmp_20 = rob_uop_15_stale_pdst;
      5'b10000:
        casez_tmp_20 = rob_uop_16_stale_pdst;
      5'b10001:
        casez_tmp_20 = rob_uop_17_stale_pdst;
      5'b10010:
        casez_tmp_20 = rob_uop_18_stale_pdst;
      5'b10011:
        casez_tmp_20 = rob_uop_19_stale_pdst;
      5'b10100:
        casez_tmp_20 = rob_uop_20_stale_pdst;
      5'b10101:
        casez_tmp_20 = rob_uop_21_stale_pdst;
      5'b10110:
        casez_tmp_20 = rob_uop_22_stale_pdst;
      5'b10111:
        casez_tmp_20 = rob_uop_23_stale_pdst;
      5'b11000:
        casez_tmp_20 = rob_uop_24_stale_pdst;
      5'b11001:
        casez_tmp_20 = rob_uop_25_stale_pdst;
      5'b11010:
        casez_tmp_20 = rob_uop_26_stale_pdst;
      5'b11011:
        casez_tmp_20 = rob_uop_27_stale_pdst;
      5'b11100:
        casez_tmp_20 = rob_uop_28_stale_pdst;
      5'b11101:
        casez_tmp_20 = rob_uop_29_stale_pdst;
      5'b11110:
        casez_tmp_20 = rob_uop_30_stale_pdst;
      default:
        casez_tmp_20 = rob_uop_31_stale_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_21;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_21 = rob_uop_0_is_fencei;
      5'b00001:
        casez_tmp_21 = rob_uop_1_is_fencei;
      5'b00010:
        casez_tmp_21 = rob_uop_2_is_fencei;
      5'b00011:
        casez_tmp_21 = rob_uop_3_is_fencei;
      5'b00100:
        casez_tmp_21 = rob_uop_4_is_fencei;
      5'b00101:
        casez_tmp_21 = rob_uop_5_is_fencei;
      5'b00110:
        casez_tmp_21 = rob_uop_6_is_fencei;
      5'b00111:
        casez_tmp_21 = rob_uop_7_is_fencei;
      5'b01000:
        casez_tmp_21 = rob_uop_8_is_fencei;
      5'b01001:
        casez_tmp_21 = rob_uop_9_is_fencei;
      5'b01010:
        casez_tmp_21 = rob_uop_10_is_fencei;
      5'b01011:
        casez_tmp_21 = rob_uop_11_is_fencei;
      5'b01100:
        casez_tmp_21 = rob_uop_12_is_fencei;
      5'b01101:
        casez_tmp_21 = rob_uop_13_is_fencei;
      5'b01110:
        casez_tmp_21 = rob_uop_14_is_fencei;
      5'b01111:
        casez_tmp_21 = rob_uop_15_is_fencei;
      5'b10000:
        casez_tmp_21 = rob_uop_16_is_fencei;
      5'b10001:
        casez_tmp_21 = rob_uop_17_is_fencei;
      5'b10010:
        casez_tmp_21 = rob_uop_18_is_fencei;
      5'b10011:
        casez_tmp_21 = rob_uop_19_is_fencei;
      5'b10100:
        casez_tmp_21 = rob_uop_20_is_fencei;
      5'b10101:
        casez_tmp_21 = rob_uop_21_is_fencei;
      5'b10110:
        casez_tmp_21 = rob_uop_22_is_fencei;
      5'b10111:
        casez_tmp_21 = rob_uop_23_is_fencei;
      5'b11000:
        casez_tmp_21 = rob_uop_24_is_fencei;
      5'b11001:
        casez_tmp_21 = rob_uop_25_is_fencei;
      5'b11010:
        casez_tmp_21 = rob_uop_26_is_fencei;
      5'b11011:
        casez_tmp_21 = rob_uop_27_is_fencei;
      5'b11100:
        casez_tmp_21 = rob_uop_28_is_fencei;
      5'b11101:
        casez_tmp_21 = rob_uop_29_is_fencei;
      5'b11110:
        casez_tmp_21 = rob_uop_30_is_fencei;
      default:
        casez_tmp_21 = rob_uop_31_is_fencei;
    endcase
  end // always @(*)
  reg         casez_tmp_22;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_22 = rob_uop_0_uses_ldq;
      5'b00001:
        casez_tmp_22 = rob_uop_1_uses_ldq;
      5'b00010:
        casez_tmp_22 = rob_uop_2_uses_ldq;
      5'b00011:
        casez_tmp_22 = rob_uop_3_uses_ldq;
      5'b00100:
        casez_tmp_22 = rob_uop_4_uses_ldq;
      5'b00101:
        casez_tmp_22 = rob_uop_5_uses_ldq;
      5'b00110:
        casez_tmp_22 = rob_uop_6_uses_ldq;
      5'b00111:
        casez_tmp_22 = rob_uop_7_uses_ldq;
      5'b01000:
        casez_tmp_22 = rob_uop_8_uses_ldq;
      5'b01001:
        casez_tmp_22 = rob_uop_9_uses_ldq;
      5'b01010:
        casez_tmp_22 = rob_uop_10_uses_ldq;
      5'b01011:
        casez_tmp_22 = rob_uop_11_uses_ldq;
      5'b01100:
        casez_tmp_22 = rob_uop_12_uses_ldq;
      5'b01101:
        casez_tmp_22 = rob_uop_13_uses_ldq;
      5'b01110:
        casez_tmp_22 = rob_uop_14_uses_ldq;
      5'b01111:
        casez_tmp_22 = rob_uop_15_uses_ldq;
      5'b10000:
        casez_tmp_22 = rob_uop_16_uses_ldq;
      5'b10001:
        casez_tmp_22 = rob_uop_17_uses_ldq;
      5'b10010:
        casez_tmp_22 = rob_uop_18_uses_ldq;
      5'b10011:
        casez_tmp_22 = rob_uop_19_uses_ldq;
      5'b10100:
        casez_tmp_22 = rob_uop_20_uses_ldq;
      5'b10101:
        casez_tmp_22 = rob_uop_21_uses_ldq;
      5'b10110:
        casez_tmp_22 = rob_uop_22_uses_ldq;
      5'b10111:
        casez_tmp_22 = rob_uop_23_uses_ldq;
      5'b11000:
        casez_tmp_22 = rob_uop_24_uses_ldq;
      5'b11001:
        casez_tmp_22 = rob_uop_25_uses_ldq;
      5'b11010:
        casez_tmp_22 = rob_uop_26_uses_ldq;
      5'b11011:
        casez_tmp_22 = rob_uop_27_uses_ldq;
      5'b11100:
        casez_tmp_22 = rob_uop_28_uses_ldq;
      5'b11101:
        casez_tmp_22 = rob_uop_29_uses_ldq;
      5'b11110:
        casez_tmp_22 = rob_uop_30_uses_ldq;
      default:
        casez_tmp_22 = rob_uop_31_uses_ldq;
    endcase
  end // always @(*)
  reg         casez_tmp_23;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_23 = rob_uop_0_uses_stq;
      5'b00001:
        casez_tmp_23 = rob_uop_1_uses_stq;
      5'b00010:
        casez_tmp_23 = rob_uop_2_uses_stq;
      5'b00011:
        casez_tmp_23 = rob_uop_3_uses_stq;
      5'b00100:
        casez_tmp_23 = rob_uop_4_uses_stq;
      5'b00101:
        casez_tmp_23 = rob_uop_5_uses_stq;
      5'b00110:
        casez_tmp_23 = rob_uop_6_uses_stq;
      5'b00111:
        casez_tmp_23 = rob_uop_7_uses_stq;
      5'b01000:
        casez_tmp_23 = rob_uop_8_uses_stq;
      5'b01001:
        casez_tmp_23 = rob_uop_9_uses_stq;
      5'b01010:
        casez_tmp_23 = rob_uop_10_uses_stq;
      5'b01011:
        casez_tmp_23 = rob_uop_11_uses_stq;
      5'b01100:
        casez_tmp_23 = rob_uop_12_uses_stq;
      5'b01101:
        casez_tmp_23 = rob_uop_13_uses_stq;
      5'b01110:
        casez_tmp_23 = rob_uop_14_uses_stq;
      5'b01111:
        casez_tmp_23 = rob_uop_15_uses_stq;
      5'b10000:
        casez_tmp_23 = rob_uop_16_uses_stq;
      5'b10001:
        casez_tmp_23 = rob_uop_17_uses_stq;
      5'b10010:
        casez_tmp_23 = rob_uop_18_uses_stq;
      5'b10011:
        casez_tmp_23 = rob_uop_19_uses_stq;
      5'b10100:
        casez_tmp_23 = rob_uop_20_uses_stq;
      5'b10101:
        casez_tmp_23 = rob_uop_21_uses_stq;
      5'b10110:
        casez_tmp_23 = rob_uop_22_uses_stq;
      5'b10111:
        casez_tmp_23 = rob_uop_23_uses_stq;
      5'b11000:
        casez_tmp_23 = rob_uop_24_uses_stq;
      5'b11001:
        casez_tmp_23 = rob_uop_25_uses_stq;
      5'b11010:
        casez_tmp_23 = rob_uop_26_uses_stq;
      5'b11011:
        casez_tmp_23 = rob_uop_27_uses_stq;
      5'b11100:
        casez_tmp_23 = rob_uop_28_uses_stq;
      5'b11101:
        casez_tmp_23 = rob_uop_29_uses_stq;
      5'b11110:
        casez_tmp_23 = rob_uop_30_uses_stq;
      default:
        casez_tmp_23 = rob_uop_31_uses_stq;
    endcase
  end // always @(*)
  reg         casez_tmp_24;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_24 = rob_uop_0_is_sys_pc2epc;
      5'b00001:
        casez_tmp_24 = rob_uop_1_is_sys_pc2epc;
      5'b00010:
        casez_tmp_24 = rob_uop_2_is_sys_pc2epc;
      5'b00011:
        casez_tmp_24 = rob_uop_3_is_sys_pc2epc;
      5'b00100:
        casez_tmp_24 = rob_uop_4_is_sys_pc2epc;
      5'b00101:
        casez_tmp_24 = rob_uop_5_is_sys_pc2epc;
      5'b00110:
        casez_tmp_24 = rob_uop_6_is_sys_pc2epc;
      5'b00111:
        casez_tmp_24 = rob_uop_7_is_sys_pc2epc;
      5'b01000:
        casez_tmp_24 = rob_uop_8_is_sys_pc2epc;
      5'b01001:
        casez_tmp_24 = rob_uop_9_is_sys_pc2epc;
      5'b01010:
        casez_tmp_24 = rob_uop_10_is_sys_pc2epc;
      5'b01011:
        casez_tmp_24 = rob_uop_11_is_sys_pc2epc;
      5'b01100:
        casez_tmp_24 = rob_uop_12_is_sys_pc2epc;
      5'b01101:
        casez_tmp_24 = rob_uop_13_is_sys_pc2epc;
      5'b01110:
        casez_tmp_24 = rob_uop_14_is_sys_pc2epc;
      5'b01111:
        casez_tmp_24 = rob_uop_15_is_sys_pc2epc;
      5'b10000:
        casez_tmp_24 = rob_uop_16_is_sys_pc2epc;
      5'b10001:
        casez_tmp_24 = rob_uop_17_is_sys_pc2epc;
      5'b10010:
        casez_tmp_24 = rob_uop_18_is_sys_pc2epc;
      5'b10011:
        casez_tmp_24 = rob_uop_19_is_sys_pc2epc;
      5'b10100:
        casez_tmp_24 = rob_uop_20_is_sys_pc2epc;
      5'b10101:
        casez_tmp_24 = rob_uop_21_is_sys_pc2epc;
      5'b10110:
        casez_tmp_24 = rob_uop_22_is_sys_pc2epc;
      5'b10111:
        casez_tmp_24 = rob_uop_23_is_sys_pc2epc;
      5'b11000:
        casez_tmp_24 = rob_uop_24_is_sys_pc2epc;
      5'b11001:
        casez_tmp_24 = rob_uop_25_is_sys_pc2epc;
      5'b11010:
        casez_tmp_24 = rob_uop_26_is_sys_pc2epc;
      5'b11011:
        casez_tmp_24 = rob_uop_27_is_sys_pc2epc;
      5'b11100:
        casez_tmp_24 = rob_uop_28_is_sys_pc2epc;
      5'b11101:
        casez_tmp_24 = rob_uop_29_is_sys_pc2epc;
      5'b11110:
        casez_tmp_24 = rob_uop_30_is_sys_pc2epc;
      default:
        casez_tmp_24 = rob_uop_31_is_sys_pc2epc;
    endcase
  end // always @(*)
  reg         casez_tmp_25;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_25 = rob_uop_0_flush_on_commit;
      5'b00001:
        casez_tmp_25 = rob_uop_1_flush_on_commit;
      5'b00010:
        casez_tmp_25 = rob_uop_2_flush_on_commit;
      5'b00011:
        casez_tmp_25 = rob_uop_3_flush_on_commit;
      5'b00100:
        casez_tmp_25 = rob_uop_4_flush_on_commit;
      5'b00101:
        casez_tmp_25 = rob_uop_5_flush_on_commit;
      5'b00110:
        casez_tmp_25 = rob_uop_6_flush_on_commit;
      5'b00111:
        casez_tmp_25 = rob_uop_7_flush_on_commit;
      5'b01000:
        casez_tmp_25 = rob_uop_8_flush_on_commit;
      5'b01001:
        casez_tmp_25 = rob_uop_9_flush_on_commit;
      5'b01010:
        casez_tmp_25 = rob_uop_10_flush_on_commit;
      5'b01011:
        casez_tmp_25 = rob_uop_11_flush_on_commit;
      5'b01100:
        casez_tmp_25 = rob_uop_12_flush_on_commit;
      5'b01101:
        casez_tmp_25 = rob_uop_13_flush_on_commit;
      5'b01110:
        casez_tmp_25 = rob_uop_14_flush_on_commit;
      5'b01111:
        casez_tmp_25 = rob_uop_15_flush_on_commit;
      5'b10000:
        casez_tmp_25 = rob_uop_16_flush_on_commit;
      5'b10001:
        casez_tmp_25 = rob_uop_17_flush_on_commit;
      5'b10010:
        casez_tmp_25 = rob_uop_18_flush_on_commit;
      5'b10011:
        casez_tmp_25 = rob_uop_19_flush_on_commit;
      5'b10100:
        casez_tmp_25 = rob_uop_20_flush_on_commit;
      5'b10101:
        casez_tmp_25 = rob_uop_21_flush_on_commit;
      5'b10110:
        casez_tmp_25 = rob_uop_22_flush_on_commit;
      5'b10111:
        casez_tmp_25 = rob_uop_23_flush_on_commit;
      5'b11000:
        casez_tmp_25 = rob_uop_24_flush_on_commit;
      5'b11001:
        casez_tmp_25 = rob_uop_25_flush_on_commit;
      5'b11010:
        casez_tmp_25 = rob_uop_26_flush_on_commit;
      5'b11011:
        casez_tmp_25 = rob_uop_27_flush_on_commit;
      5'b11100:
        casez_tmp_25 = rob_uop_28_flush_on_commit;
      5'b11101:
        casez_tmp_25 = rob_uop_29_flush_on_commit;
      5'b11110:
        casez_tmp_25 = rob_uop_30_flush_on_commit;
      default:
        casez_tmp_25 = rob_uop_31_flush_on_commit;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_26;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_26 = rob_uop_0_ldst;
      5'b00001:
        casez_tmp_26 = rob_uop_1_ldst;
      5'b00010:
        casez_tmp_26 = rob_uop_2_ldst;
      5'b00011:
        casez_tmp_26 = rob_uop_3_ldst;
      5'b00100:
        casez_tmp_26 = rob_uop_4_ldst;
      5'b00101:
        casez_tmp_26 = rob_uop_5_ldst;
      5'b00110:
        casez_tmp_26 = rob_uop_6_ldst;
      5'b00111:
        casez_tmp_26 = rob_uop_7_ldst;
      5'b01000:
        casez_tmp_26 = rob_uop_8_ldst;
      5'b01001:
        casez_tmp_26 = rob_uop_9_ldst;
      5'b01010:
        casez_tmp_26 = rob_uop_10_ldst;
      5'b01011:
        casez_tmp_26 = rob_uop_11_ldst;
      5'b01100:
        casez_tmp_26 = rob_uop_12_ldst;
      5'b01101:
        casez_tmp_26 = rob_uop_13_ldst;
      5'b01110:
        casez_tmp_26 = rob_uop_14_ldst;
      5'b01111:
        casez_tmp_26 = rob_uop_15_ldst;
      5'b10000:
        casez_tmp_26 = rob_uop_16_ldst;
      5'b10001:
        casez_tmp_26 = rob_uop_17_ldst;
      5'b10010:
        casez_tmp_26 = rob_uop_18_ldst;
      5'b10011:
        casez_tmp_26 = rob_uop_19_ldst;
      5'b10100:
        casez_tmp_26 = rob_uop_20_ldst;
      5'b10101:
        casez_tmp_26 = rob_uop_21_ldst;
      5'b10110:
        casez_tmp_26 = rob_uop_22_ldst;
      5'b10111:
        casez_tmp_26 = rob_uop_23_ldst;
      5'b11000:
        casez_tmp_26 = rob_uop_24_ldst;
      5'b11001:
        casez_tmp_26 = rob_uop_25_ldst;
      5'b11010:
        casez_tmp_26 = rob_uop_26_ldst;
      5'b11011:
        casez_tmp_26 = rob_uop_27_ldst;
      5'b11100:
        casez_tmp_26 = rob_uop_28_ldst;
      5'b11101:
        casez_tmp_26 = rob_uop_29_ldst;
      5'b11110:
        casez_tmp_26 = rob_uop_30_ldst;
      default:
        casez_tmp_26 = rob_uop_31_ldst;
    endcase
  end // always @(*)
  reg         casez_tmp_27;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_27 = rob_uop_0_ldst_val;
      5'b00001:
        casez_tmp_27 = rob_uop_1_ldst_val;
      5'b00010:
        casez_tmp_27 = rob_uop_2_ldst_val;
      5'b00011:
        casez_tmp_27 = rob_uop_3_ldst_val;
      5'b00100:
        casez_tmp_27 = rob_uop_4_ldst_val;
      5'b00101:
        casez_tmp_27 = rob_uop_5_ldst_val;
      5'b00110:
        casez_tmp_27 = rob_uop_6_ldst_val;
      5'b00111:
        casez_tmp_27 = rob_uop_7_ldst_val;
      5'b01000:
        casez_tmp_27 = rob_uop_8_ldst_val;
      5'b01001:
        casez_tmp_27 = rob_uop_9_ldst_val;
      5'b01010:
        casez_tmp_27 = rob_uop_10_ldst_val;
      5'b01011:
        casez_tmp_27 = rob_uop_11_ldst_val;
      5'b01100:
        casez_tmp_27 = rob_uop_12_ldst_val;
      5'b01101:
        casez_tmp_27 = rob_uop_13_ldst_val;
      5'b01110:
        casez_tmp_27 = rob_uop_14_ldst_val;
      5'b01111:
        casez_tmp_27 = rob_uop_15_ldst_val;
      5'b10000:
        casez_tmp_27 = rob_uop_16_ldst_val;
      5'b10001:
        casez_tmp_27 = rob_uop_17_ldst_val;
      5'b10010:
        casez_tmp_27 = rob_uop_18_ldst_val;
      5'b10011:
        casez_tmp_27 = rob_uop_19_ldst_val;
      5'b10100:
        casez_tmp_27 = rob_uop_20_ldst_val;
      5'b10101:
        casez_tmp_27 = rob_uop_21_ldst_val;
      5'b10110:
        casez_tmp_27 = rob_uop_22_ldst_val;
      5'b10111:
        casez_tmp_27 = rob_uop_23_ldst_val;
      5'b11000:
        casez_tmp_27 = rob_uop_24_ldst_val;
      5'b11001:
        casez_tmp_27 = rob_uop_25_ldst_val;
      5'b11010:
        casez_tmp_27 = rob_uop_26_ldst_val;
      5'b11011:
        casez_tmp_27 = rob_uop_27_ldst_val;
      5'b11100:
        casez_tmp_27 = rob_uop_28_ldst_val;
      5'b11101:
        casez_tmp_27 = rob_uop_29_ldst_val;
      5'b11110:
        casez_tmp_27 = rob_uop_30_ldst_val;
      default:
        casez_tmp_27 = rob_uop_31_ldst_val;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_28;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_28 = rob_uop_0_dst_rtype;
      5'b00001:
        casez_tmp_28 = rob_uop_1_dst_rtype;
      5'b00010:
        casez_tmp_28 = rob_uop_2_dst_rtype;
      5'b00011:
        casez_tmp_28 = rob_uop_3_dst_rtype;
      5'b00100:
        casez_tmp_28 = rob_uop_4_dst_rtype;
      5'b00101:
        casez_tmp_28 = rob_uop_5_dst_rtype;
      5'b00110:
        casez_tmp_28 = rob_uop_6_dst_rtype;
      5'b00111:
        casez_tmp_28 = rob_uop_7_dst_rtype;
      5'b01000:
        casez_tmp_28 = rob_uop_8_dst_rtype;
      5'b01001:
        casez_tmp_28 = rob_uop_9_dst_rtype;
      5'b01010:
        casez_tmp_28 = rob_uop_10_dst_rtype;
      5'b01011:
        casez_tmp_28 = rob_uop_11_dst_rtype;
      5'b01100:
        casez_tmp_28 = rob_uop_12_dst_rtype;
      5'b01101:
        casez_tmp_28 = rob_uop_13_dst_rtype;
      5'b01110:
        casez_tmp_28 = rob_uop_14_dst_rtype;
      5'b01111:
        casez_tmp_28 = rob_uop_15_dst_rtype;
      5'b10000:
        casez_tmp_28 = rob_uop_16_dst_rtype;
      5'b10001:
        casez_tmp_28 = rob_uop_17_dst_rtype;
      5'b10010:
        casez_tmp_28 = rob_uop_18_dst_rtype;
      5'b10011:
        casez_tmp_28 = rob_uop_19_dst_rtype;
      5'b10100:
        casez_tmp_28 = rob_uop_20_dst_rtype;
      5'b10101:
        casez_tmp_28 = rob_uop_21_dst_rtype;
      5'b10110:
        casez_tmp_28 = rob_uop_22_dst_rtype;
      5'b10111:
        casez_tmp_28 = rob_uop_23_dst_rtype;
      5'b11000:
        casez_tmp_28 = rob_uop_24_dst_rtype;
      5'b11001:
        casez_tmp_28 = rob_uop_25_dst_rtype;
      5'b11010:
        casez_tmp_28 = rob_uop_26_dst_rtype;
      5'b11011:
        casez_tmp_28 = rob_uop_27_dst_rtype;
      5'b11100:
        casez_tmp_28 = rob_uop_28_dst_rtype;
      5'b11101:
        casez_tmp_28 = rob_uop_29_dst_rtype;
      5'b11110:
        casez_tmp_28 = rob_uop_30_dst_rtype;
      default:
        casez_tmp_28 = rob_uop_31_dst_rtype;
    endcase
  end // always @(*)
  reg         casez_tmp_29;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_29 = rob_uop_0_fp_val;
      5'b00001:
        casez_tmp_29 = rob_uop_1_fp_val;
      5'b00010:
        casez_tmp_29 = rob_uop_2_fp_val;
      5'b00011:
        casez_tmp_29 = rob_uop_3_fp_val;
      5'b00100:
        casez_tmp_29 = rob_uop_4_fp_val;
      5'b00101:
        casez_tmp_29 = rob_uop_5_fp_val;
      5'b00110:
        casez_tmp_29 = rob_uop_6_fp_val;
      5'b00111:
        casez_tmp_29 = rob_uop_7_fp_val;
      5'b01000:
        casez_tmp_29 = rob_uop_8_fp_val;
      5'b01001:
        casez_tmp_29 = rob_uop_9_fp_val;
      5'b01010:
        casez_tmp_29 = rob_uop_10_fp_val;
      5'b01011:
        casez_tmp_29 = rob_uop_11_fp_val;
      5'b01100:
        casez_tmp_29 = rob_uop_12_fp_val;
      5'b01101:
        casez_tmp_29 = rob_uop_13_fp_val;
      5'b01110:
        casez_tmp_29 = rob_uop_14_fp_val;
      5'b01111:
        casez_tmp_29 = rob_uop_15_fp_val;
      5'b10000:
        casez_tmp_29 = rob_uop_16_fp_val;
      5'b10001:
        casez_tmp_29 = rob_uop_17_fp_val;
      5'b10010:
        casez_tmp_29 = rob_uop_18_fp_val;
      5'b10011:
        casez_tmp_29 = rob_uop_19_fp_val;
      5'b10100:
        casez_tmp_29 = rob_uop_20_fp_val;
      5'b10101:
        casez_tmp_29 = rob_uop_21_fp_val;
      5'b10110:
        casez_tmp_29 = rob_uop_22_fp_val;
      5'b10111:
        casez_tmp_29 = rob_uop_23_fp_val;
      5'b11000:
        casez_tmp_29 = rob_uop_24_fp_val;
      5'b11001:
        casez_tmp_29 = rob_uop_25_fp_val;
      5'b11010:
        casez_tmp_29 = rob_uop_26_fp_val;
      5'b11011:
        casez_tmp_29 = rob_uop_27_fp_val;
      5'b11100:
        casez_tmp_29 = rob_uop_28_fp_val;
      5'b11101:
        casez_tmp_29 = rob_uop_29_fp_val;
      5'b11110:
        casez_tmp_29 = rob_uop_30_fp_val;
      default:
        casez_tmp_29 = rob_uop_31_fp_val;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_30;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_30 = rob_uop_0_debug_fsrc;
      5'b00001:
        casez_tmp_30 = rob_uop_1_debug_fsrc;
      5'b00010:
        casez_tmp_30 = rob_uop_2_debug_fsrc;
      5'b00011:
        casez_tmp_30 = rob_uop_3_debug_fsrc;
      5'b00100:
        casez_tmp_30 = rob_uop_4_debug_fsrc;
      5'b00101:
        casez_tmp_30 = rob_uop_5_debug_fsrc;
      5'b00110:
        casez_tmp_30 = rob_uop_6_debug_fsrc;
      5'b00111:
        casez_tmp_30 = rob_uop_7_debug_fsrc;
      5'b01000:
        casez_tmp_30 = rob_uop_8_debug_fsrc;
      5'b01001:
        casez_tmp_30 = rob_uop_9_debug_fsrc;
      5'b01010:
        casez_tmp_30 = rob_uop_10_debug_fsrc;
      5'b01011:
        casez_tmp_30 = rob_uop_11_debug_fsrc;
      5'b01100:
        casez_tmp_30 = rob_uop_12_debug_fsrc;
      5'b01101:
        casez_tmp_30 = rob_uop_13_debug_fsrc;
      5'b01110:
        casez_tmp_30 = rob_uop_14_debug_fsrc;
      5'b01111:
        casez_tmp_30 = rob_uop_15_debug_fsrc;
      5'b10000:
        casez_tmp_30 = rob_uop_16_debug_fsrc;
      5'b10001:
        casez_tmp_30 = rob_uop_17_debug_fsrc;
      5'b10010:
        casez_tmp_30 = rob_uop_18_debug_fsrc;
      5'b10011:
        casez_tmp_30 = rob_uop_19_debug_fsrc;
      5'b10100:
        casez_tmp_30 = rob_uop_20_debug_fsrc;
      5'b10101:
        casez_tmp_30 = rob_uop_21_debug_fsrc;
      5'b10110:
        casez_tmp_30 = rob_uop_22_debug_fsrc;
      5'b10111:
        casez_tmp_30 = rob_uop_23_debug_fsrc;
      5'b11000:
        casez_tmp_30 = rob_uop_24_debug_fsrc;
      5'b11001:
        casez_tmp_30 = rob_uop_25_debug_fsrc;
      5'b11010:
        casez_tmp_30 = rob_uop_26_debug_fsrc;
      5'b11011:
        casez_tmp_30 = rob_uop_27_debug_fsrc;
      5'b11100:
        casez_tmp_30 = rob_uop_28_debug_fsrc;
      5'b11101:
        casez_tmp_30 = rob_uop_29_debug_fsrc;
      5'b11110:
        casez_tmp_30 = rob_uop_30_debug_fsrc;
      default:
        casez_tmp_30 = rob_uop_31_debug_fsrc;
    endcase
  end // always @(*)
  wire        _GEN_15 = io_brupdate_b2_mispredict & io_brupdate_b2_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_16 = io_brupdate_b2_uop_rob_idx[6:2] == com_idx;
  wire        rbk_row = _io_commit_rollback_T_3 & ~full;
  reg         casez_tmp_31;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_31 = rob_val_0;
      5'b00001:
        casez_tmp_31 = rob_val_1;
      5'b00010:
        casez_tmp_31 = rob_val_2;
      5'b00011:
        casez_tmp_31 = rob_val_3;
      5'b00100:
        casez_tmp_31 = rob_val_4;
      5'b00101:
        casez_tmp_31 = rob_val_5;
      5'b00110:
        casez_tmp_31 = rob_val_6;
      5'b00111:
        casez_tmp_31 = rob_val_7;
      5'b01000:
        casez_tmp_31 = rob_val_8;
      5'b01001:
        casez_tmp_31 = rob_val_9;
      5'b01010:
        casez_tmp_31 = rob_val_10;
      5'b01011:
        casez_tmp_31 = rob_val_11;
      5'b01100:
        casez_tmp_31 = rob_val_12;
      5'b01101:
        casez_tmp_31 = rob_val_13;
      5'b01110:
        casez_tmp_31 = rob_val_14;
      5'b01111:
        casez_tmp_31 = rob_val_15;
      5'b10000:
        casez_tmp_31 = rob_val_16;
      5'b10001:
        casez_tmp_31 = rob_val_17;
      5'b10010:
        casez_tmp_31 = rob_val_18;
      5'b10011:
        casez_tmp_31 = rob_val_19;
      5'b10100:
        casez_tmp_31 = rob_val_20;
      5'b10101:
        casez_tmp_31 = rob_val_21;
      5'b10110:
        casez_tmp_31 = rob_val_22;
      5'b10111:
        casez_tmp_31 = rob_val_23;
      5'b11000:
        casez_tmp_31 = rob_val_24;
      5'b11001:
        casez_tmp_31 = rob_val_25;
      5'b11010:
        casez_tmp_31 = rob_val_26;
      5'b11011:
        casez_tmp_31 = rob_val_27;
      5'b11100:
        casez_tmp_31 = rob_val_28;
      5'b11101:
        casez_tmp_31 = rob_val_29;
      5'b11110:
        casez_tmp_31 = rob_val_30;
      default:
        casez_tmp_31 = rob_val_31;
    endcase
  end // always @(*)
  wire        _io_commit_rbk_valids_0_output = rbk_row & casez_tmp_31;
  reg  [4:0]  casez_tmp_32;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_32 = rob_fflags_0_0;
      5'b00001:
        casez_tmp_32 = rob_fflags_0_1;
      5'b00010:
        casez_tmp_32 = rob_fflags_0_2;
      5'b00011:
        casez_tmp_32 = rob_fflags_0_3;
      5'b00100:
        casez_tmp_32 = rob_fflags_0_4;
      5'b00101:
        casez_tmp_32 = rob_fflags_0_5;
      5'b00110:
        casez_tmp_32 = rob_fflags_0_6;
      5'b00111:
        casez_tmp_32 = rob_fflags_0_7;
      5'b01000:
        casez_tmp_32 = rob_fflags_0_8;
      5'b01001:
        casez_tmp_32 = rob_fflags_0_9;
      5'b01010:
        casez_tmp_32 = rob_fflags_0_10;
      5'b01011:
        casez_tmp_32 = rob_fflags_0_11;
      5'b01100:
        casez_tmp_32 = rob_fflags_0_12;
      5'b01101:
        casez_tmp_32 = rob_fflags_0_13;
      5'b01110:
        casez_tmp_32 = rob_fflags_0_14;
      5'b01111:
        casez_tmp_32 = rob_fflags_0_15;
      5'b10000:
        casez_tmp_32 = rob_fflags_0_16;
      5'b10001:
        casez_tmp_32 = rob_fflags_0_17;
      5'b10010:
        casez_tmp_32 = rob_fflags_0_18;
      5'b10011:
        casez_tmp_32 = rob_fflags_0_19;
      5'b10100:
        casez_tmp_32 = rob_fflags_0_20;
      5'b10101:
        casez_tmp_32 = rob_fflags_0_21;
      5'b10110:
        casez_tmp_32 = rob_fflags_0_22;
      5'b10111:
        casez_tmp_32 = rob_fflags_0_23;
      5'b11000:
        casez_tmp_32 = rob_fflags_0_24;
      5'b11001:
        casez_tmp_32 = rob_fflags_0_25;
      5'b11010:
        casez_tmp_32 = rob_fflags_0_26;
      5'b11011:
        casez_tmp_32 = rob_fflags_0_27;
      5'b11100:
        casez_tmp_32 = rob_fflags_0_28;
      5'b11101:
        casez_tmp_32 = rob_fflags_0_29;
      5'b11110:
        casez_tmp_32 = rob_fflags_0_30;
      default:
        casez_tmp_32 = rob_fflags_0_31;
    endcase
  end // always @(*)
  reg         casez_tmp_33;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_33 = rob_uop_0_uses_ldq;
      5'b00001:
        casez_tmp_33 = rob_uop_1_uses_ldq;
      5'b00010:
        casez_tmp_33 = rob_uop_2_uses_ldq;
      5'b00011:
        casez_tmp_33 = rob_uop_3_uses_ldq;
      5'b00100:
        casez_tmp_33 = rob_uop_4_uses_ldq;
      5'b00101:
        casez_tmp_33 = rob_uop_5_uses_ldq;
      5'b00110:
        casez_tmp_33 = rob_uop_6_uses_ldq;
      5'b00111:
        casez_tmp_33 = rob_uop_7_uses_ldq;
      5'b01000:
        casez_tmp_33 = rob_uop_8_uses_ldq;
      5'b01001:
        casez_tmp_33 = rob_uop_9_uses_ldq;
      5'b01010:
        casez_tmp_33 = rob_uop_10_uses_ldq;
      5'b01011:
        casez_tmp_33 = rob_uop_11_uses_ldq;
      5'b01100:
        casez_tmp_33 = rob_uop_12_uses_ldq;
      5'b01101:
        casez_tmp_33 = rob_uop_13_uses_ldq;
      5'b01110:
        casez_tmp_33 = rob_uop_14_uses_ldq;
      5'b01111:
        casez_tmp_33 = rob_uop_15_uses_ldq;
      5'b10000:
        casez_tmp_33 = rob_uop_16_uses_ldq;
      5'b10001:
        casez_tmp_33 = rob_uop_17_uses_ldq;
      5'b10010:
        casez_tmp_33 = rob_uop_18_uses_ldq;
      5'b10011:
        casez_tmp_33 = rob_uop_19_uses_ldq;
      5'b10100:
        casez_tmp_33 = rob_uop_20_uses_ldq;
      5'b10101:
        casez_tmp_33 = rob_uop_21_uses_ldq;
      5'b10110:
        casez_tmp_33 = rob_uop_22_uses_ldq;
      5'b10111:
        casez_tmp_33 = rob_uop_23_uses_ldq;
      5'b11000:
        casez_tmp_33 = rob_uop_24_uses_ldq;
      5'b11001:
        casez_tmp_33 = rob_uop_25_uses_ldq;
      5'b11010:
        casez_tmp_33 = rob_uop_26_uses_ldq;
      5'b11011:
        casez_tmp_33 = rob_uop_27_uses_ldq;
      5'b11100:
        casez_tmp_33 = rob_uop_28_uses_ldq;
      5'b11101:
        casez_tmp_33 = rob_uop_29_uses_ldq;
      5'b11110:
        casez_tmp_33 = rob_uop_30_uses_ldq;
      default:
        casez_tmp_33 = rob_uop_31_uses_ldq;
    endcase
  end // always @(*)
  reg         casez_tmp_34;
  always @(*) begin
    casez (rob_pnr)
      5'b00000:
        casez_tmp_34 = rob_unsafe_0;
      5'b00001:
        casez_tmp_34 = rob_unsafe_1;
      5'b00010:
        casez_tmp_34 = rob_unsafe_2;
      5'b00011:
        casez_tmp_34 = rob_unsafe_3;
      5'b00100:
        casez_tmp_34 = rob_unsafe_4;
      5'b00101:
        casez_tmp_34 = rob_unsafe_5;
      5'b00110:
        casez_tmp_34 = rob_unsafe_6;
      5'b00111:
        casez_tmp_34 = rob_unsafe_7;
      5'b01000:
        casez_tmp_34 = rob_unsafe_8;
      5'b01001:
        casez_tmp_34 = rob_unsafe_9;
      5'b01010:
        casez_tmp_34 = rob_unsafe_10;
      5'b01011:
        casez_tmp_34 = rob_unsafe_11;
      5'b01100:
        casez_tmp_34 = rob_unsafe_12;
      5'b01101:
        casez_tmp_34 = rob_unsafe_13;
      5'b01110:
        casez_tmp_34 = rob_unsafe_14;
      5'b01111:
        casez_tmp_34 = rob_unsafe_15;
      5'b10000:
        casez_tmp_34 = rob_unsafe_16;
      5'b10001:
        casez_tmp_34 = rob_unsafe_17;
      5'b10010:
        casez_tmp_34 = rob_unsafe_18;
      5'b10011:
        casez_tmp_34 = rob_unsafe_19;
      5'b10100:
        casez_tmp_34 = rob_unsafe_20;
      5'b10101:
        casez_tmp_34 = rob_unsafe_21;
      5'b10110:
        casez_tmp_34 = rob_unsafe_22;
      5'b10111:
        casez_tmp_34 = rob_unsafe_23;
      5'b11000:
        casez_tmp_34 = rob_unsafe_24;
      5'b11001:
        casez_tmp_34 = rob_unsafe_25;
      5'b11010:
        casez_tmp_34 = rob_unsafe_26;
      5'b11011:
        casez_tmp_34 = rob_unsafe_27;
      5'b11100:
        casez_tmp_34 = rob_unsafe_28;
      5'b11101:
        casez_tmp_34 = rob_unsafe_29;
      5'b11110:
        casez_tmp_34 = rob_unsafe_30;
      default:
        casez_tmp_34 = rob_unsafe_31;
    endcase
  end // always @(*)
  reg         casez_tmp_35;
  always @(*) begin
    casez (rob_pnr)
      5'b00000:
        casez_tmp_35 = rob_exception_0;
      5'b00001:
        casez_tmp_35 = rob_exception_1;
      5'b00010:
        casez_tmp_35 = rob_exception_2;
      5'b00011:
        casez_tmp_35 = rob_exception_3;
      5'b00100:
        casez_tmp_35 = rob_exception_4;
      5'b00101:
        casez_tmp_35 = rob_exception_5;
      5'b00110:
        casez_tmp_35 = rob_exception_6;
      5'b00111:
        casez_tmp_35 = rob_exception_7;
      5'b01000:
        casez_tmp_35 = rob_exception_8;
      5'b01001:
        casez_tmp_35 = rob_exception_9;
      5'b01010:
        casez_tmp_35 = rob_exception_10;
      5'b01011:
        casez_tmp_35 = rob_exception_11;
      5'b01100:
        casez_tmp_35 = rob_exception_12;
      5'b01101:
        casez_tmp_35 = rob_exception_13;
      5'b01110:
        casez_tmp_35 = rob_exception_14;
      5'b01111:
        casez_tmp_35 = rob_exception_15;
      5'b10000:
        casez_tmp_35 = rob_exception_16;
      5'b10001:
        casez_tmp_35 = rob_exception_17;
      5'b10010:
        casez_tmp_35 = rob_exception_18;
      5'b10011:
        casez_tmp_35 = rob_exception_19;
      5'b10100:
        casez_tmp_35 = rob_exception_20;
      5'b10101:
        casez_tmp_35 = rob_exception_21;
      5'b10110:
        casez_tmp_35 = rob_exception_22;
      5'b10111:
        casez_tmp_35 = rob_exception_23;
      5'b11000:
        casez_tmp_35 = rob_exception_24;
      5'b11001:
        casez_tmp_35 = rob_exception_25;
      5'b11010:
        casez_tmp_35 = rob_exception_26;
      5'b11011:
        casez_tmp_35 = rob_exception_27;
      5'b11100:
        casez_tmp_35 = rob_exception_28;
      5'b11101:
        casez_tmp_35 = rob_exception_29;
      5'b11110:
        casez_tmp_35 = rob_exception_30;
      default:
        casez_tmp_35 = rob_exception_31;
    endcase
  end // always @(*)
  reg         casez_tmp_36;
  always @(*) begin
    casez (rob_pnr)
      5'b00000:
        casez_tmp_36 = rob_val_0;
      5'b00001:
        casez_tmp_36 = rob_val_1;
      5'b00010:
        casez_tmp_36 = rob_val_2;
      5'b00011:
        casez_tmp_36 = rob_val_3;
      5'b00100:
        casez_tmp_36 = rob_val_4;
      5'b00101:
        casez_tmp_36 = rob_val_5;
      5'b00110:
        casez_tmp_36 = rob_val_6;
      5'b00111:
        casez_tmp_36 = rob_val_7;
      5'b01000:
        casez_tmp_36 = rob_val_8;
      5'b01001:
        casez_tmp_36 = rob_val_9;
      5'b01010:
        casez_tmp_36 = rob_val_10;
      5'b01011:
        casez_tmp_36 = rob_val_11;
      5'b01100:
        casez_tmp_36 = rob_val_12;
      5'b01101:
        casez_tmp_36 = rob_val_13;
      5'b01110:
        casez_tmp_36 = rob_val_14;
      5'b01111:
        casez_tmp_36 = rob_val_15;
      5'b10000:
        casez_tmp_36 = rob_val_16;
      5'b10001:
        casez_tmp_36 = rob_val_17;
      5'b10010:
        casez_tmp_36 = rob_val_18;
      5'b10011:
        casez_tmp_36 = rob_val_19;
      5'b10100:
        casez_tmp_36 = rob_val_20;
      5'b10101:
        casez_tmp_36 = rob_val_21;
      5'b10110:
        casez_tmp_36 = rob_val_22;
      5'b10111:
        casez_tmp_36 = rob_val_23;
      5'b11000:
        casez_tmp_36 = rob_val_24;
      5'b11001:
        casez_tmp_36 = rob_val_25;
      5'b11010:
        casez_tmp_36 = rob_val_26;
      5'b11011:
        casez_tmp_36 = rob_val_27;
      5'b11100:
        casez_tmp_36 = rob_val_28;
      5'b11101:
        casez_tmp_36 = rob_val_29;
      5'b11110:
        casez_tmp_36 = rob_val_30;
      default:
        casez_tmp_36 = rob_val_31;
    endcase
  end // always @(*)
  reg         casez_tmp_37;
  always @(*) begin
    casez (io_wb_resps_0_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_37 = rob_val_0;
      5'b00001:
        casez_tmp_37 = rob_val_1;
      5'b00010:
        casez_tmp_37 = rob_val_2;
      5'b00011:
        casez_tmp_37 = rob_val_3;
      5'b00100:
        casez_tmp_37 = rob_val_4;
      5'b00101:
        casez_tmp_37 = rob_val_5;
      5'b00110:
        casez_tmp_37 = rob_val_6;
      5'b00111:
        casez_tmp_37 = rob_val_7;
      5'b01000:
        casez_tmp_37 = rob_val_8;
      5'b01001:
        casez_tmp_37 = rob_val_9;
      5'b01010:
        casez_tmp_37 = rob_val_10;
      5'b01011:
        casez_tmp_37 = rob_val_11;
      5'b01100:
        casez_tmp_37 = rob_val_12;
      5'b01101:
        casez_tmp_37 = rob_val_13;
      5'b01110:
        casez_tmp_37 = rob_val_14;
      5'b01111:
        casez_tmp_37 = rob_val_15;
      5'b10000:
        casez_tmp_37 = rob_val_16;
      5'b10001:
        casez_tmp_37 = rob_val_17;
      5'b10010:
        casez_tmp_37 = rob_val_18;
      5'b10011:
        casez_tmp_37 = rob_val_19;
      5'b10100:
        casez_tmp_37 = rob_val_20;
      5'b10101:
        casez_tmp_37 = rob_val_21;
      5'b10110:
        casez_tmp_37 = rob_val_22;
      5'b10111:
        casez_tmp_37 = rob_val_23;
      5'b11000:
        casez_tmp_37 = rob_val_24;
      5'b11001:
        casez_tmp_37 = rob_val_25;
      5'b11010:
        casez_tmp_37 = rob_val_26;
      5'b11011:
        casez_tmp_37 = rob_val_27;
      5'b11100:
        casez_tmp_37 = rob_val_28;
      5'b11101:
        casez_tmp_37 = rob_val_29;
      5'b11110:
        casez_tmp_37 = rob_val_30;
      default:
        casez_tmp_37 = rob_val_31;
    endcase
  end // always @(*)
  reg         casez_tmp_38;
  always @(*) begin
    casez (io_wb_resps_0_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_38 = rob_bsy_0;
      5'b00001:
        casez_tmp_38 = rob_bsy_1;
      5'b00010:
        casez_tmp_38 = rob_bsy_2;
      5'b00011:
        casez_tmp_38 = rob_bsy_3;
      5'b00100:
        casez_tmp_38 = rob_bsy_4;
      5'b00101:
        casez_tmp_38 = rob_bsy_5;
      5'b00110:
        casez_tmp_38 = rob_bsy_6;
      5'b00111:
        casez_tmp_38 = rob_bsy_7;
      5'b01000:
        casez_tmp_38 = rob_bsy_8;
      5'b01001:
        casez_tmp_38 = rob_bsy_9;
      5'b01010:
        casez_tmp_38 = rob_bsy_10;
      5'b01011:
        casez_tmp_38 = rob_bsy_11;
      5'b01100:
        casez_tmp_38 = rob_bsy_12;
      5'b01101:
        casez_tmp_38 = rob_bsy_13;
      5'b01110:
        casez_tmp_38 = rob_bsy_14;
      5'b01111:
        casez_tmp_38 = rob_bsy_15;
      5'b10000:
        casez_tmp_38 = rob_bsy_16;
      5'b10001:
        casez_tmp_38 = rob_bsy_17;
      5'b10010:
        casez_tmp_38 = rob_bsy_18;
      5'b10011:
        casez_tmp_38 = rob_bsy_19;
      5'b10100:
        casez_tmp_38 = rob_bsy_20;
      5'b10101:
        casez_tmp_38 = rob_bsy_21;
      5'b10110:
        casez_tmp_38 = rob_bsy_22;
      5'b10111:
        casez_tmp_38 = rob_bsy_23;
      5'b11000:
        casez_tmp_38 = rob_bsy_24;
      5'b11001:
        casez_tmp_38 = rob_bsy_25;
      5'b11010:
        casez_tmp_38 = rob_bsy_26;
      5'b11011:
        casez_tmp_38 = rob_bsy_27;
      5'b11100:
        casez_tmp_38 = rob_bsy_28;
      5'b11101:
        casez_tmp_38 = rob_bsy_29;
      5'b11110:
        casez_tmp_38 = rob_bsy_30;
      default:
        casez_tmp_38 = rob_bsy_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_39;
  always @(*) begin
    casez (io_wb_resps_0_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_39 = rob_uop_0_pdst;
      5'b00001:
        casez_tmp_39 = rob_uop_1_pdst;
      5'b00010:
        casez_tmp_39 = rob_uop_2_pdst;
      5'b00011:
        casez_tmp_39 = rob_uop_3_pdst;
      5'b00100:
        casez_tmp_39 = rob_uop_4_pdst;
      5'b00101:
        casez_tmp_39 = rob_uop_5_pdst;
      5'b00110:
        casez_tmp_39 = rob_uop_6_pdst;
      5'b00111:
        casez_tmp_39 = rob_uop_7_pdst;
      5'b01000:
        casez_tmp_39 = rob_uop_8_pdst;
      5'b01001:
        casez_tmp_39 = rob_uop_9_pdst;
      5'b01010:
        casez_tmp_39 = rob_uop_10_pdst;
      5'b01011:
        casez_tmp_39 = rob_uop_11_pdst;
      5'b01100:
        casez_tmp_39 = rob_uop_12_pdst;
      5'b01101:
        casez_tmp_39 = rob_uop_13_pdst;
      5'b01110:
        casez_tmp_39 = rob_uop_14_pdst;
      5'b01111:
        casez_tmp_39 = rob_uop_15_pdst;
      5'b10000:
        casez_tmp_39 = rob_uop_16_pdst;
      5'b10001:
        casez_tmp_39 = rob_uop_17_pdst;
      5'b10010:
        casez_tmp_39 = rob_uop_18_pdst;
      5'b10011:
        casez_tmp_39 = rob_uop_19_pdst;
      5'b10100:
        casez_tmp_39 = rob_uop_20_pdst;
      5'b10101:
        casez_tmp_39 = rob_uop_21_pdst;
      5'b10110:
        casez_tmp_39 = rob_uop_22_pdst;
      5'b10111:
        casez_tmp_39 = rob_uop_23_pdst;
      5'b11000:
        casez_tmp_39 = rob_uop_24_pdst;
      5'b11001:
        casez_tmp_39 = rob_uop_25_pdst;
      5'b11010:
        casez_tmp_39 = rob_uop_26_pdst;
      5'b11011:
        casez_tmp_39 = rob_uop_27_pdst;
      5'b11100:
        casez_tmp_39 = rob_uop_28_pdst;
      5'b11101:
        casez_tmp_39 = rob_uop_29_pdst;
      5'b11110:
        casez_tmp_39 = rob_uop_30_pdst;
      default:
        casez_tmp_39 = rob_uop_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_40;
  always @(*) begin
    casez (io_wb_resps_0_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_40 = rob_uop_0_ldst_val;
      5'b00001:
        casez_tmp_40 = rob_uop_1_ldst_val;
      5'b00010:
        casez_tmp_40 = rob_uop_2_ldst_val;
      5'b00011:
        casez_tmp_40 = rob_uop_3_ldst_val;
      5'b00100:
        casez_tmp_40 = rob_uop_4_ldst_val;
      5'b00101:
        casez_tmp_40 = rob_uop_5_ldst_val;
      5'b00110:
        casez_tmp_40 = rob_uop_6_ldst_val;
      5'b00111:
        casez_tmp_40 = rob_uop_7_ldst_val;
      5'b01000:
        casez_tmp_40 = rob_uop_8_ldst_val;
      5'b01001:
        casez_tmp_40 = rob_uop_9_ldst_val;
      5'b01010:
        casez_tmp_40 = rob_uop_10_ldst_val;
      5'b01011:
        casez_tmp_40 = rob_uop_11_ldst_val;
      5'b01100:
        casez_tmp_40 = rob_uop_12_ldst_val;
      5'b01101:
        casez_tmp_40 = rob_uop_13_ldst_val;
      5'b01110:
        casez_tmp_40 = rob_uop_14_ldst_val;
      5'b01111:
        casez_tmp_40 = rob_uop_15_ldst_val;
      5'b10000:
        casez_tmp_40 = rob_uop_16_ldst_val;
      5'b10001:
        casez_tmp_40 = rob_uop_17_ldst_val;
      5'b10010:
        casez_tmp_40 = rob_uop_18_ldst_val;
      5'b10011:
        casez_tmp_40 = rob_uop_19_ldst_val;
      5'b10100:
        casez_tmp_40 = rob_uop_20_ldst_val;
      5'b10101:
        casez_tmp_40 = rob_uop_21_ldst_val;
      5'b10110:
        casez_tmp_40 = rob_uop_22_ldst_val;
      5'b10111:
        casez_tmp_40 = rob_uop_23_ldst_val;
      5'b11000:
        casez_tmp_40 = rob_uop_24_ldst_val;
      5'b11001:
        casez_tmp_40 = rob_uop_25_ldst_val;
      5'b11010:
        casez_tmp_40 = rob_uop_26_ldst_val;
      5'b11011:
        casez_tmp_40 = rob_uop_27_ldst_val;
      5'b11100:
        casez_tmp_40 = rob_uop_28_ldst_val;
      5'b11101:
        casez_tmp_40 = rob_uop_29_ldst_val;
      5'b11110:
        casez_tmp_40 = rob_uop_30_ldst_val;
      default:
        casez_tmp_40 = rob_uop_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_41;
  always @(*) begin
    casez (io_wb_resps_1_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_41 = rob_val_0;
      5'b00001:
        casez_tmp_41 = rob_val_1;
      5'b00010:
        casez_tmp_41 = rob_val_2;
      5'b00011:
        casez_tmp_41 = rob_val_3;
      5'b00100:
        casez_tmp_41 = rob_val_4;
      5'b00101:
        casez_tmp_41 = rob_val_5;
      5'b00110:
        casez_tmp_41 = rob_val_6;
      5'b00111:
        casez_tmp_41 = rob_val_7;
      5'b01000:
        casez_tmp_41 = rob_val_8;
      5'b01001:
        casez_tmp_41 = rob_val_9;
      5'b01010:
        casez_tmp_41 = rob_val_10;
      5'b01011:
        casez_tmp_41 = rob_val_11;
      5'b01100:
        casez_tmp_41 = rob_val_12;
      5'b01101:
        casez_tmp_41 = rob_val_13;
      5'b01110:
        casez_tmp_41 = rob_val_14;
      5'b01111:
        casez_tmp_41 = rob_val_15;
      5'b10000:
        casez_tmp_41 = rob_val_16;
      5'b10001:
        casez_tmp_41 = rob_val_17;
      5'b10010:
        casez_tmp_41 = rob_val_18;
      5'b10011:
        casez_tmp_41 = rob_val_19;
      5'b10100:
        casez_tmp_41 = rob_val_20;
      5'b10101:
        casez_tmp_41 = rob_val_21;
      5'b10110:
        casez_tmp_41 = rob_val_22;
      5'b10111:
        casez_tmp_41 = rob_val_23;
      5'b11000:
        casez_tmp_41 = rob_val_24;
      5'b11001:
        casez_tmp_41 = rob_val_25;
      5'b11010:
        casez_tmp_41 = rob_val_26;
      5'b11011:
        casez_tmp_41 = rob_val_27;
      5'b11100:
        casez_tmp_41 = rob_val_28;
      5'b11101:
        casez_tmp_41 = rob_val_29;
      5'b11110:
        casez_tmp_41 = rob_val_30;
      default:
        casez_tmp_41 = rob_val_31;
    endcase
  end // always @(*)
  reg         casez_tmp_42;
  always @(*) begin
    casez (io_wb_resps_1_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_42 = rob_bsy_0;
      5'b00001:
        casez_tmp_42 = rob_bsy_1;
      5'b00010:
        casez_tmp_42 = rob_bsy_2;
      5'b00011:
        casez_tmp_42 = rob_bsy_3;
      5'b00100:
        casez_tmp_42 = rob_bsy_4;
      5'b00101:
        casez_tmp_42 = rob_bsy_5;
      5'b00110:
        casez_tmp_42 = rob_bsy_6;
      5'b00111:
        casez_tmp_42 = rob_bsy_7;
      5'b01000:
        casez_tmp_42 = rob_bsy_8;
      5'b01001:
        casez_tmp_42 = rob_bsy_9;
      5'b01010:
        casez_tmp_42 = rob_bsy_10;
      5'b01011:
        casez_tmp_42 = rob_bsy_11;
      5'b01100:
        casez_tmp_42 = rob_bsy_12;
      5'b01101:
        casez_tmp_42 = rob_bsy_13;
      5'b01110:
        casez_tmp_42 = rob_bsy_14;
      5'b01111:
        casez_tmp_42 = rob_bsy_15;
      5'b10000:
        casez_tmp_42 = rob_bsy_16;
      5'b10001:
        casez_tmp_42 = rob_bsy_17;
      5'b10010:
        casez_tmp_42 = rob_bsy_18;
      5'b10011:
        casez_tmp_42 = rob_bsy_19;
      5'b10100:
        casez_tmp_42 = rob_bsy_20;
      5'b10101:
        casez_tmp_42 = rob_bsy_21;
      5'b10110:
        casez_tmp_42 = rob_bsy_22;
      5'b10111:
        casez_tmp_42 = rob_bsy_23;
      5'b11000:
        casez_tmp_42 = rob_bsy_24;
      5'b11001:
        casez_tmp_42 = rob_bsy_25;
      5'b11010:
        casez_tmp_42 = rob_bsy_26;
      5'b11011:
        casez_tmp_42 = rob_bsy_27;
      5'b11100:
        casez_tmp_42 = rob_bsy_28;
      5'b11101:
        casez_tmp_42 = rob_bsy_29;
      5'b11110:
        casez_tmp_42 = rob_bsy_30;
      default:
        casez_tmp_42 = rob_bsy_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_43;
  always @(*) begin
    casez (io_wb_resps_1_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_43 = rob_uop_0_pdst;
      5'b00001:
        casez_tmp_43 = rob_uop_1_pdst;
      5'b00010:
        casez_tmp_43 = rob_uop_2_pdst;
      5'b00011:
        casez_tmp_43 = rob_uop_3_pdst;
      5'b00100:
        casez_tmp_43 = rob_uop_4_pdst;
      5'b00101:
        casez_tmp_43 = rob_uop_5_pdst;
      5'b00110:
        casez_tmp_43 = rob_uop_6_pdst;
      5'b00111:
        casez_tmp_43 = rob_uop_7_pdst;
      5'b01000:
        casez_tmp_43 = rob_uop_8_pdst;
      5'b01001:
        casez_tmp_43 = rob_uop_9_pdst;
      5'b01010:
        casez_tmp_43 = rob_uop_10_pdst;
      5'b01011:
        casez_tmp_43 = rob_uop_11_pdst;
      5'b01100:
        casez_tmp_43 = rob_uop_12_pdst;
      5'b01101:
        casez_tmp_43 = rob_uop_13_pdst;
      5'b01110:
        casez_tmp_43 = rob_uop_14_pdst;
      5'b01111:
        casez_tmp_43 = rob_uop_15_pdst;
      5'b10000:
        casez_tmp_43 = rob_uop_16_pdst;
      5'b10001:
        casez_tmp_43 = rob_uop_17_pdst;
      5'b10010:
        casez_tmp_43 = rob_uop_18_pdst;
      5'b10011:
        casez_tmp_43 = rob_uop_19_pdst;
      5'b10100:
        casez_tmp_43 = rob_uop_20_pdst;
      5'b10101:
        casez_tmp_43 = rob_uop_21_pdst;
      5'b10110:
        casez_tmp_43 = rob_uop_22_pdst;
      5'b10111:
        casez_tmp_43 = rob_uop_23_pdst;
      5'b11000:
        casez_tmp_43 = rob_uop_24_pdst;
      5'b11001:
        casez_tmp_43 = rob_uop_25_pdst;
      5'b11010:
        casez_tmp_43 = rob_uop_26_pdst;
      5'b11011:
        casez_tmp_43 = rob_uop_27_pdst;
      5'b11100:
        casez_tmp_43 = rob_uop_28_pdst;
      5'b11101:
        casez_tmp_43 = rob_uop_29_pdst;
      5'b11110:
        casez_tmp_43 = rob_uop_30_pdst;
      default:
        casez_tmp_43 = rob_uop_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_44;
  always @(*) begin
    casez (io_wb_resps_1_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_44 = rob_uop_0_ldst_val;
      5'b00001:
        casez_tmp_44 = rob_uop_1_ldst_val;
      5'b00010:
        casez_tmp_44 = rob_uop_2_ldst_val;
      5'b00011:
        casez_tmp_44 = rob_uop_3_ldst_val;
      5'b00100:
        casez_tmp_44 = rob_uop_4_ldst_val;
      5'b00101:
        casez_tmp_44 = rob_uop_5_ldst_val;
      5'b00110:
        casez_tmp_44 = rob_uop_6_ldst_val;
      5'b00111:
        casez_tmp_44 = rob_uop_7_ldst_val;
      5'b01000:
        casez_tmp_44 = rob_uop_8_ldst_val;
      5'b01001:
        casez_tmp_44 = rob_uop_9_ldst_val;
      5'b01010:
        casez_tmp_44 = rob_uop_10_ldst_val;
      5'b01011:
        casez_tmp_44 = rob_uop_11_ldst_val;
      5'b01100:
        casez_tmp_44 = rob_uop_12_ldst_val;
      5'b01101:
        casez_tmp_44 = rob_uop_13_ldst_val;
      5'b01110:
        casez_tmp_44 = rob_uop_14_ldst_val;
      5'b01111:
        casez_tmp_44 = rob_uop_15_ldst_val;
      5'b10000:
        casez_tmp_44 = rob_uop_16_ldst_val;
      5'b10001:
        casez_tmp_44 = rob_uop_17_ldst_val;
      5'b10010:
        casez_tmp_44 = rob_uop_18_ldst_val;
      5'b10011:
        casez_tmp_44 = rob_uop_19_ldst_val;
      5'b10100:
        casez_tmp_44 = rob_uop_20_ldst_val;
      5'b10101:
        casez_tmp_44 = rob_uop_21_ldst_val;
      5'b10110:
        casez_tmp_44 = rob_uop_22_ldst_val;
      5'b10111:
        casez_tmp_44 = rob_uop_23_ldst_val;
      5'b11000:
        casez_tmp_44 = rob_uop_24_ldst_val;
      5'b11001:
        casez_tmp_44 = rob_uop_25_ldst_val;
      5'b11010:
        casez_tmp_44 = rob_uop_26_ldst_val;
      5'b11011:
        casez_tmp_44 = rob_uop_27_ldst_val;
      5'b11100:
        casez_tmp_44 = rob_uop_28_ldst_val;
      5'b11101:
        casez_tmp_44 = rob_uop_29_ldst_val;
      5'b11110:
        casez_tmp_44 = rob_uop_30_ldst_val;
      default:
        casez_tmp_44 = rob_uop_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_45;
  always @(*) begin
    casez (io_wb_resps_2_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_45 = rob_val_0;
      5'b00001:
        casez_tmp_45 = rob_val_1;
      5'b00010:
        casez_tmp_45 = rob_val_2;
      5'b00011:
        casez_tmp_45 = rob_val_3;
      5'b00100:
        casez_tmp_45 = rob_val_4;
      5'b00101:
        casez_tmp_45 = rob_val_5;
      5'b00110:
        casez_tmp_45 = rob_val_6;
      5'b00111:
        casez_tmp_45 = rob_val_7;
      5'b01000:
        casez_tmp_45 = rob_val_8;
      5'b01001:
        casez_tmp_45 = rob_val_9;
      5'b01010:
        casez_tmp_45 = rob_val_10;
      5'b01011:
        casez_tmp_45 = rob_val_11;
      5'b01100:
        casez_tmp_45 = rob_val_12;
      5'b01101:
        casez_tmp_45 = rob_val_13;
      5'b01110:
        casez_tmp_45 = rob_val_14;
      5'b01111:
        casez_tmp_45 = rob_val_15;
      5'b10000:
        casez_tmp_45 = rob_val_16;
      5'b10001:
        casez_tmp_45 = rob_val_17;
      5'b10010:
        casez_tmp_45 = rob_val_18;
      5'b10011:
        casez_tmp_45 = rob_val_19;
      5'b10100:
        casez_tmp_45 = rob_val_20;
      5'b10101:
        casez_tmp_45 = rob_val_21;
      5'b10110:
        casez_tmp_45 = rob_val_22;
      5'b10111:
        casez_tmp_45 = rob_val_23;
      5'b11000:
        casez_tmp_45 = rob_val_24;
      5'b11001:
        casez_tmp_45 = rob_val_25;
      5'b11010:
        casez_tmp_45 = rob_val_26;
      5'b11011:
        casez_tmp_45 = rob_val_27;
      5'b11100:
        casez_tmp_45 = rob_val_28;
      5'b11101:
        casez_tmp_45 = rob_val_29;
      5'b11110:
        casez_tmp_45 = rob_val_30;
      default:
        casez_tmp_45 = rob_val_31;
    endcase
  end // always @(*)
  reg         casez_tmp_46;
  always @(*) begin
    casez (io_wb_resps_2_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_46 = rob_bsy_0;
      5'b00001:
        casez_tmp_46 = rob_bsy_1;
      5'b00010:
        casez_tmp_46 = rob_bsy_2;
      5'b00011:
        casez_tmp_46 = rob_bsy_3;
      5'b00100:
        casez_tmp_46 = rob_bsy_4;
      5'b00101:
        casez_tmp_46 = rob_bsy_5;
      5'b00110:
        casez_tmp_46 = rob_bsy_6;
      5'b00111:
        casez_tmp_46 = rob_bsy_7;
      5'b01000:
        casez_tmp_46 = rob_bsy_8;
      5'b01001:
        casez_tmp_46 = rob_bsy_9;
      5'b01010:
        casez_tmp_46 = rob_bsy_10;
      5'b01011:
        casez_tmp_46 = rob_bsy_11;
      5'b01100:
        casez_tmp_46 = rob_bsy_12;
      5'b01101:
        casez_tmp_46 = rob_bsy_13;
      5'b01110:
        casez_tmp_46 = rob_bsy_14;
      5'b01111:
        casez_tmp_46 = rob_bsy_15;
      5'b10000:
        casez_tmp_46 = rob_bsy_16;
      5'b10001:
        casez_tmp_46 = rob_bsy_17;
      5'b10010:
        casez_tmp_46 = rob_bsy_18;
      5'b10011:
        casez_tmp_46 = rob_bsy_19;
      5'b10100:
        casez_tmp_46 = rob_bsy_20;
      5'b10101:
        casez_tmp_46 = rob_bsy_21;
      5'b10110:
        casez_tmp_46 = rob_bsy_22;
      5'b10111:
        casez_tmp_46 = rob_bsy_23;
      5'b11000:
        casez_tmp_46 = rob_bsy_24;
      5'b11001:
        casez_tmp_46 = rob_bsy_25;
      5'b11010:
        casez_tmp_46 = rob_bsy_26;
      5'b11011:
        casez_tmp_46 = rob_bsy_27;
      5'b11100:
        casez_tmp_46 = rob_bsy_28;
      5'b11101:
        casez_tmp_46 = rob_bsy_29;
      5'b11110:
        casez_tmp_46 = rob_bsy_30;
      default:
        casez_tmp_46 = rob_bsy_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_47;
  always @(*) begin
    casez (io_wb_resps_2_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_47 = rob_uop_0_pdst;
      5'b00001:
        casez_tmp_47 = rob_uop_1_pdst;
      5'b00010:
        casez_tmp_47 = rob_uop_2_pdst;
      5'b00011:
        casez_tmp_47 = rob_uop_3_pdst;
      5'b00100:
        casez_tmp_47 = rob_uop_4_pdst;
      5'b00101:
        casez_tmp_47 = rob_uop_5_pdst;
      5'b00110:
        casez_tmp_47 = rob_uop_6_pdst;
      5'b00111:
        casez_tmp_47 = rob_uop_7_pdst;
      5'b01000:
        casez_tmp_47 = rob_uop_8_pdst;
      5'b01001:
        casez_tmp_47 = rob_uop_9_pdst;
      5'b01010:
        casez_tmp_47 = rob_uop_10_pdst;
      5'b01011:
        casez_tmp_47 = rob_uop_11_pdst;
      5'b01100:
        casez_tmp_47 = rob_uop_12_pdst;
      5'b01101:
        casez_tmp_47 = rob_uop_13_pdst;
      5'b01110:
        casez_tmp_47 = rob_uop_14_pdst;
      5'b01111:
        casez_tmp_47 = rob_uop_15_pdst;
      5'b10000:
        casez_tmp_47 = rob_uop_16_pdst;
      5'b10001:
        casez_tmp_47 = rob_uop_17_pdst;
      5'b10010:
        casez_tmp_47 = rob_uop_18_pdst;
      5'b10011:
        casez_tmp_47 = rob_uop_19_pdst;
      5'b10100:
        casez_tmp_47 = rob_uop_20_pdst;
      5'b10101:
        casez_tmp_47 = rob_uop_21_pdst;
      5'b10110:
        casez_tmp_47 = rob_uop_22_pdst;
      5'b10111:
        casez_tmp_47 = rob_uop_23_pdst;
      5'b11000:
        casez_tmp_47 = rob_uop_24_pdst;
      5'b11001:
        casez_tmp_47 = rob_uop_25_pdst;
      5'b11010:
        casez_tmp_47 = rob_uop_26_pdst;
      5'b11011:
        casez_tmp_47 = rob_uop_27_pdst;
      5'b11100:
        casez_tmp_47 = rob_uop_28_pdst;
      5'b11101:
        casez_tmp_47 = rob_uop_29_pdst;
      5'b11110:
        casez_tmp_47 = rob_uop_30_pdst;
      default:
        casez_tmp_47 = rob_uop_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_48;
  always @(*) begin
    casez (io_wb_resps_2_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_48 = rob_uop_0_ldst_val;
      5'b00001:
        casez_tmp_48 = rob_uop_1_ldst_val;
      5'b00010:
        casez_tmp_48 = rob_uop_2_ldst_val;
      5'b00011:
        casez_tmp_48 = rob_uop_3_ldst_val;
      5'b00100:
        casez_tmp_48 = rob_uop_4_ldst_val;
      5'b00101:
        casez_tmp_48 = rob_uop_5_ldst_val;
      5'b00110:
        casez_tmp_48 = rob_uop_6_ldst_val;
      5'b00111:
        casez_tmp_48 = rob_uop_7_ldst_val;
      5'b01000:
        casez_tmp_48 = rob_uop_8_ldst_val;
      5'b01001:
        casez_tmp_48 = rob_uop_9_ldst_val;
      5'b01010:
        casez_tmp_48 = rob_uop_10_ldst_val;
      5'b01011:
        casez_tmp_48 = rob_uop_11_ldst_val;
      5'b01100:
        casez_tmp_48 = rob_uop_12_ldst_val;
      5'b01101:
        casez_tmp_48 = rob_uop_13_ldst_val;
      5'b01110:
        casez_tmp_48 = rob_uop_14_ldst_val;
      5'b01111:
        casez_tmp_48 = rob_uop_15_ldst_val;
      5'b10000:
        casez_tmp_48 = rob_uop_16_ldst_val;
      5'b10001:
        casez_tmp_48 = rob_uop_17_ldst_val;
      5'b10010:
        casez_tmp_48 = rob_uop_18_ldst_val;
      5'b10011:
        casez_tmp_48 = rob_uop_19_ldst_val;
      5'b10100:
        casez_tmp_48 = rob_uop_20_ldst_val;
      5'b10101:
        casez_tmp_48 = rob_uop_21_ldst_val;
      5'b10110:
        casez_tmp_48 = rob_uop_22_ldst_val;
      5'b10111:
        casez_tmp_48 = rob_uop_23_ldst_val;
      5'b11000:
        casez_tmp_48 = rob_uop_24_ldst_val;
      5'b11001:
        casez_tmp_48 = rob_uop_25_ldst_val;
      5'b11010:
        casez_tmp_48 = rob_uop_26_ldst_val;
      5'b11011:
        casez_tmp_48 = rob_uop_27_ldst_val;
      5'b11100:
        casez_tmp_48 = rob_uop_28_ldst_val;
      5'b11101:
        casez_tmp_48 = rob_uop_29_ldst_val;
      5'b11110:
        casez_tmp_48 = rob_uop_30_ldst_val;
      default:
        casez_tmp_48 = rob_uop_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_49;
  always @(*) begin
    casez (io_wb_resps_3_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_49 = rob_val_0;
      5'b00001:
        casez_tmp_49 = rob_val_1;
      5'b00010:
        casez_tmp_49 = rob_val_2;
      5'b00011:
        casez_tmp_49 = rob_val_3;
      5'b00100:
        casez_tmp_49 = rob_val_4;
      5'b00101:
        casez_tmp_49 = rob_val_5;
      5'b00110:
        casez_tmp_49 = rob_val_6;
      5'b00111:
        casez_tmp_49 = rob_val_7;
      5'b01000:
        casez_tmp_49 = rob_val_8;
      5'b01001:
        casez_tmp_49 = rob_val_9;
      5'b01010:
        casez_tmp_49 = rob_val_10;
      5'b01011:
        casez_tmp_49 = rob_val_11;
      5'b01100:
        casez_tmp_49 = rob_val_12;
      5'b01101:
        casez_tmp_49 = rob_val_13;
      5'b01110:
        casez_tmp_49 = rob_val_14;
      5'b01111:
        casez_tmp_49 = rob_val_15;
      5'b10000:
        casez_tmp_49 = rob_val_16;
      5'b10001:
        casez_tmp_49 = rob_val_17;
      5'b10010:
        casez_tmp_49 = rob_val_18;
      5'b10011:
        casez_tmp_49 = rob_val_19;
      5'b10100:
        casez_tmp_49 = rob_val_20;
      5'b10101:
        casez_tmp_49 = rob_val_21;
      5'b10110:
        casez_tmp_49 = rob_val_22;
      5'b10111:
        casez_tmp_49 = rob_val_23;
      5'b11000:
        casez_tmp_49 = rob_val_24;
      5'b11001:
        casez_tmp_49 = rob_val_25;
      5'b11010:
        casez_tmp_49 = rob_val_26;
      5'b11011:
        casez_tmp_49 = rob_val_27;
      5'b11100:
        casez_tmp_49 = rob_val_28;
      5'b11101:
        casez_tmp_49 = rob_val_29;
      5'b11110:
        casez_tmp_49 = rob_val_30;
      default:
        casez_tmp_49 = rob_val_31;
    endcase
  end // always @(*)
  reg         casez_tmp_50;
  always @(*) begin
    casez (io_wb_resps_3_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_50 = rob_bsy_0;
      5'b00001:
        casez_tmp_50 = rob_bsy_1;
      5'b00010:
        casez_tmp_50 = rob_bsy_2;
      5'b00011:
        casez_tmp_50 = rob_bsy_3;
      5'b00100:
        casez_tmp_50 = rob_bsy_4;
      5'b00101:
        casez_tmp_50 = rob_bsy_5;
      5'b00110:
        casez_tmp_50 = rob_bsy_6;
      5'b00111:
        casez_tmp_50 = rob_bsy_7;
      5'b01000:
        casez_tmp_50 = rob_bsy_8;
      5'b01001:
        casez_tmp_50 = rob_bsy_9;
      5'b01010:
        casez_tmp_50 = rob_bsy_10;
      5'b01011:
        casez_tmp_50 = rob_bsy_11;
      5'b01100:
        casez_tmp_50 = rob_bsy_12;
      5'b01101:
        casez_tmp_50 = rob_bsy_13;
      5'b01110:
        casez_tmp_50 = rob_bsy_14;
      5'b01111:
        casez_tmp_50 = rob_bsy_15;
      5'b10000:
        casez_tmp_50 = rob_bsy_16;
      5'b10001:
        casez_tmp_50 = rob_bsy_17;
      5'b10010:
        casez_tmp_50 = rob_bsy_18;
      5'b10011:
        casez_tmp_50 = rob_bsy_19;
      5'b10100:
        casez_tmp_50 = rob_bsy_20;
      5'b10101:
        casez_tmp_50 = rob_bsy_21;
      5'b10110:
        casez_tmp_50 = rob_bsy_22;
      5'b10111:
        casez_tmp_50 = rob_bsy_23;
      5'b11000:
        casez_tmp_50 = rob_bsy_24;
      5'b11001:
        casez_tmp_50 = rob_bsy_25;
      5'b11010:
        casez_tmp_50 = rob_bsy_26;
      5'b11011:
        casez_tmp_50 = rob_bsy_27;
      5'b11100:
        casez_tmp_50 = rob_bsy_28;
      5'b11101:
        casez_tmp_50 = rob_bsy_29;
      5'b11110:
        casez_tmp_50 = rob_bsy_30;
      default:
        casez_tmp_50 = rob_bsy_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_51;
  always @(*) begin
    casez (io_wb_resps_3_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_51 = rob_uop_0_pdst;
      5'b00001:
        casez_tmp_51 = rob_uop_1_pdst;
      5'b00010:
        casez_tmp_51 = rob_uop_2_pdst;
      5'b00011:
        casez_tmp_51 = rob_uop_3_pdst;
      5'b00100:
        casez_tmp_51 = rob_uop_4_pdst;
      5'b00101:
        casez_tmp_51 = rob_uop_5_pdst;
      5'b00110:
        casez_tmp_51 = rob_uop_6_pdst;
      5'b00111:
        casez_tmp_51 = rob_uop_7_pdst;
      5'b01000:
        casez_tmp_51 = rob_uop_8_pdst;
      5'b01001:
        casez_tmp_51 = rob_uop_9_pdst;
      5'b01010:
        casez_tmp_51 = rob_uop_10_pdst;
      5'b01011:
        casez_tmp_51 = rob_uop_11_pdst;
      5'b01100:
        casez_tmp_51 = rob_uop_12_pdst;
      5'b01101:
        casez_tmp_51 = rob_uop_13_pdst;
      5'b01110:
        casez_tmp_51 = rob_uop_14_pdst;
      5'b01111:
        casez_tmp_51 = rob_uop_15_pdst;
      5'b10000:
        casez_tmp_51 = rob_uop_16_pdst;
      5'b10001:
        casez_tmp_51 = rob_uop_17_pdst;
      5'b10010:
        casez_tmp_51 = rob_uop_18_pdst;
      5'b10011:
        casez_tmp_51 = rob_uop_19_pdst;
      5'b10100:
        casez_tmp_51 = rob_uop_20_pdst;
      5'b10101:
        casez_tmp_51 = rob_uop_21_pdst;
      5'b10110:
        casez_tmp_51 = rob_uop_22_pdst;
      5'b10111:
        casez_tmp_51 = rob_uop_23_pdst;
      5'b11000:
        casez_tmp_51 = rob_uop_24_pdst;
      5'b11001:
        casez_tmp_51 = rob_uop_25_pdst;
      5'b11010:
        casez_tmp_51 = rob_uop_26_pdst;
      5'b11011:
        casez_tmp_51 = rob_uop_27_pdst;
      5'b11100:
        casez_tmp_51 = rob_uop_28_pdst;
      5'b11101:
        casez_tmp_51 = rob_uop_29_pdst;
      5'b11110:
        casez_tmp_51 = rob_uop_30_pdst;
      default:
        casez_tmp_51 = rob_uop_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_52;
  always @(*) begin
    casez (io_wb_resps_3_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_52 = rob_uop_0_ldst_val;
      5'b00001:
        casez_tmp_52 = rob_uop_1_ldst_val;
      5'b00010:
        casez_tmp_52 = rob_uop_2_ldst_val;
      5'b00011:
        casez_tmp_52 = rob_uop_3_ldst_val;
      5'b00100:
        casez_tmp_52 = rob_uop_4_ldst_val;
      5'b00101:
        casez_tmp_52 = rob_uop_5_ldst_val;
      5'b00110:
        casez_tmp_52 = rob_uop_6_ldst_val;
      5'b00111:
        casez_tmp_52 = rob_uop_7_ldst_val;
      5'b01000:
        casez_tmp_52 = rob_uop_8_ldst_val;
      5'b01001:
        casez_tmp_52 = rob_uop_9_ldst_val;
      5'b01010:
        casez_tmp_52 = rob_uop_10_ldst_val;
      5'b01011:
        casez_tmp_52 = rob_uop_11_ldst_val;
      5'b01100:
        casez_tmp_52 = rob_uop_12_ldst_val;
      5'b01101:
        casez_tmp_52 = rob_uop_13_ldst_val;
      5'b01110:
        casez_tmp_52 = rob_uop_14_ldst_val;
      5'b01111:
        casez_tmp_52 = rob_uop_15_ldst_val;
      5'b10000:
        casez_tmp_52 = rob_uop_16_ldst_val;
      5'b10001:
        casez_tmp_52 = rob_uop_17_ldst_val;
      5'b10010:
        casez_tmp_52 = rob_uop_18_ldst_val;
      5'b10011:
        casez_tmp_52 = rob_uop_19_ldst_val;
      5'b10100:
        casez_tmp_52 = rob_uop_20_ldst_val;
      5'b10101:
        casez_tmp_52 = rob_uop_21_ldst_val;
      5'b10110:
        casez_tmp_52 = rob_uop_22_ldst_val;
      5'b10111:
        casez_tmp_52 = rob_uop_23_ldst_val;
      5'b11000:
        casez_tmp_52 = rob_uop_24_ldst_val;
      5'b11001:
        casez_tmp_52 = rob_uop_25_ldst_val;
      5'b11010:
        casez_tmp_52 = rob_uop_26_ldst_val;
      5'b11011:
        casez_tmp_52 = rob_uop_27_ldst_val;
      5'b11100:
        casez_tmp_52 = rob_uop_28_ldst_val;
      5'b11101:
        casez_tmp_52 = rob_uop_29_ldst_val;
      5'b11110:
        casez_tmp_52 = rob_uop_30_ldst_val;
      default:
        casez_tmp_52 = rob_uop_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_53;
  always @(*) begin
    casez (io_wb_resps_4_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_53 = rob_val_0;
      5'b00001:
        casez_tmp_53 = rob_val_1;
      5'b00010:
        casez_tmp_53 = rob_val_2;
      5'b00011:
        casez_tmp_53 = rob_val_3;
      5'b00100:
        casez_tmp_53 = rob_val_4;
      5'b00101:
        casez_tmp_53 = rob_val_5;
      5'b00110:
        casez_tmp_53 = rob_val_6;
      5'b00111:
        casez_tmp_53 = rob_val_7;
      5'b01000:
        casez_tmp_53 = rob_val_8;
      5'b01001:
        casez_tmp_53 = rob_val_9;
      5'b01010:
        casez_tmp_53 = rob_val_10;
      5'b01011:
        casez_tmp_53 = rob_val_11;
      5'b01100:
        casez_tmp_53 = rob_val_12;
      5'b01101:
        casez_tmp_53 = rob_val_13;
      5'b01110:
        casez_tmp_53 = rob_val_14;
      5'b01111:
        casez_tmp_53 = rob_val_15;
      5'b10000:
        casez_tmp_53 = rob_val_16;
      5'b10001:
        casez_tmp_53 = rob_val_17;
      5'b10010:
        casez_tmp_53 = rob_val_18;
      5'b10011:
        casez_tmp_53 = rob_val_19;
      5'b10100:
        casez_tmp_53 = rob_val_20;
      5'b10101:
        casez_tmp_53 = rob_val_21;
      5'b10110:
        casez_tmp_53 = rob_val_22;
      5'b10111:
        casez_tmp_53 = rob_val_23;
      5'b11000:
        casez_tmp_53 = rob_val_24;
      5'b11001:
        casez_tmp_53 = rob_val_25;
      5'b11010:
        casez_tmp_53 = rob_val_26;
      5'b11011:
        casez_tmp_53 = rob_val_27;
      5'b11100:
        casez_tmp_53 = rob_val_28;
      5'b11101:
        casez_tmp_53 = rob_val_29;
      5'b11110:
        casez_tmp_53 = rob_val_30;
      default:
        casez_tmp_53 = rob_val_31;
    endcase
  end // always @(*)
  reg         casez_tmp_54;
  always @(*) begin
    casez (io_wb_resps_4_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_54 = rob_bsy_0;
      5'b00001:
        casez_tmp_54 = rob_bsy_1;
      5'b00010:
        casez_tmp_54 = rob_bsy_2;
      5'b00011:
        casez_tmp_54 = rob_bsy_3;
      5'b00100:
        casez_tmp_54 = rob_bsy_4;
      5'b00101:
        casez_tmp_54 = rob_bsy_5;
      5'b00110:
        casez_tmp_54 = rob_bsy_6;
      5'b00111:
        casez_tmp_54 = rob_bsy_7;
      5'b01000:
        casez_tmp_54 = rob_bsy_8;
      5'b01001:
        casez_tmp_54 = rob_bsy_9;
      5'b01010:
        casez_tmp_54 = rob_bsy_10;
      5'b01011:
        casez_tmp_54 = rob_bsy_11;
      5'b01100:
        casez_tmp_54 = rob_bsy_12;
      5'b01101:
        casez_tmp_54 = rob_bsy_13;
      5'b01110:
        casez_tmp_54 = rob_bsy_14;
      5'b01111:
        casez_tmp_54 = rob_bsy_15;
      5'b10000:
        casez_tmp_54 = rob_bsy_16;
      5'b10001:
        casez_tmp_54 = rob_bsy_17;
      5'b10010:
        casez_tmp_54 = rob_bsy_18;
      5'b10011:
        casez_tmp_54 = rob_bsy_19;
      5'b10100:
        casez_tmp_54 = rob_bsy_20;
      5'b10101:
        casez_tmp_54 = rob_bsy_21;
      5'b10110:
        casez_tmp_54 = rob_bsy_22;
      5'b10111:
        casez_tmp_54 = rob_bsy_23;
      5'b11000:
        casez_tmp_54 = rob_bsy_24;
      5'b11001:
        casez_tmp_54 = rob_bsy_25;
      5'b11010:
        casez_tmp_54 = rob_bsy_26;
      5'b11011:
        casez_tmp_54 = rob_bsy_27;
      5'b11100:
        casez_tmp_54 = rob_bsy_28;
      5'b11101:
        casez_tmp_54 = rob_bsy_29;
      5'b11110:
        casez_tmp_54 = rob_bsy_30;
      default:
        casez_tmp_54 = rob_bsy_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_55;
  always @(*) begin
    casez (io_wb_resps_4_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_55 = rob_uop_0_pdst;
      5'b00001:
        casez_tmp_55 = rob_uop_1_pdst;
      5'b00010:
        casez_tmp_55 = rob_uop_2_pdst;
      5'b00011:
        casez_tmp_55 = rob_uop_3_pdst;
      5'b00100:
        casez_tmp_55 = rob_uop_4_pdst;
      5'b00101:
        casez_tmp_55 = rob_uop_5_pdst;
      5'b00110:
        casez_tmp_55 = rob_uop_6_pdst;
      5'b00111:
        casez_tmp_55 = rob_uop_7_pdst;
      5'b01000:
        casez_tmp_55 = rob_uop_8_pdst;
      5'b01001:
        casez_tmp_55 = rob_uop_9_pdst;
      5'b01010:
        casez_tmp_55 = rob_uop_10_pdst;
      5'b01011:
        casez_tmp_55 = rob_uop_11_pdst;
      5'b01100:
        casez_tmp_55 = rob_uop_12_pdst;
      5'b01101:
        casez_tmp_55 = rob_uop_13_pdst;
      5'b01110:
        casez_tmp_55 = rob_uop_14_pdst;
      5'b01111:
        casez_tmp_55 = rob_uop_15_pdst;
      5'b10000:
        casez_tmp_55 = rob_uop_16_pdst;
      5'b10001:
        casez_tmp_55 = rob_uop_17_pdst;
      5'b10010:
        casez_tmp_55 = rob_uop_18_pdst;
      5'b10011:
        casez_tmp_55 = rob_uop_19_pdst;
      5'b10100:
        casez_tmp_55 = rob_uop_20_pdst;
      5'b10101:
        casez_tmp_55 = rob_uop_21_pdst;
      5'b10110:
        casez_tmp_55 = rob_uop_22_pdst;
      5'b10111:
        casez_tmp_55 = rob_uop_23_pdst;
      5'b11000:
        casez_tmp_55 = rob_uop_24_pdst;
      5'b11001:
        casez_tmp_55 = rob_uop_25_pdst;
      5'b11010:
        casez_tmp_55 = rob_uop_26_pdst;
      5'b11011:
        casez_tmp_55 = rob_uop_27_pdst;
      5'b11100:
        casez_tmp_55 = rob_uop_28_pdst;
      5'b11101:
        casez_tmp_55 = rob_uop_29_pdst;
      5'b11110:
        casez_tmp_55 = rob_uop_30_pdst;
      default:
        casez_tmp_55 = rob_uop_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_56;
  always @(*) begin
    casez (io_wb_resps_4_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_56 = rob_uop_0_ldst_val;
      5'b00001:
        casez_tmp_56 = rob_uop_1_ldst_val;
      5'b00010:
        casez_tmp_56 = rob_uop_2_ldst_val;
      5'b00011:
        casez_tmp_56 = rob_uop_3_ldst_val;
      5'b00100:
        casez_tmp_56 = rob_uop_4_ldst_val;
      5'b00101:
        casez_tmp_56 = rob_uop_5_ldst_val;
      5'b00110:
        casez_tmp_56 = rob_uop_6_ldst_val;
      5'b00111:
        casez_tmp_56 = rob_uop_7_ldst_val;
      5'b01000:
        casez_tmp_56 = rob_uop_8_ldst_val;
      5'b01001:
        casez_tmp_56 = rob_uop_9_ldst_val;
      5'b01010:
        casez_tmp_56 = rob_uop_10_ldst_val;
      5'b01011:
        casez_tmp_56 = rob_uop_11_ldst_val;
      5'b01100:
        casez_tmp_56 = rob_uop_12_ldst_val;
      5'b01101:
        casez_tmp_56 = rob_uop_13_ldst_val;
      5'b01110:
        casez_tmp_56 = rob_uop_14_ldst_val;
      5'b01111:
        casez_tmp_56 = rob_uop_15_ldst_val;
      5'b10000:
        casez_tmp_56 = rob_uop_16_ldst_val;
      5'b10001:
        casez_tmp_56 = rob_uop_17_ldst_val;
      5'b10010:
        casez_tmp_56 = rob_uop_18_ldst_val;
      5'b10011:
        casez_tmp_56 = rob_uop_19_ldst_val;
      5'b10100:
        casez_tmp_56 = rob_uop_20_ldst_val;
      5'b10101:
        casez_tmp_56 = rob_uop_21_ldst_val;
      5'b10110:
        casez_tmp_56 = rob_uop_22_ldst_val;
      5'b10111:
        casez_tmp_56 = rob_uop_23_ldst_val;
      5'b11000:
        casez_tmp_56 = rob_uop_24_ldst_val;
      5'b11001:
        casez_tmp_56 = rob_uop_25_ldst_val;
      5'b11010:
        casez_tmp_56 = rob_uop_26_ldst_val;
      5'b11011:
        casez_tmp_56 = rob_uop_27_ldst_val;
      5'b11100:
        casez_tmp_56 = rob_uop_28_ldst_val;
      5'b11101:
        casez_tmp_56 = rob_uop_29_ldst_val;
      5'b11110:
        casez_tmp_56 = rob_uop_30_ldst_val;
      default:
        casez_tmp_56 = rob_uop_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_57;
  always @(*) begin
    casez (io_wb_resps_5_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_57 = rob_val_0;
      5'b00001:
        casez_tmp_57 = rob_val_1;
      5'b00010:
        casez_tmp_57 = rob_val_2;
      5'b00011:
        casez_tmp_57 = rob_val_3;
      5'b00100:
        casez_tmp_57 = rob_val_4;
      5'b00101:
        casez_tmp_57 = rob_val_5;
      5'b00110:
        casez_tmp_57 = rob_val_6;
      5'b00111:
        casez_tmp_57 = rob_val_7;
      5'b01000:
        casez_tmp_57 = rob_val_8;
      5'b01001:
        casez_tmp_57 = rob_val_9;
      5'b01010:
        casez_tmp_57 = rob_val_10;
      5'b01011:
        casez_tmp_57 = rob_val_11;
      5'b01100:
        casez_tmp_57 = rob_val_12;
      5'b01101:
        casez_tmp_57 = rob_val_13;
      5'b01110:
        casez_tmp_57 = rob_val_14;
      5'b01111:
        casez_tmp_57 = rob_val_15;
      5'b10000:
        casez_tmp_57 = rob_val_16;
      5'b10001:
        casez_tmp_57 = rob_val_17;
      5'b10010:
        casez_tmp_57 = rob_val_18;
      5'b10011:
        casez_tmp_57 = rob_val_19;
      5'b10100:
        casez_tmp_57 = rob_val_20;
      5'b10101:
        casez_tmp_57 = rob_val_21;
      5'b10110:
        casez_tmp_57 = rob_val_22;
      5'b10111:
        casez_tmp_57 = rob_val_23;
      5'b11000:
        casez_tmp_57 = rob_val_24;
      5'b11001:
        casez_tmp_57 = rob_val_25;
      5'b11010:
        casez_tmp_57 = rob_val_26;
      5'b11011:
        casez_tmp_57 = rob_val_27;
      5'b11100:
        casez_tmp_57 = rob_val_28;
      5'b11101:
        casez_tmp_57 = rob_val_29;
      5'b11110:
        casez_tmp_57 = rob_val_30;
      default:
        casez_tmp_57 = rob_val_31;
    endcase
  end // always @(*)
  reg         casez_tmp_58;
  always @(*) begin
    casez (io_wb_resps_5_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_58 = rob_bsy_0;
      5'b00001:
        casez_tmp_58 = rob_bsy_1;
      5'b00010:
        casez_tmp_58 = rob_bsy_2;
      5'b00011:
        casez_tmp_58 = rob_bsy_3;
      5'b00100:
        casez_tmp_58 = rob_bsy_4;
      5'b00101:
        casez_tmp_58 = rob_bsy_5;
      5'b00110:
        casez_tmp_58 = rob_bsy_6;
      5'b00111:
        casez_tmp_58 = rob_bsy_7;
      5'b01000:
        casez_tmp_58 = rob_bsy_8;
      5'b01001:
        casez_tmp_58 = rob_bsy_9;
      5'b01010:
        casez_tmp_58 = rob_bsy_10;
      5'b01011:
        casez_tmp_58 = rob_bsy_11;
      5'b01100:
        casez_tmp_58 = rob_bsy_12;
      5'b01101:
        casez_tmp_58 = rob_bsy_13;
      5'b01110:
        casez_tmp_58 = rob_bsy_14;
      5'b01111:
        casez_tmp_58 = rob_bsy_15;
      5'b10000:
        casez_tmp_58 = rob_bsy_16;
      5'b10001:
        casez_tmp_58 = rob_bsy_17;
      5'b10010:
        casez_tmp_58 = rob_bsy_18;
      5'b10011:
        casez_tmp_58 = rob_bsy_19;
      5'b10100:
        casez_tmp_58 = rob_bsy_20;
      5'b10101:
        casez_tmp_58 = rob_bsy_21;
      5'b10110:
        casez_tmp_58 = rob_bsy_22;
      5'b10111:
        casez_tmp_58 = rob_bsy_23;
      5'b11000:
        casez_tmp_58 = rob_bsy_24;
      5'b11001:
        casez_tmp_58 = rob_bsy_25;
      5'b11010:
        casez_tmp_58 = rob_bsy_26;
      5'b11011:
        casez_tmp_58 = rob_bsy_27;
      5'b11100:
        casez_tmp_58 = rob_bsy_28;
      5'b11101:
        casez_tmp_58 = rob_bsy_29;
      5'b11110:
        casez_tmp_58 = rob_bsy_30;
      default:
        casez_tmp_58 = rob_bsy_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_59;
  always @(*) begin
    casez (io_wb_resps_5_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_59 = rob_uop_0_pdst;
      5'b00001:
        casez_tmp_59 = rob_uop_1_pdst;
      5'b00010:
        casez_tmp_59 = rob_uop_2_pdst;
      5'b00011:
        casez_tmp_59 = rob_uop_3_pdst;
      5'b00100:
        casez_tmp_59 = rob_uop_4_pdst;
      5'b00101:
        casez_tmp_59 = rob_uop_5_pdst;
      5'b00110:
        casez_tmp_59 = rob_uop_6_pdst;
      5'b00111:
        casez_tmp_59 = rob_uop_7_pdst;
      5'b01000:
        casez_tmp_59 = rob_uop_8_pdst;
      5'b01001:
        casez_tmp_59 = rob_uop_9_pdst;
      5'b01010:
        casez_tmp_59 = rob_uop_10_pdst;
      5'b01011:
        casez_tmp_59 = rob_uop_11_pdst;
      5'b01100:
        casez_tmp_59 = rob_uop_12_pdst;
      5'b01101:
        casez_tmp_59 = rob_uop_13_pdst;
      5'b01110:
        casez_tmp_59 = rob_uop_14_pdst;
      5'b01111:
        casez_tmp_59 = rob_uop_15_pdst;
      5'b10000:
        casez_tmp_59 = rob_uop_16_pdst;
      5'b10001:
        casez_tmp_59 = rob_uop_17_pdst;
      5'b10010:
        casez_tmp_59 = rob_uop_18_pdst;
      5'b10011:
        casez_tmp_59 = rob_uop_19_pdst;
      5'b10100:
        casez_tmp_59 = rob_uop_20_pdst;
      5'b10101:
        casez_tmp_59 = rob_uop_21_pdst;
      5'b10110:
        casez_tmp_59 = rob_uop_22_pdst;
      5'b10111:
        casez_tmp_59 = rob_uop_23_pdst;
      5'b11000:
        casez_tmp_59 = rob_uop_24_pdst;
      5'b11001:
        casez_tmp_59 = rob_uop_25_pdst;
      5'b11010:
        casez_tmp_59 = rob_uop_26_pdst;
      5'b11011:
        casez_tmp_59 = rob_uop_27_pdst;
      5'b11100:
        casez_tmp_59 = rob_uop_28_pdst;
      5'b11101:
        casez_tmp_59 = rob_uop_29_pdst;
      5'b11110:
        casez_tmp_59 = rob_uop_30_pdst;
      default:
        casez_tmp_59 = rob_uop_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_60;
  always @(*) begin
    casez (io_wb_resps_5_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_60 = rob_uop_0_ldst_val;
      5'b00001:
        casez_tmp_60 = rob_uop_1_ldst_val;
      5'b00010:
        casez_tmp_60 = rob_uop_2_ldst_val;
      5'b00011:
        casez_tmp_60 = rob_uop_3_ldst_val;
      5'b00100:
        casez_tmp_60 = rob_uop_4_ldst_val;
      5'b00101:
        casez_tmp_60 = rob_uop_5_ldst_val;
      5'b00110:
        casez_tmp_60 = rob_uop_6_ldst_val;
      5'b00111:
        casez_tmp_60 = rob_uop_7_ldst_val;
      5'b01000:
        casez_tmp_60 = rob_uop_8_ldst_val;
      5'b01001:
        casez_tmp_60 = rob_uop_9_ldst_val;
      5'b01010:
        casez_tmp_60 = rob_uop_10_ldst_val;
      5'b01011:
        casez_tmp_60 = rob_uop_11_ldst_val;
      5'b01100:
        casez_tmp_60 = rob_uop_12_ldst_val;
      5'b01101:
        casez_tmp_60 = rob_uop_13_ldst_val;
      5'b01110:
        casez_tmp_60 = rob_uop_14_ldst_val;
      5'b01111:
        casez_tmp_60 = rob_uop_15_ldst_val;
      5'b10000:
        casez_tmp_60 = rob_uop_16_ldst_val;
      5'b10001:
        casez_tmp_60 = rob_uop_17_ldst_val;
      5'b10010:
        casez_tmp_60 = rob_uop_18_ldst_val;
      5'b10011:
        casez_tmp_60 = rob_uop_19_ldst_val;
      5'b10100:
        casez_tmp_60 = rob_uop_20_ldst_val;
      5'b10101:
        casez_tmp_60 = rob_uop_21_ldst_val;
      5'b10110:
        casez_tmp_60 = rob_uop_22_ldst_val;
      5'b10111:
        casez_tmp_60 = rob_uop_23_ldst_val;
      5'b11000:
        casez_tmp_60 = rob_uop_24_ldst_val;
      5'b11001:
        casez_tmp_60 = rob_uop_25_ldst_val;
      5'b11010:
        casez_tmp_60 = rob_uop_26_ldst_val;
      5'b11011:
        casez_tmp_60 = rob_uop_27_ldst_val;
      5'b11100:
        casez_tmp_60 = rob_uop_28_ldst_val;
      5'b11101:
        casez_tmp_60 = rob_uop_29_ldst_val;
      5'b11110:
        casez_tmp_60 = rob_uop_30_ldst_val;
      default:
        casez_tmp_60 = rob_uop_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_61;
  always @(*) begin
    casez (io_wb_resps_6_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_61 = rob_val_0;
      5'b00001:
        casez_tmp_61 = rob_val_1;
      5'b00010:
        casez_tmp_61 = rob_val_2;
      5'b00011:
        casez_tmp_61 = rob_val_3;
      5'b00100:
        casez_tmp_61 = rob_val_4;
      5'b00101:
        casez_tmp_61 = rob_val_5;
      5'b00110:
        casez_tmp_61 = rob_val_6;
      5'b00111:
        casez_tmp_61 = rob_val_7;
      5'b01000:
        casez_tmp_61 = rob_val_8;
      5'b01001:
        casez_tmp_61 = rob_val_9;
      5'b01010:
        casez_tmp_61 = rob_val_10;
      5'b01011:
        casez_tmp_61 = rob_val_11;
      5'b01100:
        casez_tmp_61 = rob_val_12;
      5'b01101:
        casez_tmp_61 = rob_val_13;
      5'b01110:
        casez_tmp_61 = rob_val_14;
      5'b01111:
        casez_tmp_61 = rob_val_15;
      5'b10000:
        casez_tmp_61 = rob_val_16;
      5'b10001:
        casez_tmp_61 = rob_val_17;
      5'b10010:
        casez_tmp_61 = rob_val_18;
      5'b10011:
        casez_tmp_61 = rob_val_19;
      5'b10100:
        casez_tmp_61 = rob_val_20;
      5'b10101:
        casez_tmp_61 = rob_val_21;
      5'b10110:
        casez_tmp_61 = rob_val_22;
      5'b10111:
        casez_tmp_61 = rob_val_23;
      5'b11000:
        casez_tmp_61 = rob_val_24;
      5'b11001:
        casez_tmp_61 = rob_val_25;
      5'b11010:
        casez_tmp_61 = rob_val_26;
      5'b11011:
        casez_tmp_61 = rob_val_27;
      5'b11100:
        casez_tmp_61 = rob_val_28;
      5'b11101:
        casez_tmp_61 = rob_val_29;
      5'b11110:
        casez_tmp_61 = rob_val_30;
      default:
        casez_tmp_61 = rob_val_31;
    endcase
  end // always @(*)
  reg         casez_tmp_62;
  always @(*) begin
    casez (io_wb_resps_6_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_62 = rob_bsy_0;
      5'b00001:
        casez_tmp_62 = rob_bsy_1;
      5'b00010:
        casez_tmp_62 = rob_bsy_2;
      5'b00011:
        casez_tmp_62 = rob_bsy_3;
      5'b00100:
        casez_tmp_62 = rob_bsy_4;
      5'b00101:
        casez_tmp_62 = rob_bsy_5;
      5'b00110:
        casez_tmp_62 = rob_bsy_6;
      5'b00111:
        casez_tmp_62 = rob_bsy_7;
      5'b01000:
        casez_tmp_62 = rob_bsy_8;
      5'b01001:
        casez_tmp_62 = rob_bsy_9;
      5'b01010:
        casez_tmp_62 = rob_bsy_10;
      5'b01011:
        casez_tmp_62 = rob_bsy_11;
      5'b01100:
        casez_tmp_62 = rob_bsy_12;
      5'b01101:
        casez_tmp_62 = rob_bsy_13;
      5'b01110:
        casez_tmp_62 = rob_bsy_14;
      5'b01111:
        casez_tmp_62 = rob_bsy_15;
      5'b10000:
        casez_tmp_62 = rob_bsy_16;
      5'b10001:
        casez_tmp_62 = rob_bsy_17;
      5'b10010:
        casez_tmp_62 = rob_bsy_18;
      5'b10011:
        casez_tmp_62 = rob_bsy_19;
      5'b10100:
        casez_tmp_62 = rob_bsy_20;
      5'b10101:
        casez_tmp_62 = rob_bsy_21;
      5'b10110:
        casez_tmp_62 = rob_bsy_22;
      5'b10111:
        casez_tmp_62 = rob_bsy_23;
      5'b11000:
        casez_tmp_62 = rob_bsy_24;
      5'b11001:
        casez_tmp_62 = rob_bsy_25;
      5'b11010:
        casez_tmp_62 = rob_bsy_26;
      5'b11011:
        casez_tmp_62 = rob_bsy_27;
      5'b11100:
        casez_tmp_62 = rob_bsy_28;
      5'b11101:
        casez_tmp_62 = rob_bsy_29;
      5'b11110:
        casez_tmp_62 = rob_bsy_30;
      default:
        casez_tmp_62 = rob_bsy_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_63;
  always @(*) begin
    casez (io_wb_resps_6_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_63 = rob_uop_0_pdst;
      5'b00001:
        casez_tmp_63 = rob_uop_1_pdst;
      5'b00010:
        casez_tmp_63 = rob_uop_2_pdst;
      5'b00011:
        casez_tmp_63 = rob_uop_3_pdst;
      5'b00100:
        casez_tmp_63 = rob_uop_4_pdst;
      5'b00101:
        casez_tmp_63 = rob_uop_5_pdst;
      5'b00110:
        casez_tmp_63 = rob_uop_6_pdst;
      5'b00111:
        casez_tmp_63 = rob_uop_7_pdst;
      5'b01000:
        casez_tmp_63 = rob_uop_8_pdst;
      5'b01001:
        casez_tmp_63 = rob_uop_9_pdst;
      5'b01010:
        casez_tmp_63 = rob_uop_10_pdst;
      5'b01011:
        casez_tmp_63 = rob_uop_11_pdst;
      5'b01100:
        casez_tmp_63 = rob_uop_12_pdst;
      5'b01101:
        casez_tmp_63 = rob_uop_13_pdst;
      5'b01110:
        casez_tmp_63 = rob_uop_14_pdst;
      5'b01111:
        casez_tmp_63 = rob_uop_15_pdst;
      5'b10000:
        casez_tmp_63 = rob_uop_16_pdst;
      5'b10001:
        casez_tmp_63 = rob_uop_17_pdst;
      5'b10010:
        casez_tmp_63 = rob_uop_18_pdst;
      5'b10011:
        casez_tmp_63 = rob_uop_19_pdst;
      5'b10100:
        casez_tmp_63 = rob_uop_20_pdst;
      5'b10101:
        casez_tmp_63 = rob_uop_21_pdst;
      5'b10110:
        casez_tmp_63 = rob_uop_22_pdst;
      5'b10111:
        casez_tmp_63 = rob_uop_23_pdst;
      5'b11000:
        casez_tmp_63 = rob_uop_24_pdst;
      5'b11001:
        casez_tmp_63 = rob_uop_25_pdst;
      5'b11010:
        casez_tmp_63 = rob_uop_26_pdst;
      5'b11011:
        casez_tmp_63 = rob_uop_27_pdst;
      5'b11100:
        casez_tmp_63 = rob_uop_28_pdst;
      5'b11101:
        casez_tmp_63 = rob_uop_29_pdst;
      5'b11110:
        casez_tmp_63 = rob_uop_30_pdst;
      default:
        casez_tmp_63 = rob_uop_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_64;
  always @(*) begin
    casez (io_wb_resps_6_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_64 = rob_uop_0_ldst_val;
      5'b00001:
        casez_tmp_64 = rob_uop_1_ldst_val;
      5'b00010:
        casez_tmp_64 = rob_uop_2_ldst_val;
      5'b00011:
        casez_tmp_64 = rob_uop_3_ldst_val;
      5'b00100:
        casez_tmp_64 = rob_uop_4_ldst_val;
      5'b00101:
        casez_tmp_64 = rob_uop_5_ldst_val;
      5'b00110:
        casez_tmp_64 = rob_uop_6_ldst_val;
      5'b00111:
        casez_tmp_64 = rob_uop_7_ldst_val;
      5'b01000:
        casez_tmp_64 = rob_uop_8_ldst_val;
      5'b01001:
        casez_tmp_64 = rob_uop_9_ldst_val;
      5'b01010:
        casez_tmp_64 = rob_uop_10_ldst_val;
      5'b01011:
        casez_tmp_64 = rob_uop_11_ldst_val;
      5'b01100:
        casez_tmp_64 = rob_uop_12_ldst_val;
      5'b01101:
        casez_tmp_64 = rob_uop_13_ldst_val;
      5'b01110:
        casez_tmp_64 = rob_uop_14_ldst_val;
      5'b01111:
        casez_tmp_64 = rob_uop_15_ldst_val;
      5'b10000:
        casez_tmp_64 = rob_uop_16_ldst_val;
      5'b10001:
        casez_tmp_64 = rob_uop_17_ldst_val;
      5'b10010:
        casez_tmp_64 = rob_uop_18_ldst_val;
      5'b10011:
        casez_tmp_64 = rob_uop_19_ldst_val;
      5'b10100:
        casez_tmp_64 = rob_uop_20_ldst_val;
      5'b10101:
        casez_tmp_64 = rob_uop_21_ldst_val;
      5'b10110:
        casez_tmp_64 = rob_uop_22_ldst_val;
      5'b10111:
        casez_tmp_64 = rob_uop_23_ldst_val;
      5'b11000:
        casez_tmp_64 = rob_uop_24_ldst_val;
      5'b11001:
        casez_tmp_64 = rob_uop_25_ldst_val;
      5'b11010:
        casez_tmp_64 = rob_uop_26_ldst_val;
      5'b11011:
        casez_tmp_64 = rob_uop_27_ldst_val;
      5'b11100:
        casez_tmp_64 = rob_uop_28_ldst_val;
      5'b11101:
        casez_tmp_64 = rob_uop_29_ldst_val;
      5'b11110:
        casez_tmp_64 = rob_uop_30_ldst_val;
      default:
        casez_tmp_64 = rob_uop_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_65;
  always @(*) begin
    casez (io_wb_resps_7_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_65 = rob_val_0;
      5'b00001:
        casez_tmp_65 = rob_val_1;
      5'b00010:
        casez_tmp_65 = rob_val_2;
      5'b00011:
        casez_tmp_65 = rob_val_3;
      5'b00100:
        casez_tmp_65 = rob_val_4;
      5'b00101:
        casez_tmp_65 = rob_val_5;
      5'b00110:
        casez_tmp_65 = rob_val_6;
      5'b00111:
        casez_tmp_65 = rob_val_7;
      5'b01000:
        casez_tmp_65 = rob_val_8;
      5'b01001:
        casez_tmp_65 = rob_val_9;
      5'b01010:
        casez_tmp_65 = rob_val_10;
      5'b01011:
        casez_tmp_65 = rob_val_11;
      5'b01100:
        casez_tmp_65 = rob_val_12;
      5'b01101:
        casez_tmp_65 = rob_val_13;
      5'b01110:
        casez_tmp_65 = rob_val_14;
      5'b01111:
        casez_tmp_65 = rob_val_15;
      5'b10000:
        casez_tmp_65 = rob_val_16;
      5'b10001:
        casez_tmp_65 = rob_val_17;
      5'b10010:
        casez_tmp_65 = rob_val_18;
      5'b10011:
        casez_tmp_65 = rob_val_19;
      5'b10100:
        casez_tmp_65 = rob_val_20;
      5'b10101:
        casez_tmp_65 = rob_val_21;
      5'b10110:
        casez_tmp_65 = rob_val_22;
      5'b10111:
        casez_tmp_65 = rob_val_23;
      5'b11000:
        casez_tmp_65 = rob_val_24;
      5'b11001:
        casez_tmp_65 = rob_val_25;
      5'b11010:
        casez_tmp_65 = rob_val_26;
      5'b11011:
        casez_tmp_65 = rob_val_27;
      5'b11100:
        casez_tmp_65 = rob_val_28;
      5'b11101:
        casez_tmp_65 = rob_val_29;
      5'b11110:
        casez_tmp_65 = rob_val_30;
      default:
        casez_tmp_65 = rob_val_31;
    endcase
  end // always @(*)
  reg         casez_tmp_66;
  always @(*) begin
    casez (io_wb_resps_7_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_66 = rob_bsy_0;
      5'b00001:
        casez_tmp_66 = rob_bsy_1;
      5'b00010:
        casez_tmp_66 = rob_bsy_2;
      5'b00011:
        casez_tmp_66 = rob_bsy_3;
      5'b00100:
        casez_tmp_66 = rob_bsy_4;
      5'b00101:
        casez_tmp_66 = rob_bsy_5;
      5'b00110:
        casez_tmp_66 = rob_bsy_6;
      5'b00111:
        casez_tmp_66 = rob_bsy_7;
      5'b01000:
        casez_tmp_66 = rob_bsy_8;
      5'b01001:
        casez_tmp_66 = rob_bsy_9;
      5'b01010:
        casez_tmp_66 = rob_bsy_10;
      5'b01011:
        casez_tmp_66 = rob_bsy_11;
      5'b01100:
        casez_tmp_66 = rob_bsy_12;
      5'b01101:
        casez_tmp_66 = rob_bsy_13;
      5'b01110:
        casez_tmp_66 = rob_bsy_14;
      5'b01111:
        casez_tmp_66 = rob_bsy_15;
      5'b10000:
        casez_tmp_66 = rob_bsy_16;
      5'b10001:
        casez_tmp_66 = rob_bsy_17;
      5'b10010:
        casez_tmp_66 = rob_bsy_18;
      5'b10011:
        casez_tmp_66 = rob_bsy_19;
      5'b10100:
        casez_tmp_66 = rob_bsy_20;
      5'b10101:
        casez_tmp_66 = rob_bsy_21;
      5'b10110:
        casez_tmp_66 = rob_bsy_22;
      5'b10111:
        casez_tmp_66 = rob_bsy_23;
      5'b11000:
        casez_tmp_66 = rob_bsy_24;
      5'b11001:
        casez_tmp_66 = rob_bsy_25;
      5'b11010:
        casez_tmp_66 = rob_bsy_26;
      5'b11011:
        casez_tmp_66 = rob_bsy_27;
      5'b11100:
        casez_tmp_66 = rob_bsy_28;
      5'b11101:
        casez_tmp_66 = rob_bsy_29;
      5'b11110:
        casez_tmp_66 = rob_bsy_30;
      default:
        casez_tmp_66 = rob_bsy_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_67;
  always @(*) begin
    casez (io_wb_resps_7_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_67 = rob_uop_0_pdst;
      5'b00001:
        casez_tmp_67 = rob_uop_1_pdst;
      5'b00010:
        casez_tmp_67 = rob_uop_2_pdst;
      5'b00011:
        casez_tmp_67 = rob_uop_3_pdst;
      5'b00100:
        casez_tmp_67 = rob_uop_4_pdst;
      5'b00101:
        casez_tmp_67 = rob_uop_5_pdst;
      5'b00110:
        casez_tmp_67 = rob_uop_6_pdst;
      5'b00111:
        casez_tmp_67 = rob_uop_7_pdst;
      5'b01000:
        casez_tmp_67 = rob_uop_8_pdst;
      5'b01001:
        casez_tmp_67 = rob_uop_9_pdst;
      5'b01010:
        casez_tmp_67 = rob_uop_10_pdst;
      5'b01011:
        casez_tmp_67 = rob_uop_11_pdst;
      5'b01100:
        casez_tmp_67 = rob_uop_12_pdst;
      5'b01101:
        casez_tmp_67 = rob_uop_13_pdst;
      5'b01110:
        casez_tmp_67 = rob_uop_14_pdst;
      5'b01111:
        casez_tmp_67 = rob_uop_15_pdst;
      5'b10000:
        casez_tmp_67 = rob_uop_16_pdst;
      5'b10001:
        casez_tmp_67 = rob_uop_17_pdst;
      5'b10010:
        casez_tmp_67 = rob_uop_18_pdst;
      5'b10011:
        casez_tmp_67 = rob_uop_19_pdst;
      5'b10100:
        casez_tmp_67 = rob_uop_20_pdst;
      5'b10101:
        casez_tmp_67 = rob_uop_21_pdst;
      5'b10110:
        casez_tmp_67 = rob_uop_22_pdst;
      5'b10111:
        casez_tmp_67 = rob_uop_23_pdst;
      5'b11000:
        casez_tmp_67 = rob_uop_24_pdst;
      5'b11001:
        casez_tmp_67 = rob_uop_25_pdst;
      5'b11010:
        casez_tmp_67 = rob_uop_26_pdst;
      5'b11011:
        casez_tmp_67 = rob_uop_27_pdst;
      5'b11100:
        casez_tmp_67 = rob_uop_28_pdst;
      5'b11101:
        casez_tmp_67 = rob_uop_29_pdst;
      5'b11110:
        casez_tmp_67 = rob_uop_30_pdst;
      default:
        casez_tmp_67 = rob_uop_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_68;
  always @(*) begin
    casez (io_wb_resps_7_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_68 = rob_uop_0_ldst_val;
      5'b00001:
        casez_tmp_68 = rob_uop_1_ldst_val;
      5'b00010:
        casez_tmp_68 = rob_uop_2_ldst_val;
      5'b00011:
        casez_tmp_68 = rob_uop_3_ldst_val;
      5'b00100:
        casez_tmp_68 = rob_uop_4_ldst_val;
      5'b00101:
        casez_tmp_68 = rob_uop_5_ldst_val;
      5'b00110:
        casez_tmp_68 = rob_uop_6_ldst_val;
      5'b00111:
        casez_tmp_68 = rob_uop_7_ldst_val;
      5'b01000:
        casez_tmp_68 = rob_uop_8_ldst_val;
      5'b01001:
        casez_tmp_68 = rob_uop_9_ldst_val;
      5'b01010:
        casez_tmp_68 = rob_uop_10_ldst_val;
      5'b01011:
        casez_tmp_68 = rob_uop_11_ldst_val;
      5'b01100:
        casez_tmp_68 = rob_uop_12_ldst_val;
      5'b01101:
        casez_tmp_68 = rob_uop_13_ldst_val;
      5'b01110:
        casez_tmp_68 = rob_uop_14_ldst_val;
      5'b01111:
        casez_tmp_68 = rob_uop_15_ldst_val;
      5'b10000:
        casez_tmp_68 = rob_uop_16_ldst_val;
      5'b10001:
        casez_tmp_68 = rob_uop_17_ldst_val;
      5'b10010:
        casez_tmp_68 = rob_uop_18_ldst_val;
      5'b10011:
        casez_tmp_68 = rob_uop_19_ldst_val;
      5'b10100:
        casez_tmp_68 = rob_uop_20_ldst_val;
      5'b10101:
        casez_tmp_68 = rob_uop_21_ldst_val;
      5'b10110:
        casez_tmp_68 = rob_uop_22_ldst_val;
      5'b10111:
        casez_tmp_68 = rob_uop_23_ldst_val;
      5'b11000:
        casez_tmp_68 = rob_uop_24_ldst_val;
      5'b11001:
        casez_tmp_68 = rob_uop_25_ldst_val;
      5'b11010:
        casez_tmp_68 = rob_uop_26_ldst_val;
      5'b11011:
        casez_tmp_68 = rob_uop_27_ldst_val;
      5'b11100:
        casez_tmp_68 = rob_uop_28_ldst_val;
      5'b11101:
        casez_tmp_68 = rob_uop_29_ldst_val;
      5'b11110:
        casez_tmp_68 = rob_uop_30_ldst_val;
      default:
        casez_tmp_68 = rob_uop_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_69;
  always @(*) begin
    casez (io_wb_resps_8_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_69 = rob_val_0;
      5'b00001:
        casez_tmp_69 = rob_val_1;
      5'b00010:
        casez_tmp_69 = rob_val_2;
      5'b00011:
        casez_tmp_69 = rob_val_3;
      5'b00100:
        casez_tmp_69 = rob_val_4;
      5'b00101:
        casez_tmp_69 = rob_val_5;
      5'b00110:
        casez_tmp_69 = rob_val_6;
      5'b00111:
        casez_tmp_69 = rob_val_7;
      5'b01000:
        casez_tmp_69 = rob_val_8;
      5'b01001:
        casez_tmp_69 = rob_val_9;
      5'b01010:
        casez_tmp_69 = rob_val_10;
      5'b01011:
        casez_tmp_69 = rob_val_11;
      5'b01100:
        casez_tmp_69 = rob_val_12;
      5'b01101:
        casez_tmp_69 = rob_val_13;
      5'b01110:
        casez_tmp_69 = rob_val_14;
      5'b01111:
        casez_tmp_69 = rob_val_15;
      5'b10000:
        casez_tmp_69 = rob_val_16;
      5'b10001:
        casez_tmp_69 = rob_val_17;
      5'b10010:
        casez_tmp_69 = rob_val_18;
      5'b10011:
        casez_tmp_69 = rob_val_19;
      5'b10100:
        casez_tmp_69 = rob_val_20;
      5'b10101:
        casez_tmp_69 = rob_val_21;
      5'b10110:
        casez_tmp_69 = rob_val_22;
      5'b10111:
        casez_tmp_69 = rob_val_23;
      5'b11000:
        casez_tmp_69 = rob_val_24;
      5'b11001:
        casez_tmp_69 = rob_val_25;
      5'b11010:
        casez_tmp_69 = rob_val_26;
      5'b11011:
        casez_tmp_69 = rob_val_27;
      5'b11100:
        casez_tmp_69 = rob_val_28;
      5'b11101:
        casez_tmp_69 = rob_val_29;
      5'b11110:
        casez_tmp_69 = rob_val_30;
      default:
        casez_tmp_69 = rob_val_31;
    endcase
  end // always @(*)
  reg         casez_tmp_70;
  always @(*) begin
    casez (io_wb_resps_8_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_70 = rob_bsy_0;
      5'b00001:
        casez_tmp_70 = rob_bsy_1;
      5'b00010:
        casez_tmp_70 = rob_bsy_2;
      5'b00011:
        casez_tmp_70 = rob_bsy_3;
      5'b00100:
        casez_tmp_70 = rob_bsy_4;
      5'b00101:
        casez_tmp_70 = rob_bsy_5;
      5'b00110:
        casez_tmp_70 = rob_bsy_6;
      5'b00111:
        casez_tmp_70 = rob_bsy_7;
      5'b01000:
        casez_tmp_70 = rob_bsy_8;
      5'b01001:
        casez_tmp_70 = rob_bsy_9;
      5'b01010:
        casez_tmp_70 = rob_bsy_10;
      5'b01011:
        casez_tmp_70 = rob_bsy_11;
      5'b01100:
        casez_tmp_70 = rob_bsy_12;
      5'b01101:
        casez_tmp_70 = rob_bsy_13;
      5'b01110:
        casez_tmp_70 = rob_bsy_14;
      5'b01111:
        casez_tmp_70 = rob_bsy_15;
      5'b10000:
        casez_tmp_70 = rob_bsy_16;
      5'b10001:
        casez_tmp_70 = rob_bsy_17;
      5'b10010:
        casez_tmp_70 = rob_bsy_18;
      5'b10011:
        casez_tmp_70 = rob_bsy_19;
      5'b10100:
        casez_tmp_70 = rob_bsy_20;
      5'b10101:
        casez_tmp_70 = rob_bsy_21;
      5'b10110:
        casez_tmp_70 = rob_bsy_22;
      5'b10111:
        casez_tmp_70 = rob_bsy_23;
      5'b11000:
        casez_tmp_70 = rob_bsy_24;
      5'b11001:
        casez_tmp_70 = rob_bsy_25;
      5'b11010:
        casez_tmp_70 = rob_bsy_26;
      5'b11011:
        casez_tmp_70 = rob_bsy_27;
      5'b11100:
        casez_tmp_70 = rob_bsy_28;
      5'b11101:
        casez_tmp_70 = rob_bsy_29;
      5'b11110:
        casez_tmp_70 = rob_bsy_30;
      default:
        casez_tmp_70 = rob_bsy_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_71;
  always @(*) begin
    casez (io_wb_resps_8_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_71 = rob_uop_0_pdst;
      5'b00001:
        casez_tmp_71 = rob_uop_1_pdst;
      5'b00010:
        casez_tmp_71 = rob_uop_2_pdst;
      5'b00011:
        casez_tmp_71 = rob_uop_3_pdst;
      5'b00100:
        casez_tmp_71 = rob_uop_4_pdst;
      5'b00101:
        casez_tmp_71 = rob_uop_5_pdst;
      5'b00110:
        casez_tmp_71 = rob_uop_6_pdst;
      5'b00111:
        casez_tmp_71 = rob_uop_7_pdst;
      5'b01000:
        casez_tmp_71 = rob_uop_8_pdst;
      5'b01001:
        casez_tmp_71 = rob_uop_9_pdst;
      5'b01010:
        casez_tmp_71 = rob_uop_10_pdst;
      5'b01011:
        casez_tmp_71 = rob_uop_11_pdst;
      5'b01100:
        casez_tmp_71 = rob_uop_12_pdst;
      5'b01101:
        casez_tmp_71 = rob_uop_13_pdst;
      5'b01110:
        casez_tmp_71 = rob_uop_14_pdst;
      5'b01111:
        casez_tmp_71 = rob_uop_15_pdst;
      5'b10000:
        casez_tmp_71 = rob_uop_16_pdst;
      5'b10001:
        casez_tmp_71 = rob_uop_17_pdst;
      5'b10010:
        casez_tmp_71 = rob_uop_18_pdst;
      5'b10011:
        casez_tmp_71 = rob_uop_19_pdst;
      5'b10100:
        casez_tmp_71 = rob_uop_20_pdst;
      5'b10101:
        casez_tmp_71 = rob_uop_21_pdst;
      5'b10110:
        casez_tmp_71 = rob_uop_22_pdst;
      5'b10111:
        casez_tmp_71 = rob_uop_23_pdst;
      5'b11000:
        casez_tmp_71 = rob_uop_24_pdst;
      5'b11001:
        casez_tmp_71 = rob_uop_25_pdst;
      5'b11010:
        casez_tmp_71 = rob_uop_26_pdst;
      5'b11011:
        casez_tmp_71 = rob_uop_27_pdst;
      5'b11100:
        casez_tmp_71 = rob_uop_28_pdst;
      5'b11101:
        casez_tmp_71 = rob_uop_29_pdst;
      5'b11110:
        casez_tmp_71 = rob_uop_30_pdst;
      default:
        casez_tmp_71 = rob_uop_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_72;
  always @(*) begin
    casez (io_wb_resps_8_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_72 = rob_uop_0_ldst_val;
      5'b00001:
        casez_tmp_72 = rob_uop_1_ldst_val;
      5'b00010:
        casez_tmp_72 = rob_uop_2_ldst_val;
      5'b00011:
        casez_tmp_72 = rob_uop_3_ldst_val;
      5'b00100:
        casez_tmp_72 = rob_uop_4_ldst_val;
      5'b00101:
        casez_tmp_72 = rob_uop_5_ldst_val;
      5'b00110:
        casez_tmp_72 = rob_uop_6_ldst_val;
      5'b00111:
        casez_tmp_72 = rob_uop_7_ldst_val;
      5'b01000:
        casez_tmp_72 = rob_uop_8_ldst_val;
      5'b01001:
        casez_tmp_72 = rob_uop_9_ldst_val;
      5'b01010:
        casez_tmp_72 = rob_uop_10_ldst_val;
      5'b01011:
        casez_tmp_72 = rob_uop_11_ldst_val;
      5'b01100:
        casez_tmp_72 = rob_uop_12_ldst_val;
      5'b01101:
        casez_tmp_72 = rob_uop_13_ldst_val;
      5'b01110:
        casez_tmp_72 = rob_uop_14_ldst_val;
      5'b01111:
        casez_tmp_72 = rob_uop_15_ldst_val;
      5'b10000:
        casez_tmp_72 = rob_uop_16_ldst_val;
      5'b10001:
        casez_tmp_72 = rob_uop_17_ldst_val;
      5'b10010:
        casez_tmp_72 = rob_uop_18_ldst_val;
      5'b10011:
        casez_tmp_72 = rob_uop_19_ldst_val;
      5'b10100:
        casez_tmp_72 = rob_uop_20_ldst_val;
      5'b10101:
        casez_tmp_72 = rob_uop_21_ldst_val;
      5'b10110:
        casez_tmp_72 = rob_uop_22_ldst_val;
      5'b10111:
        casez_tmp_72 = rob_uop_23_ldst_val;
      5'b11000:
        casez_tmp_72 = rob_uop_24_ldst_val;
      5'b11001:
        casez_tmp_72 = rob_uop_25_ldst_val;
      5'b11010:
        casez_tmp_72 = rob_uop_26_ldst_val;
      5'b11011:
        casez_tmp_72 = rob_uop_27_ldst_val;
      5'b11100:
        casez_tmp_72 = rob_uop_28_ldst_val;
      5'b11101:
        casez_tmp_72 = rob_uop_29_ldst_val;
      5'b11110:
        casez_tmp_72 = rob_uop_30_ldst_val;
      default:
        casez_tmp_72 = rob_uop_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_73;
  always @(*) begin
    casez (io_wb_resps_9_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_73 = rob_val_0;
      5'b00001:
        casez_tmp_73 = rob_val_1;
      5'b00010:
        casez_tmp_73 = rob_val_2;
      5'b00011:
        casez_tmp_73 = rob_val_3;
      5'b00100:
        casez_tmp_73 = rob_val_4;
      5'b00101:
        casez_tmp_73 = rob_val_5;
      5'b00110:
        casez_tmp_73 = rob_val_6;
      5'b00111:
        casez_tmp_73 = rob_val_7;
      5'b01000:
        casez_tmp_73 = rob_val_8;
      5'b01001:
        casez_tmp_73 = rob_val_9;
      5'b01010:
        casez_tmp_73 = rob_val_10;
      5'b01011:
        casez_tmp_73 = rob_val_11;
      5'b01100:
        casez_tmp_73 = rob_val_12;
      5'b01101:
        casez_tmp_73 = rob_val_13;
      5'b01110:
        casez_tmp_73 = rob_val_14;
      5'b01111:
        casez_tmp_73 = rob_val_15;
      5'b10000:
        casez_tmp_73 = rob_val_16;
      5'b10001:
        casez_tmp_73 = rob_val_17;
      5'b10010:
        casez_tmp_73 = rob_val_18;
      5'b10011:
        casez_tmp_73 = rob_val_19;
      5'b10100:
        casez_tmp_73 = rob_val_20;
      5'b10101:
        casez_tmp_73 = rob_val_21;
      5'b10110:
        casez_tmp_73 = rob_val_22;
      5'b10111:
        casez_tmp_73 = rob_val_23;
      5'b11000:
        casez_tmp_73 = rob_val_24;
      5'b11001:
        casez_tmp_73 = rob_val_25;
      5'b11010:
        casez_tmp_73 = rob_val_26;
      5'b11011:
        casez_tmp_73 = rob_val_27;
      5'b11100:
        casez_tmp_73 = rob_val_28;
      5'b11101:
        casez_tmp_73 = rob_val_29;
      5'b11110:
        casez_tmp_73 = rob_val_30;
      default:
        casez_tmp_73 = rob_val_31;
    endcase
  end // always @(*)
  reg         casez_tmp_74;
  always @(*) begin
    casez (io_wb_resps_9_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_74 = rob_bsy_0;
      5'b00001:
        casez_tmp_74 = rob_bsy_1;
      5'b00010:
        casez_tmp_74 = rob_bsy_2;
      5'b00011:
        casez_tmp_74 = rob_bsy_3;
      5'b00100:
        casez_tmp_74 = rob_bsy_4;
      5'b00101:
        casez_tmp_74 = rob_bsy_5;
      5'b00110:
        casez_tmp_74 = rob_bsy_6;
      5'b00111:
        casez_tmp_74 = rob_bsy_7;
      5'b01000:
        casez_tmp_74 = rob_bsy_8;
      5'b01001:
        casez_tmp_74 = rob_bsy_9;
      5'b01010:
        casez_tmp_74 = rob_bsy_10;
      5'b01011:
        casez_tmp_74 = rob_bsy_11;
      5'b01100:
        casez_tmp_74 = rob_bsy_12;
      5'b01101:
        casez_tmp_74 = rob_bsy_13;
      5'b01110:
        casez_tmp_74 = rob_bsy_14;
      5'b01111:
        casez_tmp_74 = rob_bsy_15;
      5'b10000:
        casez_tmp_74 = rob_bsy_16;
      5'b10001:
        casez_tmp_74 = rob_bsy_17;
      5'b10010:
        casez_tmp_74 = rob_bsy_18;
      5'b10011:
        casez_tmp_74 = rob_bsy_19;
      5'b10100:
        casez_tmp_74 = rob_bsy_20;
      5'b10101:
        casez_tmp_74 = rob_bsy_21;
      5'b10110:
        casez_tmp_74 = rob_bsy_22;
      5'b10111:
        casez_tmp_74 = rob_bsy_23;
      5'b11000:
        casez_tmp_74 = rob_bsy_24;
      5'b11001:
        casez_tmp_74 = rob_bsy_25;
      5'b11010:
        casez_tmp_74 = rob_bsy_26;
      5'b11011:
        casez_tmp_74 = rob_bsy_27;
      5'b11100:
        casez_tmp_74 = rob_bsy_28;
      5'b11101:
        casez_tmp_74 = rob_bsy_29;
      5'b11110:
        casez_tmp_74 = rob_bsy_30;
      default:
        casez_tmp_74 = rob_bsy_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_75;
  always @(*) begin
    casez (io_wb_resps_9_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_75 = rob_uop_0_pdst;
      5'b00001:
        casez_tmp_75 = rob_uop_1_pdst;
      5'b00010:
        casez_tmp_75 = rob_uop_2_pdst;
      5'b00011:
        casez_tmp_75 = rob_uop_3_pdst;
      5'b00100:
        casez_tmp_75 = rob_uop_4_pdst;
      5'b00101:
        casez_tmp_75 = rob_uop_5_pdst;
      5'b00110:
        casez_tmp_75 = rob_uop_6_pdst;
      5'b00111:
        casez_tmp_75 = rob_uop_7_pdst;
      5'b01000:
        casez_tmp_75 = rob_uop_8_pdst;
      5'b01001:
        casez_tmp_75 = rob_uop_9_pdst;
      5'b01010:
        casez_tmp_75 = rob_uop_10_pdst;
      5'b01011:
        casez_tmp_75 = rob_uop_11_pdst;
      5'b01100:
        casez_tmp_75 = rob_uop_12_pdst;
      5'b01101:
        casez_tmp_75 = rob_uop_13_pdst;
      5'b01110:
        casez_tmp_75 = rob_uop_14_pdst;
      5'b01111:
        casez_tmp_75 = rob_uop_15_pdst;
      5'b10000:
        casez_tmp_75 = rob_uop_16_pdst;
      5'b10001:
        casez_tmp_75 = rob_uop_17_pdst;
      5'b10010:
        casez_tmp_75 = rob_uop_18_pdst;
      5'b10011:
        casez_tmp_75 = rob_uop_19_pdst;
      5'b10100:
        casez_tmp_75 = rob_uop_20_pdst;
      5'b10101:
        casez_tmp_75 = rob_uop_21_pdst;
      5'b10110:
        casez_tmp_75 = rob_uop_22_pdst;
      5'b10111:
        casez_tmp_75 = rob_uop_23_pdst;
      5'b11000:
        casez_tmp_75 = rob_uop_24_pdst;
      5'b11001:
        casez_tmp_75 = rob_uop_25_pdst;
      5'b11010:
        casez_tmp_75 = rob_uop_26_pdst;
      5'b11011:
        casez_tmp_75 = rob_uop_27_pdst;
      5'b11100:
        casez_tmp_75 = rob_uop_28_pdst;
      5'b11101:
        casez_tmp_75 = rob_uop_29_pdst;
      5'b11110:
        casez_tmp_75 = rob_uop_30_pdst;
      default:
        casez_tmp_75 = rob_uop_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_76;
  always @(*) begin
    casez (io_wb_resps_9_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_76 = rob_uop_0_ldst_val;
      5'b00001:
        casez_tmp_76 = rob_uop_1_ldst_val;
      5'b00010:
        casez_tmp_76 = rob_uop_2_ldst_val;
      5'b00011:
        casez_tmp_76 = rob_uop_3_ldst_val;
      5'b00100:
        casez_tmp_76 = rob_uop_4_ldst_val;
      5'b00101:
        casez_tmp_76 = rob_uop_5_ldst_val;
      5'b00110:
        casez_tmp_76 = rob_uop_6_ldst_val;
      5'b00111:
        casez_tmp_76 = rob_uop_7_ldst_val;
      5'b01000:
        casez_tmp_76 = rob_uop_8_ldst_val;
      5'b01001:
        casez_tmp_76 = rob_uop_9_ldst_val;
      5'b01010:
        casez_tmp_76 = rob_uop_10_ldst_val;
      5'b01011:
        casez_tmp_76 = rob_uop_11_ldst_val;
      5'b01100:
        casez_tmp_76 = rob_uop_12_ldst_val;
      5'b01101:
        casez_tmp_76 = rob_uop_13_ldst_val;
      5'b01110:
        casez_tmp_76 = rob_uop_14_ldst_val;
      5'b01111:
        casez_tmp_76 = rob_uop_15_ldst_val;
      5'b10000:
        casez_tmp_76 = rob_uop_16_ldst_val;
      5'b10001:
        casez_tmp_76 = rob_uop_17_ldst_val;
      5'b10010:
        casez_tmp_76 = rob_uop_18_ldst_val;
      5'b10011:
        casez_tmp_76 = rob_uop_19_ldst_val;
      5'b10100:
        casez_tmp_76 = rob_uop_20_ldst_val;
      5'b10101:
        casez_tmp_76 = rob_uop_21_ldst_val;
      5'b10110:
        casez_tmp_76 = rob_uop_22_ldst_val;
      5'b10111:
        casez_tmp_76 = rob_uop_23_ldst_val;
      5'b11000:
        casez_tmp_76 = rob_uop_24_ldst_val;
      5'b11001:
        casez_tmp_76 = rob_uop_25_ldst_val;
      5'b11010:
        casez_tmp_76 = rob_uop_26_ldst_val;
      5'b11011:
        casez_tmp_76 = rob_uop_27_ldst_val;
      5'b11100:
        casez_tmp_76 = rob_uop_28_ldst_val;
      5'b11101:
        casez_tmp_76 = rob_uop_29_ldst_val;
      5'b11110:
        casez_tmp_76 = rob_uop_30_ldst_val;
      default:
        casez_tmp_76 = rob_uop_31_ldst_val;
    endcase
  end // always @(*)
  reg         rob_val_1_0;
  reg         rob_val_1_1;
  reg         rob_val_1_2;
  reg         rob_val_1_3;
  reg         rob_val_1_4;
  reg         rob_val_1_5;
  reg         rob_val_1_6;
  reg         rob_val_1_7;
  reg         rob_val_1_8;
  reg         rob_val_1_9;
  reg         rob_val_1_10;
  reg         rob_val_1_11;
  reg         rob_val_1_12;
  reg         rob_val_1_13;
  reg         rob_val_1_14;
  reg         rob_val_1_15;
  reg         rob_val_1_16;
  reg         rob_val_1_17;
  reg         rob_val_1_18;
  reg         rob_val_1_19;
  reg         rob_val_1_20;
  reg         rob_val_1_21;
  reg         rob_val_1_22;
  reg         rob_val_1_23;
  reg         rob_val_1_24;
  reg         rob_val_1_25;
  reg         rob_val_1_26;
  reg         rob_val_1_27;
  reg         rob_val_1_28;
  reg         rob_val_1_29;
  reg         rob_val_1_30;
  reg         rob_val_1_31;
  reg         rob_bsy_1_0;
  reg         rob_bsy_1_1;
  reg         rob_bsy_1_2;
  reg         rob_bsy_1_3;
  reg         rob_bsy_1_4;
  reg         rob_bsy_1_5;
  reg         rob_bsy_1_6;
  reg         rob_bsy_1_7;
  reg         rob_bsy_1_8;
  reg         rob_bsy_1_9;
  reg         rob_bsy_1_10;
  reg         rob_bsy_1_11;
  reg         rob_bsy_1_12;
  reg         rob_bsy_1_13;
  reg         rob_bsy_1_14;
  reg         rob_bsy_1_15;
  reg         rob_bsy_1_16;
  reg         rob_bsy_1_17;
  reg         rob_bsy_1_18;
  reg         rob_bsy_1_19;
  reg         rob_bsy_1_20;
  reg         rob_bsy_1_21;
  reg         rob_bsy_1_22;
  reg         rob_bsy_1_23;
  reg         rob_bsy_1_24;
  reg         rob_bsy_1_25;
  reg         rob_bsy_1_26;
  reg         rob_bsy_1_27;
  reg         rob_bsy_1_28;
  reg         rob_bsy_1_29;
  reg         rob_bsy_1_30;
  reg         rob_bsy_1_31;
  reg         rob_unsafe_1_0;
  reg         rob_unsafe_1_1;
  reg         rob_unsafe_1_2;
  reg         rob_unsafe_1_3;
  reg         rob_unsafe_1_4;
  reg         rob_unsafe_1_5;
  reg         rob_unsafe_1_6;
  reg         rob_unsafe_1_7;
  reg         rob_unsafe_1_8;
  reg         rob_unsafe_1_9;
  reg         rob_unsafe_1_10;
  reg         rob_unsafe_1_11;
  reg         rob_unsafe_1_12;
  reg         rob_unsafe_1_13;
  reg         rob_unsafe_1_14;
  reg         rob_unsafe_1_15;
  reg         rob_unsafe_1_16;
  reg         rob_unsafe_1_17;
  reg         rob_unsafe_1_18;
  reg         rob_unsafe_1_19;
  reg         rob_unsafe_1_20;
  reg         rob_unsafe_1_21;
  reg         rob_unsafe_1_22;
  reg         rob_unsafe_1_23;
  reg         rob_unsafe_1_24;
  reg         rob_unsafe_1_25;
  reg         rob_unsafe_1_26;
  reg         rob_unsafe_1_27;
  reg         rob_unsafe_1_28;
  reg         rob_unsafe_1_29;
  reg         rob_unsafe_1_30;
  reg         rob_unsafe_1_31;
  reg  [6:0]  rob_uop_1_0_uopc;
  reg         rob_uop_1_0_is_rvc;
  reg         rob_uop_1_0_is_br;
  reg         rob_uop_1_0_is_jalr;
  reg         rob_uop_1_0_is_jal;
  reg  [19:0] rob_uop_1_0_br_mask;
  reg  [5:0]  rob_uop_1_0_ftq_idx;
  reg         rob_uop_1_0_edge_inst;
  reg  [5:0]  rob_uop_1_0_pc_lob;
  reg  [6:0]  rob_uop_1_0_pdst;
  reg  [6:0]  rob_uop_1_0_stale_pdst;
  reg         rob_uop_1_0_is_fencei;
  reg         rob_uop_1_0_uses_ldq;
  reg         rob_uop_1_0_uses_stq;
  reg         rob_uop_1_0_is_sys_pc2epc;
  reg         rob_uop_1_0_flush_on_commit;
  reg  [5:0]  rob_uop_1_0_ldst;
  reg         rob_uop_1_0_ldst_val;
  reg  [1:0]  rob_uop_1_0_dst_rtype;
  reg         rob_uop_1_0_fp_val;
  reg  [1:0]  rob_uop_1_0_debug_fsrc;
  reg  [6:0]  rob_uop_1_1_uopc;
  reg         rob_uop_1_1_is_rvc;
  reg         rob_uop_1_1_is_br;
  reg         rob_uop_1_1_is_jalr;
  reg         rob_uop_1_1_is_jal;
  reg  [19:0] rob_uop_1_1_br_mask;
  reg  [5:0]  rob_uop_1_1_ftq_idx;
  reg         rob_uop_1_1_edge_inst;
  reg  [5:0]  rob_uop_1_1_pc_lob;
  reg  [6:0]  rob_uop_1_1_pdst;
  reg  [6:0]  rob_uop_1_1_stale_pdst;
  reg         rob_uop_1_1_is_fencei;
  reg         rob_uop_1_1_uses_ldq;
  reg         rob_uop_1_1_uses_stq;
  reg         rob_uop_1_1_is_sys_pc2epc;
  reg         rob_uop_1_1_flush_on_commit;
  reg  [5:0]  rob_uop_1_1_ldst;
  reg         rob_uop_1_1_ldst_val;
  reg  [1:0]  rob_uop_1_1_dst_rtype;
  reg         rob_uop_1_1_fp_val;
  reg  [1:0]  rob_uop_1_1_debug_fsrc;
  reg  [6:0]  rob_uop_1_2_uopc;
  reg         rob_uop_1_2_is_rvc;
  reg         rob_uop_1_2_is_br;
  reg         rob_uop_1_2_is_jalr;
  reg         rob_uop_1_2_is_jal;
  reg  [19:0] rob_uop_1_2_br_mask;
  reg  [5:0]  rob_uop_1_2_ftq_idx;
  reg         rob_uop_1_2_edge_inst;
  reg  [5:0]  rob_uop_1_2_pc_lob;
  reg  [6:0]  rob_uop_1_2_pdst;
  reg  [6:0]  rob_uop_1_2_stale_pdst;
  reg         rob_uop_1_2_is_fencei;
  reg         rob_uop_1_2_uses_ldq;
  reg         rob_uop_1_2_uses_stq;
  reg         rob_uop_1_2_is_sys_pc2epc;
  reg         rob_uop_1_2_flush_on_commit;
  reg  [5:0]  rob_uop_1_2_ldst;
  reg         rob_uop_1_2_ldst_val;
  reg  [1:0]  rob_uop_1_2_dst_rtype;
  reg         rob_uop_1_2_fp_val;
  reg  [1:0]  rob_uop_1_2_debug_fsrc;
  reg  [6:0]  rob_uop_1_3_uopc;
  reg         rob_uop_1_3_is_rvc;
  reg         rob_uop_1_3_is_br;
  reg         rob_uop_1_3_is_jalr;
  reg         rob_uop_1_3_is_jal;
  reg  [19:0] rob_uop_1_3_br_mask;
  reg  [5:0]  rob_uop_1_3_ftq_idx;
  reg         rob_uop_1_3_edge_inst;
  reg  [5:0]  rob_uop_1_3_pc_lob;
  reg  [6:0]  rob_uop_1_3_pdst;
  reg  [6:0]  rob_uop_1_3_stale_pdst;
  reg         rob_uop_1_3_is_fencei;
  reg         rob_uop_1_3_uses_ldq;
  reg         rob_uop_1_3_uses_stq;
  reg         rob_uop_1_3_is_sys_pc2epc;
  reg         rob_uop_1_3_flush_on_commit;
  reg  [5:0]  rob_uop_1_3_ldst;
  reg         rob_uop_1_3_ldst_val;
  reg  [1:0]  rob_uop_1_3_dst_rtype;
  reg         rob_uop_1_3_fp_val;
  reg  [1:0]  rob_uop_1_3_debug_fsrc;
  reg  [6:0]  rob_uop_1_4_uopc;
  reg         rob_uop_1_4_is_rvc;
  reg         rob_uop_1_4_is_br;
  reg         rob_uop_1_4_is_jalr;
  reg         rob_uop_1_4_is_jal;
  reg  [19:0] rob_uop_1_4_br_mask;
  reg  [5:0]  rob_uop_1_4_ftq_idx;
  reg         rob_uop_1_4_edge_inst;
  reg  [5:0]  rob_uop_1_4_pc_lob;
  reg  [6:0]  rob_uop_1_4_pdst;
  reg  [6:0]  rob_uop_1_4_stale_pdst;
  reg         rob_uop_1_4_is_fencei;
  reg         rob_uop_1_4_uses_ldq;
  reg         rob_uop_1_4_uses_stq;
  reg         rob_uop_1_4_is_sys_pc2epc;
  reg         rob_uop_1_4_flush_on_commit;
  reg  [5:0]  rob_uop_1_4_ldst;
  reg         rob_uop_1_4_ldst_val;
  reg  [1:0]  rob_uop_1_4_dst_rtype;
  reg         rob_uop_1_4_fp_val;
  reg  [1:0]  rob_uop_1_4_debug_fsrc;
  reg  [6:0]  rob_uop_1_5_uopc;
  reg         rob_uop_1_5_is_rvc;
  reg         rob_uop_1_5_is_br;
  reg         rob_uop_1_5_is_jalr;
  reg         rob_uop_1_5_is_jal;
  reg  [19:0] rob_uop_1_5_br_mask;
  reg  [5:0]  rob_uop_1_5_ftq_idx;
  reg         rob_uop_1_5_edge_inst;
  reg  [5:0]  rob_uop_1_5_pc_lob;
  reg  [6:0]  rob_uop_1_5_pdst;
  reg  [6:0]  rob_uop_1_5_stale_pdst;
  reg         rob_uop_1_5_is_fencei;
  reg         rob_uop_1_5_uses_ldq;
  reg         rob_uop_1_5_uses_stq;
  reg         rob_uop_1_5_is_sys_pc2epc;
  reg         rob_uop_1_5_flush_on_commit;
  reg  [5:0]  rob_uop_1_5_ldst;
  reg         rob_uop_1_5_ldst_val;
  reg  [1:0]  rob_uop_1_5_dst_rtype;
  reg         rob_uop_1_5_fp_val;
  reg  [1:0]  rob_uop_1_5_debug_fsrc;
  reg  [6:0]  rob_uop_1_6_uopc;
  reg         rob_uop_1_6_is_rvc;
  reg         rob_uop_1_6_is_br;
  reg         rob_uop_1_6_is_jalr;
  reg         rob_uop_1_6_is_jal;
  reg  [19:0] rob_uop_1_6_br_mask;
  reg  [5:0]  rob_uop_1_6_ftq_idx;
  reg         rob_uop_1_6_edge_inst;
  reg  [5:0]  rob_uop_1_6_pc_lob;
  reg  [6:0]  rob_uop_1_6_pdst;
  reg  [6:0]  rob_uop_1_6_stale_pdst;
  reg         rob_uop_1_6_is_fencei;
  reg         rob_uop_1_6_uses_ldq;
  reg         rob_uop_1_6_uses_stq;
  reg         rob_uop_1_6_is_sys_pc2epc;
  reg         rob_uop_1_6_flush_on_commit;
  reg  [5:0]  rob_uop_1_6_ldst;
  reg         rob_uop_1_6_ldst_val;
  reg  [1:0]  rob_uop_1_6_dst_rtype;
  reg         rob_uop_1_6_fp_val;
  reg  [1:0]  rob_uop_1_6_debug_fsrc;
  reg  [6:0]  rob_uop_1_7_uopc;
  reg         rob_uop_1_7_is_rvc;
  reg         rob_uop_1_7_is_br;
  reg         rob_uop_1_7_is_jalr;
  reg         rob_uop_1_7_is_jal;
  reg  [19:0] rob_uop_1_7_br_mask;
  reg  [5:0]  rob_uop_1_7_ftq_idx;
  reg         rob_uop_1_7_edge_inst;
  reg  [5:0]  rob_uop_1_7_pc_lob;
  reg  [6:0]  rob_uop_1_7_pdst;
  reg  [6:0]  rob_uop_1_7_stale_pdst;
  reg         rob_uop_1_7_is_fencei;
  reg         rob_uop_1_7_uses_ldq;
  reg         rob_uop_1_7_uses_stq;
  reg         rob_uop_1_7_is_sys_pc2epc;
  reg         rob_uop_1_7_flush_on_commit;
  reg  [5:0]  rob_uop_1_7_ldst;
  reg         rob_uop_1_7_ldst_val;
  reg  [1:0]  rob_uop_1_7_dst_rtype;
  reg         rob_uop_1_7_fp_val;
  reg  [1:0]  rob_uop_1_7_debug_fsrc;
  reg  [6:0]  rob_uop_1_8_uopc;
  reg         rob_uop_1_8_is_rvc;
  reg         rob_uop_1_8_is_br;
  reg         rob_uop_1_8_is_jalr;
  reg         rob_uop_1_8_is_jal;
  reg  [19:0] rob_uop_1_8_br_mask;
  reg  [5:0]  rob_uop_1_8_ftq_idx;
  reg         rob_uop_1_8_edge_inst;
  reg  [5:0]  rob_uop_1_8_pc_lob;
  reg  [6:0]  rob_uop_1_8_pdst;
  reg  [6:0]  rob_uop_1_8_stale_pdst;
  reg         rob_uop_1_8_is_fencei;
  reg         rob_uop_1_8_uses_ldq;
  reg         rob_uop_1_8_uses_stq;
  reg         rob_uop_1_8_is_sys_pc2epc;
  reg         rob_uop_1_8_flush_on_commit;
  reg  [5:0]  rob_uop_1_8_ldst;
  reg         rob_uop_1_8_ldst_val;
  reg  [1:0]  rob_uop_1_8_dst_rtype;
  reg         rob_uop_1_8_fp_val;
  reg  [1:0]  rob_uop_1_8_debug_fsrc;
  reg  [6:0]  rob_uop_1_9_uopc;
  reg         rob_uop_1_9_is_rvc;
  reg         rob_uop_1_9_is_br;
  reg         rob_uop_1_9_is_jalr;
  reg         rob_uop_1_9_is_jal;
  reg  [19:0] rob_uop_1_9_br_mask;
  reg  [5:0]  rob_uop_1_9_ftq_idx;
  reg         rob_uop_1_9_edge_inst;
  reg  [5:0]  rob_uop_1_9_pc_lob;
  reg  [6:0]  rob_uop_1_9_pdst;
  reg  [6:0]  rob_uop_1_9_stale_pdst;
  reg         rob_uop_1_9_is_fencei;
  reg         rob_uop_1_9_uses_ldq;
  reg         rob_uop_1_9_uses_stq;
  reg         rob_uop_1_9_is_sys_pc2epc;
  reg         rob_uop_1_9_flush_on_commit;
  reg  [5:0]  rob_uop_1_9_ldst;
  reg         rob_uop_1_9_ldst_val;
  reg  [1:0]  rob_uop_1_9_dst_rtype;
  reg         rob_uop_1_9_fp_val;
  reg  [1:0]  rob_uop_1_9_debug_fsrc;
  reg  [6:0]  rob_uop_1_10_uopc;
  reg         rob_uop_1_10_is_rvc;
  reg         rob_uop_1_10_is_br;
  reg         rob_uop_1_10_is_jalr;
  reg         rob_uop_1_10_is_jal;
  reg  [19:0] rob_uop_1_10_br_mask;
  reg  [5:0]  rob_uop_1_10_ftq_idx;
  reg         rob_uop_1_10_edge_inst;
  reg  [5:0]  rob_uop_1_10_pc_lob;
  reg  [6:0]  rob_uop_1_10_pdst;
  reg  [6:0]  rob_uop_1_10_stale_pdst;
  reg         rob_uop_1_10_is_fencei;
  reg         rob_uop_1_10_uses_ldq;
  reg         rob_uop_1_10_uses_stq;
  reg         rob_uop_1_10_is_sys_pc2epc;
  reg         rob_uop_1_10_flush_on_commit;
  reg  [5:0]  rob_uop_1_10_ldst;
  reg         rob_uop_1_10_ldst_val;
  reg  [1:0]  rob_uop_1_10_dst_rtype;
  reg         rob_uop_1_10_fp_val;
  reg  [1:0]  rob_uop_1_10_debug_fsrc;
  reg  [6:0]  rob_uop_1_11_uopc;
  reg         rob_uop_1_11_is_rvc;
  reg         rob_uop_1_11_is_br;
  reg         rob_uop_1_11_is_jalr;
  reg         rob_uop_1_11_is_jal;
  reg  [19:0] rob_uop_1_11_br_mask;
  reg  [5:0]  rob_uop_1_11_ftq_idx;
  reg         rob_uop_1_11_edge_inst;
  reg  [5:0]  rob_uop_1_11_pc_lob;
  reg  [6:0]  rob_uop_1_11_pdst;
  reg  [6:0]  rob_uop_1_11_stale_pdst;
  reg         rob_uop_1_11_is_fencei;
  reg         rob_uop_1_11_uses_ldq;
  reg         rob_uop_1_11_uses_stq;
  reg         rob_uop_1_11_is_sys_pc2epc;
  reg         rob_uop_1_11_flush_on_commit;
  reg  [5:0]  rob_uop_1_11_ldst;
  reg         rob_uop_1_11_ldst_val;
  reg  [1:0]  rob_uop_1_11_dst_rtype;
  reg         rob_uop_1_11_fp_val;
  reg  [1:0]  rob_uop_1_11_debug_fsrc;
  reg  [6:0]  rob_uop_1_12_uopc;
  reg         rob_uop_1_12_is_rvc;
  reg         rob_uop_1_12_is_br;
  reg         rob_uop_1_12_is_jalr;
  reg         rob_uop_1_12_is_jal;
  reg  [19:0] rob_uop_1_12_br_mask;
  reg  [5:0]  rob_uop_1_12_ftq_idx;
  reg         rob_uop_1_12_edge_inst;
  reg  [5:0]  rob_uop_1_12_pc_lob;
  reg  [6:0]  rob_uop_1_12_pdst;
  reg  [6:0]  rob_uop_1_12_stale_pdst;
  reg         rob_uop_1_12_is_fencei;
  reg         rob_uop_1_12_uses_ldq;
  reg         rob_uop_1_12_uses_stq;
  reg         rob_uop_1_12_is_sys_pc2epc;
  reg         rob_uop_1_12_flush_on_commit;
  reg  [5:0]  rob_uop_1_12_ldst;
  reg         rob_uop_1_12_ldst_val;
  reg  [1:0]  rob_uop_1_12_dst_rtype;
  reg         rob_uop_1_12_fp_val;
  reg  [1:0]  rob_uop_1_12_debug_fsrc;
  reg  [6:0]  rob_uop_1_13_uopc;
  reg         rob_uop_1_13_is_rvc;
  reg         rob_uop_1_13_is_br;
  reg         rob_uop_1_13_is_jalr;
  reg         rob_uop_1_13_is_jal;
  reg  [19:0] rob_uop_1_13_br_mask;
  reg  [5:0]  rob_uop_1_13_ftq_idx;
  reg         rob_uop_1_13_edge_inst;
  reg  [5:0]  rob_uop_1_13_pc_lob;
  reg  [6:0]  rob_uop_1_13_pdst;
  reg  [6:0]  rob_uop_1_13_stale_pdst;
  reg         rob_uop_1_13_is_fencei;
  reg         rob_uop_1_13_uses_ldq;
  reg         rob_uop_1_13_uses_stq;
  reg         rob_uop_1_13_is_sys_pc2epc;
  reg         rob_uop_1_13_flush_on_commit;
  reg  [5:0]  rob_uop_1_13_ldst;
  reg         rob_uop_1_13_ldst_val;
  reg  [1:0]  rob_uop_1_13_dst_rtype;
  reg         rob_uop_1_13_fp_val;
  reg  [1:0]  rob_uop_1_13_debug_fsrc;
  reg  [6:0]  rob_uop_1_14_uopc;
  reg         rob_uop_1_14_is_rvc;
  reg         rob_uop_1_14_is_br;
  reg         rob_uop_1_14_is_jalr;
  reg         rob_uop_1_14_is_jal;
  reg  [19:0] rob_uop_1_14_br_mask;
  reg  [5:0]  rob_uop_1_14_ftq_idx;
  reg         rob_uop_1_14_edge_inst;
  reg  [5:0]  rob_uop_1_14_pc_lob;
  reg  [6:0]  rob_uop_1_14_pdst;
  reg  [6:0]  rob_uop_1_14_stale_pdst;
  reg         rob_uop_1_14_is_fencei;
  reg         rob_uop_1_14_uses_ldq;
  reg         rob_uop_1_14_uses_stq;
  reg         rob_uop_1_14_is_sys_pc2epc;
  reg         rob_uop_1_14_flush_on_commit;
  reg  [5:0]  rob_uop_1_14_ldst;
  reg         rob_uop_1_14_ldst_val;
  reg  [1:0]  rob_uop_1_14_dst_rtype;
  reg         rob_uop_1_14_fp_val;
  reg  [1:0]  rob_uop_1_14_debug_fsrc;
  reg  [6:0]  rob_uop_1_15_uopc;
  reg         rob_uop_1_15_is_rvc;
  reg         rob_uop_1_15_is_br;
  reg         rob_uop_1_15_is_jalr;
  reg         rob_uop_1_15_is_jal;
  reg  [19:0] rob_uop_1_15_br_mask;
  reg  [5:0]  rob_uop_1_15_ftq_idx;
  reg         rob_uop_1_15_edge_inst;
  reg  [5:0]  rob_uop_1_15_pc_lob;
  reg  [6:0]  rob_uop_1_15_pdst;
  reg  [6:0]  rob_uop_1_15_stale_pdst;
  reg         rob_uop_1_15_is_fencei;
  reg         rob_uop_1_15_uses_ldq;
  reg         rob_uop_1_15_uses_stq;
  reg         rob_uop_1_15_is_sys_pc2epc;
  reg         rob_uop_1_15_flush_on_commit;
  reg  [5:0]  rob_uop_1_15_ldst;
  reg         rob_uop_1_15_ldst_val;
  reg  [1:0]  rob_uop_1_15_dst_rtype;
  reg         rob_uop_1_15_fp_val;
  reg  [1:0]  rob_uop_1_15_debug_fsrc;
  reg  [6:0]  rob_uop_1_16_uopc;
  reg         rob_uop_1_16_is_rvc;
  reg         rob_uop_1_16_is_br;
  reg         rob_uop_1_16_is_jalr;
  reg         rob_uop_1_16_is_jal;
  reg  [19:0] rob_uop_1_16_br_mask;
  reg  [5:0]  rob_uop_1_16_ftq_idx;
  reg         rob_uop_1_16_edge_inst;
  reg  [5:0]  rob_uop_1_16_pc_lob;
  reg  [6:0]  rob_uop_1_16_pdst;
  reg  [6:0]  rob_uop_1_16_stale_pdst;
  reg         rob_uop_1_16_is_fencei;
  reg         rob_uop_1_16_uses_ldq;
  reg         rob_uop_1_16_uses_stq;
  reg         rob_uop_1_16_is_sys_pc2epc;
  reg         rob_uop_1_16_flush_on_commit;
  reg  [5:0]  rob_uop_1_16_ldst;
  reg         rob_uop_1_16_ldst_val;
  reg  [1:0]  rob_uop_1_16_dst_rtype;
  reg         rob_uop_1_16_fp_val;
  reg  [1:0]  rob_uop_1_16_debug_fsrc;
  reg  [6:0]  rob_uop_1_17_uopc;
  reg         rob_uop_1_17_is_rvc;
  reg         rob_uop_1_17_is_br;
  reg         rob_uop_1_17_is_jalr;
  reg         rob_uop_1_17_is_jal;
  reg  [19:0] rob_uop_1_17_br_mask;
  reg  [5:0]  rob_uop_1_17_ftq_idx;
  reg         rob_uop_1_17_edge_inst;
  reg  [5:0]  rob_uop_1_17_pc_lob;
  reg  [6:0]  rob_uop_1_17_pdst;
  reg  [6:0]  rob_uop_1_17_stale_pdst;
  reg         rob_uop_1_17_is_fencei;
  reg         rob_uop_1_17_uses_ldq;
  reg         rob_uop_1_17_uses_stq;
  reg         rob_uop_1_17_is_sys_pc2epc;
  reg         rob_uop_1_17_flush_on_commit;
  reg  [5:0]  rob_uop_1_17_ldst;
  reg         rob_uop_1_17_ldst_val;
  reg  [1:0]  rob_uop_1_17_dst_rtype;
  reg         rob_uop_1_17_fp_val;
  reg  [1:0]  rob_uop_1_17_debug_fsrc;
  reg  [6:0]  rob_uop_1_18_uopc;
  reg         rob_uop_1_18_is_rvc;
  reg         rob_uop_1_18_is_br;
  reg         rob_uop_1_18_is_jalr;
  reg         rob_uop_1_18_is_jal;
  reg  [19:0] rob_uop_1_18_br_mask;
  reg  [5:0]  rob_uop_1_18_ftq_idx;
  reg         rob_uop_1_18_edge_inst;
  reg  [5:0]  rob_uop_1_18_pc_lob;
  reg  [6:0]  rob_uop_1_18_pdst;
  reg  [6:0]  rob_uop_1_18_stale_pdst;
  reg         rob_uop_1_18_is_fencei;
  reg         rob_uop_1_18_uses_ldq;
  reg         rob_uop_1_18_uses_stq;
  reg         rob_uop_1_18_is_sys_pc2epc;
  reg         rob_uop_1_18_flush_on_commit;
  reg  [5:0]  rob_uop_1_18_ldst;
  reg         rob_uop_1_18_ldst_val;
  reg  [1:0]  rob_uop_1_18_dst_rtype;
  reg         rob_uop_1_18_fp_val;
  reg  [1:0]  rob_uop_1_18_debug_fsrc;
  reg  [6:0]  rob_uop_1_19_uopc;
  reg         rob_uop_1_19_is_rvc;
  reg         rob_uop_1_19_is_br;
  reg         rob_uop_1_19_is_jalr;
  reg         rob_uop_1_19_is_jal;
  reg  [19:0] rob_uop_1_19_br_mask;
  reg  [5:0]  rob_uop_1_19_ftq_idx;
  reg         rob_uop_1_19_edge_inst;
  reg  [5:0]  rob_uop_1_19_pc_lob;
  reg  [6:0]  rob_uop_1_19_pdst;
  reg  [6:0]  rob_uop_1_19_stale_pdst;
  reg         rob_uop_1_19_is_fencei;
  reg         rob_uop_1_19_uses_ldq;
  reg         rob_uop_1_19_uses_stq;
  reg         rob_uop_1_19_is_sys_pc2epc;
  reg         rob_uop_1_19_flush_on_commit;
  reg  [5:0]  rob_uop_1_19_ldst;
  reg         rob_uop_1_19_ldst_val;
  reg  [1:0]  rob_uop_1_19_dst_rtype;
  reg         rob_uop_1_19_fp_val;
  reg  [1:0]  rob_uop_1_19_debug_fsrc;
  reg  [6:0]  rob_uop_1_20_uopc;
  reg         rob_uop_1_20_is_rvc;
  reg         rob_uop_1_20_is_br;
  reg         rob_uop_1_20_is_jalr;
  reg         rob_uop_1_20_is_jal;
  reg  [19:0] rob_uop_1_20_br_mask;
  reg  [5:0]  rob_uop_1_20_ftq_idx;
  reg         rob_uop_1_20_edge_inst;
  reg  [5:0]  rob_uop_1_20_pc_lob;
  reg  [6:0]  rob_uop_1_20_pdst;
  reg  [6:0]  rob_uop_1_20_stale_pdst;
  reg         rob_uop_1_20_is_fencei;
  reg         rob_uop_1_20_uses_ldq;
  reg         rob_uop_1_20_uses_stq;
  reg         rob_uop_1_20_is_sys_pc2epc;
  reg         rob_uop_1_20_flush_on_commit;
  reg  [5:0]  rob_uop_1_20_ldst;
  reg         rob_uop_1_20_ldst_val;
  reg  [1:0]  rob_uop_1_20_dst_rtype;
  reg         rob_uop_1_20_fp_val;
  reg  [1:0]  rob_uop_1_20_debug_fsrc;
  reg  [6:0]  rob_uop_1_21_uopc;
  reg         rob_uop_1_21_is_rvc;
  reg         rob_uop_1_21_is_br;
  reg         rob_uop_1_21_is_jalr;
  reg         rob_uop_1_21_is_jal;
  reg  [19:0] rob_uop_1_21_br_mask;
  reg  [5:0]  rob_uop_1_21_ftq_idx;
  reg         rob_uop_1_21_edge_inst;
  reg  [5:0]  rob_uop_1_21_pc_lob;
  reg  [6:0]  rob_uop_1_21_pdst;
  reg  [6:0]  rob_uop_1_21_stale_pdst;
  reg         rob_uop_1_21_is_fencei;
  reg         rob_uop_1_21_uses_ldq;
  reg         rob_uop_1_21_uses_stq;
  reg         rob_uop_1_21_is_sys_pc2epc;
  reg         rob_uop_1_21_flush_on_commit;
  reg  [5:0]  rob_uop_1_21_ldst;
  reg         rob_uop_1_21_ldst_val;
  reg  [1:0]  rob_uop_1_21_dst_rtype;
  reg         rob_uop_1_21_fp_val;
  reg  [1:0]  rob_uop_1_21_debug_fsrc;
  reg  [6:0]  rob_uop_1_22_uopc;
  reg         rob_uop_1_22_is_rvc;
  reg         rob_uop_1_22_is_br;
  reg         rob_uop_1_22_is_jalr;
  reg         rob_uop_1_22_is_jal;
  reg  [19:0] rob_uop_1_22_br_mask;
  reg  [5:0]  rob_uop_1_22_ftq_idx;
  reg         rob_uop_1_22_edge_inst;
  reg  [5:0]  rob_uop_1_22_pc_lob;
  reg  [6:0]  rob_uop_1_22_pdst;
  reg  [6:0]  rob_uop_1_22_stale_pdst;
  reg         rob_uop_1_22_is_fencei;
  reg         rob_uop_1_22_uses_ldq;
  reg         rob_uop_1_22_uses_stq;
  reg         rob_uop_1_22_is_sys_pc2epc;
  reg         rob_uop_1_22_flush_on_commit;
  reg  [5:0]  rob_uop_1_22_ldst;
  reg         rob_uop_1_22_ldst_val;
  reg  [1:0]  rob_uop_1_22_dst_rtype;
  reg         rob_uop_1_22_fp_val;
  reg  [1:0]  rob_uop_1_22_debug_fsrc;
  reg  [6:0]  rob_uop_1_23_uopc;
  reg         rob_uop_1_23_is_rvc;
  reg         rob_uop_1_23_is_br;
  reg         rob_uop_1_23_is_jalr;
  reg         rob_uop_1_23_is_jal;
  reg  [19:0] rob_uop_1_23_br_mask;
  reg  [5:0]  rob_uop_1_23_ftq_idx;
  reg         rob_uop_1_23_edge_inst;
  reg  [5:0]  rob_uop_1_23_pc_lob;
  reg  [6:0]  rob_uop_1_23_pdst;
  reg  [6:0]  rob_uop_1_23_stale_pdst;
  reg         rob_uop_1_23_is_fencei;
  reg         rob_uop_1_23_uses_ldq;
  reg         rob_uop_1_23_uses_stq;
  reg         rob_uop_1_23_is_sys_pc2epc;
  reg         rob_uop_1_23_flush_on_commit;
  reg  [5:0]  rob_uop_1_23_ldst;
  reg         rob_uop_1_23_ldst_val;
  reg  [1:0]  rob_uop_1_23_dst_rtype;
  reg         rob_uop_1_23_fp_val;
  reg  [1:0]  rob_uop_1_23_debug_fsrc;
  reg  [6:0]  rob_uop_1_24_uopc;
  reg         rob_uop_1_24_is_rvc;
  reg         rob_uop_1_24_is_br;
  reg         rob_uop_1_24_is_jalr;
  reg         rob_uop_1_24_is_jal;
  reg  [19:0] rob_uop_1_24_br_mask;
  reg  [5:0]  rob_uop_1_24_ftq_idx;
  reg         rob_uop_1_24_edge_inst;
  reg  [5:0]  rob_uop_1_24_pc_lob;
  reg  [6:0]  rob_uop_1_24_pdst;
  reg  [6:0]  rob_uop_1_24_stale_pdst;
  reg         rob_uop_1_24_is_fencei;
  reg         rob_uop_1_24_uses_ldq;
  reg         rob_uop_1_24_uses_stq;
  reg         rob_uop_1_24_is_sys_pc2epc;
  reg         rob_uop_1_24_flush_on_commit;
  reg  [5:0]  rob_uop_1_24_ldst;
  reg         rob_uop_1_24_ldst_val;
  reg  [1:0]  rob_uop_1_24_dst_rtype;
  reg         rob_uop_1_24_fp_val;
  reg  [1:0]  rob_uop_1_24_debug_fsrc;
  reg  [6:0]  rob_uop_1_25_uopc;
  reg         rob_uop_1_25_is_rvc;
  reg         rob_uop_1_25_is_br;
  reg         rob_uop_1_25_is_jalr;
  reg         rob_uop_1_25_is_jal;
  reg  [19:0] rob_uop_1_25_br_mask;
  reg  [5:0]  rob_uop_1_25_ftq_idx;
  reg         rob_uop_1_25_edge_inst;
  reg  [5:0]  rob_uop_1_25_pc_lob;
  reg  [6:0]  rob_uop_1_25_pdst;
  reg  [6:0]  rob_uop_1_25_stale_pdst;
  reg         rob_uop_1_25_is_fencei;
  reg         rob_uop_1_25_uses_ldq;
  reg         rob_uop_1_25_uses_stq;
  reg         rob_uop_1_25_is_sys_pc2epc;
  reg         rob_uop_1_25_flush_on_commit;
  reg  [5:0]  rob_uop_1_25_ldst;
  reg         rob_uop_1_25_ldst_val;
  reg  [1:0]  rob_uop_1_25_dst_rtype;
  reg         rob_uop_1_25_fp_val;
  reg  [1:0]  rob_uop_1_25_debug_fsrc;
  reg  [6:0]  rob_uop_1_26_uopc;
  reg         rob_uop_1_26_is_rvc;
  reg         rob_uop_1_26_is_br;
  reg         rob_uop_1_26_is_jalr;
  reg         rob_uop_1_26_is_jal;
  reg  [19:0] rob_uop_1_26_br_mask;
  reg  [5:0]  rob_uop_1_26_ftq_idx;
  reg         rob_uop_1_26_edge_inst;
  reg  [5:0]  rob_uop_1_26_pc_lob;
  reg  [6:0]  rob_uop_1_26_pdst;
  reg  [6:0]  rob_uop_1_26_stale_pdst;
  reg         rob_uop_1_26_is_fencei;
  reg         rob_uop_1_26_uses_ldq;
  reg         rob_uop_1_26_uses_stq;
  reg         rob_uop_1_26_is_sys_pc2epc;
  reg         rob_uop_1_26_flush_on_commit;
  reg  [5:0]  rob_uop_1_26_ldst;
  reg         rob_uop_1_26_ldst_val;
  reg  [1:0]  rob_uop_1_26_dst_rtype;
  reg         rob_uop_1_26_fp_val;
  reg  [1:0]  rob_uop_1_26_debug_fsrc;
  reg  [6:0]  rob_uop_1_27_uopc;
  reg         rob_uop_1_27_is_rvc;
  reg         rob_uop_1_27_is_br;
  reg         rob_uop_1_27_is_jalr;
  reg         rob_uop_1_27_is_jal;
  reg  [19:0] rob_uop_1_27_br_mask;
  reg  [5:0]  rob_uop_1_27_ftq_idx;
  reg         rob_uop_1_27_edge_inst;
  reg  [5:0]  rob_uop_1_27_pc_lob;
  reg  [6:0]  rob_uop_1_27_pdst;
  reg  [6:0]  rob_uop_1_27_stale_pdst;
  reg         rob_uop_1_27_is_fencei;
  reg         rob_uop_1_27_uses_ldq;
  reg         rob_uop_1_27_uses_stq;
  reg         rob_uop_1_27_is_sys_pc2epc;
  reg         rob_uop_1_27_flush_on_commit;
  reg  [5:0]  rob_uop_1_27_ldst;
  reg         rob_uop_1_27_ldst_val;
  reg  [1:0]  rob_uop_1_27_dst_rtype;
  reg         rob_uop_1_27_fp_val;
  reg  [1:0]  rob_uop_1_27_debug_fsrc;
  reg  [6:0]  rob_uop_1_28_uopc;
  reg         rob_uop_1_28_is_rvc;
  reg         rob_uop_1_28_is_br;
  reg         rob_uop_1_28_is_jalr;
  reg         rob_uop_1_28_is_jal;
  reg  [19:0] rob_uop_1_28_br_mask;
  reg  [5:0]  rob_uop_1_28_ftq_idx;
  reg         rob_uop_1_28_edge_inst;
  reg  [5:0]  rob_uop_1_28_pc_lob;
  reg  [6:0]  rob_uop_1_28_pdst;
  reg  [6:0]  rob_uop_1_28_stale_pdst;
  reg         rob_uop_1_28_is_fencei;
  reg         rob_uop_1_28_uses_ldq;
  reg         rob_uop_1_28_uses_stq;
  reg         rob_uop_1_28_is_sys_pc2epc;
  reg         rob_uop_1_28_flush_on_commit;
  reg  [5:0]  rob_uop_1_28_ldst;
  reg         rob_uop_1_28_ldst_val;
  reg  [1:0]  rob_uop_1_28_dst_rtype;
  reg         rob_uop_1_28_fp_val;
  reg  [1:0]  rob_uop_1_28_debug_fsrc;
  reg  [6:0]  rob_uop_1_29_uopc;
  reg         rob_uop_1_29_is_rvc;
  reg         rob_uop_1_29_is_br;
  reg         rob_uop_1_29_is_jalr;
  reg         rob_uop_1_29_is_jal;
  reg  [19:0] rob_uop_1_29_br_mask;
  reg  [5:0]  rob_uop_1_29_ftq_idx;
  reg         rob_uop_1_29_edge_inst;
  reg  [5:0]  rob_uop_1_29_pc_lob;
  reg  [6:0]  rob_uop_1_29_pdst;
  reg  [6:0]  rob_uop_1_29_stale_pdst;
  reg         rob_uop_1_29_is_fencei;
  reg         rob_uop_1_29_uses_ldq;
  reg         rob_uop_1_29_uses_stq;
  reg         rob_uop_1_29_is_sys_pc2epc;
  reg         rob_uop_1_29_flush_on_commit;
  reg  [5:0]  rob_uop_1_29_ldst;
  reg         rob_uop_1_29_ldst_val;
  reg  [1:0]  rob_uop_1_29_dst_rtype;
  reg         rob_uop_1_29_fp_val;
  reg  [1:0]  rob_uop_1_29_debug_fsrc;
  reg  [6:0]  rob_uop_1_30_uopc;
  reg         rob_uop_1_30_is_rvc;
  reg         rob_uop_1_30_is_br;
  reg         rob_uop_1_30_is_jalr;
  reg         rob_uop_1_30_is_jal;
  reg  [19:0] rob_uop_1_30_br_mask;
  reg  [5:0]  rob_uop_1_30_ftq_idx;
  reg         rob_uop_1_30_edge_inst;
  reg  [5:0]  rob_uop_1_30_pc_lob;
  reg  [6:0]  rob_uop_1_30_pdst;
  reg  [6:0]  rob_uop_1_30_stale_pdst;
  reg         rob_uop_1_30_is_fencei;
  reg         rob_uop_1_30_uses_ldq;
  reg         rob_uop_1_30_uses_stq;
  reg         rob_uop_1_30_is_sys_pc2epc;
  reg         rob_uop_1_30_flush_on_commit;
  reg  [5:0]  rob_uop_1_30_ldst;
  reg         rob_uop_1_30_ldst_val;
  reg  [1:0]  rob_uop_1_30_dst_rtype;
  reg         rob_uop_1_30_fp_val;
  reg  [1:0]  rob_uop_1_30_debug_fsrc;
  reg  [6:0]  rob_uop_1_31_uopc;
  reg         rob_uop_1_31_is_rvc;
  reg         rob_uop_1_31_is_br;
  reg         rob_uop_1_31_is_jalr;
  reg         rob_uop_1_31_is_jal;
  reg  [19:0] rob_uop_1_31_br_mask;
  reg  [5:0]  rob_uop_1_31_ftq_idx;
  reg         rob_uop_1_31_edge_inst;
  reg  [5:0]  rob_uop_1_31_pc_lob;
  reg  [6:0]  rob_uop_1_31_pdst;
  reg  [6:0]  rob_uop_1_31_stale_pdst;
  reg         rob_uop_1_31_is_fencei;
  reg         rob_uop_1_31_uses_ldq;
  reg         rob_uop_1_31_uses_stq;
  reg         rob_uop_1_31_is_sys_pc2epc;
  reg         rob_uop_1_31_flush_on_commit;
  reg  [5:0]  rob_uop_1_31_ldst;
  reg         rob_uop_1_31_ldst_val;
  reg  [1:0]  rob_uop_1_31_dst_rtype;
  reg         rob_uop_1_31_fp_val;
  reg  [1:0]  rob_uop_1_31_debug_fsrc;
  reg         rob_exception_1_0;
  reg         rob_exception_1_1;
  reg         rob_exception_1_2;
  reg         rob_exception_1_3;
  reg         rob_exception_1_4;
  reg         rob_exception_1_5;
  reg         rob_exception_1_6;
  reg         rob_exception_1_7;
  reg         rob_exception_1_8;
  reg         rob_exception_1_9;
  reg         rob_exception_1_10;
  reg         rob_exception_1_11;
  reg         rob_exception_1_12;
  reg         rob_exception_1_13;
  reg         rob_exception_1_14;
  reg         rob_exception_1_15;
  reg         rob_exception_1_16;
  reg         rob_exception_1_17;
  reg         rob_exception_1_18;
  reg         rob_exception_1_19;
  reg         rob_exception_1_20;
  reg         rob_exception_1_21;
  reg         rob_exception_1_22;
  reg         rob_exception_1_23;
  reg         rob_exception_1_24;
  reg         rob_exception_1_25;
  reg         rob_exception_1_26;
  reg         rob_exception_1_27;
  reg         rob_exception_1_28;
  reg         rob_exception_1_29;
  reg         rob_exception_1_30;
  reg         rob_exception_1_31;
  reg         rob_predicated_1_0;
  reg         rob_predicated_1_1;
  reg         rob_predicated_1_2;
  reg         rob_predicated_1_3;
  reg         rob_predicated_1_4;
  reg         rob_predicated_1_5;
  reg         rob_predicated_1_6;
  reg         rob_predicated_1_7;
  reg         rob_predicated_1_8;
  reg         rob_predicated_1_9;
  reg         rob_predicated_1_10;
  reg         rob_predicated_1_11;
  reg         rob_predicated_1_12;
  reg         rob_predicated_1_13;
  reg         rob_predicated_1_14;
  reg         rob_predicated_1_15;
  reg         rob_predicated_1_16;
  reg         rob_predicated_1_17;
  reg         rob_predicated_1_18;
  reg         rob_predicated_1_19;
  reg         rob_predicated_1_20;
  reg         rob_predicated_1_21;
  reg         rob_predicated_1_22;
  reg         rob_predicated_1_23;
  reg         rob_predicated_1_24;
  reg         rob_predicated_1_25;
  reg         rob_predicated_1_26;
  reg         rob_predicated_1_27;
  reg         rob_predicated_1_28;
  reg         rob_predicated_1_29;
  reg         rob_predicated_1_30;
  reg         rob_predicated_1_31;
  reg         casez_tmp_77;
  always @(*) begin
    casez (rob_tail)
      5'b00000:
        casez_tmp_77 = rob_val_1_0;
      5'b00001:
        casez_tmp_77 = rob_val_1_1;
      5'b00010:
        casez_tmp_77 = rob_val_1_2;
      5'b00011:
        casez_tmp_77 = rob_val_1_3;
      5'b00100:
        casez_tmp_77 = rob_val_1_4;
      5'b00101:
        casez_tmp_77 = rob_val_1_5;
      5'b00110:
        casez_tmp_77 = rob_val_1_6;
      5'b00111:
        casez_tmp_77 = rob_val_1_7;
      5'b01000:
        casez_tmp_77 = rob_val_1_8;
      5'b01001:
        casez_tmp_77 = rob_val_1_9;
      5'b01010:
        casez_tmp_77 = rob_val_1_10;
      5'b01011:
        casez_tmp_77 = rob_val_1_11;
      5'b01100:
        casez_tmp_77 = rob_val_1_12;
      5'b01101:
        casez_tmp_77 = rob_val_1_13;
      5'b01110:
        casez_tmp_77 = rob_val_1_14;
      5'b01111:
        casez_tmp_77 = rob_val_1_15;
      5'b10000:
        casez_tmp_77 = rob_val_1_16;
      5'b10001:
        casez_tmp_77 = rob_val_1_17;
      5'b10010:
        casez_tmp_77 = rob_val_1_18;
      5'b10011:
        casez_tmp_77 = rob_val_1_19;
      5'b10100:
        casez_tmp_77 = rob_val_1_20;
      5'b10101:
        casez_tmp_77 = rob_val_1_21;
      5'b10110:
        casez_tmp_77 = rob_val_1_22;
      5'b10111:
        casez_tmp_77 = rob_val_1_23;
      5'b11000:
        casez_tmp_77 = rob_val_1_24;
      5'b11001:
        casez_tmp_77 = rob_val_1_25;
      5'b11010:
        casez_tmp_77 = rob_val_1_26;
      5'b11011:
        casez_tmp_77 = rob_val_1_27;
      5'b11100:
        casez_tmp_77 = rob_val_1_28;
      5'b11101:
        casez_tmp_77 = rob_val_1_29;
      5'b11110:
        casez_tmp_77 = rob_val_1_30;
      default:
        casez_tmp_77 = rob_val_1_31;
    endcase
  end // always @(*)
  wire        _GEN_17 = io_wb_resps_0_valid & io_wb_resps_0_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_18 = io_wb_resps_1_valid & io_wb_resps_1_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_19 = io_wb_resps_2_valid & io_wb_resps_2_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_20 = io_wb_resps_3_valid & io_wb_resps_3_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_21 = io_wb_resps_4_valid & io_wb_resps_4_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_22 = io_wb_resps_5_valid & io_wb_resps_5_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_23 = io_wb_resps_6_valid & io_wb_resps_6_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_24 = io_wb_resps_7_valid & io_wb_resps_7_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_25 = io_wb_resps_8_valid & io_wb_resps_8_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_26 = io_wb_resps_9_valid & io_wb_resps_9_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_27 = io_lsu_clr_bsy_0_valid & io_lsu_clr_bsy_0_bits[1:0] == 2'h1;
  reg         casez_tmp_78;
  always @(*) begin
    casez (io_lsu_clr_bsy_0_bits[6:2])
      5'b00000:
        casez_tmp_78 = rob_val_1_0;
      5'b00001:
        casez_tmp_78 = rob_val_1_1;
      5'b00010:
        casez_tmp_78 = rob_val_1_2;
      5'b00011:
        casez_tmp_78 = rob_val_1_3;
      5'b00100:
        casez_tmp_78 = rob_val_1_4;
      5'b00101:
        casez_tmp_78 = rob_val_1_5;
      5'b00110:
        casez_tmp_78 = rob_val_1_6;
      5'b00111:
        casez_tmp_78 = rob_val_1_7;
      5'b01000:
        casez_tmp_78 = rob_val_1_8;
      5'b01001:
        casez_tmp_78 = rob_val_1_9;
      5'b01010:
        casez_tmp_78 = rob_val_1_10;
      5'b01011:
        casez_tmp_78 = rob_val_1_11;
      5'b01100:
        casez_tmp_78 = rob_val_1_12;
      5'b01101:
        casez_tmp_78 = rob_val_1_13;
      5'b01110:
        casez_tmp_78 = rob_val_1_14;
      5'b01111:
        casez_tmp_78 = rob_val_1_15;
      5'b10000:
        casez_tmp_78 = rob_val_1_16;
      5'b10001:
        casez_tmp_78 = rob_val_1_17;
      5'b10010:
        casez_tmp_78 = rob_val_1_18;
      5'b10011:
        casez_tmp_78 = rob_val_1_19;
      5'b10100:
        casez_tmp_78 = rob_val_1_20;
      5'b10101:
        casez_tmp_78 = rob_val_1_21;
      5'b10110:
        casez_tmp_78 = rob_val_1_22;
      5'b10111:
        casez_tmp_78 = rob_val_1_23;
      5'b11000:
        casez_tmp_78 = rob_val_1_24;
      5'b11001:
        casez_tmp_78 = rob_val_1_25;
      5'b11010:
        casez_tmp_78 = rob_val_1_26;
      5'b11011:
        casez_tmp_78 = rob_val_1_27;
      5'b11100:
        casez_tmp_78 = rob_val_1_28;
      5'b11101:
        casez_tmp_78 = rob_val_1_29;
      5'b11110:
        casez_tmp_78 = rob_val_1_30;
      default:
        casez_tmp_78 = rob_val_1_31;
    endcase
  end // always @(*)
  reg         casez_tmp_79;
  always @(*) begin
    casez (io_lsu_clr_bsy_0_bits[6:2])
      5'b00000:
        casez_tmp_79 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_79 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_79 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_79 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_79 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_79 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_79 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_79 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_79 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_79 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_79 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_79 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_79 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_79 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_79 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_79 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_79 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_79 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_79 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_79 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_79 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_79 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_79 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_79 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_79 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_79 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_79 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_79 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_79 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_79 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_79 = rob_bsy_1_30;
      default:
        casez_tmp_79 = rob_bsy_1_31;
    endcase
  end // always @(*)
  wire        _GEN_28 = io_lsu_clr_bsy_1_valid & io_lsu_clr_bsy_1_bits[1:0] == 2'h1;
  reg         casez_tmp_80;
  always @(*) begin
    casez (io_lsu_clr_bsy_1_bits[6:2])
      5'b00000:
        casez_tmp_80 = rob_val_1_0;
      5'b00001:
        casez_tmp_80 = rob_val_1_1;
      5'b00010:
        casez_tmp_80 = rob_val_1_2;
      5'b00011:
        casez_tmp_80 = rob_val_1_3;
      5'b00100:
        casez_tmp_80 = rob_val_1_4;
      5'b00101:
        casez_tmp_80 = rob_val_1_5;
      5'b00110:
        casez_tmp_80 = rob_val_1_6;
      5'b00111:
        casez_tmp_80 = rob_val_1_7;
      5'b01000:
        casez_tmp_80 = rob_val_1_8;
      5'b01001:
        casez_tmp_80 = rob_val_1_9;
      5'b01010:
        casez_tmp_80 = rob_val_1_10;
      5'b01011:
        casez_tmp_80 = rob_val_1_11;
      5'b01100:
        casez_tmp_80 = rob_val_1_12;
      5'b01101:
        casez_tmp_80 = rob_val_1_13;
      5'b01110:
        casez_tmp_80 = rob_val_1_14;
      5'b01111:
        casez_tmp_80 = rob_val_1_15;
      5'b10000:
        casez_tmp_80 = rob_val_1_16;
      5'b10001:
        casez_tmp_80 = rob_val_1_17;
      5'b10010:
        casez_tmp_80 = rob_val_1_18;
      5'b10011:
        casez_tmp_80 = rob_val_1_19;
      5'b10100:
        casez_tmp_80 = rob_val_1_20;
      5'b10101:
        casez_tmp_80 = rob_val_1_21;
      5'b10110:
        casez_tmp_80 = rob_val_1_22;
      5'b10111:
        casez_tmp_80 = rob_val_1_23;
      5'b11000:
        casez_tmp_80 = rob_val_1_24;
      5'b11001:
        casez_tmp_80 = rob_val_1_25;
      5'b11010:
        casez_tmp_80 = rob_val_1_26;
      5'b11011:
        casez_tmp_80 = rob_val_1_27;
      5'b11100:
        casez_tmp_80 = rob_val_1_28;
      5'b11101:
        casez_tmp_80 = rob_val_1_29;
      5'b11110:
        casez_tmp_80 = rob_val_1_30;
      default:
        casez_tmp_80 = rob_val_1_31;
    endcase
  end // always @(*)
  reg         casez_tmp_81;
  always @(*) begin
    casez (io_lsu_clr_bsy_1_bits[6:2])
      5'b00000:
        casez_tmp_81 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_81 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_81 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_81 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_81 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_81 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_81 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_81 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_81 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_81 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_81 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_81 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_81 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_81 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_81 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_81 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_81 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_81 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_81 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_81 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_81 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_81 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_81 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_81 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_81 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_81 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_81 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_81 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_81 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_81 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_81 = rob_bsy_1_30;
      default:
        casez_tmp_81 = rob_bsy_1_31;
    endcase
  end // always @(*)
  wire        _GEN_29 = io_lsu_clr_bsy_2_valid & io_lsu_clr_bsy_2_bits[1:0] == 2'h1;
  reg         casez_tmp_82;
  always @(*) begin
    casez (io_lsu_clr_bsy_2_bits[6:2])
      5'b00000:
        casez_tmp_82 = rob_val_1_0;
      5'b00001:
        casez_tmp_82 = rob_val_1_1;
      5'b00010:
        casez_tmp_82 = rob_val_1_2;
      5'b00011:
        casez_tmp_82 = rob_val_1_3;
      5'b00100:
        casez_tmp_82 = rob_val_1_4;
      5'b00101:
        casez_tmp_82 = rob_val_1_5;
      5'b00110:
        casez_tmp_82 = rob_val_1_6;
      5'b00111:
        casez_tmp_82 = rob_val_1_7;
      5'b01000:
        casez_tmp_82 = rob_val_1_8;
      5'b01001:
        casez_tmp_82 = rob_val_1_9;
      5'b01010:
        casez_tmp_82 = rob_val_1_10;
      5'b01011:
        casez_tmp_82 = rob_val_1_11;
      5'b01100:
        casez_tmp_82 = rob_val_1_12;
      5'b01101:
        casez_tmp_82 = rob_val_1_13;
      5'b01110:
        casez_tmp_82 = rob_val_1_14;
      5'b01111:
        casez_tmp_82 = rob_val_1_15;
      5'b10000:
        casez_tmp_82 = rob_val_1_16;
      5'b10001:
        casez_tmp_82 = rob_val_1_17;
      5'b10010:
        casez_tmp_82 = rob_val_1_18;
      5'b10011:
        casez_tmp_82 = rob_val_1_19;
      5'b10100:
        casez_tmp_82 = rob_val_1_20;
      5'b10101:
        casez_tmp_82 = rob_val_1_21;
      5'b10110:
        casez_tmp_82 = rob_val_1_22;
      5'b10111:
        casez_tmp_82 = rob_val_1_23;
      5'b11000:
        casez_tmp_82 = rob_val_1_24;
      5'b11001:
        casez_tmp_82 = rob_val_1_25;
      5'b11010:
        casez_tmp_82 = rob_val_1_26;
      5'b11011:
        casez_tmp_82 = rob_val_1_27;
      5'b11100:
        casez_tmp_82 = rob_val_1_28;
      5'b11101:
        casez_tmp_82 = rob_val_1_29;
      5'b11110:
        casez_tmp_82 = rob_val_1_30;
      default:
        casez_tmp_82 = rob_val_1_31;
    endcase
  end // always @(*)
  reg         casez_tmp_83;
  always @(*) begin
    casez (io_lsu_clr_bsy_2_bits[6:2])
      5'b00000:
        casez_tmp_83 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_83 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_83 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_83 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_83 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_83 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_83 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_83 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_83 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_83 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_83 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_83 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_83 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_83 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_83 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_83 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_83 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_83 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_83 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_83 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_83 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_83 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_83 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_83 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_83 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_83 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_83 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_83 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_83 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_83 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_83 = rob_bsy_1_30;
      default:
        casez_tmp_83 = rob_bsy_1_31;
    endcase
  end // always @(*)
  wire        _GEN_30 = io_lxcpt_valid & io_lxcpt_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_31 = _GEN_30 & _GEN_13 & ~reset;
  reg         casez_tmp_84;
  always @(*) begin
    casez (io_lxcpt_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_84 = rob_unsafe_1_0;
      5'b00001:
        casez_tmp_84 = rob_unsafe_1_1;
      5'b00010:
        casez_tmp_84 = rob_unsafe_1_2;
      5'b00011:
        casez_tmp_84 = rob_unsafe_1_3;
      5'b00100:
        casez_tmp_84 = rob_unsafe_1_4;
      5'b00101:
        casez_tmp_84 = rob_unsafe_1_5;
      5'b00110:
        casez_tmp_84 = rob_unsafe_1_6;
      5'b00111:
        casez_tmp_84 = rob_unsafe_1_7;
      5'b01000:
        casez_tmp_84 = rob_unsafe_1_8;
      5'b01001:
        casez_tmp_84 = rob_unsafe_1_9;
      5'b01010:
        casez_tmp_84 = rob_unsafe_1_10;
      5'b01011:
        casez_tmp_84 = rob_unsafe_1_11;
      5'b01100:
        casez_tmp_84 = rob_unsafe_1_12;
      5'b01101:
        casez_tmp_84 = rob_unsafe_1_13;
      5'b01110:
        casez_tmp_84 = rob_unsafe_1_14;
      5'b01111:
        casez_tmp_84 = rob_unsafe_1_15;
      5'b10000:
        casez_tmp_84 = rob_unsafe_1_16;
      5'b10001:
        casez_tmp_84 = rob_unsafe_1_17;
      5'b10010:
        casez_tmp_84 = rob_unsafe_1_18;
      5'b10011:
        casez_tmp_84 = rob_unsafe_1_19;
      5'b10100:
        casez_tmp_84 = rob_unsafe_1_20;
      5'b10101:
        casez_tmp_84 = rob_unsafe_1_21;
      5'b10110:
        casez_tmp_84 = rob_unsafe_1_22;
      5'b10111:
        casez_tmp_84 = rob_unsafe_1_23;
      5'b11000:
        casez_tmp_84 = rob_unsafe_1_24;
      5'b11001:
        casez_tmp_84 = rob_unsafe_1_25;
      5'b11010:
        casez_tmp_84 = rob_unsafe_1_26;
      5'b11011:
        casez_tmp_84 = rob_unsafe_1_27;
      5'b11100:
        casez_tmp_84 = rob_unsafe_1_28;
      5'b11101:
        casez_tmp_84 = rob_unsafe_1_29;
      5'b11110:
        casez_tmp_84 = rob_unsafe_1_30;
      default:
        casez_tmp_84 = rob_unsafe_1_31;
    endcase
  end // always @(*)
  reg         casez_tmp_85;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_85 = rob_val_1_0;
      5'b00001:
        casez_tmp_85 = rob_val_1_1;
      5'b00010:
        casez_tmp_85 = rob_val_1_2;
      5'b00011:
        casez_tmp_85 = rob_val_1_3;
      5'b00100:
        casez_tmp_85 = rob_val_1_4;
      5'b00101:
        casez_tmp_85 = rob_val_1_5;
      5'b00110:
        casez_tmp_85 = rob_val_1_6;
      5'b00111:
        casez_tmp_85 = rob_val_1_7;
      5'b01000:
        casez_tmp_85 = rob_val_1_8;
      5'b01001:
        casez_tmp_85 = rob_val_1_9;
      5'b01010:
        casez_tmp_85 = rob_val_1_10;
      5'b01011:
        casez_tmp_85 = rob_val_1_11;
      5'b01100:
        casez_tmp_85 = rob_val_1_12;
      5'b01101:
        casez_tmp_85 = rob_val_1_13;
      5'b01110:
        casez_tmp_85 = rob_val_1_14;
      5'b01111:
        casez_tmp_85 = rob_val_1_15;
      5'b10000:
        casez_tmp_85 = rob_val_1_16;
      5'b10001:
        casez_tmp_85 = rob_val_1_17;
      5'b10010:
        casez_tmp_85 = rob_val_1_18;
      5'b10011:
        casez_tmp_85 = rob_val_1_19;
      5'b10100:
        casez_tmp_85 = rob_val_1_20;
      5'b10101:
        casez_tmp_85 = rob_val_1_21;
      5'b10110:
        casez_tmp_85 = rob_val_1_22;
      5'b10111:
        casez_tmp_85 = rob_val_1_23;
      5'b11000:
        casez_tmp_85 = rob_val_1_24;
      5'b11001:
        casez_tmp_85 = rob_val_1_25;
      5'b11010:
        casez_tmp_85 = rob_val_1_26;
      5'b11011:
        casez_tmp_85 = rob_val_1_27;
      5'b11100:
        casez_tmp_85 = rob_val_1_28;
      5'b11101:
        casez_tmp_85 = rob_val_1_29;
      5'b11110:
        casez_tmp_85 = rob_val_1_30;
      default:
        casez_tmp_85 = rob_val_1_31;
    endcase
  end // always @(*)
  reg         casez_tmp_86;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_86 = rob_exception_1_0;
      5'b00001:
        casez_tmp_86 = rob_exception_1_1;
      5'b00010:
        casez_tmp_86 = rob_exception_1_2;
      5'b00011:
        casez_tmp_86 = rob_exception_1_3;
      5'b00100:
        casez_tmp_86 = rob_exception_1_4;
      5'b00101:
        casez_tmp_86 = rob_exception_1_5;
      5'b00110:
        casez_tmp_86 = rob_exception_1_6;
      5'b00111:
        casez_tmp_86 = rob_exception_1_7;
      5'b01000:
        casez_tmp_86 = rob_exception_1_8;
      5'b01001:
        casez_tmp_86 = rob_exception_1_9;
      5'b01010:
        casez_tmp_86 = rob_exception_1_10;
      5'b01011:
        casez_tmp_86 = rob_exception_1_11;
      5'b01100:
        casez_tmp_86 = rob_exception_1_12;
      5'b01101:
        casez_tmp_86 = rob_exception_1_13;
      5'b01110:
        casez_tmp_86 = rob_exception_1_14;
      5'b01111:
        casez_tmp_86 = rob_exception_1_15;
      5'b10000:
        casez_tmp_86 = rob_exception_1_16;
      5'b10001:
        casez_tmp_86 = rob_exception_1_17;
      5'b10010:
        casez_tmp_86 = rob_exception_1_18;
      5'b10011:
        casez_tmp_86 = rob_exception_1_19;
      5'b10100:
        casez_tmp_86 = rob_exception_1_20;
      5'b10101:
        casez_tmp_86 = rob_exception_1_21;
      5'b10110:
        casez_tmp_86 = rob_exception_1_22;
      5'b10111:
        casez_tmp_86 = rob_exception_1_23;
      5'b11000:
        casez_tmp_86 = rob_exception_1_24;
      5'b11001:
        casez_tmp_86 = rob_exception_1_25;
      5'b11010:
        casez_tmp_86 = rob_exception_1_26;
      5'b11011:
        casez_tmp_86 = rob_exception_1_27;
      5'b11100:
        casez_tmp_86 = rob_exception_1_28;
      5'b11101:
        casez_tmp_86 = rob_exception_1_29;
      5'b11110:
        casez_tmp_86 = rob_exception_1_30;
      default:
        casez_tmp_86 = rob_exception_1_31;
    endcase
  end // always @(*)
  wire        can_throw_exception_1 = casez_tmp_85 & casez_tmp_86;
  reg         casez_tmp_87;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_87 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_87 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_87 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_87 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_87 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_87 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_87 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_87 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_87 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_87 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_87 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_87 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_87 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_87 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_87 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_87 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_87 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_87 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_87 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_87 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_87 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_87 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_87 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_87 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_87 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_87 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_87 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_87 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_87 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_87 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_87 = rob_bsy_1_30;
      default:
        casez_tmp_87 = rob_bsy_1_31;
    endcase
  end // always @(*)
  wire        can_commit_1 = casez_tmp_85 & ~casez_tmp_87 & ~io_csr_stall;
  reg         casez_tmp_88;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_88 = rob_predicated_1_0;
      5'b00001:
        casez_tmp_88 = rob_predicated_1_1;
      5'b00010:
        casez_tmp_88 = rob_predicated_1_2;
      5'b00011:
        casez_tmp_88 = rob_predicated_1_3;
      5'b00100:
        casez_tmp_88 = rob_predicated_1_4;
      5'b00101:
        casez_tmp_88 = rob_predicated_1_5;
      5'b00110:
        casez_tmp_88 = rob_predicated_1_6;
      5'b00111:
        casez_tmp_88 = rob_predicated_1_7;
      5'b01000:
        casez_tmp_88 = rob_predicated_1_8;
      5'b01001:
        casez_tmp_88 = rob_predicated_1_9;
      5'b01010:
        casez_tmp_88 = rob_predicated_1_10;
      5'b01011:
        casez_tmp_88 = rob_predicated_1_11;
      5'b01100:
        casez_tmp_88 = rob_predicated_1_12;
      5'b01101:
        casez_tmp_88 = rob_predicated_1_13;
      5'b01110:
        casez_tmp_88 = rob_predicated_1_14;
      5'b01111:
        casez_tmp_88 = rob_predicated_1_15;
      5'b10000:
        casez_tmp_88 = rob_predicated_1_16;
      5'b10001:
        casez_tmp_88 = rob_predicated_1_17;
      5'b10010:
        casez_tmp_88 = rob_predicated_1_18;
      5'b10011:
        casez_tmp_88 = rob_predicated_1_19;
      5'b10100:
        casez_tmp_88 = rob_predicated_1_20;
      5'b10101:
        casez_tmp_88 = rob_predicated_1_21;
      5'b10110:
        casez_tmp_88 = rob_predicated_1_22;
      5'b10111:
        casez_tmp_88 = rob_predicated_1_23;
      5'b11000:
        casez_tmp_88 = rob_predicated_1_24;
      5'b11001:
        casez_tmp_88 = rob_predicated_1_25;
      5'b11010:
        casez_tmp_88 = rob_predicated_1_26;
      5'b11011:
        casez_tmp_88 = rob_predicated_1_27;
      5'b11100:
        casez_tmp_88 = rob_predicated_1_28;
      5'b11101:
        casez_tmp_88 = rob_predicated_1_29;
      5'b11110:
        casez_tmp_88 = rob_predicated_1_30;
      default:
        casez_tmp_88 = rob_predicated_1_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_89;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_89 = rob_uop_1_0_uopc;
      5'b00001:
        casez_tmp_89 = rob_uop_1_1_uopc;
      5'b00010:
        casez_tmp_89 = rob_uop_1_2_uopc;
      5'b00011:
        casez_tmp_89 = rob_uop_1_3_uopc;
      5'b00100:
        casez_tmp_89 = rob_uop_1_4_uopc;
      5'b00101:
        casez_tmp_89 = rob_uop_1_5_uopc;
      5'b00110:
        casez_tmp_89 = rob_uop_1_6_uopc;
      5'b00111:
        casez_tmp_89 = rob_uop_1_7_uopc;
      5'b01000:
        casez_tmp_89 = rob_uop_1_8_uopc;
      5'b01001:
        casez_tmp_89 = rob_uop_1_9_uopc;
      5'b01010:
        casez_tmp_89 = rob_uop_1_10_uopc;
      5'b01011:
        casez_tmp_89 = rob_uop_1_11_uopc;
      5'b01100:
        casez_tmp_89 = rob_uop_1_12_uopc;
      5'b01101:
        casez_tmp_89 = rob_uop_1_13_uopc;
      5'b01110:
        casez_tmp_89 = rob_uop_1_14_uopc;
      5'b01111:
        casez_tmp_89 = rob_uop_1_15_uopc;
      5'b10000:
        casez_tmp_89 = rob_uop_1_16_uopc;
      5'b10001:
        casez_tmp_89 = rob_uop_1_17_uopc;
      5'b10010:
        casez_tmp_89 = rob_uop_1_18_uopc;
      5'b10011:
        casez_tmp_89 = rob_uop_1_19_uopc;
      5'b10100:
        casez_tmp_89 = rob_uop_1_20_uopc;
      5'b10101:
        casez_tmp_89 = rob_uop_1_21_uopc;
      5'b10110:
        casez_tmp_89 = rob_uop_1_22_uopc;
      5'b10111:
        casez_tmp_89 = rob_uop_1_23_uopc;
      5'b11000:
        casez_tmp_89 = rob_uop_1_24_uopc;
      5'b11001:
        casez_tmp_89 = rob_uop_1_25_uopc;
      5'b11010:
        casez_tmp_89 = rob_uop_1_26_uopc;
      5'b11011:
        casez_tmp_89 = rob_uop_1_27_uopc;
      5'b11100:
        casez_tmp_89 = rob_uop_1_28_uopc;
      5'b11101:
        casez_tmp_89 = rob_uop_1_29_uopc;
      5'b11110:
        casez_tmp_89 = rob_uop_1_30_uopc;
      default:
        casez_tmp_89 = rob_uop_1_31_uopc;
    endcase
  end // always @(*)
  reg         casez_tmp_90;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_90 = rob_uop_1_0_is_rvc;
      5'b00001:
        casez_tmp_90 = rob_uop_1_1_is_rvc;
      5'b00010:
        casez_tmp_90 = rob_uop_1_2_is_rvc;
      5'b00011:
        casez_tmp_90 = rob_uop_1_3_is_rvc;
      5'b00100:
        casez_tmp_90 = rob_uop_1_4_is_rvc;
      5'b00101:
        casez_tmp_90 = rob_uop_1_5_is_rvc;
      5'b00110:
        casez_tmp_90 = rob_uop_1_6_is_rvc;
      5'b00111:
        casez_tmp_90 = rob_uop_1_7_is_rvc;
      5'b01000:
        casez_tmp_90 = rob_uop_1_8_is_rvc;
      5'b01001:
        casez_tmp_90 = rob_uop_1_9_is_rvc;
      5'b01010:
        casez_tmp_90 = rob_uop_1_10_is_rvc;
      5'b01011:
        casez_tmp_90 = rob_uop_1_11_is_rvc;
      5'b01100:
        casez_tmp_90 = rob_uop_1_12_is_rvc;
      5'b01101:
        casez_tmp_90 = rob_uop_1_13_is_rvc;
      5'b01110:
        casez_tmp_90 = rob_uop_1_14_is_rvc;
      5'b01111:
        casez_tmp_90 = rob_uop_1_15_is_rvc;
      5'b10000:
        casez_tmp_90 = rob_uop_1_16_is_rvc;
      5'b10001:
        casez_tmp_90 = rob_uop_1_17_is_rvc;
      5'b10010:
        casez_tmp_90 = rob_uop_1_18_is_rvc;
      5'b10011:
        casez_tmp_90 = rob_uop_1_19_is_rvc;
      5'b10100:
        casez_tmp_90 = rob_uop_1_20_is_rvc;
      5'b10101:
        casez_tmp_90 = rob_uop_1_21_is_rvc;
      5'b10110:
        casez_tmp_90 = rob_uop_1_22_is_rvc;
      5'b10111:
        casez_tmp_90 = rob_uop_1_23_is_rvc;
      5'b11000:
        casez_tmp_90 = rob_uop_1_24_is_rvc;
      5'b11001:
        casez_tmp_90 = rob_uop_1_25_is_rvc;
      5'b11010:
        casez_tmp_90 = rob_uop_1_26_is_rvc;
      5'b11011:
        casez_tmp_90 = rob_uop_1_27_is_rvc;
      5'b11100:
        casez_tmp_90 = rob_uop_1_28_is_rvc;
      5'b11101:
        casez_tmp_90 = rob_uop_1_29_is_rvc;
      5'b11110:
        casez_tmp_90 = rob_uop_1_30_is_rvc;
      default:
        casez_tmp_90 = rob_uop_1_31_is_rvc;
    endcase
  end // always @(*)
  reg         casez_tmp_91;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_91 = rob_uop_1_0_is_br;
      5'b00001:
        casez_tmp_91 = rob_uop_1_1_is_br;
      5'b00010:
        casez_tmp_91 = rob_uop_1_2_is_br;
      5'b00011:
        casez_tmp_91 = rob_uop_1_3_is_br;
      5'b00100:
        casez_tmp_91 = rob_uop_1_4_is_br;
      5'b00101:
        casez_tmp_91 = rob_uop_1_5_is_br;
      5'b00110:
        casez_tmp_91 = rob_uop_1_6_is_br;
      5'b00111:
        casez_tmp_91 = rob_uop_1_7_is_br;
      5'b01000:
        casez_tmp_91 = rob_uop_1_8_is_br;
      5'b01001:
        casez_tmp_91 = rob_uop_1_9_is_br;
      5'b01010:
        casez_tmp_91 = rob_uop_1_10_is_br;
      5'b01011:
        casez_tmp_91 = rob_uop_1_11_is_br;
      5'b01100:
        casez_tmp_91 = rob_uop_1_12_is_br;
      5'b01101:
        casez_tmp_91 = rob_uop_1_13_is_br;
      5'b01110:
        casez_tmp_91 = rob_uop_1_14_is_br;
      5'b01111:
        casez_tmp_91 = rob_uop_1_15_is_br;
      5'b10000:
        casez_tmp_91 = rob_uop_1_16_is_br;
      5'b10001:
        casez_tmp_91 = rob_uop_1_17_is_br;
      5'b10010:
        casez_tmp_91 = rob_uop_1_18_is_br;
      5'b10011:
        casez_tmp_91 = rob_uop_1_19_is_br;
      5'b10100:
        casez_tmp_91 = rob_uop_1_20_is_br;
      5'b10101:
        casez_tmp_91 = rob_uop_1_21_is_br;
      5'b10110:
        casez_tmp_91 = rob_uop_1_22_is_br;
      5'b10111:
        casez_tmp_91 = rob_uop_1_23_is_br;
      5'b11000:
        casez_tmp_91 = rob_uop_1_24_is_br;
      5'b11001:
        casez_tmp_91 = rob_uop_1_25_is_br;
      5'b11010:
        casez_tmp_91 = rob_uop_1_26_is_br;
      5'b11011:
        casez_tmp_91 = rob_uop_1_27_is_br;
      5'b11100:
        casez_tmp_91 = rob_uop_1_28_is_br;
      5'b11101:
        casez_tmp_91 = rob_uop_1_29_is_br;
      5'b11110:
        casez_tmp_91 = rob_uop_1_30_is_br;
      default:
        casez_tmp_91 = rob_uop_1_31_is_br;
    endcase
  end // always @(*)
  reg         casez_tmp_92;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_92 = rob_uop_1_0_is_jalr;
      5'b00001:
        casez_tmp_92 = rob_uop_1_1_is_jalr;
      5'b00010:
        casez_tmp_92 = rob_uop_1_2_is_jalr;
      5'b00011:
        casez_tmp_92 = rob_uop_1_3_is_jalr;
      5'b00100:
        casez_tmp_92 = rob_uop_1_4_is_jalr;
      5'b00101:
        casez_tmp_92 = rob_uop_1_5_is_jalr;
      5'b00110:
        casez_tmp_92 = rob_uop_1_6_is_jalr;
      5'b00111:
        casez_tmp_92 = rob_uop_1_7_is_jalr;
      5'b01000:
        casez_tmp_92 = rob_uop_1_8_is_jalr;
      5'b01001:
        casez_tmp_92 = rob_uop_1_9_is_jalr;
      5'b01010:
        casez_tmp_92 = rob_uop_1_10_is_jalr;
      5'b01011:
        casez_tmp_92 = rob_uop_1_11_is_jalr;
      5'b01100:
        casez_tmp_92 = rob_uop_1_12_is_jalr;
      5'b01101:
        casez_tmp_92 = rob_uop_1_13_is_jalr;
      5'b01110:
        casez_tmp_92 = rob_uop_1_14_is_jalr;
      5'b01111:
        casez_tmp_92 = rob_uop_1_15_is_jalr;
      5'b10000:
        casez_tmp_92 = rob_uop_1_16_is_jalr;
      5'b10001:
        casez_tmp_92 = rob_uop_1_17_is_jalr;
      5'b10010:
        casez_tmp_92 = rob_uop_1_18_is_jalr;
      5'b10011:
        casez_tmp_92 = rob_uop_1_19_is_jalr;
      5'b10100:
        casez_tmp_92 = rob_uop_1_20_is_jalr;
      5'b10101:
        casez_tmp_92 = rob_uop_1_21_is_jalr;
      5'b10110:
        casez_tmp_92 = rob_uop_1_22_is_jalr;
      5'b10111:
        casez_tmp_92 = rob_uop_1_23_is_jalr;
      5'b11000:
        casez_tmp_92 = rob_uop_1_24_is_jalr;
      5'b11001:
        casez_tmp_92 = rob_uop_1_25_is_jalr;
      5'b11010:
        casez_tmp_92 = rob_uop_1_26_is_jalr;
      5'b11011:
        casez_tmp_92 = rob_uop_1_27_is_jalr;
      5'b11100:
        casez_tmp_92 = rob_uop_1_28_is_jalr;
      5'b11101:
        casez_tmp_92 = rob_uop_1_29_is_jalr;
      5'b11110:
        casez_tmp_92 = rob_uop_1_30_is_jalr;
      default:
        casez_tmp_92 = rob_uop_1_31_is_jalr;
    endcase
  end // always @(*)
  reg         casez_tmp_93;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_93 = rob_uop_1_0_is_jal;
      5'b00001:
        casez_tmp_93 = rob_uop_1_1_is_jal;
      5'b00010:
        casez_tmp_93 = rob_uop_1_2_is_jal;
      5'b00011:
        casez_tmp_93 = rob_uop_1_3_is_jal;
      5'b00100:
        casez_tmp_93 = rob_uop_1_4_is_jal;
      5'b00101:
        casez_tmp_93 = rob_uop_1_5_is_jal;
      5'b00110:
        casez_tmp_93 = rob_uop_1_6_is_jal;
      5'b00111:
        casez_tmp_93 = rob_uop_1_7_is_jal;
      5'b01000:
        casez_tmp_93 = rob_uop_1_8_is_jal;
      5'b01001:
        casez_tmp_93 = rob_uop_1_9_is_jal;
      5'b01010:
        casez_tmp_93 = rob_uop_1_10_is_jal;
      5'b01011:
        casez_tmp_93 = rob_uop_1_11_is_jal;
      5'b01100:
        casez_tmp_93 = rob_uop_1_12_is_jal;
      5'b01101:
        casez_tmp_93 = rob_uop_1_13_is_jal;
      5'b01110:
        casez_tmp_93 = rob_uop_1_14_is_jal;
      5'b01111:
        casez_tmp_93 = rob_uop_1_15_is_jal;
      5'b10000:
        casez_tmp_93 = rob_uop_1_16_is_jal;
      5'b10001:
        casez_tmp_93 = rob_uop_1_17_is_jal;
      5'b10010:
        casez_tmp_93 = rob_uop_1_18_is_jal;
      5'b10011:
        casez_tmp_93 = rob_uop_1_19_is_jal;
      5'b10100:
        casez_tmp_93 = rob_uop_1_20_is_jal;
      5'b10101:
        casez_tmp_93 = rob_uop_1_21_is_jal;
      5'b10110:
        casez_tmp_93 = rob_uop_1_22_is_jal;
      5'b10111:
        casez_tmp_93 = rob_uop_1_23_is_jal;
      5'b11000:
        casez_tmp_93 = rob_uop_1_24_is_jal;
      5'b11001:
        casez_tmp_93 = rob_uop_1_25_is_jal;
      5'b11010:
        casez_tmp_93 = rob_uop_1_26_is_jal;
      5'b11011:
        casez_tmp_93 = rob_uop_1_27_is_jal;
      5'b11100:
        casez_tmp_93 = rob_uop_1_28_is_jal;
      5'b11101:
        casez_tmp_93 = rob_uop_1_29_is_jal;
      5'b11110:
        casez_tmp_93 = rob_uop_1_30_is_jal;
      default:
        casez_tmp_93 = rob_uop_1_31_is_jal;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_94;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_94 = rob_uop_1_0_ftq_idx;
      5'b00001:
        casez_tmp_94 = rob_uop_1_1_ftq_idx;
      5'b00010:
        casez_tmp_94 = rob_uop_1_2_ftq_idx;
      5'b00011:
        casez_tmp_94 = rob_uop_1_3_ftq_idx;
      5'b00100:
        casez_tmp_94 = rob_uop_1_4_ftq_idx;
      5'b00101:
        casez_tmp_94 = rob_uop_1_5_ftq_idx;
      5'b00110:
        casez_tmp_94 = rob_uop_1_6_ftq_idx;
      5'b00111:
        casez_tmp_94 = rob_uop_1_7_ftq_idx;
      5'b01000:
        casez_tmp_94 = rob_uop_1_8_ftq_idx;
      5'b01001:
        casez_tmp_94 = rob_uop_1_9_ftq_idx;
      5'b01010:
        casez_tmp_94 = rob_uop_1_10_ftq_idx;
      5'b01011:
        casez_tmp_94 = rob_uop_1_11_ftq_idx;
      5'b01100:
        casez_tmp_94 = rob_uop_1_12_ftq_idx;
      5'b01101:
        casez_tmp_94 = rob_uop_1_13_ftq_idx;
      5'b01110:
        casez_tmp_94 = rob_uop_1_14_ftq_idx;
      5'b01111:
        casez_tmp_94 = rob_uop_1_15_ftq_idx;
      5'b10000:
        casez_tmp_94 = rob_uop_1_16_ftq_idx;
      5'b10001:
        casez_tmp_94 = rob_uop_1_17_ftq_idx;
      5'b10010:
        casez_tmp_94 = rob_uop_1_18_ftq_idx;
      5'b10011:
        casez_tmp_94 = rob_uop_1_19_ftq_idx;
      5'b10100:
        casez_tmp_94 = rob_uop_1_20_ftq_idx;
      5'b10101:
        casez_tmp_94 = rob_uop_1_21_ftq_idx;
      5'b10110:
        casez_tmp_94 = rob_uop_1_22_ftq_idx;
      5'b10111:
        casez_tmp_94 = rob_uop_1_23_ftq_idx;
      5'b11000:
        casez_tmp_94 = rob_uop_1_24_ftq_idx;
      5'b11001:
        casez_tmp_94 = rob_uop_1_25_ftq_idx;
      5'b11010:
        casez_tmp_94 = rob_uop_1_26_ftq_idx;
      5'b11011:
        casez_tmp_94 = rob_uop_1_27_ftq_idx;
      5'b11100:
        casez_tmp_94 = rob_uop_1_28_ftq_idx;
      5'b11101:
        casez_tmp_94 = rob_uop_1_29_ftq_idx;
      5'b11110:
        casez_tmp_94 = rob_uop_1_30_ftq_idx;
      default:
        casez_tmp_94 = rob_uop_1_31_ftq_idx;
    endcase
  end // always @(*)
  reg         casez_tmp_95;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_95 = rob_uop_1_0_edge_inst;
      5'b00001:
        casez_tmp_95 = rob_uop_1_1_edge_inst;
      5'b00010:
        casez_tmp_95 = rob_uop_1_2_edge_inst;
      5'b00011:
        casez_tmp_95 = rob_uop_1_3_edge_inst;
      5'b00100:
        casez_tmp_95 = rob_uop_1_4_edge_inst;
      5'b00101:
        casez_tmp_95 = rob_uop_1_5_edge_inst;
      5'b00110:
        casez_tmp_95 = rob_uop_1_6_edge_inst;
      5'b00111:
        casez_tmp_95 = rob_uop_1_7_edge_inst;
      5'b01000:
        casez_tmp_95 = rob_uop_1_8_edge_inst;
      5'b01001:
        casez_tmp_95 = rob_uop_1_9_edge_inst;
      5'b01010:
        casez_tmp_95 = rob_uop_1_10_edge_inst;
      5'b01011:
        casez_tmp_95 = rob_uop_1_11_edge_inst;
      5'b01100:
        casez_tmp_95 = rob_uop_1_12_edge_inst;
      5'b01101:
        casez_tmp_95 = rob_uop_1_13_edge_inst;
      5'b01110:
        casez_tmp_95 = rob_uop_1_14_edge_inst;
      5'b01111:
        casez_tmp_95 = rob_uop_1_15_edge_inst;
      5'b10000:
        casez_tmp_95 = rob_uop_1_16_edge_inst;
      5'b10001:
        casez_tmp_95 = rob_uop_1_17_edge_inst;
      5'b10010:
        casez_tmp_95 = rob_uop_1_18_edge_inst;
      5'b10011:
        casez_tmp_95 = rob_uop_1_19_edge_inst;
      5'b10100:
        casez_tmp_95 = rob_uop_1_20_edge_inst;
      5'b10101:
        casez_tmp_95 = rob_uop_1_21_edge_inst;
      5'b10110:
        casez_tmp_95 = rob_uop_1_22_edge_inst;
      5'b10111:
        casez_tmp_95 = rob_uop_1_23_edge_inst;
      5'b11000:
        casez_tmp_95 = rob_uop_1_24_edge_inst;
      5'b11001:
        casez_tmp_95 = rob_uop_1_25_edge_inst;
      5'b11010:
        casez_tmp_95 = rob_uop_1_26_edge_inst;
      5'b11011:
        casez_tmp_95 = rob_uop_1_27_edge_inst;
      5'b11100:
        casez_tmp_95 = rob_uop_1_28_edge_inst;
      5'b11101:
        casez_tmp_95 = rob_uop_1_29_edge_inst;
      5'b11110:
        casez_tmp_95 = rob_uop_1_30_edge_inst;
      default:
        casez_tmp_95 = rob_uop_1_31_edge_inst;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_96;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_96 = rob_uop_1_0_pc_lob;
      5'b00001:
        casez_tmp_96 = rob_uop_1_1_pc_lob;
      5'b00010:
        casez_tmp_96 = rob_uop_1_2_pc_lob;
      5'b00011:
        casez_tmp_96 = rob_uop_1_3_pc_lob;
      5'b00100:
        casez_tmp_96 = rob_uop_1_4_pc_lob;
      5'b00101:
        casez_tmp_96 = rob_uop_1_5_pc_lob;
      5'b00110:
        casez_tmp_96 = rob_uop_1_6_pc_lob;
      5'b00111:
        casez_tmp_96 = rob_uop_1_7_pc_lob;
      5'b01000:
        casez_tmp_96 = rob_uop_1_8_pc_lob;
      5'b01001:
        casez_tmp_96 = rob_uop_1_9_pc_lob;
      5'b01010:
        casez_tmp_96 = rob_uop_1_10_pc_lob;
      5'b01011:
        casez_tmp_96 = rob_uop_1_11_pc_lob;
      5'b01100:
        casez_tmp_96 = rob_uop_1_12_pc_lob;
      5'b01101:
        casez_tmp_96 = rob_uop_1_13_pc_lob;
      5'b01110:
        casez_tmp_96 = rob_uop_1_14_pc_lob;
      5'b01111:
        casez_tmp_96 = rob_uop_1_15_pc_lob;
      5'b10000:
        casez_tmp_96 = rob_uop_1_16_pc_lob;
      5'b10001:
        casez_tmp_96 = rob_uop_1_17_pc_lob;
      5'b10010:
        casez_tmp_96 = rob_uop_1_18_pc_lob;
      5'b10011:
        casez_tmp_96 = rob_uop_1_19_pc_lob;
      5'b10100:
        casez_tmp_96 = rob_uop_1_20_pc_lob;
      5'b10101:
        casez_tmp_96 = rob_uop_1_21_pc_lob;
      5'b10110:
        casez_tmp_96 = rob_uop_1_22_pc_lob;
      5'b10111:
        casez_tmp_96 = rob_uop_1_23_pc_lob;
      5'b11000:
        casez_tmp_96 = rob_uop_1_24_pc_lob;
      5'b11001:
        casez_tmp_96 = rob_uop_1_25_pc_lob;
      5'b11010:
        casez_tmp_96 = rob_uop_1_26_pc_lob;
      5'b11011:
        casez_tmp_96 = rob_uop_1_27_pc_lob;
      5'b11100:
        casez_tmp_96 = rob_uop_1_28_pc_lob;
      5'b11101:
        casez_tmp_96 = rob_uop_1_29_pc_lob;
      5'b11110:
        casez_tmp_96 = rob_uop_1_30_pc_lob;
      default:
        casez_tmp_96 = rob_uop_1_31_pc_lob;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_97;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_97 = rob_uop_1_0_pdst;
      5'b00001:
        casez_tmp_97 = rob_uop_1_1_pdst;
      5'b00010:
        casez_tmp_97 = rob_uop_1_2_pdst;
      5'b00011:
        casez_tmp_97 = rob_uop_1_3_pdst;
      5'b00100:
        casez_tmp_97 = rob_uop_1_4_pdst;
      5'b00101:
        casez_tmp_97 = rob_uop_1_5_pdst;
      5'b00110:
        casez_tmp_97 = rob_uop_1_6_pdst;
      5'b00111:
        casez_tmp_97 = rob_uop_1_7_pdst;
      5'b01000:
        casez_tmp_97 = rob_uop_1_8_pdst;
      5'b01001:
        casez_tmp_97 = rob_uop_1_9_pdst;
      5'b01010:
        casez_tmp_97 = rob_uop_1_10_pdst;
      5'b01011:
        casez_tmp_97 = rob_uop_1_11_pdst;
      5'b01100:
        casez_tmp_97 = rob_uop_1_12_pdst;
      5'b01101:
        casez_tmp_97 = rob_uop_1_13_pdst;
      5'b01110:
        casez_tmp_97 = rob_uop_1_14_pdst;
      5'b01111:
        casez_tmp_97 = rob_uop_1_15_pdst;
      5'b10000:
        casez_tmp_97 = rob_uop_1_16_pdst;
      5'b10001:
        casez_tmp_97 = rob_uop_1_17_pdst;
      5'b10010:
        casez_tmp_97 = rob_uop_1_18_pdst;
      5'b10011:
        casez_tmp_97 = rob_uop_1_19_pdst;
      5'b10100:
        casez_tmp_97 = rob_uop_1_20_pdst;
      5'b10101:
        casez_tmp_97 = rob_uop_1_21_pdst;
      5'b10110:
        casez_tmp_97 = rob_uop_1_22_pdst;
      5'b10111:
        casez_tmp_97 = rob_uop_1_23_pdst;
      5'b11000:
        casez_tmp_97 = rob_uop_1_24_pdst;
      5'b11001:
        casez_tmp_97 = rob_uop_1_25_pdst;
      5'b11010:
        casez_tmp_97 = rob_uop_1_26_pdst;
      5'b11011:
        casez_tmp_97 = rob_uop_1_27_pdst;
      5'b11100:
        casez_tmp_97 = rob_uop_1_28_pdst;
      5'b11101:
        casez_tmp_97 = rob_uop_1_29_pdst;
      5'b11110:
        casez_tmp_97 = rob_uop_1_30_pdst;
      default:
        casez_tmp_97 = rob_uop_1_31_pdst;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_98;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_98 = rob_uop_1_0_stale_pdst;
      5'b00001:
        casez_tmp_98 = rob_uop_1_1_stale_pdst;
      5'b00010:
        casez_tmp_98 = rob_uop_1_2_stale_pdst;
      5'b00011:
        casez_tmp_98 = rob_uop_1_3_stale_pdst;
      5'b00100:
        casez_tmp_98 = rob_uop_1_4_stale_pdst;
      5'b00101:
        casez_tmp_98 = rob_uop_1_5_stale_pdst;
      5'b00110:
        casez_tmp_98 = rob_uop_1_6_stale_pdst;
      5'b00111:
        casez_tmp_98 = rob_uop_1_7_stale_pdst;
      5'b01000:
        casez_tmp_98 = rob_uop_1_8_stale_pdst;
      5'b01001:
        casez_tmp_98 = rob_uop_1_9_stale_pdst;
      5'b01010:
        casez_tmp_98 = rob_uop_1_10_stale_pdst;
      5'b01011:
        casez_tmp_98 = rob_uop_1_11_stale_pdst;
      5'b01100:
        casez_tmp_98 = rob_uop_1_12_stale_pdst;
      5'b01101:
        casez_tmp_98 = rob_uop_1_13_stale_pdst;
      5'b01110:
        casez_tmp_98 = rob_uop_1_14_stale_pdst;
      5'b01111:
        casez_tmp_98 = rob_uop_1_15_stale_pdst;
      5'b10000:
        casez_tmp_98 = rob_uop_1_16_stale_pdst;
      5'b10001:
        casez_tmp_98 = rob_uop_1_17_stale_pdst;
      5'b10010:
        casez_tmp_98 = rob_uop_1_18_stale_pdst;
      5'b10011:
        casez_tmp_98 = rob_uop_1_19_stale_pdst;
      5'b10100:
        casez_tmp_98 = rob_uop_1_20_stale_pdst;
      5'b10101:
        casez_tmp_98 = rob_uop_1_21_stale_pdst;
      5'b10110:
        casez_tmp_98 = rob_uop_1_22_stale_pdst;
      5'b10111:
        casez_tmp_98 = rob_uop_1_23_stale_pdst;
      5'b11000:
        casez_tmp_98 = rob_uop_1_24_stale_pdst;
      5'b11001:
        casez_tmp_98 = rob_uop_1_25_stale_pdst;
      5'b11010:
        casez_tmp_98 = rob_uop_1_26_stale_pdst;
      5'b11011:
        casez_tmp_98 = rob_uop_1_27_stale_pdst;
      5'b11100:
        casez_tmp_98 = rob_uop_1_28_stale_pdst;
      5'b11101:
        casez_tmp_98 = rob_uop_1_29_stale_pdst;
      5'b11110:
        casez_tmp_98 = rob_uop_1_30_stale_pdst;
      default:
        casez_tmp_98 = rob_uop_1_31_stale_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_99;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_99 = rob_uop_1_0_is_fencei;
      5'b00001:
        casez_tmp_99 = rob_uop_1_1_is_fencei;
      5'b00010:
        casez_tmp_99 = rob_uop_1_2_is_fencei;
      5'b00011:
        casez_tmp_99 = rob_uop_1_3_is_fencei;
      5'b00100:
        casez_tmp_99 = rob_uop_1_4_is_fencei;
      5'b00101:
        casez_tmp_99 = rob_uop_1_5_is_fencei;
      5'b00110:
        casez_tmp_99 = rob_uop_1_6_is_fencei;
      5'b00111:
        casez_tmp_99 = rob_uop_1_7_is_fencei;
      5'b01000:
        casez_tmp_99 = rob_uop_1_8_is_fencei;
      5'b01001:
        casez_tmp_99 = rob_uop_1_9_is_fencei;
      5'b01010:
        casez_tmp_99 = rob_uop_1_10_is_fencei;
      5'b01011:
        casez_tmp_99 = rob_uop_1_11_is_fencei;
      5'b01100:
        casez_tmp_99 = rob_uop_1_12_is_fencei;
      5'b01101:
        casez_tmp_99 = rob_uop_1_13_is_fencei;
      5'b01110:
        casez_tmp_99 = rob_uop_1_14_is_fencei;
      5'b01111:
        casez_tmp_99 = rob_uop_1_15_is_fencei;
      5'b10000:
        casez_tmp_99 = rob_uop_1_16_is_fencei;
      5'b10001:
        casez_tmp_99 = rob_uop_1_17_is_fencei;
      5'b10010:
        casez_tmp_99 = rob_uop_1_18_is_fencei;
      5'b10011:
        casez_tmp_99 = rob_uop_1_19_is_fencei;
      5'b10100:
        casez_tmp_99 = rob_uop_1_20_is_fencei;
      5'b10101:
        casez_tmp_99 = rob_uop_1_21_is_fencei;
      5'b10110:
        casez_tmp_99 = rob_uop_1_22_is_fencei;
      5'b10111:
        casez_tmp_99 = rob_uop_1_23_is_fencei;
      5'b11000:
        casez_tmp_99 = rob_uop_1_24_is_fencei;
      5'b11001:
        casez_tmp_99 = rob_uop_1_25_is_fencei;
      5'b11010:
        casez_tmp_99 = rob_uop_1_26_is_fencei;
      5'b11011:
        casez_tmp_99 = rob_uop_1_27_is_fencei;
      5'b11100:
        casez_tmp_99 = rob_uop_1_28_is_fencei;
      5'b11101:
        casez_tmp_99 = rob_uop_1_29_is_fencei;
      5'b11110:
        casez_tmp_99 = rob_uop_1_30_is_fencei;
      default:
        casez_tmp_99 = rob_uop_1_31_is_fencei;
    endcase
  end // always @(*)
  reg         casez_tmp_100;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_100 = rob_uop_1_0_uses_ldq;
      5'b00001:
        casez_tmp_100 = rob_uop_1_1_uses_ldq;
      5'b00010:
        casez_tmp_100 = rob_uop_1_2_uses_ldq;
      5'b00011:
        casez_tmp_100 = rob_uop_1_3_uses_ldq;
      5'b00100:
        casez_tmp_100 = rob_uop_1_4_uses_ldq;
      5'b00101:
        casez_tmp_100 = rob_uop_1_5_uses_ldq;
      5'b00110:
        casez_tmp_100 = rob_uop_1_6_uses_ldq;
      5'b00111:
        casez_tmp_100 = rob_uop_1_7_uses_ldq;
      5'b01000:
        casez_tmp_100 = rob_uop_1_8_uses_ldq;
      5'b01001:
        casez_tmp_100 = rob_uop_1_9_uses_ldq;
      5'b01010:
        casez_tmp_100 = rob_uop_1_10_uses_ldq;
      5'b01011:
        casez_tmp_100 = rob_uop_1_11_uses_ldq;
      5'b01100:
        casez_tmp_100 = rob_uop_1_12_uses_ldq;
      5'b01101:
        casez_tmp_100 = rob_uop_1_13_uses_ldq;
      5'b01110:
        casez_tmp_100 = rob_uop_1_14_uses_ldq;
      5'b01111:
        casez_tmp_100 = rob_uop_1_15_uses_ldq;
      5'b10000:
        casez_tmp_100 = rob_uop_1_16_uses_ldq;
      5'b10001:
        casez_tmp_100 = rob_uop_1_17_uses_ldq;
      5'b10010:
        casez_tmp_100 = rob_uop_1_18_uses_ldq;
      5'b10011:
        casez_tmp_100 = rob_uop_1_19_uses_ldq;
      5'b10100:
        casez_tmp_100 = rob_uop_1_20_uses_ldq;
      5'b10101:
        casez_tmp_100 = rob_uop_1_21_uses_ldq;
      5'b10110:
        casez_tmp_100 = rob_uop_1_22_uses_ldq;
      5'b10111:
        casez_tmp_100 = rob_uop_1_23_uses_ldq;
      5'b11000:
        casez_tmp_100 = rob_uop_1_24_uses_ldq;
      5'b11001:
        casez_tmp_100 = rob_uop_1_25_uses_ldq;
      5'b11010:
        casez_tmp_100 = rob_uop_1_26_uses_ldq;
      5'b11011:
        casez_tmp_100 = rob_uop_1_27_uses_ldq;
      5'b11100:
        casez_tmp_100 = rob_uop_1_28_uses_ldq;
      5'b11101:
        casez_tmp_100 = rob_uop_1_29_uses_ldq;
      5'b11110:
        casez_tmp_100 = rob_uop_1_30_uses_ldq;
      default:
        casez_tmp_100 = rob_uop_1_31_uses_ldq;
    endcase
  end // always @(*)
  reg         casez_tmp_101;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_101 = rob_uop_1_0_uses_stq;
      5'b00001:
        casez_tmp_101 = rob_uop_1_1_uses_stq;
      5'b00010:
        casez_tmp_101 = rob_uop_1_2_uses_stq;
      5'b00011:
        casez_tmp_101 = rob_uop_1_3_uses_stq;
      5'b00100:
        casez_tmp_101 = rob_uop_1_4_uses_stq;
      5'b00101:
        casez_tmp_101 = rob_uop_1_5_uses_stq;
      5'b00110:
        casez_tmp_101 = rob_uop_1_6_uses_stq;
      5'b00111:
        casez_tmp_101 = rob_uop_1_7_uses_stq;
      5'b01000:
        casez_tmp_101 = rob_uop_1_8_uses_stq;
      5'b01001:
        casez_tmp_101 = rob_uop_1_9_uses_stq;
      5'b01010:
        casez_tmp_101 = rob_uop_1_10_uses_stq;
      5'b01011:
        casez_tmp_101 = rob_uop_1_11_uses_stq;
      5'b01100:
        casez_tmp_101 = rob_uop_1_12_uses_stq;
      5'b01101:
        casez_tmp_101 = rob_uop_1_13_uses_stq;
      5'b01110:
        casez_tmp_101 = rob_uop_1_14_uses_stq;
      5'b01111:
        casez_tmp_101 = rob_uop_1_15_uses_stq;
      5'b10000:
        casez_tmp_101 = rob_uop_1_16_uses_stq;
      5'b10001:
        casez_tmp_101 = rob_uop_1_17_uses_stq;
      5'b10010:
        casez_tmp_101 = rob_uop_1_18_uses_stq;
      5'b10011:
        casez_tmp_101 = rob_uop_1_19_uses_stq;
      5'b10100:
        casez_tmp_101 = rob_uop_1_20_uses_stq;
      5'b10101:
        casez_tmp_101 = rob_uop_1_21_uses_stq;
      5'b10110:
        casez_tmp_101 = rob_uop_1_22_uses_stq;
      5'b10111:
        casez_tmp_101 = rob_uop_1_23_uses_stq;
      5'b11000:
        casez_tmp_101 = rob_uop_1_24_uses_stq;
      5'b11001:
        casez_tmp_101 = rob_uop_1_25_uses_stq;
      5'b11010:
        casez_tmp_101 = rob_uop_1_26_uses_stq;
      5'b11011:
        casez_tmp_101 = rob_uop_1_27_uses_stq;
      5'b11100:
        casez_tmp_101 = rob_uop_1_28_uses_stq;
      5'b11101:
        casez_tmp_101 = rob_uop_1_29_uses_stq;
      5'b11110:
        casez_tmp_101 = rob_uop_1_30_uses_stq;
      default:
        casez_tmp_101 = rob_uop_1_31_uses_stq;
    endcase
  end // always @(*)
  reg         casez_tmp_102;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_102 = rob_uop_1_0_is_sys_pc2epc;
      5'b00001:
        casez_tmp_102 = rob_uop_1_1_is_sys_pc2epc;
      5'b00010:
        casez_tmp_102 = rob_uop_1_2_is_sys_pc2epc;
      5'b00011:
        casez_tmp_102 = rob_uop_1_3_is_sys_pc2epc;
      5'b00100:
        casez_tmp_102 = rob_uop_1_4_is_sys_pc2epc;
      5'b00101:
        casez_tmp_102 = rob_uop_1_5_is_sys_pc2epc;
      5'b00110:
        casez_tmp_102 = rob_uop_1_6_is_sys_pc2epc;
      5'b00111:
        casez_tmp_102 = rob_uop_1_7_is_sys_pc2epc;
      5'b01000:
        casez_tmp_102 = rob_uop_1_8_is_sys_pc2epc;
      5'b01001:
        casez_tmp_102 = rob_uop_1_9_is_sys_pc2epc;
      5'b01010:
        casez_tmp_102 = rob_uop_1_10_is_sys_pc2epc;
      5'b01011:
        casez_tmp_102 = rob_uop_1_11_is_sys_pc2epc;
      5'b01100:
        casez_tmp_102 = rob_uop_1_12_is_sys_pc2epc;
      5'b01101:
        casez_tmp_102 = rob_uop_1_13_is_sys_pc2epc;
      5'b01110:
        casez_tmp_102 = rob_uop_1_14_is_sys_pc2epc;
      5'b01111:
        casez_tmp_102 = rob_uop_1_15_is_sys_pc2epc;
      5'b10000:
        casez_tmp_102 = rob_uop_1_16_is_sys_pc2epc;
      5'b10001:
        casez_tmp_102 = rob_uop_1_17_is_sys_pc2epc;
      5'b10010:
        casez_tmp_102 = rob_uop_1_18_is_sys_pc2epc;
      5'b10011:
        casez_tmp_102 = rob_uop_1_19_is_sys_pc2epc;
      5'b10100:
        casez_tmp_102 = rob_uop_1_20_is_sys_pc2epc;
      5'b10101:
        casez_tmp_102 = rob_uop_1_21_is_sys_pc2epc;
      5'b10110:
        casez_tmp_102 = rob_uop_1_22_is_sys_pc2epc;
      5'b10111:
        casez_tmp_102 = rob_uop_1_23_is_sys_pc2epc;
      5'b11000:
        casez_tmp_102 = rob_uop_1_24_is_sys_pc2epc;
      5'b11001:
        casez_tmp_102 = rob_uop_1_25_is_sys_pc2epc;
      5'b11010:
        casez_tmp_102 = rob_uop_1_26_is_sys_pc2epc;
      5'b11011:
        casez_tmp_102 = rob_uop_1_27_is_sys_pc2epc;
      5'b11100:
        casez_tmp_102 = rob_uop_1_28_is_sys_pc2epc;
      5'b11101:
        casez_tmp_102 = rob_uop_1_29_is_sys_pc2epc;
      5'b11110:
        casez_tmp_102 = rob_uop_1_30_is_sys_pc2epc;
      default:
        casez_tmp_102 = rob_uop_1_31_is_sys_pc2epc;
    endcase
  end // always @(*)
  reg         casez_tmp_103;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_103 = rob_uop_1_0_flush_on_commit;
      5'b00001:
        casez_tmp_103 = rob_uop_1_1_flush_on_commit;
      5'b00010:
        casez_tmp_103 = rob_uop_1_2_flush_on_commit;
      5'b00011:
        casez_tmp_103 = rob_uop_1_3_flush_on_commit;
      5'b00100:
        casez_tmp_103 = rob_uop_1_4_flush_on_commit;
      5'b00101:
        casez_tmp_103 = rob_uop_1_5_flush_on_commit;
      5'b00110:
        casez_tmp_103 = rob_uop_1_6_flush_on_commit;
      5'b00111:
        casez_tmp_103 = rob_uop_1_7_flush_on_commit;
      5'b01000:
        casez_tmp_103 = rob_uop_1_8_flush_on_commit;
      5'b01001:
        casez_tmp_103 = rob_uop_1_9_flush_on_commit;
      5'b01010:
        casez_tmp_103 = rob_uop_1_10_flush_on_commit;
      5'b01011:
        casez_tmp_103 = rob_uop_1_11_flush_on_commit;
      5'b01100:
        casez_tmp_103 = rob_uop_1_12_flush_on_commit;
      5'b01101:
        casez_tmp_103 = rob_uop_1_13_flush_on_commit;
      5'b01110:
        casez_tmp_103 = rob_uop_1_14_flush_on_commit;
      5'b01111:
        casez_tmp_103 = rob_uop_1_15_flush_on_commit;
      5'b10000:
        casez_tmp_103 = rob_uop_1_16_flush_on_commit;
      5'b10001:
        casez_tmp_103 = rob_uop_1_17_flush_on_commit;
      5'b10010:
        casez_tmp_103 = rob_uop_1_18_flush_on_commit;
      5'b10011:
        casez_tmp_103 = rob_uop_1_19_flush_on_commit;
      5'b10100:
        casez_tmp_103 = rob_uop_1_20_flush_on_commit;
      5'b10101:
        casez_tmp_103 = rob_uop_1_21_flush_on_commit;
      5'b10110:
        casez_tmp_103 = rob_uop_1_22_flush_on_commit;
      5'b10111:
        casez_tmp_103 = rob_uop_1_23_flush_on_commit;
      5'b11000:
        casez_tmp_103 = rob_uop_1_24_flush_on_commit;
      5'b11001:
        casez_tmp_103 = rob_uop_1_25_flush_on_commit;
      5'b11010:
        casez_tmp_103 = rob_uop_1_26_flush_on_commit;
      5'b11011:
        casez_tmp_103 = rob_uop_1_27_flush_on_commit;
      5'b11100:
        casez_tmp_103 = rob_uop_1_28_flush_on_commit;
      5'b11101:
        casez_tmp_103 = rob_uop_1_29_flush_on_commit;
      5'b11110:
        casez_tmp_103 = rob_uop_1_30_flush_on_commit;
      default:
        casez_tmp_103 = rob_uop_1_31_flush_on_commit;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_104;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_104 = rob_uop_1_0_ldst;
      5'b00001:
        casez_tmp_104 = rob_uop_1_1_ldst;
      5'b00010:
        casez_tmp_104 = rob_uop_1_2_ldst;
      5'b00011:
        casez_tmp_104 = rob_uop_1_3_ldst;
      5'b00100:
        casez_tmp_104 = rob_uop_1_4_ldst;
      5'b00101:
        casez_tmp_104 = rob_uop_1_5_ldst;
      5'b00110:
        casez_tmp_104 = rob_uop_1_6_ldst;
      5'b00111:
        casez_tmp_104 = rob_uop_1_7_ldst;
      5'b01000:
        casez_tmp_104 = rob_uop_1_8_ldst;
      5'b01001:
        casez_tmp_104 = rob_uop_1_9_ldst;
      5'b01010:
        casez_tmp_104 = rob_uop_1_10_ldst;
      5'b01011:
        casez_tmp_104 = rob_uop_1_11_ldst;
      5'b01100:
        casez_tmp_104 = rob_uop_1_12_ldst;
      5'b01101:
        casez_tmp_104 = rob_uop_1_13_ldst;
      5'b01110:
        casez_tmp_104 = rob_uop_1_14_ldst;
      5'b01111:
        casez_tmp_104 = rob_uop_1_15_ldst;
      5'b10000:
        casez_tmp_104 = rob_uop_1_16_ldst;
      5'b10001:
        casez_tmp_104 = rob_uop_1_17_ldst;
      5'b10010:
        casez_tmp_104 = rob_uop_1_18_ldst;
      5'b10011:
        casez_tmp_104 = rob_uop_1_19_ldst;
      5'b10100:
        casez_tmp_104 = rob_uop_1_20_ldst;
      5'b10101:
        casez_tmp_104 = rob_uop_1_21_ldst;
      5'b10110:
        casez_tmp_104 = rob_uop_1_22_ldst;
      5'b10111:
        casez_tmp_104 = rob_uop_1_23_ldst;
      5'b11000:
        casez_tmp_104 = rob_uop_1_24_ldst;
      5'b11001:
        casez_tmp_104 = rob_uop_1_25_ldst;
      5'b11010:
        casez_tmp_104 = rob_uop_1_26_ldst;
      5'b11011:
        casez_tmp_104 = rob_uop_1_27_ldst;
      5'b11100:
        casez_tmp_104 = rob_uop_1_28_ldst;
      5'b11101:
        casez_tmp_104 = rob_uop_1_29_ldst;
      5'b11110:
        casez_tmp_104 = rob_uop_1_30_ldst;
      default:
        casez_tmp_104 = rob_uop_1_31_ldst;
    endcase
  end // always @(*)
  reg         casez_tmp_105;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_105 = rob_uop_1_0_ldst_val;
      5'b00001:
        casez_tmp_105 = rob_uop_1_1_ldst_val;
      5'b00010:
        casez_tmp_105 = rob_uop_1_2_ldst_val;
      5'b00011:
        casez_tmp_105 = rob_uop_1_3_ldst_val;
      5'b00100:
        casez_tmp_105 = rob_uop_1_4_ldst_val;
      5'b00101:
        casez_tmp_105 = rob_uop_1_5_ldst_val;
      5'b00110:
        casez_tmp_105 = rob_uop_1_6_ldst_val;
      5'b00111:
        casez_tmp_105 = rob_uop_1_7_ldst_val;
      5'b01000:
        casez_tmp_105 = rob_uop_1_8_ldst_val;
      5'b01001:
        casez_tmp_105 = rob_uop_1_9_ldst_val;
      5'b01010:
        casez_tmp_105 = rob_uop_1_10_ldst_val;
      5'b01011:
        casez_tmp_105 = rob_uop_1_11_ldst_val;
      5'b01100:
        casez_tmp_105 = rob_uop_1_12_ldst_val;
      5'b01101:
        casez_tmp_105 = rob_uop_1_13_ldst_val;
      5'b01110:
        casez_tmp_105 = rob_uop_1_14_ldst_val;
      5'b01111:
        casez_tmp_105 = rob_uop_1_15_ldst_val;
      5'b10000:
        casez_tmp_105 = rob_uop_1_16_ldst_val;
      5'b10001:
        casez_tmp_105 = rob_uop_1_17_ldst_val;
      5'b10010:
        casez_tmp_105 = rob_uop_1_18_ldst_val;
      5'b10011:
        casez_tmp_105 = rob_uop_1_19_ldst_val;
      5'b10100:
        casez_tmp_105 = rob_uop_1_20_ldst_val;
      5'b10101:
        casez_tmp_105 = rob_uop_1_21_ldst_val;
      5'b10110:
        casez_tmp_105 = rob_uop_1_22_ldst_val;
      5'b10111:
        casez_tmp_105 = rob_uop_1_23_ldst_val;
      5'b11000:
        casez_tmp_105 = rob_uop_1_24_ldst_val;
      5'b11001:
        casez_tmp_105 = rob_uop_1_25_ldst_val;
      5'b11010:
        casez_tmp_105 = rob_uop_1_26_ldst_val;
      5'b11011:
        casez_tmp_105 = rob_uop_1_27_ldst_val;
      5'b11100:
        casez_tmp_105 = rob_uop_1_28_ldst_val;
      5'b11101:
        casez_tmp_105 = rob_uop_1_29_ldst_val;
      5'b11110:
        casez_tmp_105 = rob_uop_1_30_ldst_val;
      default:
        casez_tmp_105 = rob_uop_1_31_ldst_val;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_106;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_106 = rob_uop_1_0_dst_rtype;
      5'b00001:
        casez_tmp_106 = rob_uop_1_1_dst_rtype;
      5'b00010:
        casez_tmp_106 = rob_uop_1_2_dst_rtype;
      5'b00011:
        casez_tmp_106 = rob_uop_1_3_dst_rtype;
      5'b00100:
        casez_tmp_106 = rob_uop_1_4_dst_rtype;
      5'b00101:
        casez_tmp_106 = rob_uop_1_5_dst_rtype;
      5'b00110:
        casez_tmp_106 = rob_uop_1_6_dst_rtype;
      5'b00111:
        casez_tmp_106 = rob_uop_1_7_dst_rtype;
      5'b01000:
        casez_tmp_106 = rob_uop_1_8_dst_rtype;
      5'b01001:
        casez_tmp_106 = rob_uop_1_9_dst_rtype;
      5'b01010:
        casez_tmp_106 = rob_uop_1_10_dst_rtype;
      5'b01011:
        casez_tmp_106 = rob_uop_1_11_dst_rtype;
      5'b01100:
        casez_tmp_106 = rob_uop_1_12_dst_rtype;
      5'b01101:
        casez_tmp_106 = rob_uop_1_13_dst_rtype;
      5'b01110:
        casez_tmp_106 = rob_uop_1_14_dst_rtype;
      5'b01111:
        casez_tmp_106 = rob_uop_1_15_dst_rtype;
      5'b10000:
        casez_tmp_106 = rob_uop_1_16_dst_rtype;
      5'b10001:
        casez_tmp_106 = rob_uop_1_17_dst_rtype;
      5'b10010:
        casez_tmp_106 = rob_uop_1_18_dst_rtype;
      5'b10011:
        casez_tmp_106 = rob_uop_1_19_dst_rtype;
      5'b10100:
        casez_tmp_106 = rob_uop_1_20_dst_rtype;
      5'b10101:
        casez_tmp_106 = rob_uop_1_21_dst_rtype;
      5'b10110:
        casez_tmp_106 = rob_uop_1_22_dst_rtype;
      5'b10111:
        casez_tmp_106 = rob_uop_1_23_dst_rtype;
      5'b11000:
        casez_tmp_106 = rob_uop_1_24_dst_rtype;
      5'b11001:
        casez_tmp_106 = rob_uop_1_25_dst_rtype;
      5'b11010:
        casez_tmp_106 = rob_uop_1_26_dst_rtype;
      5'b11011:
        casez_tmp_106 = rob_uop_1_27_dst_rtype;
      5'b11100:
        casez_tmp_106 = rob_uop_1_28_dst_rtype;
      5'b11101:
        casez_tmp_106 = rob_uop_1_29_dst_rtype;
      5'b11110:
        casez_tmp_106 = rob_uop_1_30_dst_rtype;
      default:
        casez_tmp_106 = rob_uop_1_31_dst_rtype;
    endcase
  end // always @(*)
  reg         casez_tmp_107;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_107 = rob_uop_1_0_fp_val;
      5'b00001:
        casez_tmp_107 = rob_uop_1_1_fp_val;
      5'b00010:
        casez_tmp_107 = rob_uop_1_2_fp_val;
      5'b00011:
        casez_tmp_107 = rob_uop_1_3_fp_val;
      5'b00100:
        casez_tmp_107 = rob_uop_1_4_fp_val;
      5'b00101:
        casez_tmp_107 = rob_uop_1_5_fp_val;
      5'b00110:
        casez_tmp_107 = rob_uop_1_6_fp_val;
      5'b00111:
        casez_tmp_107 = rob_uop_1_7_fp_val;
      5'b01000:
        casez_tmp_107 = rob_uop_1_8_fp_val;
      5'b01001:
        casez_tmp_107 = rob_uop_1_9_fp_val;
      5'b01010:
        casez_tmp_107 = rob_uop_1_10_fp_val;
      5'b01011:
        casez_tmp_107 = rob_uop_1_11_fp_val;
      5'b01100:
        casez_tmp_107 = rob_uop_1_12_fp_val;
      5'b01101:
        casez_tmp_107 = rob_uop_1_13_fp_val;
      5'b01110:
        casez_tmp_107 = rob_uop_1_14_fp_val;
      5'b01111:
        casez_tmp_107 = rob_uop_1_15_fp_val;
      5'b10000:
        casez_tmp_107 = rob_uop_1_16_fp_val;
      5'b10001:
        casez_tmp_107 = rob_uop_1_17_fp_val;
      5'b10010:
        casez_tmp_107 = rob_uop_1_18_fp_val;
      5'b10011:
        casez_tmp_107 = rob_uop_1_19_fp_val;
      5'b10100:
        casez_tmp_107 = rob_uop_1_20_fp_val;
      5'b10101:
        casez_tmp_107 = rob_uop_1_21_fp_val;
      5'b10110:
        casez_tmp_107 = rob_uop_1_22_fp_val;
      5'b10111:
        casez_tmp_107 = rob_uop_1_23_fp_val;
      5'b11000:
        casez_tmp_107 = rob_uop_1_24_fp_val;
      5'b11001:
        casez_tmp_107 = rob_uop_1_25_fp_val;
      5'b11010:
        casez_tmp_107 = rob_uop_1_26_fp_val;
      5'b11011:
        casez_tmp_107 = rob_uop_1_27_fp_val;
      5'b11100:
        casez_tmp_107 = rob_uop_1_28_fp_val;
      5'b11101:
        casez_tmp_107 = rob_uop_1_29_fp_val;
      5'b11110:
        casez_tmp_107 = rob_uop_1_30_fp_val;
      default:
        casez_tmp_107 = rob_uop_1_31_fp_val;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_108;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_108 = rob_uop_1_0_debug_fsrc;
      5'b00001:
        casez_tmp_108 = rob_uop_1_1_debug_fsrc;
      5'b00010:
        casez_tmp_108 = rob_uop_1_2_debug_fsrc;
      5'b00011:
        casez_tmp_108 = rob_uop_1_3_debug_fsrc;
      5'b00100:
        casez_tmp_108 = rob_uop_1_4_debug_fsrc;
      5'b00101:
        casez_tmp_108 = rob_uop_1_5_debug_fsrc;
      5'b00110:
        casez_tmp_108 = rob_uop_1_6_debug_fsrc;
      5'b00111:
        casez_tmp_108 = rob_uop_1_7_debug_fsrc;
      5'b01000:
        casez_tmp_108 = rob_uop_1_8_debug_fsrc;
      5'b01001:
        casez_tmp_108 = rob_uop_1_9_debug_fsrc;
      5'b01010:
        casez_tmp_108 = rob_uop_1_10_debug_fsrc;
      5'b01011:
        casez_tmp_108 = rob_uop_1_11_debug_fsrc;
      5'b01100:
        casez_tmp_108 = rob_uop_1_12_debug_fsrc;
      5'b01101:
        casez_tmp_108 = rob_uop_1_13_debug_fsrc;
      5'b01110:
        casez_tmp_108 = rob_uop_1_14_debug_fsrc;
      5'b01111:
        casez_tmp_108 = rob_uop_1_15_debug_fsrc;
      5'b10000:
        casez_tmp_108 = rob_uop_1_16_debug_fsrc;
      5'b10001:
        casez_tmp_108 = rob_uop_1_17_debug_fsrc;
      5'b10010:
        casez_tmp_108 = rob_uop_1_18_debug_fsrc;
      5'b10011:
        casez_tmp_108 = rob_uop_1_19_debug_fsrc;
      5'b10100:
        casez_tmp_108 = rob_uop_1_20_debug_fsrc;
      5'b10101:
        casez_tmp_108 = rob_uop_1_21_debug_fsrc;
      5'b10110:
        casez_tmp_108 = rob_uop_1_22_debug_fsrc;
      5'b10111:
        casez_tmp_108 = rob_uop_1_23_debug_fsrc;
      5'b11000:
        casez_tmp_108 = rob_uop_1_24_debug_fsrc;
      5'b11001:
        casez_tmp_108 = rob_uop_1_25_debug_fsrc;
      5'b11010:
        casez_tmp_108 = rob_uop_1_26_debug_fsrc;
      5'b11011:
        casez_tmp_108 = rob_uop_1_27_debug_fsrc;
      5'b11100:
        casez_tmp_108 = rob_uop_1_28_debug_fsrc;
      5'b11101:
        casez_tmp_108 = rob_uop_1_29_debug_fsrc;
      5'b11110:
        casez_tmp_108 = rob_uop_1_30_debug_fsrc;
      default:
        casez_tmp_108 = rob_uop_1_31_debug_fsrc;
    endcase
  end // always @(*)
  wire        _GEN_32 = io_brupdate_b2_mispredict & io_brupdate_b2_uop_rob_idx[1:0] == 2'h1;
  wire        rbk_row_1 = _io_commit_rollback_T_3 & ~full;
  reg         casez_tmp_109;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_109 = rob_val_1_0;
      5'b00001:
        casez_tmp_109 = rob_val_1_1;
      5'b00010:
        casez_tmp_109 = rob_val_1_2;
      5'b00011:
        casez_tmp_109 = rob_val_1_3;
      5'b00100:
        casez_tmp_109 = rob_val_1_4;
      5'b00101:
        casez_tmp_109 = rob_val_1_5;
      5'b00110:
        casez_tmp_109 = rob_val_1_6;
      5'b00111:
        casez_tmp_109 = rob_val_1_7;
      5'b01000:
        casez_tmp_109 = rob_val_1_8;
      5'b01001:
        casez_tmp_109 = rob_val_1_9;
      5'b01010:
        casez_tmp_109 = rob_val_1_10;
      5'b01011:
        casez_tmp_109 = rob_val_1_11;
      5'b01100:
        casez_tmp_109 = rob_val_1_12;
      5'b01101:
        casez_tmp_109 = rob_val_1_13;
      5'b01110:
        casez_tmp_109 = rob_val_1_14;
      5'b01111:
        casez_tmp_109 = rob_val_1_15;
      5'b10000:
        casez_tmp_109 = rob_val_1_16;
      5'b10001:
        casez_tmp_109 = rob_val_1_17;
      5'b10010:
        casez_tmp_109 = rob_val_1_18;
      5'b10011:
        casez_tmp_109 = rob_val_1_19;
      5'b10100:
        casez_tmp_109 = rob_val_1_20;
      5'b10101:
        casez_tmp_109 = rob_val_1_21;
      5'b10110:
        casez_tmp_109 = rob_val_1_22;
      5'b10111:
        casez_tmp_109 = rob_val_1_23;
      5'b11000:
        casez_tmp_109 = rob_val_1_24;
      5'b11001:
        casez_tmp_109 = rob_val_1_25;
      5'b11010:
        casez_tmp_109 = rob_val_1_26;
      5'b11011:
        casez_tmp_109 = rob_val_1_27;
      5'b11100:
        casez_tmp_109 = rob_val_1_28;
      5'b11101:
        casez_tmp_109 = rob_val_1_29;
      5'b11110:
        casez_tmp_109 = rob_val_1_30;
      default:
        casez_tmp_109 = rob_val_1_31;
    endcase
  end // always @(*)
  wire        _io_commit_rbk_valids_1_output = rbk_row_1 & casez_tmp_109;
  reg  [4:0]  casez_tmp_110;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_110 = rob_fflags_1_0;
      5'b00001:
        casez_tmp_110 = rob_fflags_1_1;
      5'b00010:
        casez_tmp_110 = rob_fflags_1_2;
      5'b00011:
        casez_tmp_110 = rob_fflags_1_3;
      5'b00100:
        casez_tmp_110 = rob_fflags_1_4;
      5'b00101:
        casez_tmp_110 = rob_fflags_1_5;
      5'b00110:
        casez_tmp_110 = rob_fflags_1_6;
      5'b00111:
        casez_tmp_110 = rob_fflags_1_7;
      5'b01000:
        casez_tmp_110 = rob_fflags_1_8;
      5'b01001:
        casez_tmp_110 = rob_fflags_1_9;
      5'b01010:
        casez_tmp_110 = rob_fflags_1_10;
      5'b01011:
        casez_tmp_110 = rob_fflags_1_11;
      5'b01100:
        casez_tmp_110 = rob_fflags_1_12;
      5'b01101:
        casez_tmp_110 = rob_fflags_1_13;
      5'b01110:
        casez_tmp_110 = rob_fflags_1_14;
      5'b01111:
        casez_tmp_110 = rob_fflags_1_15;
      5'b10000:
        casez_tmp_110 = rob_fflags_1_16;
      5'b10001:
        casez_tmp_110 = rob_fflags_1_17;
      5'b10010:
        casez_tmp_110 = rob_fflags_1_18;
      5'b10011:
        casez_tmp_110 = rob_fflags_1_19;
      5'b10100:
        casez_tmp_110 = rob_fflags_1_20;
      5'b10101:
        casez_tmp_110 = rob_fflags_1_21;
      5'b10110:
        casez_tmp_110 = rob_fflags_1_22;
      5'b10111:
        casez_tmp_110 = rob_fflags_1_23;
      5'b11000:
        casez_tmp_110 = rob_fflags_1_24;
      5'b11001:
        casez_tmp_110 = rob_fflags_1_25;
      5'b11010:
        casez_tmp_110 = rob_fflags_1_26;
      5'b11011:
        casez_tmp_110 = rob_fflags_1_27;
      5'b11100:
        casez_tmp_110 = rob_fflags_1_28;
      5'b11101:
        casez_tmp_110 = rob_fflags_1_29;
      5'b11110:
        casez_tmp_110 = rob_fflags_1_30;
      default:
        casez_tmp_110 = rob_fflags_1_31;
    endcase
  end // always @(*)
  reg         casez_tmp_111;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_111 = rob_uop_1_0_uses_ldq;
      5'b00001:
        casez_tmp_111 = rob_uop_1_1_uses_ldq;
      5'b00010:
        casez_tmp_111 = rob_uop_1_2_uses_ldq;
      5'b00011:
        casez_tmp_111 = rob_uop_1_3_uses_ldq;
      5'b00100:
        casez_tmp_111 = rob_uop_1_4_uses_ldq;
      5'b00101:
        casez_tmp_111 = rob_uop_1_5_uses_ldq;
      5'b00110:
        casez_tmp_111 = rob_uop_1_6_uses_ldq;
      5'b00111:
        casez_tmp_111 = rob_uop_1_7_uses_ldq;
      5'b01000:
        casez_tmp_111 = rob_uop_1_8_uses_ldq;
      5'b01001:
        casez_tmp_111 = rob_uop_1_9_uses_ldq;
      5'b01010:
        casez_tmp_111 = rob_uop_1_10_uses_ldq;
      5'b01011:
        casez_tmp_111 = rob_uop_1_11_uses_ldq;
      5'b01100:
        casez_tmp_111 = rob_uop_1_12_uses_ldq;
      5'b01101:
        casez_tmp_111 = rob_uop_1_13_uses_ldq;
      5'b01110:
        casez_tmp_111 = rob_uop_1_14_uses_ldq;
      5'b01111:
        casez_tmp_111 = rob_uop_1_15_uses_ldq;
      5'b10000:
        casez_tmp_111 = rob_uop_1_16_uses_ldq;
      5'b10001:
        casez_tmp_111 = rob_uop_1_17_uses_ldq;
      5'b10010:
        casez_tmp_111 = rob_uop_1_18_uses_ldq;
      5'b10011:
        casez_tmp_111 = rob_uop_1_19_uses_ldq;
      5'b10100:
        casez_tmp_111 = rob_uop_1_20_uses_ldq;
      5'b10101:
        casez_tmp_111 = rob_uop_1_21_uses_ldq;
      5'b10110:
        casez_tmp_111 = rob_uop_1_22_uses_ldq;
      5'b10111:
        casez_tmp_111 = rob_uop_1_23_uses_ldq;
      5'b11000:
        casez_tmp_111 = rob_uop_1_24_uses_ldq;
      5'b11001:
        casez_tmp_111 = rob_uop_1_25_uses_ldq;
      5'b11010:
        casez_tmp_111 = rob_uop_1_26_uses_ldq;
      5'b11011:
        casez_tmp_111 = rob_uop_1_27_uses_ldq;
      5'b11100:
        casez_tmp_111 = rob_uop_1_28_uses_ldq;
      5'b11101:
        casez_tmp_111 = rob_uop_1_29_uses_ldq;
      5'b11110:
        casez_tmp_111 = rob_uop_1_30_uses_ldq;
      default:
        casez_tmp_111 = rob_uop_1_31_uses_ldq;
    endcase
  end // always @(*)
  reg         casez_tmp_112;
  always @(*) begin
    casez (rob_pnr)
      5'b00000:
        casez_tmp_112 = rob_unsafe_1_0;
      5'b00001:
        casez_tmp_112 = rob_unsafe_1_1;
      5'b00010:
        casez_tmp_112 = rob_unsafe_1_2;
      5'b00011:
        casez_tmp_112 = rob_unsafe_1_3;
      5'b00100:
        casez_tmp_112 = rob_unsafe_1_4;
      5'b00101:
        casez_tmp_112 = rob_unsafe_1_5;
      5'b00110:
        casez_tmp_112 = rob_unsafe_1_6;
      5'b00111:
        casez_tmp_112 = rob_unsafe_1_7;
      5'b01000:
        casez_tmp_112 = rob_unsafe_1_8;
      5'b01001:
        casez_tmp_112 = rob_unsafe_1_9;
      5'b01010:
        casez_tmp_112 = rob_unsafe_1_10;
      5'b01011:
        casez_tmp_112 = rob_unsafe_1_11;
      5'b01100:
        casez_tmp_112 = rob_unsafe_1_12;
      5'b01101:
        casez_tmp_112 = rob_unsafe_1_13;
      5'b01110:
        casez_tmp_112 = rob_unsafe_1_14;
      5'b01111:
        casez_tmp_112 = rob_unsafe_1_15;
      5'b10000:
        casez_tmp_112 = rob_unsafe_1_16;
      5'b10001:
        casez_tmp_112 = rob_unsafe_1_17;
      5'b10010:
        casez_tmp_112 = rob_unsafe_1_18;
      5'b10011:
        casez_tmp_112 = rob_unsafe_1_19;
      5'b10100:
        casez_tmp_112 = rob_unsafe_1_20;
      5'b10101:
        casez_tmp_112 = rob_unsafe_1_21;
      5'b10110:
        casez_tmp_112 = rob_unsafe_1_22;
      5'b10111:
        casez_tmp_112 = rob_unsafe_1_23;
      5'b11000:
        casez_tmp_112 = rob_unsafe_1_24;
      5'b11001:
        casez_tmp_112 = rob_unsafe_1_25;
      5'b11010:
        casez_tmp_112 = rob_unsafe_1_26;
      5'b11011:
        casez_tmp_112 = rob_unsafe_1_27;
      5'b11100:
        casez_tmp_112 = rob_unsafe_1_28;
      5'b11101:
        casez_tmp_112 = rob_unsafe_1_29;
      5'b11110:
        casez_tmp_112 = rob_unsafe_1_30;
      default:
        casez_tmp_112 = rob_unsafe_1_31;
    endcase
  end // always @(*)
  reg         casez_tmp_113;
  always @(*) begin
    casez (rob_pnr)
      5'b00000:
        casez_tmp_113 = rob_exception_1_0;
      5'b00001:
        casez_tmp_113 = rob_exception_1_1;
      5'b00010:
        casez_tmp_113 = rob_exception_1_2;
      5'b00011:
        casez_tmp_113 = rob_exception_1_3;
      5'b00100:
        casez_tmp_113 = rob_exception_1_4;
      5'b00101:
        casez_tmp_113 = rob_exception_1_5;
      5'b00110:
        casez_tmp_113 = rob_exception_1_6;
      5'b00111:
        casez_tmp_113 = rob_exception_1_7;
      5'b01000:
        casez_tmp_113 = rob_exception_1_8;
      5'b01001:
        casez_tmp_113 = rob_exception_1_9;
      5'b01010:
        casez_tmp_113 = rob_exception_1_10;
      5'b01011:
        casez_tmp_113 = rob_exception_1_11;
      5'b01100:
        casez_tmp_113 = rob_exception_1_12;
      5'b01101:
        casez_tmp_113 = rob_exception_1_13;
      5'b01110:
        casez_tmp_113 = rob_exception_1_14;
      5'b01111:
        casez_tmp_113 = rob_exception_1_15;
      5'b10000:
        casez_tmp_113 = rob_exception_1_16;
      5'b10001:
        casez_tmp_113 = rob_exception_1_17;
      5'b10010:
        casez_tmp_113 = rob_exception_1_18;
      5'b10011:
        casez_tmp_113 = rob_exception_1_19;
      5'b10100:
        casez_tmp_113 = rob_exception_1_20;
      5'b10101:
        casez_tmp_113 = rob_exception_1_21;
      5'b10110:
        casez_tmp_113 = rob_exception_1_22;
      5'b10111:
        casez_tmp_113 = rob_exception_1_23;
      5'b11000:
        casez_tmp_113 = rob_exception_1_24;
      5'b11001:
        casez_tmp_113 = rob_exception_1_25;
      5'b11010:
        casez_tmp_113 = rob_exception_1_26;
      5'b11011:
        casez_tmp_113 = rob_exception_1_27;
      5'b11100:
        casez_tmp_113 = rob_exception_1_28;
      5'b11101:
        casez_tmp_113 = rob_exception_1_29;
      5'b11110:
        casez_tmp_113 = rob_exception_1_30;
      default:
        casez_tmp_113 = rob_exception_1_31;
    endcase
  end // always @(*)
  reg         casez_tmp_114;
  always @(*) begin
    casez (rob_pnr)
      5'b00000:
        casez_tmp_114 = rob_val_1_0;
      5'b00001:
        casez_tmp_114 = rob_val_1_1;
      5'b00010:
        casez_tmp_114 = rob_val_1_2;
      5'b00011:
        casez_tmp_114 = rob_val_1_3;
      5'b00100:
        casez_tmp_114 = rob_val_1_4;
      5'b00101:
        casez_tmp_114 = rob_val_1_5;
      5'b00110:
        casez_tmp_114 = rob_val_1_6;
      5'b00111:
        casez_tmp_114 = rob_val_1_7;
      5'b01000:
        casez_tmp_114 = rob_val_1_8;
      5'b01001:
        casez_tmp_114 = rob_val_1_9;
      5'b01010:
        casez_tmp_114 = rob_val_1_10;
      5'b01011:
        casez_tmp_114 = rob_val_1_11;
      5'b01100:
        casez_tmp_114 = rob_val_1_12;
      5'b01101:
        casez_tmp_114 = rob_val_1_13;
      5'b01110:
        casez_tmp_114 = rob_val_1_14;
      5'b01111:
        casez_tmp_114 = rob_val_1_15;
      5'b10000:
        casez_tmp_114 = rob_val_1_16;
      5'b10001:
        casez_tmp_114 = rob_val_1_17;
      5'b10010:
        casez_tmp_114 = rob_val_1_18;
      5'b10011:
        casez_tmp_114 = rob_val_1_19;
      5'b10100:
        casez_tmp_114 = rob_val_1_20;
      5'b10101:
        casez_tmp_114 = rob_val_1_21;
      5'b10110:
        casez_tmp_114 = rob_val_1_22;
      5'b10111:
        casez_tmp_114 = rob_val_1_23;
      5'b11000:
        casez_tmp_114 = rob_val_1_24;
      5'b11001:
        casez_tmp_114 = rob_val_1_25;
      5'b11010:
        casez_tmp_114 = rob_val_1_26;
      5'b11011:
        casez_tmp_114 = rob_val_1_27;
      5'b11100:
        casez_tmp_114 = rob_val_1_28;
      5'b11101:
        casez_tmp_114 = rob_val_1_29;
      5'b11110:
        casez_tmp_114 = rob_val_1_30;
      default:
        casez_tmp_114 = rob_val_1_31;
    endcase
  end // always @(*)
  reg         casez_tmp_115;
  always @(*) begin
    casez (io_wb_resps_0_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_115 = rob_val_1_0;
      5'b00001:
        casez_tmp_115 = rob_val_1_1;
      5'b00010:
        casez_tmp_115 = rob_val_1_2;
      5'b00011:
        casez_tmp_115 = rob_val_1_3;
      5'b00100:
        casez_tmp_115 = rob_val_1_4;
      5'b00101:
        casez_tmp_115 = rob_val_1_5;
      5'b00110:
        casez_tmp_115 = rob_val_1_6;
      5'b00111:
        casez_tmp_115 = rob_val_1_7;
      5'b01000:
        casez_tmp_115 = rob_val_1_8;
      5'b01001:
        casez_tmp_115 = rob_val_1_9;
      5'b01010:
        casez_tmp_115 = rob_val_1_10;
      5'b01011:
        casez_tmp_115 = rob_val_1_11;
      5'b01100:
        casez_tmp_115 = rob_val_1_12;
      5'b01101:
        casez_tmp_115 = rob_val_1_13;
      5'b01110:
        casez_tmp_115 = rob_val_1_14;
      5'b01111:
        casez_tmp_115 = rob_val_1_15;
      5'b10000:
        casez_tmp_115 = rob_val_1_16;
      5'b10001:
        casez_tmp_115 = rob_val_1_17;
      5'b10010:
        casez_tmp_115 = rob_val_1_18;
      5'b10011:
        casez_tmp_115 = rob_val_1_19;
      5'b10100:
        casez_tmp_115 = rob_val_1_20;
      5'b10101:
        casez_tmp_115 = rob_val_1_21;
      5'b10110:
        casez_tmp_115 = rob_val_1_22;
      5'b10111:
        casez_tmp_115 = rob_val_1_23;
      5'b11000:
        casez_tmp_115 = rob_val_1_24;
      5'b11001:
        casez_tmp_115 = rob_val_1_25;
      5'b11010:
        casez_tmp_115 = rob_val_1_26;
      5'b11011:
        casez_tmp_115 = rob_val_1_27;
      5'b11100:
        casez_tmp_115 = rob_val_1_28;
      5'b11101:
        casez_tmp_115 = rob_val_1_29;
      5'b11110:
        casez_tmp_115 = rob_val_1_30;
      default:
        casez_tmp_115 = rob_val_1_31;
    endcase
  end // always @(*)
  reg         casez_tmp_116;
  always @(*) begin
    casez (io_wb_resps_0_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_116 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_116 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_116 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_116 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_116 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_116 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_116 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_116 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_116 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_116 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_116 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_116 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_116 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_116 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_116 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_116 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_116 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_116 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_116 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_116 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_116 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_116 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_116 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_116 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_116 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_116 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_116 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_116 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_116 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_116 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_116 = rob_bsy_1_30;
      default:
        casez_tmp_116 = rob_bsy_1_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_117;
  always @(*) begin
    casez (io_wb_resps_0_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_117 = rob_uop_1_0_pdst;
      5'b00001:
        casez_tmp_117 = rob_uop_1_1_pdst;
      5'b00010:
        casez_tmp_117 = rob_uop_1_2_pdst;
      5'b00011:
        casez_tmp_117 = rob_uop_1_3_pdst;
      5'b00100:
        casez_tmp_117 = rob_uop_1_4_pdst;
      5'b00101:
        casez_tmp_117 = rob_uop_1_5_pdst;
      5'b00110:
        casez_tmp_117 = rob_uop_1_6_pdst;
      5'b00111:
        casez_tmp_117 = rob_uop_1_7_pdst;
      5'b01000:
        casez_tmp_117 = rob_uop_1_8_pdst;
      5'b01001:
        casez_tmp_117 = rob_uop_1_9_pdst;
      5'b01010:
        casez_tmp_117 = rob_uop_1_10_pdst;
      5'b01011:
        casez_tmp_117 = rob_uop_1_11_pdst;
      5'b01100:
        casez_tmp_117 = rob_uop_1_12_pdst;
      5'b01101:
        casez_tmp_117 = rob_uop_1_13_pdst;
      5'b01110:
        casez_tmp_117 = rob_uop_1_14_pdst;
      5'b01111:
        casez_tmp_117 = rob_uop_1_15_pdst;
      5'b10000:
        casez_tmp_117 = rob_uop_1_16_pdst;
      5'b10001:
        casez_tmp_117 = rob_uop_1_17_pdst;
      5'b10010:
        casez_tmp_117 = rob_uop_1_18_pdst;
      5'b10011:
        casez_tmp_117 = rob_uop_1_19_pdst;
      5'b10100:
        casez_tmp_117 = rob_uop_1_20_pdst;
      5'b10101:
        casez_tmp_117 = rob_uop_1_21_pdst;
      5'b10110:
        casez_tmp_117 = rob_uop_1_22_pdst;
      5'b10111:
        casez_tmp_117 = rob_uop_1_23_pdst;
      5'b11000:
        casez_tmp_117 = rob_uop_1_24_pdst;
      5'b11001:
        casez_tmp_117 = rob_uop_1_25_pdst;
      5'b11010:
        casez_tmp_117 = rob_uop_1_26_pdst;
      5'b11011:
        casez_tmp_117 = rob_uop_1_27_pdst;
      5'b11100:
        casez_tmp_117 = rob_uop_1_28_pdst;
      5'b11101:
        casez_tmp_117 = rob_uop_1_29_pdst;
      5'b11110:
        casez_tmp_117 = rob_uop_1_30_pdst;
      default:
        casez_tmp_117 = rob_uop_1_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_118;
  always @(*) begin
    casez (io_wb_resps_0_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_118 = rob_uop_1_0_ldst_val;
      5'b00001:
        casez_tmp_118 = rob_uop_1_1_ldst_val;
      5'b00010:
        casez_tmp_118 = rob_uop_1_2_ldst_val;
      5'b00011:
        casez_tmp_118 = rob_uop_1_3_ldst_val;
      5'b00100:
        casez_tmp_118 = rob_uop_1_4_ldst_val;
      5'b00101:
        casez_tmp_118 = rob_uop_1_5_ldst_val;
      5'b00110:
        casez_tmp_118 = rob_uop_1_6_ldst_val;
      5'b00111:
        casez_tmp_118 = rob_uop_1_7_ldst_val;
      5'b01000:
        casez_tmp_118 = rob_uop_1_8_ldst_val;
      5'b01001:
        casez_tmp_118 = rob_uop_1_9_ldst_val;
      5'b01010:
        casez_tmp_118 = rob_uop_1_10_ldst_val;
      5'b01011:
        casez_tmp_118 = rob_uop_1_11_ldst_val;
      5'b01100:
        casez_tmp_118 = rob_uop_1_12_ldst_val;
      5'b01101:
        casez_tmp_118 = rob_uop_1_13_ldst_val;
      5'b01110:
        casez_tmp_118 = rob_uop_1_14_ldst_val;
      5'b01111:
        casez_tmp_118 = rob_uop_1_15_ldst_val;
      5'b10000:
        casez_tmp_118 = rob_uop_1_16_ldst_val;
      5'b10001:
        casez_tmp_118 = rob_uop_1_17_ldst_val;
      5'b10010:
        casez_tmp_118 = rob_uop_1_18_ldst_val;
      5'b10011:
        casez_tmp_118 = rob_uop_1_19_ldst_val;
      5'b10100:
        casez_tmp_118 = rob_uop_1_20_ldst_val;
      5'b10101:
        casez_tmp_118 = rob_uop_1_21_ldst_val;
      5'b10110:
        casez_tmp_118 = rob_uop_1_22_ldst_val;
      5'b10111:
        casez_tmp_118 = rob_uop_1_23_ldst_val;
      5'b11000:
        casez_tmp_118 = rob_uop_1_24_ldst_val;
      5'b11001:
        casez_tmp_118 = rob_uop_1_25_ldst_val;
      5'b11010:
        casez_tmp_118 = rob_uop_1_26_ldst_val;
      5'b11011:
        casez_tmp_118 = rob_uop_1_27_ldst_val;
      5'b11100:
        casez_tmp_118 = rob_uop_1_28_ldst_val;
      5'b11101:
        casez_tmp_118 = rob_uop_1_29_ldst_val;
      5'b11110:
        casez_tmp_118 = rob_uop_1_30_ldst_val;
      default:
        casez_tmp_118 = rob_uop_1_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_119;
  always @(*) begin
    casez (io_wb_resps_1_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_119 = rob_val_1_0;
      5'b00001:
        casez_tmp_119 = rob_val_1_1;
      5'b00010:
        casez_tmp_119 = rob_val_1_2;
      5'b00011:
        casez_tmp_119 = rob_val_1_3;
      5'b00100:
        casez_tmp_119 = rob_val_1_4;
      5'b00101:
        casez_tmp_119 = rob_val_1_5;
      5'b00110:
        casez_tmp_119 = rob_val_1_6;
      5'b00111:
        casez_tmp_119 = rob_val_1_7;
      5'b01000:
        casez_tmp_119 = rob_val_1_8;
      5'b01001:
        casez_tmp_119 = rob_val_1_9;
      5'b01010:
        casez_tmp_119 = rob_val_1_10;
      5'b01011:
        casez_tmp_119 = rob_val_1_11;
      5'b01100:
        casez_tmp_119 = rob_val_1_12;
      5'b01101:
        casez_tmp_119 = rob_val_1_13;
      5'b01110:
        casez_tmp_119 = rob_val_1_14;
      5'b01111:
        casez_tmp_119 = rob_val_1_15;
      5'b10000:
        casez_tmp_119 = rob_val_1_16;
      5'b10001:
        casez_tmp_119 = rob_val_1_17;
      5'b10010:
        casez_tmp_119 = rob_val_1_18;
      5'b10011:
        casez_tmp_119 = rob_val_1_19;
      5'b10100:
        casez_tmp_119 = rob_val_1_20;
      5'b10101:
        casez_tmp_119 = rob_val_1_21;
      5'b10110:
        casez_tmp_119 = rob_val_1_22;
      5'b10111:
        casez_tmp_119 = rob_val_1_23;
      5'b11000:
        casez_tmp_119 = rob_val_1_24;
      5'b11001:
        casez_tmp_119 = rob_val_1_25;
      5'b11010:
        casez_tmp_119 = rob_val_1_26;
      5'b11011:
        casez_tmp_119 = rob_val_1_27;
      5'b11100:
        casez_tmp_119 = rob_val_1_28;
      5'b11101:
        casez_tmp_119 = rob_val_1_29;
      5'b11110:
        casez_tmp_119 = rob_val_1_30;
      default:
        casez_tmp_119 = rob_val_1_31;
    endcase
  end // always @(*)
  reg         casez_tmp_120;
  always @(*) begin
    casez (io_wb_resps_1_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_120 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_120 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_120 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_120 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_120 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_120 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_120 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_120 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_120 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_120 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_120 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_120 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_120 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_120 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_120 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_120 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_120 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_120 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_120 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_120 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_120 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_120 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_120 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_120 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_120 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_120 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_120 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_120 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_120 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_120 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_120 = rob_bsy_1_30;
      default:
        casez_tmp_120 = rob_bsy_1_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_121;
  always @(*) begin
    casez (io_wb_resps_1_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_121 = rob_uop_1_0_pdst;
      5'b00001:
        casez_tmp_121 = rob_uop_1_1_pdst;
      5'b00010:
        casez_tmp_121 = rob_uop_1_2_pdst;
      5'b00011:
        casez_tmp_121 = rob_uop_1_3_pdst;
      5'b00100:
        casez_tmp_121 = rob_uop_1_4_pdst;
      5'b00101:
        casez_tmp_121 = rob_uop_1_5_pdst;
      5'b00110:
        casez_tmp_121 = rob_uop_1_6_pdst;
      5'b00111:
        casez_tmp_121 = rob_uop_1_7_pdst;
      5'b01000:
        casez_tmp_121 = rob_uop_1_8_pdst;
      5'b01001:
        casez_tmp_121 = rob_uop_1_9_pdst;
      5'b01010:
        casez_tmp_121 = rob_uop_1_10_pdst;
      5'b01011:
        casez_tmp_121 = rob_uop_1_11_pdst;
      5'b01100:
        casez_tmp_121 = rob_uop_1_12_pdst;
      5'b01101:
        casez_tmp_121 = rob_uop_1_13_pdst;
      5'b01110:
        casez_tmp_121 = rob_uop_1_14_pdst;
      5'b01111:
        casez_tmp_121 = rob_uop_1_15_pdst;
      5'b10000:
        casez_tmp_121 = rob_uop_1_16_pdst;
      5'b10001:
        casez_tmp_121 = rob_uop_1_17_pdst;
      5'b10010:
        casez_tmp_121 = rob_uop_1_18_pdst;
      5'b10011:
        casez_tmp_121 = rob_uop_1_19_pdst;
      5'b10100:
        casez_tmp_121 = rob_uop_1_20_pdst;
      5'b10101:
        casez_tmp_121 = rob_uop_1_21_pdst;
      5'b10110:
        casez_tmp_121 = rob_uop_1_22_pdst;
      5'b10111:
        casez_tmp_121 = rob_uop_1_23_pdst;
      5'b11000:
        casez_tmp_121 = rob_uop_1_24_pdst;
      5'b11001:
        casez_tmp_121 = rob_uop_1_25_pdst;
      5'b11010:
        casez_tmp_121 = rob_uop_1_26_pdst;
      5'b11011:
        casez_tmp_121 = rob_uop_1_27_pdst;
      5'b11100:
        casez_tmp_121 = rob_uop_1_28_pdst;
      5'b11101:
        casez_tmp_121 = rob_uop_1_29_pdst;
      5'b11110:
        casez_tmp_121 = rob_uop_1_30_pdst;
      default:
        casez_tmp_121 = rob_uop_1_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_122;
  always @(*) begin
    casez (io_wb_resps_1_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_122 = rob_uop_1_0_ldst_val;
      5'b00001:
        casez_tmp_122 = rob_uop_1_1_ldst_val;
      5'b00010:
        casez_tmp_122 = rob_uop_1_2_ldst_val;
      5'b00011:
        casez_tmp_122 = rob_uop_1_3_ldst_val;
      5'b00100:
        casez_tmp_122 = rob_uop_1_4_ldst_val;
      5'b00101:
        casez_tmp_122 = rob_uop_1_5_ldst_val;
      5'b00110:
        casez_tmp_122 = rob_uop_1_6_ldst_val;
      5'b00111:
        casez_tmp_122 = rob_uop_1_7_ldst_val;
      5'b01000:
        casez_tmp_122 = rob_uop_1_8_ldst_val;
      5'b01001:
        casez_tmp_122 = rob_uop_1_9_ldst_val;
      5'b01010:
        casez_tmp_122 = rob_uop_1_10_ldst_val;
      5'b01011:
        casez_tmp_122 = rob_uop_1_11_ldst_val;
      5'b01100:
        casez_tmp_122 = rob_uop_1_12_ldst_val;
      5'b01101:
        casez_tmp_122 = rob_uop_1_13_ldst_val;
      5'b01110:
        casez_tmp_122 = rob_uop_1_14_ldst_val;
      5'b01111:
        casez_tmp_122 = rob_uop_1_15_ldst_val;
      5'b10000:
        casez_tmp_122 = rob_uop_1_16_ldst_val;
      5'b10001:
        casez_tmp_122 = rob_uop_1_17_ldst_val;
      5'b10010:
        casez_tmp_122 = rob_uop_1_18_ldst_val;
      5'b10011:
        casez_tmp_122 = rob_uop_1_19_ldst_val;
      5'b10100:
        casez_tmp_122 = rob_uop_1_20_ldst_val;
      5'b10101:
        casez_tmp_122 = rob_uop_1_21_ldst_val;
      5'b10110:
        casez_tmp_122 = rob_uop_1_22_ldst_val;
      5'b10111:
        casez_tmp_122 = rob_uop_1_23_ldst_val;
      5'b11000:
        casez_tmp_122 = rob_uop_1_24_ldst_val;
      5'b11001:
        casez_tmp_122 = rob_uop_1_25_ldst_val;
      5'b11010:
        casez_tmp_122 = rob_uop_1_26_ldst_val;
      5'b11011:
        casez_tmp_122 = rob_uop_1_27_ldst_val;
      5'b11100:
        casez_tmp_122 = rob_uop_1_28_ldst_val;
      5'b11101:
        casez_tmp_122 = rob_uop_1_29_ldst_val;
      5'b11110:
        casez_tmp_122 = rob_uop_1_30_ldst_val;
      default:
        casez_tmp_122 = rob_uop_1_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_123;
  always @(*) begin
    casez (io_wb_resps_2_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_123 = rob_val_1_0;
      5'b00001:
        casez_tmp_123 = rob_val_1_1;
      5'b00010:
        casez_tmp_123 = rob_val_1_2;
      5'b00011:
        casez_tmp_123 = rob_val_1_3;
      5'b00100:
        casez_tmp_123 = rob_val_1_4;
      5'b00101:
        casez_tmp_123 = rob_val_1_5;
      5'b00110:
        casez_tmp_123 = rob_val_1_6;
      5'b00111:
        casez_tmp_123 = rob_val_1_7;
      5'b01000:
        casez_tmp_123 = rob_val_1_8;
      5'b01001:
        casez_tmp_123 = rob_val_1_9;
      5'b01010:
        casez_tmp_123 = rob_val_1_10;
      5'b01011:
        casez_tmp_123 = rob_val_1_11;
      5'b01100:
        casez_tmp_123 = rob_val_1_12;
      5'b01101:
        casez_tmp_123 = rob_val_1_13;
      5'b01110:
        casez_tmp_123 = rob_val_1_14;
      5'b01111:
        casez_tmp_123 = rob_val_1_15;
      5'b10000:
        casez_tmp_123 = rob_val_1_16;
      5'b10001:
        casez_tmp_123 = rob_val_1_17;
      5'b10010:
        casez_tmp_123 = rob_val_1_18;
      5'b10011:
        casez_tmp_123 = rob_val_1_19;
      5'b10100:
        casez_tmp_123 = rob_val_1_20;
      5'b10101:
        casez_tmp_123 = rob_val_1_21;
      5'b10110:
        casez_tmp_123 = rob_val_1_22;
      5'b10111:
        casez_tmp_123 = rob_val_1_23;
      5'b11000:
        casez_tmp_123 = rob_val_1_24;
      5'b11001:
        casez_tmp_123 = rob_val_1_25;
      5'b11010:
        casez_tmp_123 = rob_val_1_26;
      5'b11011:
        casez_tmp_123 = rob_val_1_27;
      5'b11100:
        casez_tmp_123 = rob_val_1_28;
      5'b11101:
        casez_tmp_123 = rob_val_1_29;
      5'b11110:
        casez_tmp_123 = rob_val_1_30;
      default:
        casez_tmp_123 = rob_val_1_31;
    endcase
  end // always @(*)
  reg         casez_tmp_124;
  always @(*) begin
    casez (io_wb_resps_2_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_124 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_124 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_124 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_124 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_124 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_124 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_124 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_124 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_124 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_124 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_124 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_124 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_124 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_124 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_124 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_124 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_124 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_124 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_124 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_124 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_124 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_124 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_124 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_124 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_124 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_124 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_124 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_124 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_124 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_124 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_124 = rob_bsy_1_30;
      default:
        casez_tmp_124 = rob_bsy_1_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_125;
  always @(*) begin
    casez (io_wb_resps_2_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_125 = rob_uop_1_0_pdst;
      5'b00001:
        casez_tmp_125 = rob_uop_1_1_pdst;
      5'b00010:
        casez_tmp_125 = rob_uop_1_2_pdst;
      5'b00011:
        casez_tmp_125 = rob_uop_1_3_pdst;
      5'b00100:
        casez_tmp_125 = rob_uop_1_4_pdst;
      5'b00101:
        casez_tmp_125 = rob_uop_1_5_pdst;
      5'b00110:
        casez_tmp_125 = rob_uop_1_6_pdst;
      5'b00111:
        casez_tmp_125 = rob_uop_1_7_pdst;
      5'b01000:
        casez_tmp_125 = rob_uop_1_8_pdst;
      5'b01001:
        casez_tmp_125 = rob_uop_1_9_pdst;
      5'b01010:
        casez_tmp_125 = rob_uop_1_10_pdst;
      5'b01011:
        casez_tmp_125 = rob_uop_1_11_pdst;
      5'b01100:
        casez_tmp_125 = rob_uop_1_12_pdst;
      5'b01101:
        casez_tmp_125 = rob_uop_1_13_pdst;
      5'b01110:
        casez_tmp_125 = rob_uop_1_14_pdst;
      5'b01111:
        casez_tmp_125 = rob_uop_1_15_pdst;
      5'b10000:
        casez_tmp_125 = rob_uop_1_16_pdst;
      5'b10001:
        casez_tmp_125 = rob_uop_1_17_pdst;
      5'b10010:
        casez_tmp_125 = rob_uop_1_18_pdst;
      5'b10011:
        casez_tmp_125 = rob_uop_1_19_pdst;
      5'b10100:
        casez_tmp_125 = rob_uop_1_20_pdst;
      5'b10101:
        casez_tmp_125 = rob_uop_1_21_pdst;
      5'b10110:
        casez_tmp_125 = rob_uop_1_22_pdst;
      5'b10111:
        casez_tmp_125 = rob_uop_1_23_pdst;
      5'b11000:
        casez_tmp_125 = rob_uop_1_24_pdst;
      5'b11001:
        casez_tmp_125 = rob_uop_1_25_pdst;
      5'b11010:
        casez_tmp_125 = rob_uop_1_26_pdst;
      5'b11011:
        casez_tmp_125 = rob_uop_1_27_pdst;
      5'b11100:
        casez_tmp_125 = rob_uop_1_28_pdst;
      5'b11101:
        casez_tmp_125 = rob_uop_1_29_pdst;
      5'b11110:
        casez_tmp_125 = rob_uop_1_30_pdst;
      default:
        casez_tmp_125 = rob_uop_1_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_126;
  always @(*) begin
    casez (io_wb_resps_2_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_126 = rob_uop_1_0_ldst_val;
      5'b00001:
        casez_tmp_126 = rob_uop_1_1_ldst_val;
      5'b00010:
        casez_tmp_126 = rob_uop_1_2_ldst_val;
      5'b00011:
        casez_tmp_126 = rob_uop_1_3_ldst_val;
      5'b00100:
        casez_tmp_126 = rob_uop_1_4_ldst_val;
      5'b00101:
        casez_tmp_126 = rob_uop_1_5_ldst_val;
      5'b00110:
        casez_tmp_126 = rob_uop_1_6_ldst_val;
      5'b00111:
        casez_tmp_126 = rob_uop_1_7_ldst_val;
      5'b01000:
        casez_tmp_126 = rob_uop_1_8_ldst_val;
      5'b01001:
        casez_tmp_126 = rob_uop_1_9_ldst_val;
      5'b01010:
        casez_tmp_126 = rob_uop_1_10_ldst_val;
      5'b01011:
        casez_tmp_126 = rob_uop_1_11_ldst_val;
      5'b01100:
        casez_tmp_126 = rob_uop_1_12_ldst_val;
      5'b01101:
        casez_tmp_126 = rob_uop_1_13_ldst_val;
      5'b01110:
        casez_tmp_126 = rob_uop_1_14_ldst_val;
      5'b01111:
        casez_tmp_126 = rob_uop_1_15_ldst_val;
      5'b10000:
        casez_tmp_126 = rob_uop_1_16_ldst_val;
      5'b10001:
        casez_tmp_126 = rob_uop_1_17_ldst_val;
      5'b10010:
        casez_tmp_126 = rob_uop_1_18_ldst_val;
      5'b10011:
        casez_tmp_126 = rob_uop_1_19_ldst_val;
      5'b10100:
        casez_tmp_126 = rob_uop_1_20_ldst_val;
      5'b10101:
        casez_tmp_126 = rob_uop_1_21_ldst_val;
      5'b10110:
        casez_tmp_126 = rob_uop_1_22_ldst_val;
      5'b10111:
        casez_tmp_126 = rob_uop_1_23_ldst_val;
      5'b11000:
        casez_tmp_126 = rob_uop_1_24_ldst_val;
      5'b11001:
        casez_tmp_126 = rob_uop_1_25_ldst_val;
      5'b11010:
        casez_tmp_126 = rob_uop_1_26_ldst_val;
      5'b11011:
        casez_tmp_126 = rob_uop_1_27_ldst_val;
      5'b11100:
        casez_tmp_126 = rob_uop_1_28_ldst_val;
      5'b11101:
        casez_tmp_126 = rob_uop_1_29_ldst_val;
      5'b11110:
        casez_tmp_126 = rob_uop_1_30_ldst_val;
      default:
        casez_tmp_126 = rob_uop_1_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_127;
  always @(*) begin
    casez (io_wb_resps_3_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_127 = rob_val_1_0;
      5'b00001:
        casez_tmp_127 = rob_val_1_1;
      5'b00010:
        casez_tmp_127 = rob_val_1_2;
      5'b00011:
        casez_tmp_127 = rob_val_1_3;
      5'b00100:
        casez_tmp_127 = rob_val_1_4;
      5'b00101:
        casez_tmp_127 = rob_val_1_5;
      5'b00110:
        casez_tmp_127 = rob_val_1_6;
      5'b00111:
        casez_tmp_127 = rob_val_1_7;
      5'b01000:
        casez_tmp_127 = rob_val_1_8;
      5'b01001:
        casez_tmp_127 = rob_val_1_9;
      5'b01010:
        casez_tmp_127 = rob_val_1_10;
      5'b01011:
        casez_tmp_127 = rob_val_1_11;
      5'b01100:
        casez_tmp_127 = rob_val_1_12;
      5'b01101:
        casez_tmp_127 = rob_val_1_13;
      5'b01110:
        casez_tmp_127 = rob_val_1_14;
      5'b01111:
        casez_tmp_127 = rob_val_1_15;
      5'b10000:
        casez_tmp_127 = rob_val_1_16;
      5'b10001:
        casez_tmp_127 = rob_val_1_17;
      5'b10010:
        casez_tmp_127 = rob_val_1_18;
      5'b10011:
        casez_tmp_127 = rob_val_1_19;
      5'b10100:
        casez_tmp_127 = rob_val_1_20;
      5'b10101:
        casez_tmp_127 = rob_val_1_21;
      5'b10110:
        casez_tmp_127 = rob_val_1_22;
      5'b10111:
        casez_tmp_127 = rob_val_1_23;
      5'b11000:
        casez_tmp_127 = rob_val_1_24;
      5'b11001:
        casez_tmp_127 = rob_val_1_25;
      5'b11010:
        casez_tmp_127 = rob_val_1_26;
      5'b11011:
        casez_tmp_127 = rob_val_1_27;
      5'b11100:
        casez_tmp_127 = rob_val_1_28;
      5'b11101:
        casez_tmp_127 = rob_val_1_29;
      5'b11110:
        casez_tmp_127 = rob_val_1_30;
      default:
        casez_tmp_127 = rob_val_1_31;
    endcase
  end // always @(*)
  reg         casez_tmp_128;
  always @(*) begin
    casez (io_wb_resps_3_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_128 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_128 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_128 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_128 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_128 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_128 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_128 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_128 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_128 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_128 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_128 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_128 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_128 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_128 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_128 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_128 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_128 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_128 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_128 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_128 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_128 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_128 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_128 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_128 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_128 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_128 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_128 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_128 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_128 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_128 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_128 = rob_bsy_1_30;
      default:
        casez_tmp_128 = rob_bsy_1_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_129;
  always @(*) begin
    casez (io_wb_resps_3_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_129 = rob_uop_1_0_pdst;
      5'b00001:
        casez_tmp_129 = rob_uop_1_1_pdst;
      5'b00010:
        casez_tmp_129 = rob_uop_1_2_pdst;
      5'b00011:
        casez_tmp_129 = rob_uop_1_3_pdst;
      5'b00100:
        casez_tmp_129 = rob_uop_1_4_pdst;
      5'b00101:
        casez_tmp_129 = rob_uop_1_5_pdst;
      5'b00110:
        casez_tmp_129 = rob_uop_1_6_pdst;
      5'b00111:
        casez_tmp_129 = rob_uop_1_7_pdst;
      5'b01000:
        casez_tmp_129 = rob_uop_1_8_pdst;
      5'b01001:
        casez_tmp_129 = rob_uop_1_9_pdst;
      5'b01010:
        casez_tmp_129 = rob_uop_1_10_pdst;
      5'b01011:
        casez_tmp_129 = rob_uop_1_11_pdst;
      5'b01100:
        casez_tmp_129 = rob_uop_1_12_pdst;
      5'b01101:
        casez_tmp_129 = rob_uop_1_13_pdst;
      5'b01110:
        casez_tmp_129 = rob_uop_1_14_pdst;
      5'b01111:
        casez_tmp_129 = rob_uop_1_15_pdst;
      5'b10000:
        casez_tmp_129 = rob_uop_1_16_pdst;
      5'b10001:
        casez_tmp_129 = rob_uop_1_17_pdst;
      5'b10010:
        casez_tmp_129 = rob_uop_1_18_pdst;
      5'b10011:
        casez_tmp_129 = rob_uop_1_19_pdst;
      5'b10100:
        casez_tmp_129 = rob_uop_1_20_pdst;
      5'b10101:
        casez_tmp_129 = rob_uop_1_21_pdst;
      5'b10110:
        casez_tmp_129 = rob_uop_1_22_pdst;
      5'b10111:
        casez_tmp_129 = rob_uop_1_23_pdst;
      5'b11000:
        casez_tmp_129 = rob_uop_1_24_pdst;
      5'b11001:
        casez_tmp_129 = rob_uop_1_25_pdst;
      5'b11010:
        casez_tmp_129 = rob_uop_1_26_pdst;
      5'b11011:
        casez_tmp_129 = rob_uop_1_27_pdst;
      5'b11100:
        casez_tmp_129 = rob_uop_1_28_pdst;
      5'b11101:
        casez_tmp_129 = rob_uop_1_29_pdst;
      5'b11110:
        casez_tmp_129 = rob_uop_1_30_pdst;
      default:
        casez_tmp_129 = rob_uop_1_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_130;
  always @(*) begin
    casez (io_wb_resps_3_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_130 = rob_uop_1_0_ldst_val;
      5'b00001:
        casez_tmp_130 = rob_uop_1_1_ldst_val;
      5'b00010:
        casez_tmp_130 = rob_uop_1_2_ldst_val;
      5'b00011:
        casez_tmp_130 = rob_uop_1_3_ldst_val;
      5'b00100:
        casez_tmp_130 = rob_uop_1_4_ldst_val;
      5'b00101:
        casez_tmp_130 = rob_uop_1_5_ldst_val;
      5'b00110:
        casez_tmp_130 = rob_uop_1_6_ldst_val;
      5'b00111:
        casez_tmp_130 = rob_uop_1_7_ldst_val;
      5'b01000:
        casez_tmp_130 = rob_uop_1_8_ldst_val;
      5'b01001:
        casez_tmp_130 = rob_uop_1_9_ldst_val;
      5'b01010:
        casez_tmp_130 = rob_uop_1_10_ldst_val;
      5'b01011:
        casez_tmp_130 = rob_uop_1_11_ldst_val;
      5'b01100:
        casez_tmp_130 = rob_uop_1_12_ldst_val;
      5'b01101:
        casez_tmp_130 = rob_uop_1_13_ldst_val;
      5'b01110:
        casez_tmp_130 = rob_uop_1_14_ldst_val;
      5'b01111:
        casez_tmp_130 = rob_uop_1_15_ldst_val;
      5'b10000:
        casez_tmp_130 = rob_uop_1_16_ldst_val;
      5'b10001:
        casez_tmp_130 = rob_uop_1_17_ldst_val;
      5'b10010:
        casez_tmp_130 = rob_uop_1_18_ldst_val;
      5'b10011:
        casez_tmp_130 = rob_uop_1_19_ldst_val;
      5'b10100:
        casez_tmp_130 = rob_uop_1_20_ldst_val;
      5'b10101:
        casez_tmp_130 = rob_uop_1_21_ldst_val;
      5'b10110:
        casez_tmp_130 = rob_uop_1_22_ldst_val;
      5'b10111:
        casez_tmp_130 = rob_uop_1_23_ldst_val;
      5'b11000:
        casez_tmp_130 = rob_uop_1_24_ldst_val;
      5'b11001:
        casez_tmp_130 = rob_uop_1_25_ldst_val;
      5'b11010:
        casez_tmp_130 = rob_uop_1_26_ldst_val;
      5'b11011:
        casez_tmp_130 = rob_uop_1_27_ldst_val;
      5'b11100:
        casez_tmp_130 = rob_uop_1_28_ldst_val;
      5'b11101:
        casez_tmp_130 = rob_uop_1_29_ldst_val;
      5'b11110:
        casez_tmp_130 = rob_uop_1_30_ldst_val;
      default:
        casez_tmp_130 = rob_uop_1_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_131;
  always @(*) begin
    casez (io_wb_resps_4_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_131 = rob_val_1_0;
      5'b00001:
        casez_tmp_131 = rob_val_1_1;
      5'b00010:
        casez_tmp_131 = rob_val_1_2;
      5'b00011:
        casez_tmp_131 = rob_val_1_3;
      5'b00100:
        casez_tmp_131 = rob_val_1_4;
      5'b00101:
        casez_tmp_131 = rob_val_1_5;
      5'b00110:
        casez_tmp_131 = rob_val_1_6;
      5'b00111:
        casez_tmp_131 = rob_val_1_7;
      5'b01000:
        casez_tmp_131 = rob_val_1_8;
      5'b01001:
        casez_tmp_131 = rob_val_1_9;
      5'b01010:
        casez_tmp_131 = rob_val_1_10;
      5'b01011:
        casez_tmp_131 = rob_val_1_11;
      5'b01100:
        casez_tmp_131 = rob_val_1_12;
      5'b01101:
        casez_tmp_131 = rob_val_1_13;
      5'b01110:
        casez_tmp_131 = rob_val_1_14;
      5'b01111:
        casez_tmp_131 = rob_val_1_15;
      5'b10000:
        casez_tmp_131 = rob_val_1_16;
      5'b10001:
        casez_tmp_131 = rob_val_1_17;
      5'b10010:
        casez_tmp_131 = rob_val_1_18;
      5'b10011:
        casez_tmp_131 = rob_val_1_19;
      5'b10100:
        casez_tmp_131 = rob_val_1_20;
      5'b10101:
        casez_tmp_131 = rob_val_1_21;
      5'b10110:
        casez_tmp_131 = rob_val_1_22;
      5'b10111:
        casez_tmp_131 = rob_val_1_23;
      5'b11000:
        casez_tmp_131 = rob_val_1_24;
      5'b11001:
        casez_tmp_131 = rob_val_1_25;
      5'b11010:
        casez_tmp_131 = rob_val_1_26;
      5'b11011:
        casez_tmp_131 = rob_val_1_27;
      5'b11100:
        casez_tmp_131 = rob_val_1_28;
      5'b11101:
        casez_tmp_131 = rob_val_1_29;
      5'b11110:
        casez_tmp_131 = rob_val_1_30;
      default:
        casez_tmp_131 = rob_val_1_31;
    endcase
  end // always @(*)
  reg         casez_tmp_132;
  always @(*) begin
    casez (io_wb_resps_4_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_132 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_132 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_132 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_132 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_132 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_132 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_132 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_132 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_132 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_132 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_132 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_132 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_132 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_132 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_132 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_132 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_132 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_132 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_132 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_132 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_132 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_132 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_132 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_132 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_132 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_132 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_132 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_132 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_132 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_132 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_132 = rob_bsy_1_30;
      default:
        casez_tmp_132 = rob_bsy_1_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_133;
  always @(*) begin
    casez (io_wb_resps_4_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_133 = rob_uop_1_0_pdst;
      5'b00001:
        casez_tmp_133 = rob_uop_1_1_pdst;
      5'b00010:
        casez_tmp_133 = rob_uop_1_2_pdst;
      5'b00011:
        casez_tmp_133 = rob_uop_1_3_pdst;
      5'b00100:
        casez_tmp_133 = rob_uop_1_4_pdst;
      5'b00101:
        casez_tmp_133 = rob_uop_1_5_pdst;
      5'b00110:
        casez_tmp_133 = rob_uop_1_6_pdst;
      5'b00111:
        casez_tmp_133 = rob_uop_1_7_pdst;
      5'b01000:
        casez_tmp_133 = rob_uop_1_8_pdst;
      5'b01001:
        casez_tmp_133 = rob_uop_1_9_pdst;
      5'b01010:
        casez_tmp_133 = rob_uop_1_10_pdst;
      5'b01011:
        casez_tmp_133 = rob_uop_1_11_pdst;
      5'b01100:
        casez_tmp_133 = rob_uop_1_12_pdst;
      5'b01101:
        casez_tmp_133 = rob_uop_1_13_pdst;
      5'b01110:
        casez_tmp_133 = rob_uop_1_14_pdst;
      5'b01111:
        casez_tmp_133 = rob_uop_1_15_pdst;
      5'b10000:
        casez_tmp_133 = rob_uop_1_16_pdst;
      5'b10001:
        casez_tmp_133 = rob_uop_1_17_pdst;
      5'b10010:
        casez_tmp_133 = rob_uop_1_18_pdst;
      5'b10011:
        casez_tmp_133 = rob_uop_1_19_pdst;
      5'b10100:
        casez_tmp_133 = rob_uop_1_20_pdst;
      5'b10101:
        casez_tmp_133 = rob_uop_1_21_pdst;
      5'b10110:
        casez_tmp_133 = rob_uop_1_22_pdst;
      5'b10111:
        casez_tmp_133 = rob_uop_1_23_pdst;
      5'b11000:
        casez_tmp_133 = rob_uop_1_24_pdst;
      5'b11001:
        casez_tmp_133 = rob_uop_1_25_pdst;
      5'b11010:
        casez_tmp_133 = rob_uop_1_26_pdst;
      5'b11011:
        casez_tmp_133 = rob_uop_1_27_pdst;
      5'b11100:
        casez_tmp_133 = rob_uop_1_28_pdst;
      5'b11101:
        casez_tmp_133 = rob_uop_1_29_pdst;
      5'b11110:
        casez_tmp_133 = rob_uop_1_30_pdst;
      default:
        casez_tmp_133 = rob_uop_1_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_134;
  always @(*) begin
    casez (io_wb_resps_4_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_134 = rob_uop_1_0_ldst_val;
      5'b00001:
        casez_tmp_134 = rob_uop_1_1_ldst_val;
      5'b00010:
        casez_tmp_134 = rob_uop_1_2_ldst_val;
      5'b00011:
        casez_tmp_134 = rob_uop_1_3_ldst_val;
      5'b00100:
        casez_tmp_134 = rob_uop_1_4_ldst_val;
      5'b00101:
        casez_tmp_134 = rob_uop_1_5_ldst_val;
      5'b00110:
        casez_tmp_134 = rob_uop_1_6_ldst_val;
      5'b00111:
        casez_tmp_134 = rob_uop_1_7_ldst_val;
      5'b01000:
        casez_tmp_134 = rob_uop_1_8_ldst_val;
      5'b01001:
        casez_tmp_134 = rob_uop_1_9_ldst_val;
      5'b01010:
        casez_tmp_134 = rob_uop_1_10_ldst_val;
      5'b01011:
        casez_tmp_134 = rob_uop_1_11_ldst_val;
      5'b01100:
        casez_tmp_134 = rob_uop_1_12_ldst_val;
      5'b01101:
        casez_tmp_134 = rob_uop_1_13_ldst_val;
      5'b01110:
        casez_tmp_134 = rob_uop_1_14_ldst_val;
      5'b01111:
        casez_tmp_134 = rob_uop_1_15_ldst_val;
      5'b10000:
        casez_tmp_134 = rob_uop_1_16_ldst_val;
      5'b10001:
        casez_tmp_134 = rob_uop_1_17_ldst_val;
      5'b10010:
        casez_tmp_134 = rob_uop_1_18_ldst_val;
      5'b10011:
        casez_tmp_134 = rob_uop_1_19_ldst_val;
      5'b10100:
        casez_tmp_134 = rob_uop_1_20_ldst_val;
      5'b10101:
        casez_tmp_134 = rob_uop_1_21_ldst_val;
      5'b10110:
        casez_tmp_134 = rob_uop_1_22_ldst_val;
      5'b10111:
        casez_tmp_134 = rob_uop_1_23_ldst_val;
      5'b11000:
        casez_tmp_134 = rob_uop_1_24_ldst_val;
      5'b11001:
        casez_tmp_134 = rob_uop_1_25_ldst_val;
      5'b11010:
        casez_tmp_134 = rob_uop_1_26_ldst_val;
      5'b11011:
        casez_tmp_134 = rob_uop_1_27_ldst_val;
      5'b11100:
        casez_tmp_134 = rob_uop_1_28_ldst_val;
      5'b11101:
        casez_tmp_134 = rob_uop_1_29_ldst_val;
      5'b11110:
        casez_tmp_134 = rob_uop_1_30_ldst_val;
      default:
        casez_tmp_134 = rob_uop_1_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_135;
  always @(*) begin
    casez (io_wb_resps_5_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_135 = rob_val_1_0;
      5'b00001:
        casez_tmp_135 = rob_val_1_1;
      5'b00010:
        casez_tmp_135 = rob_val_1_2;
      5'b00011:
        casez_tmp_135 = rob_val_1_3;
      5'b00100:
        casez_tmp_135 = rob_val_1_4;
      5'b00101:
        casez_tmp_135 = rob_val_1_5;
      5'b00110:
        casez_tmp_135 = rob_val_1_6;
      5'b00111:
        casez_tmp_135 = rob_val_1_7;
      5'b01000:
        casez_tmp_135 = rob_val_1_8;
      5'b01001:
        casez_tmp_135 = rob_val_1_9;
      5'b01010:
        casez_tmp_135 = rob_val_1_10;
      5'b01011:
        casez_tmp_135 = rob_val_1_11;
      5'b01100:
        casez_tmp_135 = rob_val_1_12;
      5'b01101:
        casez_tmp_135 = rob_val_1_13;
      5'b01110:
        casez_tmp_135 = rob_val_1_14;
      5'b01111:
        casez_tmp_135 = rob_val_1_15;
      5'b10000:
        casez_tmp_135 = rob_val_1_16;
      5'b10001:
        casez_tmp_135 = rob_val_1_17;
      5'b10010:
        casez_tmp_135 = rob_val_1_18;
      5'b10011:
        casez_tmp_135 = rob_val_1_19;
      5'b10100:
        casez_tmp_135 = rob_val_1_20;
      5'b10101:
        casez_tmp_135 = rob_val_1_21;
      5'b10110:
        casez_tmp_135 = rob_val_1_22;
      5'b10111:
        casez_tmp_135 = rob_val_1_23;
      5'b11000:
        casez_tmp_135 = rob_val_1_24;
      5'b11001:
        casez_tmp_135 = rob_val_1_25;
      5'b11010:
        casez_tmp_135 = rob_val_1_26;
      5'b11011:
        casez_tmp_135 = rob_val_1_27;
      5'b11100:
        casez_tmp_135 = rob_val_1_28;
      5'b11101:
        casez_tmp_135 = rob_val_1_29;
      5'b11110:
        casez_tmp_135 = rob_val_1_30;
      default:
        casez_tmp_135 = rob_val_1_31;
    endcase
  end // always @(*)
  reg         casez_tmp_136;
  always @(*) begin
    casez (io_wb_resps_5_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_136 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_136 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_136 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_136 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_136 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_136 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_136 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_136 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_136 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_136 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_136 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_136 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_136 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_136 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_136 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_136 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_136 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_136 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_136 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_136 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_136 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_136 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_136 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_136 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_136 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_136 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_136 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_136 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_136 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_136 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_136 = rob_bsy_1_30;
      default:
        casez_tmp_136 = rob_bsy_1_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_137;
  always @(*) begin
    casez (io_wb_resps_5_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_137 = rob_uop_1_0_pdst;
      5'b00001:
        casez_tmp_137 = rob_uop_1_1_pdst;
      5'b00010:
        casez_tmp_137 = rob_uop_1_2_pdst;
      5'b00011:
        casez_tmp_137 = rob_uop_1_3_pdst;
      5'b00100:
        casez_tmp_137 = rob_uop_1_4_pdst;
      5'b00101:
        casez_tmp_137 = rob_uop_1_5_pdst;
      5'b00110:
        casez_tmp_137 = rob_uop_1_6_pdst;
      5'b00111:
        casez_tmp_137 = rob_uop_1_7_pdst;
      5'b01000:
        casez_tmp_137 = rob_uop_1_8_pdst;
      5'b01001:
        casez_tmp_137 = rob_uop_1_9_pdst;
      5'b01010:
        casez_tmp_137 = rob_uop_1_10_pdst;
      5'b01011:
        casez_tmp_137 = rob_uop_1_11_pdst;
      5'b01100:
        casez_tmp_137 = rob_uop_1_12_pdst;
      5'b01101:
        casez_tmp_137 = rob_uop_1_13_pdst;
      5'b01110:
        casez_tmp_137 = rob_uop_1_14_pdst;
      5'b01111:
        casez_tmp_137 = rob_uop_1_15_pdst;
      5'b10000:
        casez_tmp_137 = rob_uop_1_16_pdst;
      5'b10001:
        casez_tmp_137 = rob_uop_1_17_pdst;
      5'b10010:
        casez_tmp_137 = rob_uop_1_18_pdst;
      5'b10011:
        casez_tmp_137 = rob_uop_1_19_pdst;
      5'b10100:
        casez_tmp_137 = rob_uop_1_20_pdst;
      5'b10101:
        casez_tmp_137 = rob_uop_1_21_pdst;
      5'b10110:
        casez_tmp_137 = rob_uop_1_22_pdst;
      5'b10111:
        casez_tmp_137 = rob_uop_1_23_pdst;
      5'b11000:
        casez_tmp_137 = rob_uop_1_24_pdst;
      5'b11001:
        casez_tmp_137 = rob_uop_1_25_pdst;
      5'b11010:
        casez_tmp_137 = rob_uop_1_26_pdst;
      5'b11011:
        casez_tmp_137 = rob_uop_1_27_pdst;
      5'b11100:
        casez_tmp_137 = rob_uop_1_28_pdst;
      5'b11101:
        casez_tmp_137 = rob_uop_1_29_pdst;
      5'b11110:
        casez_tmp_137 = rob_uop_1_30_pdst;
      default:
        casez_tmp_137 = rob_uop_1_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_138;
  always @(*) begin
    casez (io_wb_resps_5_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_138 = rob_uop_1_0_ldst_val;
      5'b00001:
        casez_tmp_138 = rob_uop_1_1_ldst_val;
      5'b00010:
        casez_tmp_138 = rob_uop_1_2_ldst_val;
      5'b00011:
        casez_tmp_138 = rob_uop_1_3_ldst_val;
      5'b00100:
        casez_tmp_138 = rob_uop_1_4_ldst_val;
      5'b00101:
        casez_tmp_138 = rob_uop_1_5_ldst_val;
      5'b00110:
        casez_tmp_138 = rob_uop_1_6_ldst_val;
      5'b00111:
        casez_tmp_138 = rob_uop_1_7_ldst_val;
      5'b01000:
        casez_tmp_138 = rob_uop_1_8_ldst_val;
      5'b01001:
        casez_tmp_138 = rob_uop_1_9_ldst_val;
      5'b01010:
        casez_tmp_138 = rob_uop_1_10_ldst_val;
      5'b01011:
        casez_tmp_138 = rob_uop_1_11_ldst_val;
      5'b01100:
        casez_tmp_138 = rob_uop_1_12_ldst_val;
      5'b01101:
        casez_tmp_138 = rob_uop_1_13_ldst_val;
      5'b01110:
        casez_tmp_138 = rob_uop_1_14_ldst_val;
      5'b01111:
        casez_tmp_138 = rob_uop_1_15_ldst_val;
      5'b10000:
        casez_tmp_138 = rob_uop_1_16_ldst_val;
      5'b10001:
        casez_tmp_138 = rob_uop_1_17_ldst_val;
      5'b10010:
        casez_tmp_138 = rob_uop_1_18_ldst_val;
      5'b10011:
        casez_tmp_138 = rob_uop_1_19_ldst_val;
      5'b10100:
        casez_tmp_138 = rob_uop_1_20_ldst_val;
      5'b10101:
        casez_tmp_138 = rob_uop_1_21_ldst_val;
      5'b10110:
        casez_tmp_138 = rob_uop_1_22_ldst_val;
      5'b10111:
        casez_tmp_138 = rob_uop_1_23_ldst_val;
      5'b11000:
        casez_tmp_138 = rob_uop_1_24_ldst_val;
      5'b11001:
        casez_tmp_138 = rob_uop_1_25_ldst_val;
      5'b11010:
        casez_tmp_138 = rob_uop_1_26_ldst_val;
      5'b11011:
        casez_tmp_138 = rob_uop_1_27_ldst_val;
      5'b11100:
        casez_tmp_138 = rob_uop_1_28_ldst_val;
      5'b11101:
        casez_tmp_138 = rob_uop_1_29_ldst_val;
      5'b11110:
        casez_tmp_138 = rob_uop_1_30_ldst_val;
      default:
        casez_tmp_138 = rob_uop_1_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_139;
  always @(*) begin
    casez (io_wb_resps_6_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_139 = rob_val_1_0;
      5'b00001:
        casez_tmp_139 = rob_val_1_1;
      5'b00010:
        casez_tmp_139 = rob_val_1_2;
      5'b00011:
        casez_tmp_139 = rob_val_1_3;
      5'b00100:
        casez_tmp_139 = rob_val_1_4;
      5'b00101:
        casez_tmp_139 = rob_val_1_5;
      5'b00110:
        casez_tmp_139 = rob_val_1_6;
      5'b00111:
        casez_tmp_139 = rob_val_1_7;
      5'b01000:
        casez_tmp_139 = rob_val_1_8;
      5'b01001:
        casez_tmp_139 = rob_val_1_9;
      5'b01010:
        casez_tmp_139 = rob_val_1_10;
      5'b01011:
        casez_tmp_139 = rob_val_1_11;
      5'b01100:
        casez_tmp_139 = rob_val_1_12;
      5'b01101:
        casez_tmp_139 = rob_val_1_13;
      5'b01110:
        casez_tmp_139 = rob_val_1_14;
      5'b01111:
        casez_tmp_139 = rob_val_1_15;
      5'b10000:
        casez_tmp_139 = rob_val_1_16;
      5'b10001:
        casez_tmp_139 = rob_val_1_17;
      5'b10010:
        casez_tmp_139 = rob_val_1_18;
      5'b10011:
        casez_tmp_139 = rob_val_1_19;
      5'b10100:
        casez_tmp_139 = rob_val_1_20;
      5'b10101:
        casez_tmp_139 = rob_val_1_21;
      5'b10110:
        casez_tmp_139 = rob_val_1_22;
      5'b10111:
        casez_tmp_139 = rob_val_1_23;
      5'b11000:
        casez_tmp_139 = rob_val_1_24;
      5'b11001:
        casez_tmp_139 = rob_val_1_25;
      5'b11010:
        casez_tmp_139 = rob_val_1_26;
      5'b11011:
        casez_tmp_139 = rob_val_1_27;
      5'b11100:
        casez_tmp_139 = rob_val_1_28;
      5'b11101:
        casez_tmp_139 = rob_val_1_29;
      5'b11110:
        casez_tmp_139 = rob_val_1_30;
      default:
        casez_tmp_139 = rob_val_1_31;
    endcase
  end // always @(*)
  reg         casez_tmp_140;
  always @(*) begin
    casez (io_wb_resps_6_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_140 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_140 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_140 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_140 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_140 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_140 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_140 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_140 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_140 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_140 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_140 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_140 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_140 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_140 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_140 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_140 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_140 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_140 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_140 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_140 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_140 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_140 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_140 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_140 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_140 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_140 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_140 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_140 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_140 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_140 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_140 = rob_bsy_1_30;
      default:
        casez_tmp_140 = rob_bsy_1_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_141;
  always @(*) begin
    casez (io_wb_resps_6_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_141 = rob_uop_1_0_pdst;
      5'b00001:
        casez_tmp_141 = rob_uop_1_1_pdst;
      5'b00010:
        casez_tmp_141 = rob_uop_1_2_pdst;
      5'b00011:
        casez_tmp_141 = rob_uop_1_3_pdst;
      5'b00100:
        casez_tmp_141 = rob_uop_1_4_pdst;
      5'b00101:
        casez_tmp_141 = rob_uop_1_5_pdst;
      5'b00110:
        casez_tmp_141 = rob_uop_1_6_pdst;
      5'b00111:
        casez_tmp_141 = rob_uop_1_7_pdst;
      5'b01000:
        casez_tmp_141 = rob_uop_1_8_pdst;
      5'b01001:
        casez_tmp_141 = rob_uop_1_9_pdst;
      5'b01010:
        casez_tmp_141 = rob_uop_1_10_pdst;
      5'b01011:
        casez_tmp_141 = rob_uop_1_11_pdst;
      5'b01100:
        casez_tmp_141 = rob_uop_1_12_pdst;
      5'b01101:
        casez_tmp_141 = rob_uop_1_13_pdst;
      5'b01110:
        casez_tmp_141 = rob_uop_1_14_pdst;
      5'b01111:
        casez_tmp_141 = rob_uop_1_15_pdst;
      5'b10000:
        casez_tmp_141 = rob_uop_1_16_pdst;
      5'b10001:
        casez_tmp_141 = rob_uop_1_17_pdst;
      5'b10010:
        casez_tmp_141 = rob_uop_1_18_pdst;
      5'b10011:
        casez_tmp_141 = rob_uop_1_19_pdst;
      5'b10100:
        casez_tmp_141 = rob_uop_1_20_pdst;
      5'b10101:
        casez_tmp_141 = rob_uop_1_21_pdst;
      5'b10110:
        casez_tmp_141 = rob_uop_1_22_pdst;
      5'b10111:
        casez_tmp_141 = rob_uop_1_23_pdst;
      5'b11000:
        casez_tmp_141 = rob_uop_1_24_pdst;
      5'b11001:
        casez_tmp_141 = rob_uop_1_25_pdst;
      5'b11010:
        casez_tmp_141 = rob_uop_1_26_pdst;
      5'b11011:
        casez_tmp_141 = rob_uop_1_27_pdst;
      5'b11100:
        casez_tmp_141 = rob_uop_1_28_pdst;
      5'b11101:
        casez_tmp_141 = rob_uop_1_29_pdst;
      5'b11110:
        casez_tmp_141 = rob_uop_1_30_pdst;
      default:
        casez_tmp_141 = rob_uop_1_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_142;
  always @(*) begin
    casez (io_wb_resps_6_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_142 = rob_uop_1_0_ldst_val;
      5'b00001:
        casez_tmp_142 = rob_uop_1_1_ldst_val;
      5'b00010:
        casez_tmp_142 = rob_uop_1_2_ldst_val;
      5'b00011:
        casez_tmp_142 = rob_uop_1_3_ldst_val;
      5'b00100:
        casez_tmp_142 = rob_uop_1_4_ldst_val;
      5'b00101:
        casez_tmp_142 = rob_uop_1_5_ldst_val;
      5'b00110:
        casez_tmp_142 = rob_uop_1_6_ldst_val;
      5'b00111:
        casez_tmp_142 = rob_uop_1_7_ldst_val;
      5'b01000:
        casez_tmp_142 = rob_uop_1_8_ldst_val;
      5'b01001:
        casez_tmp_142 = rob_uop_1_9_ldst_val;
      5'b01010:
        casez_tmp_142 = rob_uop_1_10_ldst_val;
      5'b01011:
        casez_tmp_142 = rob_uop_1_11_ldst_val;
      5'b01100:
        casez_tmp_142 = rob_uop_1_12_ldst_val;
      5'b01101:
        casez_tmp_142 = rob_uop_1_13_ldst_val;
      5'b01110:
        casez_tmp_142 = rob_uop_1_14_ldst_val;
      5'b01111:
        casez_tmp_142 = rob_uop_1_15_ldst_val;
      5'b10000:
        casez_tmp_142 = rob_uop_1_16_ldst_val;
      5'b10001:
        casez_tmp_142 = rob_uop_1_17_ldst_val;
      5'b10010:
        casez_tmp_142 = rob_uop_1_18_ldst_val;
      5'b10011:
        casez_tmp_142 = rob_uop_1_19_ldst_val;
      5'b10100:
        casez_tmp_142 = rob_uop_1_20_ldst_val;
      5'b10101:
        casez_tmp_142 = rob_uop_1_21_ldst_val;
      5'b10110:
        casez_tmp_142 = rob_uop_1_22_ldst_val;
      5'b10111:
        casez_tmp_142 = rob_uop_1_23_ldst_val;
      5'b11000:
        casez_tmp_142 = rob_uop_1_24_ldst_val;
      5'b11001:
        casez_tmp_142 = rob_uop_1_25_ldst_val;
      5'b11010:
        casez_tmp_142 = rob_uop_1_26_ldst_val;
      5'b11011:
        casez_tmp_142 = rob_uop_1_27_ldst_val;
      5'b11100:
        casez_tmp_142 = rob_uop_1_28_ldst_val;
      5'b11101:
        casez_tmp_142 = rob_uop_1_29_ldst_val;
      5'b11110:
        casez_tmp_142 = rob_uop_1_30_ldst_val;
      default:
        casez_tmp_142 = rob_uop_1_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_143;
  always @(*) begin
    casez (io_wb_resps_7_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_143 = rob_val_1_0;
      5'b00001:
        casez_tmp_143 = rob_val_1_1;
      5'b00010:
        casez_tmp_143 = rob_val_1_2;
      5'b00011:
        casez_tmp_143 = rob_val_1_3;
      5'b00100:
        casez_tmp_143 = rob_val_1_4;
      5'b00101:
        casez_tmp_143 = rob_val_1_5;
      5'b00110:
        casez_tmp_143 = rob_val_1_6;
      5'b00111:
        casez_tmp_143 = rob_val_1_7;
      5'b01000:
        casez_tmp_143 = rob_val_1_8;
      5'b01001:
        casez_tmp_143 = rob_val_1_9;
      5'b01010:
        casez_tmp_143 = rob_val_1_10;
      5'b01011:
        casez_tmp_143 = rob_val_1_11;
      5'b01100:
        casez_tmp_143 = rob_val_1_12;
      5'b01101:
        casez_tmp_143 = rob_val_1_13;
      5'b01110:
        casez_tmp_143 = rob_val_1_14;
      5'b01111:
        casez_tmp_143 = rob_val_1_15;
      5'b10000:
        casez_tmp_143 = rob_val_1_16;
      5'b10001:
        casez_tmp_143 = rob_val_1_17;
      5'b10010:
        casez_tmp_143 = rob_val_1_18;
      5'b10011:
        casez_tmp_143 = rob_val_1_19;
      5'b10100:
        casez_tmp_143 = rob_val_1_20;
      5'b10101:
        casez_tmp_143 = rob_val_1_21;
      5'b10110:
        casez_tmp_143 = rob_val_1_22;
      5'b10111:
        casez_tmp_143 = rob_val_1_23;
      5'b11000:
        casez_tmp_143 = rob_val_1_24;
      5'b11001:
        casez_tmp_143 = rob_val_1_25;
      5'b11010:
        casez_tmp_143 = rob_val_1_26;
      5'b11011:
        casez_tmp_143 = rob_val_1_27;
      5'b11100:
        casez_tmp_143 = rob_val_1_28;
      5'b11101:
        casez_tmp_143 = rob_val_1_29;
      5'b11110:
        casez_tmp_143 = rob_val_1_30;
      default:
        casez_tmp_143 = rob_val_1_31;
    endcase
  end // always @(*)
  reg         casez_tmp_144;
  always @(*) begin
    casez (io_wb_resps_7_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_144 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_144 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_144 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_144 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_144 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_144 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_144 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_144 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_144 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_144 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_144 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_144 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_144 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_144 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_144 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_144 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_144 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_144 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_144 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_144 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_144 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_144 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_144 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_144 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_144 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_144 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_144 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_144 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_144 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_144 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_144 = rob_bsy_1_30;
      default:
        casez_tmp_144 = rob_bsy_1_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_145;
  always @(*) begin
    casez (io_wb_resps_7_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_145 = rob_uop_1_0_pdst;
      5'b00001:
        casez_tmp_145 = rob_uop_1_1_pdst;
      5'b00010:
        casez_tmp_145 = rob_uop_1_2_pdst;
      5'b00011:
        casez_tmp_145 = rob_uop_1_3_pdst;
      5'b00100:
        casez_tmp_145 = rob_uop_1_4_pdst;
      5'b00101:
        casez_tmp_145 = rob_uop_1_5_pdst;
      5'b00110:
        casez_tmp_145 = rob_uop_1_6_pdst;
      5'b00111:
        casez_tmp_145 = rob_uop_1_7_pdst;
      5'b01000:
        casez_tmp_145 = rob_uop_1_8_pdst;
      5'b01001:
        casez_tmp_145 = rob_uop_1_9_pdst;
      5'b01010:
        casez_tmp_145 = rob_uop_1_10_pdst;
      5'b01011:
        casez_tmp_145 = rob_uop_1_11_pdst;
      5'b01100:
        casez_tmp_145 = rob_uop_1_12_pdst;
      5'b01101:
        casez_tmp_145 = rob_uop_1_13_pdst;
      5'b01110:
        casez_tmp_145 = rob_uop_1_14_pdst;
      5'b01111:
        casez_tmp_145 = rob_uop_1_15_pdst;
      5'b10000:
        casez_tmp_145 = rob_uop_1_16_pdst;
      5'b10001:
        casez_tmp_145 = rob_uop_1_17_pdst;
      5'b10010:
        casez_tmp_145 = rob_uop_1_18_pdst;
      5'b10011:
        casez_tmp_145 = rob_uop_1_19_pdst;
      5'b10100:
        casez_tmp_145 = rob_uop_1_20_pdst;
      5'b10101:
        casez_tmp_145 = rob_uop_1_21_pdst;
      5'b10110:
        casez_tmp_145 = rob_uop_1_22_pdst;
      5'b10111:
        casez_tmp_145 = rob_uop_1_23_pdst;
      5'b11000:
        casez_tmp_145 = rob_uop_1_24_pdst;
      5'b11001:
        casez_tmp_145 = rob_uop_1_25_pdst;
      5'b11010:
        casez_tmp_145 = rob_uop_1_26_pdst;
      5'b11011:
        casez_tmp_145 = rob_uop_1_27_pdst;
      5'b11100:
        casez_tmp_145 = rob_uop_1_28_pdst;
      5'b11101:
        casez_tmp_145 = rob_uop_1_29_pdst;
      5'b11110:
        casez_tmp_145 = rob_uop_1_30_pdst;
      default:
        casez_tmp_145 = rob_uop_1_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_146;
  always @(*) begin
    casez (io_wb_resps_7_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_146 = rob_uop_1_0_ldst_val;
      5'b00001:
        casez_tmp_146 = rob_uop_1_1_ldst_val;
      5'b00010:
        casez_tmp_146 = rob_uop_1_2_ldst_val;
      5'b00011:
        casez_tmp_146 = rob_uop_1_3_ldst_val;
      5'b00100:
        casez_tmp_146 = rob_uop_1_4_ldst_val;
      5'b00101:
        casez_tmp_146 = rob_uop_1_5_ldst_val;
      5'b00110:
        casez_tmp_146 = rob_uop_1_6_ldst_val;
      5'b00111:
        casez_tmp_146 = rob_uop_1_7_ldst_val;
      5'b01000:
        casez_tmp_146 = rob_uop_1_8_ldst_val;
      5'b01001:
        casez_tmp_146 = rob_uop_1_9_ldst_val;
      5'b01010:
        casez_tmp_146 = rob_uop_1_10_ldst_val;
      5'b01011:
        casez_tmp_146 = rob_uop_1_11_ldst_val;
      5'b01100:
        casez_tmp_146 = rob_uop_1_12_ldst_val;
      5'b01101:
        casez_tmp_146 = rob_uop_1_13_ldst_val;
      5'b01110:
        casez_tmp_146 = rob_uop_1_14_ldst_val;
      5'b01111:
        casez_tmp_146 = rob_uop_1_15_ldst_val;
      5'b10000:
        casez_tmp_146 = rob_uop_1_16_ldst_val;
      5'b10001:
        casez_tmp_146 = rob_uop_1_17_ldst_val;
      5'b10010:
        casez_tmp_146 = rob_uop_1_18_ldst_val;
      5'b10011:
        casez_tmp_146 = rob_uop_1_19_ldst_val;
      5'b10100:
        casez_tmp_146 = rob_uop_1_20_ldst_val;
      5'b10101:
        casez_tmp_146 = rob_uop_1_21_ldst_val;
      5'b10110:
        casez_tmp_146 = rob_uop_1_22_ldst_val;
      5'b10111:
        casez_tmp_146 = rob_uop_1_23_ldst_val;
      5'b11000:
        casez_tmp_146 = rob_uop_1_24_ldst_val;
      5'b11001:
        casez_tmp_146 = rob_uop_1_25_ldst_val;
      5'b11010:
        casez_tmp_146 = rob_uop_1_26_ldst_val;
      5'b11011:
        casez_tmp_146 = rob_uop_1_27_ldst_val;
      5'b11100:
        casez_tmp_146 = rob_uop_1_28_ldst_val;
      5'b11101:
        casez_tmp_146 = rob_uop_1_29_ldst_val;
      5'b11110:
        casez_tmp_146 = rob_uop_1_30_ldst_val;
      default:
        casez_tmp_146 = rob_uop_1_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_147;
  always @(*) begin
    casez (io_wb_resps_8_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_147 = rob_val_1_0;
      5'b00001:
        casez_tmp_147 = rob_val_1_1;
      5'b00010:
        casez_tmp_147 = rob_val_1_2;
      5'b00011:
        casez_tmp_147 = rob_val_1_3;
      5'b00100:
        casez_tmp_147 = rob_val_1_4;
      5'b00101:
        casez_tmp_147 = rob_val_1_5;
      5'b00110:
        casez_tmp_147 = rob_val_1_6;
      5'b00111:
        casez_tmp_147 = rob_val_1_7;
      5'b01000:
        casez_tmp_147 = rob_val_1_8;
      5'b01001:
        casez_tmp_147 = rob_val_1_9;
      5'b01010:
        casez_tmp_147 = rob_val_1_10;
      5'b01011:
        casez_tmp_147 = rob_val_1_11;
      5'b01100:
        casez_tmp_147 = rob_val_1_12;
      5'b01101:
        casez_tmp_147 = rob_val_1_13;
      5'b01110:
        casez_tmp_147 = rob_val_1_14;
      5'b01111:
        casez_tmp_147 = rob_val_1_15;
      5'b10000:
        casez_tmp_147 = rob_val_1_16;
      5'b10001:
        casez_tmp_147 = rob_val_1_17;
      5'b10010:
        casez_tmp_147 = rob_val_1_18;
      5'b10011:
        casez_tmp_147 = rob_val_1_19;
      5'b10100:
        casez_tmp_147 = rob_val_1_20;
      5'b10101:
        casez_tmp_147 = rob_val_1_21;
      5'b10110:
        casez_tmp_147 = rob_val_1_22;
      5'b10111:
        casez_tmp_147 = rob_val_1_23;
      5'b11000:
        casez_tmp_147 = rob_val_1_24;
      5'b11001:
        casez_tmp_147 = rob_val_1_25;
      5'b11010:
        casez_tmp_147 = rob_val_1_26;
      5'b11011:
        casez_tmp_147 = rob_val_1_27;
      5'b11100:
        casez_tmp_147 = rob_val_1_28;
      5'b11101:
        casez_tmp_147 = rob_val_1_29;
      5'b11110:
        casez_tmp_147 = rob_val_1_30;
      default:
        casez_tmp_147 = rob_val_1_31;
    endcase
  end // always @(*)
  reg         casez_tmp_148;
  always @(*) begin
    casez (io_wb_resps_8_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_148 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_148 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_148 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_148 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_148 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_148 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_148 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_148 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_148 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_148 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_148 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_148 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_148 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_148 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_148 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_148 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_148 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_148 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_148 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_148 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_148 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_148 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_148 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_148 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_148 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_148 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_148 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_148 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_148 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_148 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_148 = rob_bsy_1_30;
      default:
        casez_tmp_148 = rob_bsy_1_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_149;
  always @(*) begin
    casez (io_wb_resps_8_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_149 = rob_uop_1_0_pdst;
      5'b00001:
        casez_tmp_149 = rob_uop_1_1_pdst;
      5'b00010:
        casez_tmp_149 = rob_uop_1_2_pdst;
      5'b00011:
        casez_tmp_149 = rob_uop_1_3_pdst;
      5'b00100:
        casez_tmp_149 = rob_uop_1_4_pdst;
      5'b00101:
        casez_tmp_149 = rob_uop_1_5_pdst;
      5'b00110:
        casez_tmp_149 = rob_uop_1_6_pdst;
      5'b00111:
        casez_tmp_149 = rob_uop_1_7_pdst;
      5'b01000:
        casez_tmp_149 = rob_uop_1_8_pdst;
      5'b01001:
        casez_tmp_149 = rob_uop_1_9_pdst;
      5'b01010:
        casez_tmp_149 = rob_uop_1_10_pdst;
      5'b01011:
        casez_tmp_149 = rob_uop_1_11_pdst;
      5'b01100:
        casez_tmp_149 = rob_uop_1_12_pdst;
      5'b01101:
        casez_tmp_149 = rob_uop_1_13_pdst;
      5'b01110:
        casez_tmp_149 = rob_uop_1_14_pdst;
      5'b01111:
        casez_tmp_149 = rob_uop_1_15_pdst;
      5'b10000:
        casez_tmp_149 = rob_uop_1_16_pdst;
      5'b10001:
        casez_tmp_149 = rob_uop_1_17_pdst;
      5'b10010:
        casez_tmp_149 = rob_uop_1_18_pdst;
      5'b10011:
        casez_tmp_149 = rob_uop_1_19_pdst;
      5'b10100:
        casez_tmp_149 = rob_uop_1_20_pdst;
      5'b10101:
        casez_tmp_149 = rob_uop_1_21_pdst;
      5'b10110:
        casez_tmp_149 = rob_uop_1_22_pdst;
      5'b10111:
        casez_tmp_149 = rob_uop_1_23_pdst;
      5'b11000:
        casez_tmp_149 = rob_uop_1_24_pdst;
      5'b11001:
        casez_tmp_149 = rob_uop_1_25_pdst;
      5'b11010:
        casez_tmp_149 = rob_uop_1_26_pdst;
      5'b11011:
        casez_tmp_149 = rob_uop_1_27_pdst;
      5'b11100:
        casez_tmp_149 = rob_uop_1_28_pdst;
      5'b11101:
        casez_tmp_149 = rob_uop_1_29_pdst;
      5'b11110:
        casez_tmp_149 = rob_uop_1_30_pdst;
      default:
        casez_tmp_149 = rob_uop_1_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_150;
  always @(*) begin
    casez (io_wb_resps_8_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_150 = rob_uop_1_0_ldst_val;
      5'b00001:
        casez_tmp_150 = rob_uop_1_1_ldst_val;
      5'b00010:
        casez_tmp_150 = rob_uop_1_2_ldst_val;
      5'b00011:
        casez_tmp_150 = rob_uop_1_3_ldst_val;
      5'b00100:
        casez_tmp_150 = rob_uop_1_4_ldst_val;
      5'b00101:
        casez_tmp_150 = rob_uop_1_5_ldst_val;
      5'b00110:
        casez_tmp_150 = rob_uop_1_6_ldst_val;
      5'b00111:
        casez_tmp_150 = rob_uop_1_7_ldst_val;
      5'b01000:
        casez_tmp_150 = rob_uop_1_8_ldst_val;
      5'b01001:
        casez_tmp_150 = rob_uop_1_9_ldst_val;
      5'b01010:
        casez_tmp_150 = rob_uop_1_10_ldst_val;
      5'b01011:
        casez_tmp_150 = rob_uop_1_11_ldst_val;
      5'b01100:
        casez_tmp_150 = rob_uop_1_12_ldst_val;
      5'b01101:
        casez_tmp_150 = rob_uop_1_13_ldst_val;
      5'b01110:
        casez_tmp_150 = rob_uop_1_14_ldst_val;
      5'b01111:
        casez_tmp_150 = rob_uop_1_15_ldst_val;
      5'b10000:
        casez_tmp_150 = rob_uop_1_16_ldst_val;
      5'b10001:
        casez_tmp_150 = rob_uop_1_17_ldst_val;
      5'b10010:
        casez_tmp_150 = rob_uop_1_18_ldst_val;
      5'b10011:
        casez_tmp_150 = rob_uop_1_19_ldst_val;
      5'b10100:
        casez_tmp_150 = rob_uop_1_20_ldst_val;
      5'b10101:
        casez_tmp_150 = rob_uop_1_21_ldst_val;
      5'b10110:
        casez_tmp_150 = rob_uop_1_22_ldst_val;
      5'b10111:
        casez_tmp_150 = rob_uop_1_23_ldst_val;
      5'b11000:
        casez_tmp_150 = rob_uop_1_24_ldst_val;
      5'b11001:
        casez_tmp_150 = rob_uop_1_25_ldst_val;
      5'b11010:
        casez_tmp_150 = rob_uop_1_26_ldst_val;
      5'b11011:
        casez_tmp_150 = rob_uop_1_27_ldst_val;
      5'b11100:
        casez_tmp_150 = rob_uop_1_28_ldst_val;
      5'b11101:
        casez_tmp_150 = rob_uop_1_29_ldst_val;
      5'b11110:
        casez_tmp_150 = rob_uop_1_30_ldst_val;
      default:
        casez_tmp_150 = rob_uop_1_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_151;
  always @(*) begin
    casez (io_wb_resps_9_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_151 = rob_val_1_0;
      5'b00001:
        casez_tmp_151 = rob_val_1_1;
      5'b00010:
        casez_tmp_151 = rob_val_1_2;
      5'b00011:
        casez_tmp_151 = rob_val_1_3;
      5'b00100:
        casez_tmp_151 = rob_val_1_4;
      5'b00101:
        casez_tmp_151 = rob_val_1_5;
      5'b00110:
        casez_tmp_151 = rob_val_1_6;
      5'b00111:
        casez_tmp_151 = rob_val_1_7;
      5'b01000:
        casez_tmp_151 = rob_val_1_8;
      5'b01001:
        casez_tmp_151 = rob_val_1_9;
      5'b01010:
        casez_tmp_151 = rob_val_1_10;
      5'b01011:
        casez_tmp_151 = rob_val_1_11;
      5'b01100:
        casez_tmp_151 = rob_val_1_12;
      5'b01101:
        casez_tmp_151 = rob_val_1_13;
      5'b01110:
        casez_tmp_151 = rob_val_1_14;
      5'b01111:
        casez_tmp_151 = rob_val_1_15;
      5'b10000:
        casez_tmp_151 = rob_val_1_16;
      5'b10001:
        casez_tmp_151 = rob_val_1_17;
      5'b10010:
        casez_tmp_151 = rob_val_1_18;
      5'b10011:
        casez_tmp_151 = rob_val_1_19;
      5'b10100:
        casez_tmp_151 = rob_val_1_20;
      5'b10101:
        casez_tmp_151 = rob_val_1_21;
      5'b10110:
        casez_tmp_151 = rob_val_1_22;
      5'b10111:
        casez_tmp_151 = rob_val_1_23;
      5'b11000:
        casez_tmp_151 = rob_val_1_24;
      5'b11001:
        casez_tmp_151 = rob_val_1_25;
      5'b11010:
        casez_tmp_151 = rob_val_1_26;
      5'b11011:
        casez_tmp_151 = rob_val_1_27;
      5'b11100:
        casez_tmp_151 = rob_val_1_28;
      5'b11101:
        casez_tmp_151 = rob_val_1_29;
      5'b11110:
        casez_tmp_151 = rob_val_1_30;
      default:
        casez_tmp_151 = rob_val_1_31;
    endcase
  end // always @(*)
  reg         casez_tmp_152;
  always @(*) begin
    casez (io_wb_resps_9_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_152 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_152 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_152 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_152 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_152 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_152 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_152 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_152 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_152 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_152 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_152 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_152 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_152 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_152 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_152 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_152 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_152 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_152 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_152 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_152 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_152 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_152 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_152 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_152 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_152 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_152 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_152 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_152 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_152 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_152 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_152 = rob_bsy_1_30;
      default:
        casez_tmp_152 = rob_bsy_1_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_153;
  always @(*) begin
    casez (io_wb_resps_9_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_153 = rob_uop_1_0_pdst;
      5'b00001:
        casez_tmp_153 = rob_uop_1_1_pdst;
      5'b00010:
        casez_tmp_153 = rob_uop_1_2_pdst;
      5'b00011:
        casez_tmp_153 = rob_uop_1_3_pdst;
      5'b00100:
        casez_tmp_153 = rob_uop_1_4_pdst;
      5'b00101:
        casez_tmp_153 = rob_uop_1_5_pdst;
      5'b00110:
        casez_tmp_153 = rob_uop_1_6_pdst;
      5'b00111:
        casez_tmp_153 = rob_uop_1_7_pdst;
      5'b01000:
        casez_tmp_153 = rob_uop_1_8_pdst;
      5'b01001:
        casez_tmp_153 = rob_uop_1_9_pdst;
      5'b01010:
        casez_tmp_153 = rob_uop_1_10_pdst;
      5'b01011:
        casez_tmp_153 = rob_uop_1_11_pdst;
      5'b01100:
        casez_tmp_153 = rob_uop_1_12_pdst;
      5'b01101:
        casez_tmp_153 = rob_uop_1_13_pdst;
      5'b01110:
        casez_tmp_153 = rob_uop_1_14_pdst;
      5'b01111:
        casez_tmp_153 = rob_uop_1_15_pdst;
      5'b10000:
        casez_tmp_153 = rob_uop_1_16_pdst;
      5'b10001:
        casez_tmp_153 = rob_uop_1_17_pdst;
      5'b10010:
        casez_tmp_153 = rob_uop_1_18_pdst;
      5'b10011:
        casez_tmp_153 = rob_uop_1_19_pdst;
      5'b10100:
        casez_tmp_153 = rob_uop_1_20_pdst;
      5'b10101:
        casez_tmp_153 = rob_uop_1_21_pdst;
      5'b10110:
        casez_tmp_153 = rob_uop_1_22_pdst;
      5'b10111:
        casez_tmp_153 = rob_uop_1_23_pdst;
      5'b11000:
        casez_tmp_153 = rob_uop_1_24_pdst;
      5'b11001:
        casez_tmp_153 = rob_uop_1_25_pdst;
      5'b11010:
        casez_tmp_153 = rob_uop_1_26_pdst;
      5'b11011:
        casez_tmp_153 = rob_uop_1_27_pdst;
      5'b11100:
        casez_tmp_153 = rob_uop_1_28_pdst;
      5'b11101:
        casez_tmp_153 = rob_uop_1_29_pdst;
      5'b11110:
        casez_tmp_153 = rob_uop_1_30_pdst;
      default:
        casez_tmp_153 = rob_uop_1_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_154;
  always @(*) begin
    casez (io_wb_resps_9_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_154 = rob_uop_1_0_ldst_val;
      5'b00001:
        casez_tmp_154 = rob_uop_1_1_ldst_val;
      5'b00010:
        casez_tmp_154 = rob_uop_1_2_ldst_val;
      5'b00011:
        casez_tmp_154 = rob_uop_1_3_ldst_val;
      5'b00100:
        casez_tmp_154 = rob_uop_1_4_ldst_val;
      5'b00101:
        casez_tmp_154 = rob_uop_1_5_ldst_val;
      5'b00110:
        casez_tmp_154 = rob_uop_1_6_ldst_val;
      5'b00111:
        casez_tmp_154 = rob_uop_1_7_ldst_val;
      5'b01000:
        casez_tmp_154 = rob_uop_1_8_ldst_val;
      5'b01001:
        casez_tmp_154 = rob_uop_1_9_ldst_val;
      5'b01010:
        casez_tmp_154 = rob_uop_1_10_ldst_val;
      5'b01011:
        casez_tmp_154 = rob_uop_1_11_ldst_val;
      5'b01100:
        casez_tmp_154 = rob_uop_1_12_ldst_val;
      5'b01101:
        casez_tmp_154 = rob_uop_1_13_ldst_val;
      5'b01110:
        casez_tmp_154 = rob_uop_1_14_ldst_val;
      5'b01111:
        casez_tmp_154 = rob_uop_1_15_ldst_val;
      5'b10000:
        casez_tmp_154 = rob_uop_1_16_ldst_val;
      5'b10001:
        casez_tmp_154 = rob_uop_1_17_ldst_val;
      5'b10010:
        casez_tmp_154 = rob_uop_1_18_ldst_val;
      5'b10011:
        casez_tmp_154 = rob_uop_1_19_ldst_val;
      5'b10100:
        casez_tmp_154 = rob_uop_1_20_ldst_val;
      5'b10101:
        casez_tmp_154 = rob_uop_1_21_ldst_val;
      5'b10110:
        casez_tmp_154 = rob_uop_1_22_ldst_val;
      5'b10111:
        casez_tmp_154 = rob_uop_1_23_ldst_val;
      5'b11000:
        casez_tmp_154 = rob_uop_1_24_ldst_val;
      5'b11001:
        casez_tmp_154 = rob_uop_1_25_ldst_val;
      5'b11010:
        casez_tmp_154 = rob_uop_1_26_ldst_val;
      5'b11011:
        casez_tmp_154 = rob_uop_1_27_ldst_val;
      5'b11100:
        casez_tmp_154 = rob_uop_1_28_ldst_val;
      5'b11101:
        casez_tmp_154 = rob_uop_1_29_ldst_val;
      5'b11110:
        casez_tmp_154 = rob_uop_1_30_ldst_val;
      default:
        casez_tmp_154 = rob_uop_1_31_ldst_val;
    endcase
  end // always @(*)
  reg         rob_val_2_0;
  reg         rob_val_2_1;
  reg         rob_val_2_2;
  reg         rob_val_2_3;
  reg         rob_val_2_4;
  reg         rob_val_2_5;
  reg         rob_val_2_6;
  reg         rob_val_2_7;
  reg         rob_val_2_8;
  reg         rob_val_2_9;
  reg         rob_val_2_10;
  reg         rob_val_2_11;
  reg         rob_val_2_12;
  reg         rob_val_2_13;
  reg         rob_val_2_14;
  reg         rob_val_2_15;
  reg         rob_val_2_16;
  reg         rob_val_2_17;
  reg         rob_val_2_18;
  reg         rob_val_2_19;
  reg         rob_val_2_20;
  reg         rob_val_2_21;
  reg         rob_val_2_22;
  reg         rob_val_2_23;
  reg         rob_val_2_24;
  reg         rob_val_2_25;
  reg         rob_val_2_26;
  reg         rob_val_2_27;
  reg         rob_val_2_28;
  reg         rob_val_2_29;
  reg         rob_val_2_30;
  reg         rob_val_2_31;
  reg         rob_bsy_2_0;
  reg         rob_bsy_2_1;
  reg         rob_bsy_2_2;
  reg         rob_bsy_2_3;
  reg         rob_bsy_2_4;
  reg         rob_bsy_2_5;
  reg         rob_bsy_2_6;
  reg         rob_bsy_2_7;
  reg         rob_bsy_2_8;
  reg         rob_bsy_2_9;
  reg         rob_bsy_2_10;
  reg         rob_bsy_2_11;
  reg         rob_bsy_2_12;
  reg         rob_bsy_2_13;
  reg         rob_bsy_2_14;
  reg         rob_bsy_2_15;
  reg         rob_bsy_2_16;
  reg         rob_bsy_2_17;
  reg         rob_bsy_2_18;
  reg         rob_bsy_2_19;
  reg         rob_bsy_2_20;
  reg         rob_bsy_2_21;
  reg         rob_bsy_2_22;
  reg         rob_bsy_2_23;
  reg         rob_bsy_2_24;
  reg         rob_bsy_2_25;
  reg         rob_bsy_2_26;
  reg         rob_bsy_2_27;
  reg         rob_bsy_2_28;
  reg         rob_bsy_2_29;
  reg         rob_bsy_2_30;
  reg         rob_bsy_2_31;
  reg         rob_unsafe_2_0;
  reg         rob_unsafe_2_1;
  reg         rob_unsafe_2_2;
  reg         rob_unsafe_2_3;
  reg         rob_unsafe_2_4;
  reg         rob_unsafe_2_5;
  reg         rob_unsafe_2_6;
  reg         rob_unsafe_2_7;
  reg         rob_unsafe_2_8;
  reg         rob_unsafe_2_9;
  reg         rob_unsafe_2_10;
  reg         rob_unsafe_2_11;
  reg         rob_unsafe_2_12;
  reg         rob_unsafe_2_13;
  reg         rob_unsafe_2_14;
  reg         rob_unsafe_2_15;
  reg         rob_unsafe_2_16;
  reg         rob_unsafe_2_17;
  reg         rob_unsafe_2_18;
  reg         rob_unsafe_2_19;
  reg         rob_unsafe_2_20;
  reg         rob_unsafe_2_21;
  reg         rob_unsafe_2_22;
  reg         rob_unsafe_2_23;
  reg         rob_unsafe_2_24;
  reg         rob_unsafe_2_25;
  reg         rob_unsafe_2_26;
  reg         rob_unsafe_2_27;
  reg         rob_unsafe_2_28;
  reg         rob_unsafe_2_29;
  reg         rob_unsafe_2_30;
  reg         rob_unsafe_2_31;
  reg  [6:0]  rob_uop_2_0_uopc;
  reg         rob_uop_2_0_is_rvc;
  reg         rob_uop_2_0_is_br;
  reg         rob_uop_2_0_is_jalr;
  reg         rob_uop_2_0_is_jal;
  reg  [19:0] rob_uop_2_0_br_mask;
  reg  [5:0]  rob_uop_2_0_ftq_idx;
  reg         rob_uop_2_0_edge_inst;
  reg  [5:0]  rob_uop_2_0_pc_lob;
  reg  [6:0]  rob_uop_2_0_pdst;
  reg  [6:0]  rob_uop_2_0_stale_pdst;
  reg         rob_uop_2_0_is_fencei;
  reg         rob_uop_2_0_uses_ldq;
  reg         rob_uop_2_0_uses_stq;
  reg         rob_uop_2_0_is_sys_pc2epc;
  reg         rob_uop_2_0_flush_on_commit;
  reg  [5:0]  rob_uop_2_0_ldst;
  reg         rob_uop_2_0_ldst_val;
  reg  [1:0]  rob_uop_2_0_dst_rtype;
  reg         rob_uop_2_0_fp_val;
  reg  [1:0]  rob_uop_2_0_debug_fsrc;
  reg  [6:0]  rob_uop_2_1_uopc;
  reg         rob_uop_2_1_is_rvc;
  reg         rob_uop_2_1_is_br;
  reg         rob_uop_2_1_is_jalr;
  reg         rob_uop_2_1_is_jal;
  reg  [19:0] rob_uop_2_1_br_mask;
  reg  [5:0]  rob_uop_2_1_ftq_idx;
  reg         rob_uop_2_1_edge_inst;
  reg  [5:0]  rob_uop_2_1_pc_lob;
  reg  [6:0]  rob_uop_2_1_pdst;
  reg  [6:0]  rob_uop_2_1_stale_pdst;
  reg         rob_uop_2_1_is_fencei;
  reg         rob_uop_2_1_uses_ldq;
  reg         rob_uop_2_1_uses_stq;
  reg         rob_uop_2_1_is_sys_pc2epc;
  reg         rob_uop_2_1_flush_on_commit;
  reg  [5:0]  rob_uop_2_1_ldst;
  reg         rob_uop_2_1_ldst_val;
  reg  [1:0]  rob_uop_2_1_dst_rtype;
  reg         rob_uop_2_1_fp_val;
  reg  [1:0]  rob_uop_2_1_debug_fsrc;
  reg  [6:0]  rob_uop_2_2_uopc;
  reg         rob_uop_2_2_is_rvc;
  reg         rob_uop_2_2_is_br;
  reg         rob_uop_2_2_is_jalr;
  reg         rob_uop_2_2_is_jal;
  reg  [19:0] rob_uop_2_2_br_mask;
  reg  [5:0]  rob_uop_2_2_ftq_idx;
  reg         rob_uop_2_2_edge_inst;
  reg  [5:0]  rob_uop_2_2_pc_lob;
  reg  [6:0]  rob_uop_2_2_pdst;
  reg  [6:0]  rob_uop_2_2_stale_pdst;
  reg         rob_uop_2_2_is_fencei;
  reg         rob_uop_2_2_uses_ldq;
  reg         rob_uop_2_2_uses_stq;
  reg         rob_uop_2_2_is_sys_pc2epc;
  reg         rob_uop_2_2_flush_on_commit;
  reg  [5:0]  rob_uop_2_2_ldst;
  reg         rob_uop_2_2_ldst_val;
  reg  [1:0]  rob_uop_2_2_dst_rtype;
  reg         rob_uop_2_2_fp_val;
  reg  [1:0]  rob_uop_2_2_debug_fsrc;
  reg  [6:0]  rob_uop_2_3_uopc;
  reg         rob_uop_2_3_is_rvc;
  reg         rob_uop_2_3_is_br;
  reg         rob_uop_2_3_is_jalr;
  reg         rob_uop_2_3_is_jal;
  reg  [19:0] rob_uop_2_3_br_mask;
  reg  [5:0]  rob_uop_2_3_ftq_idx;
  reg         rob_uop_2_3_edge_inst;
  reg  [5:0]  rob_uop_2_3_pc_lob;
  reg  [6:0]  rob_uop_2_3_pdst;
  reg  [6:0]  rob_uop_2_3_stale_pdst;
  reg         rob_uop_2_3_is_fencei;
  reg         rob_uop_2_3_uses_ldq;
  reg         rob_uop_2_3_uses_stq;
  reg         rob_uop_2_3_is_sys_pc2epc;
  reg         rob_uop_2_3_flush_on_commit;
  reg  [5:0]  rob_uop_2_3_ldst;
  reg         rob_uop_2_3_ldst_val;
  reg  [1:0]  rob_uop_2_3_dst_rtype;
  reg         rob_uop_2_3_fp_val;
  reg  [1:0]  rob_uop_2_3_debug_fsrc;
  reg  [6:0]  rob_uop_2_4_uopc;
  reg         rob_uop_2_4_is_rvc;
  reg         rob_uop_2_4_is_br;
  reg         rob_uop_2_4_is_jalr;
  reg         rob_uop_2_4_is_jal;
  reg  [19:0] rob_uop_2_4_br_mask;
  reg  [5:0]  rob_uop_2_4_ftq_idx;
  reg         rob_uop_2_4_edge_inst;
  reg  [5:0]  rob_uop_2_4_pc_lob;
  reg  [6:0]  rob_uop_2_4_pdst;
  reg  [6:0]  rob_uop_2_4_stale_pdst;
  reg         rob_uop_2_4_is_fencei;
  reg         rob_uop_2_4_uses_ldq;
  reg         rob_uop_2_4_uses_stq;
  reg         rob_uop_2_4_is_sys_pc2epc;
  reg         rob_uop_2_4_flush_on_commit;
  reg  [5:0]  rob_uop_2_4_ldst;
  reg         rob_uop_2_4_ldst_val;
  reg  [1:0]  rob_uop_2_4_dst_rtype;
  reg         rob_uop_2_4_fp_val;
  reg  [1:0]  rob_uop_2_4_debug_fsrc;
  reg  [6:0]  rob_uop_2_5_uopc;
  reg         rob_uop_2_5_is_rvc;
  reg         rob_uop_2_5_is_br;
  reg         rob_uop_2_5_is_jalr;
  reg         rob_uop_2_5_is_jal;
  reg  [19:0] rob_uop_2_5_br_mask;
  reg  [5:0]  rob_uop_2_5_ftq_idx;
  reg         rob_uop_2_5_edge_inst;
  reg  [5:0]  rob_uop_2_5_pc_lob;
  reg  [6:0]  rob_uop_2_5_pdst;
  reg  [6:0]  rob_uop_2_5_stale_pdst;
  reg         rob_uop_2_5_is_fencei;
  reg         rob_uop_2_5_uses_ldq;
  reg         rob_uop_2_5_uses_stq;
  reg         rob_uop_2_5_is_sys_pc2epc;
  reg         rob_uop_2_5_flush_on_commit;
  reg  [5:0]  rob_uop_2_5_ldst;
  reg         rob_uop_2_5_ldst_val;
  reg  [1:0]  rob_uop_2_5_dst_rtype;
  reg         rob_uop_2_5_fp_val;
  reg  [1:0]  rob_uop_2_5_debug_fsrc;
  reg  [6:0]  rob_uop_2_6_uopc;
  reg         rob_uop_2_6_is_rvc;
  reg         rob_uop_2_6_is_br;
  reg         rob_uop_2_6_is_jalr;
  reg         rob_uop_2_6_is_jal;
  reg  [19:0] rob_uop_2_6_br_mask;
  reg  [5:0]  rob_uop_2_6_ftq_idx;
  reg         rob_uop_2_6_edge_inst;
  reg  [5:0]  rob_uop_2_6_pc_lob;
  reg  [6:0]  rob_uop_2_6_pdst;
  reg  [6:0]  rob_uop_2_6_stale_pdst;
  reg         rob_uop_2_6_is_fencei;
  reg         rob_uop_2_6_uses_ldq;
  reg         rob_uop_2_6_uses_stq;
  reg         rob_uop_2_6_is_sys_pc2epc;
  reg         rob_uop_2_6_flush_on_commit;
  reg  [5:0]  rob_uop_2_6_ldst;
  reg         rob_uop_2_6_ldst_val;
  reg  [1:0]  rob_uop_2_6_dst_rtype;
  reg         rob_uop_2_6_fp_val;
  reg  [1:0]  rob_uop_2_6_debug_fsrc;
  reg  [6:0]  rob_uop_2_7_uopc;
  reg         rob_uop_2_7_is_rvc;
  reg         rob_uop_2_7_is_br;
  reg         rob_uop_2_7_is_jalr;
  reg         rob_uop_2_7_is_jal;
  reg  [19:0] rob_uop_2_7_br_mask;
  reg  [5:0]  rob_uop_2_7_ftq_idx;
  reg         rob_uop_2_7_edge_inst;
  reg  [5:0]  rob_uop_2_7_pc_lob;
  reg  [6:0]  rob_uop_2_7_pdst;
  reg  [6:0]  rob_uop_2_7_stale_pdst;
  reg         rob_uop_2_7_is_fencei;
  reg         rob_uop_2_7_uses_ldq;
  reg         rob_uop_2_7_uses_stq;
  reg         rob_uop_2_7_is_sys_pc2epc;
  reg         rob_uop_2_7_flush_on_commit;
  reg  [5:0]  rob_uop_2_7_ldst;
  reg         rob_uop_2_7_ldst_val;
  reg  [1:0]  rob_uop_2_7_dst_rtype;
  reg         rob_uop_2_7_fp_val;
  reg  [1:0]  rob_uop_2_7_debug_fsrc;
  reg  [6:0]  rob_uop_2_8_uopc;
  reg         rob_uop_2_8_is_rvc;
  reg         rob_uop_2_8_is_br;
  reg         rob_uop_2_8_is_jalr;
  reg         rob_uop_2_8_is_jal;
  reg  [19:0] rob_uop_2_8_br_mask;
  reg  [5:0]  rob_uop_2_8_ftq_idx;
  reg         rob_uop_2_8_edge_inst;
  reg  [5:0]  rob_uop_2_8_pc_lob;
  reg  [6:0]  rob_uop_2_8_pdst;
  reg  [6:0]  rob_uop_2_8_stale_pdst;
  reg         rob_uop_2_8_is_fencei;
  reg         rob_uop_2_8_uses_ldq;
  reg         rob_uop_2_8_uses_stq;
  reg         rob_uop_2_8_is_sys_pc2epc;
  reg         rob_uop_2_8_flush_on_commit;
  reg  [5:0]  rob_uop_2_8_ldst;
  reg         rob_uop_2_8_ldst_val;
  reg  [1:0]  rob_uop_2_8_dst_rtype;
  reg         rob_uop_2_8_fp_val;
  reg  [1:0]  rob_uop_2_8_debug_fsrc;
  reg  [6:0]  rob_uop_2_9_uopc;
  reg         rob_uop_2_9_is_rvc;
  reg         rob_uop_2_9_is_br;
  reg         rob_uop_2_9_is_jalr;
  reg         rob_uop_2_9_is_jal;
  reg  [19:0] rob_uop_2_9_br_mask;
  reg  [5:0]  rob_uop_2_9_ftq_idx;
  reg         rob_uop_2_9_edge_inst;
  reg  [5:0]  rob_uop_2_9_pc_lob;
  reg  [6:0]  rob_uop_2_9_pdst;
  reg  [6:0]  rob_uop_2_9_stale_pdst;
  reg         rob_uop_2_9_is_fencei;
  reg         rob_uop_2_9_uses_ldq;
  reg         rob_uop_2_9_uses_stq;
  reg         rob_uop_2_9_is_sys_pc2epc;
  reg         rob_uop_2_9_flush_on_commit;
  reg  [5:0]  rob_uop_2_9_ldst;
  reg         rob_uop_2_9_ldst_val;
  reg  [1:0]  rob_uop_2_9_dst_rtype;
  reg         rob_uop_2_9_fp_val;
  reg  [1:0]  rob_uop_2_9_debug_fsrc;
  reg  [6:0]  rob_uop_2_10_uopc;
  reg         rob_uop_2_10_is_rvc;
  reg         rob_uop_2_10_is_br;
  reg         rob_uop_2_10_is_jalr;
  reg         rob_uop_2_10_is_jal;
  reg  [19:0] rob_uop_2_10_br_mask;
  reg  [5:0]  rob_uop_2_10_ftq_idx;
  reg         rob_uop_2_10_edge_inst;
  reg  [5:0]  rob_uop_2_10_pc_lob;
  reg  [6:0]  rob_uop_2_10_pdst;
  reg  [6:0]  rob_uop_2_10_stale_pdst;
  reg         rob_uop_2_10_is_fencei;
  reg         rob_uop_2_10_uses_ldq;
  reg         rob_uop_2_10_uses_stq;
  reg         rob_uop_2_10_is_sys_pc2epc;
  reg         rob_uop_2_10_flush_on_commit;
  reg  [5:0]  rob_uop_2_10_ldst;
  reg         rob_uop_2_10_ldst_val;
  reg  [1:0]  rob_uop_2_10_dst_rtype;
  reg         rob_uop_2_10_fp_val;
  reg  [1:0]  rob_uop_2_10_debug_fsrc;
  reg  [6:0]  rob_uop_2_11_uopc;
  reg         rob_uop_2_11_is_rvc;
  reg         rob_uop_2_11_is_br;
  reg         rob_uop_2_11_is_jalr;
  reg         rob_uop_2_11_is_jal;
  reg  [19:0] rob_uop_2_11_br_mask;
  reg  [5:0]  rob_uop_2_11_ftq_idx;
  reg         rob_uop_2_11_edge_inst;
  reg  [5:0]  rob_uop_2_11_pc_lob;
  reg  [6:0]  rob_uop_2_11_pdst;
  reg  [6:0]  rob_uop_2_11_stale_pdst;
  reg         rob_uop_2_11_is_fencei;
  reg         rob_uop_2_11_uses_ldq;
  reg         rob_uop_2_11_uses_stq;
  reg         rob_uop_2_11_is_sys_pc2epc;
  reg         rob_uop_2_11_flush_on_commit;
  reg  [5:0]  rob_uop_2_11_ldst;
  reg         rob_uop_2_11_ldst_val;
  reg  [1:0]  rob_uop_2_11_dst_rtype;
  reg         rob_uop_2_11_fp_val;
  reg  [1:0]  rob_uop_2_11_debug_fsrc;
  reg  [6:0]  rob_uop_2_12_uopc;
  reg         rob_uop_2_12_is_rvc;
  reg         rob_uop_2_12_is_br;
  reg         rob_uop_2_12_is_jalr;
  reg         rob_uop_2_12_is_jal;
  reg  [19:0] rob_uop_2_12_br_mask;
  reg  [5:0]  rob_uop_2_12_ftq_idx;
  reg         rob_uop_2_12_edge_inst;
  reg  [5:0]  rob_uop_2_12_pc_lob;
  reg  [6:0]  rob_uop_2_12_pdst;
  reg  [6:0]  rob_uop_2_12_stale_pdst;
  reg         rob_uop_2_12_is_fencei;
  reg         rob_uop_2_12_uses_ldq;
  reg         rob_uop_2_12_uses_stq;
  reg         rob_uop_2_12_is_sys_pc2epc;
  reg         rob_uop_2_12_flush_on_commit;
  reg  [5:0]  rob_uop_2_12_ldst;
  reg         rob_uop_2_12_ldst_val;
  reg  [1:0]  rob_uop_2_12_dst_rtype;
  reg         rob_uop_2_12_fp_val;
  reg  [1:0]  rob_uop_2_12_debug_fsrc;
  reg  [6:0]  rob_uop_2_13_uopc;
  reg         rob_uop_2_13_is_rvc;
  reg         rob_uop_2_13_is_br;
  reg         rob_uop_2_13_is_jalr;
  reg         rob_uop_2_13_is_jal;
  reg  [19:0] rob_uop_2_13_br_mask;
  reg  [5:0]  rob_uop_2_13_ftq_idx;
  reg         rob_uop_2_13_edge_inst;
  reg  [5:0]  rob_uop_2_13_pc_lob;
  reg  [6:0]  rob_uop_2_13_pdst;
  reg  [6:0]  rob_uop_2_13_stale_pdst;
  reg         rob_uop_2_13_is_fencei;
  reg         rob_uop_2_13_uses_ldq;
  reg         rob_uop_2_13_uses_stq;
  reg         rob_uop_2_13_is_sys_pc2epc;
  reg         rob_uop_2_13_flush_on_commit;
  reg  [5:0]  rob_uop_2_13_ldst;
  reg         rob_uop_2_13_ldst_val;
  reg  [1:0]  rob_uop_2_13_dst_rtype;
  reg         rob_uop_2_13_fp_val;
  reg  [1:0]  rob_uop_2_13_debug_fsrc;
  reg  [6:0]  rob_uop_2_14_uopc;
  reg         rob_uop_2_14_is_rvc;
  reg         rob_uop_2_14_is_br;
  reg         rob_uop_2_14_is_jalr;
  reg         rob_uop_2_14_is_jal;
  reg  [19:0] rob_uop_2_14_br_mask;
  reg  [5:0]  rob_uop_2_14_ftq_idx;
  reg         rob_uop_2_14_edge_inst;
  reg  [5:0]  rob_uop_2_14_pc_lob;
  reg  [6:0]  rob_uop_2_14_pdst;
  reg  [6:0]  rob_uop_2_14_stale_pdst;
  reg         rob_uop_2_14_is_fencei;
  reg         rob_uop_2_14_uses_ldq;
  reg         rob_uop_2_14_uses_stq;
  reg         rob_uop_2_14_is_sys_pc2epc;
  reg         rob_uop_2_14_flush_on_commit;
  reg  [5:0]  rob_uop_2_14_ldst;
  reg         rob_uop_2_14_ldst_val;
  reg  [1:0]  rob_uop_2_14_dst_rtype;
  reg         rob_uop_2_14_fp_val;
  reg  [1:0]  rob_uop_2_14_debug_fsrc;
  reg  [6:0]  rob_uop_2_15_uopc;
  reg         rob_uop_2_15_is_rvc;
  reg         rob_uop_2_15_is_br;
  reg         rob_uop_2_15_is_jalr;
  reg         rob_uop_2_15_is_jal;
  reg  [19:0] rob_uop_2_15_br_mask;
  reg  [5:0]  rob_uop_2_15_ftq_idx;
  reg         rob_uop_2_15_edge_inst;
  reg  [5:0]  rob_uop_2_15_pc_lob;
  reg  [6:0]  rob_uop_2_15_pdst;
  reg  [6:0]  rob_uop_2_15_stale_pdst;
  reg         rob_uop_2_15_is_fencei;
  reg         rob_uop_2_15_uses_ldq;
  reg         rob_uop_2_15_uses_stq;
  reg         rob_uop_2_15_is_sys_pc2epc;
  reg         rob_uop_2_15_flush_on_commit;
  reg  [5:0]  rob_uop_2_15_ldst;
  reg         rob_uop_2_15_ldst_val;
  reg  [1:0]  rob_uop_2_15_dst_rtype;
  reg         rob_uop_2_15_fp_val;
  reg  [1:0]  rob_uop_2_15_debug_fsrc;
  reg  [6:0]  rob_uop_2_16_uopc;
  reg         rob_uop_2_16_is_rvc;
  reg         rob_uop_2_16_is_br;
  reg         rob_uop_2_16_is_jalr;
  reg         rob_uop_2_16_is_jal;
  reg  [19:0] rob_uop_2_16_br_mask;
  reg  [5:0]  rob_uop_2_16_ftq_idx;
  reg         rob_uop_2_16_edge_inst;
  reg  [5:0]  rob_uop_2_16_pc_lob;
  reg  [6:0]  rob_uop_2_16_pdst;
  reg  [6:0]  rob_uop_2_16_stale_pdst;
  reg         rob_uop_2_16_is_fencei;
  reg         rob_uop_2_16_uses_ldq;
  reg         rob_uop_2_16_uses_stq;
  reg         rob_uop_2_16_is_sys_pc2epc;
  reg         rob_uop_2_16_flush_on_commit;
  reg  [5:0]  rob_uop_2_16_ldst;
  reg         rob_uop_2_16_ldst_val;
  reg  [1:0]  rob_uop_2_16_dst_rtype;
  reg         rob_uop_2_16_fp_val;
  reg  [1:0]  rob_uop_2_16_debug_fsrc;
  reg  [6:0]  rob_uop_2_17_uopc;
  reg         rob_uop_2_17_is_rvc;
  reg         rob_uop_2_17_is_br;
  reg         rob_uop_2_17_is_jalr;
  reg         rob_uop_2_17_is_jal;
  reg  [19:0] rob_uop_2_17_br_mask;
  reg  [5:0]  rob_uop_2_17_ftq_idx;
  reg         rob_uop_2_17_edge_inst;
  reg  [5:0]  rob_uop_2_17_pc_lob;
  reg  [6:0]  rob_uop_2_17_pdst;
  reg  [6:0]  rob_uop_2_17_stale_pdst;
  reg         rob_uop_2_17_is_fencei;
  reg         rob_uop_2_17_uses_ldq;
  reg         rob_uop_2_17_uses_stq;
  reg         rob_uop_2_17_is_sys_pc2epc;
  reg         rob_uop_2_17_flush_on_commit;
  reg  [5:0]  rob_uop_2_17_ldst;
  reg         rob_uop_2_17_ldst_val;
  reg  [1:0]  rob_uop_2_17_dst_rtype;
  reg         rob_uop_2_17_fp_val;
  reg  [1:0]  rob_uop_2_17_debug_fsrc;
  reg  [6:0]  rob_uop_2_18_uopc;
  reg         rob_uop_2_18_is_rvc;
  reg         rob_uop_2_18_is_br;
  reg         rob_uop_2_18_is_jalr;
  reg         rob_uop_2_18_is_jal;
  reg  [19:0] rob_uop_2_18_br_mask;
  reg  [5:0]  rob_uop_2_18_ftq_idx;
  reg         rob_uop_2_18_edge_inst;
  reg  [5:0]  rob_uop_2_18_pc_lob;
  reg  [6:0]  rob_uop_2_18_pdst;
  reg  [6:0]  rob_uop_2_18_stale_pdst;
  reg         rob_uop_2_18_is_fencei;
  reg         rob_uop_2_18_uses_ldq;
  reg         rob_uop_2_18_uses_stq;
  reg         rob_uop_2_18_is_sys_pc2epc;
  reg         rob_uop_2_18_flush_on_commit;
  reg  [5:0]  rob_uop_2_18_ldst;
  reg         rob_uop_2_18_ldst_val;
  reg  [1:0]  rob_uop_2_18_dst_rtype;
  reg         rob_uop_2_18_fp_val;
  reg  [1:0]  rob_uop_2_18_debug_fsrc;
  reg  [6:0]  rob_uop_2_19_uopc;
  reg         rob_uop_2_19_is_rvc;
  reg         rob_uop_2_19_is_br;
  reg         rob_uop_2_19_is_jalr;
  reg         rob_uop_2_19_is_jal;
  reg  [19:0] rob_uop_2_19_br_mask;
  reg  [5:0]  rob_uop_2_19_ftq_idx;
  reg         rob_uop_2_19_edge_inst;
  reg  [5:0]  rob_uop_2_19_pc_lob;
  reg  [6:0]  rob_uop_2_19_pdst;
  reg  [6:0]  rob_uop_2_19_stale_pdst;
  reg         rob_uop_2_19_is_fencei;
  reg         rob_uop_2_19_uses_ldq;
  reg         rob_uop_2_19_uses_stq;
  reg         rob_uop_2_19_is_sys_pc2epc;
  reg         rob_uop_2_19_flush_on_commit;
  reg  [5:0]  rob_uop_2_19_ldst;
  reg         rob_uop_2_19_ldst_val;
  reg  [1:0]  rob_uop_2_19_dst_rtype;
  reg         rob_uop_2_19_fp_val;
  reg  [1:0]  rob_uop_2_19_debug_fsrc;
  reg  [6:0]  rob_uop_2_20_uopc;
  reg         rob_uop_2_20_is_rvc;
  reg         rob_uop_2_20_is_br;
  reg         rob_uop_2_20_is_jalr;
  reg         rob_uop_2_20_is_jal;
  reg  [19:0] rob_uop_2_20_br_mask;
  reg  [5:0]  rob_uop_2_20_ftq_idx;
  reg         rob_uop_2_20_edge_inst;
  reg  [5:0]  rob_uop_2_20_pc_lob;
  reg  [6:0]  rob_uop_2_20_pdst;
  reg  [6:0]  rob_uop_2_20_stale_pdst;
  reg         rob_uop_2_20_is_fencei;
  reg         rob_uop_2_20_uses_ldq;
  reg         rob_uop_2_20_uses_stq;
  reg         rob_uop_2_20_is_sys_pc2epc;
  reg         rob_uop_2_20_flush_on_commit;
  reg  [5:0]  rob_uop_2_20_ldst;
  reg         rob_uop_2_20_ldst_val;
  reg  [1:0]  rob_uop_2_20_dst_rtype;
  reg         rob_uop_2_20_fp_val;
  reg  [1:0]  rob_uop_2_20_debug_fsrc;
  reg  [6:0]  rob_uop_2_21_uopc;
  reg         rob_uop_2_21_is_rvc;
  reg         rob_uop_2_21_is_br;
  reg         rob_uop_2_21_is_jalr;
  reg         rob_uop_2_21_is_jal;
  reg  [19:0] rob_uop_2_21_br_mask;
  reg  [5:0]  rob_uop_2_21_ftq_idx;
  reg         rob_uop_2_21_edge_inst;
  reg  [5:0]  rob_uop_2_21_pc_lob;
  reg  [6:0]  rob_uop_2_21_pdst;
  reg  [6:0]  rob_uop_2_21_stale_pdst;
  reg         rob_uop_2_21_is_fencei;
  reg         rob_uop_2_21_uses_ldq;
  reg         rob_uop_2_21_uses_stq;
  reg         rob_uop_2_21_is_sys_pc2epc;
  reg         rob_uop_2_21_flush_on_commit;
  reg  [5:0]  rob_uop_2_21_ldst;
  reg         rob_uop_2_21_ldst_val;
  reg  [1:0]  rob_uop_2_21_dst_rtype;
  reg         rob_uop_2_21_fp_val;
  reg  [1:0]  rob_uop_2_21_debug_fsrc;
  reg  [6:0]  rob_uop_2_22_uopc;
  reg         rob_uop_2_22_is_rvc;
  reg         rob_uop_2_22_is_br;
  reg         rob_uop_2_22_is_jalr;
  reg         rob_uop_2_22_is_jal;
  reg  [19:0] rob_uop_2_22_br_mask;
  reg  [5:0]  rob_uop_2_22_ftq_idx;
  reg         rob_uop_2_22_edge_inst;
  reg  [5:0]  rob_uop_2_22_pc_lob;
  reg  [6:0]  rob_uop_2_22_pdst;
  reg  [6:0]  rob_uop_2_22_stale_pdst;
  reg         rob_uop_2_22_is_fencei;
  reg         rob_uop_2_22_uses_ldq;
  reg         rob_uop_2_22_uses_stq;
  reg         rob_uop_2_22_is_sys_pc2epc;
  reg         rob_uop_2_22_flush_on_commit;
  reg  [5:0]  rob_uop_2_22_ldst;
  reg         rob_uop_2_22_ldst_val;
  reg  [1:0]  rob_uop_2_22_dst_rtype;
  reg         rob_uop_2_22_fp_val;
  reg  [1:0]  rob_uop_2_22_debug_fsrc;
  reg  [6:0]  rob_uop_2_23_uopc;
  reg         rob_uop_2_23_is_rvc;
  reg         rob_uop_2_23_is_br;
  reg         rob_uop_2_23_is_jalr;
  reg         rob_uop_2_23_is_jal;
  reg  [19:0] rob_uop_2_23_br_mask;
  reg  [5:0]  rob_uop_2_23_ftq_idx;
  reg         rob_uop_2_23_edge_inst;
  reg  [5:0]  rob_uop_2_23_pc_lob;
  reg  [6:0]  rob_uop_2_23_pdst;
  reg  [6:0]  rob_uop_2_23_stale_pdst;
  reg         rob_uop_2_23_is_fencei;
  reg         rob_uop_2_23_uses_ldq;
  reg         rob_uop_2_23_uses_stq;
  reg         rob_uop_2_23_is_sys_pc2epc;
  reg         rob_uop_2_23_flush_on_commit;
  reg  [5:0]  rob_uop_2_23_ldst;
  reg         rob_uop_2_23_ldst_val;
  reg  [1:0]  rob_uop_2_23_dst_rtype;
  reg         rob_uop_2_23_fp_val;
  reg  [1:0]  rob_uop_2_23_debug_fsrc;
  reg  [6:0]  rob_uop_2_24_uopc;
  reg         rob_uop_2_24_is_rvc;
  reg         rob_uop_2_24_is_br;
  reg         rob_uop_2_24_is_jalr;
  reg         rob_uop_2_24_is_jal;
  reg  [19:0] rob_uop_2_24_br_mask;
  reg  [5:0]  rob_uop_2_24_ftq_idx;
  reg         rob_uop_2_24_edge_inst;
  reg  [5:0]  rob_uop_2_24_pc_lob;
  reg  [6:0]  rob_uop_2_24_pdst;
  reg  [6:0]  rob_uop_2_24_stale_pdst;
  reg         rob_uop_2_24_is_fencei;
  reg         rob_uop_2_24_uses_ldq;
  reg         rob_uop_2_24_uses_stq;
  reg         rob_uop_2_24_is_sys_pc2epc;
  reg         rob_uop_2_24_flush_on_commit;
  reg  [5:0]  rob_uop_2_24_ldst;
  reg         rob_uop_2_24_ldst_val;
  reg  [1:0]  rob_uop_2_24_dst_rtype;
  reg         rob_uop_2_24_fp_val;
  reg  [1:0]  rob_uop_2_24_debug_fsrc;
  reg  [6:0]  rob_uop_2_25_uopc;
  reg         rob_uop_2_25_is_rvc;
  reg         rob_uop_2_25_is_br;
  reg         rob_uop_2_25_is_jalr;
  reg         rob_uop_2_25_is_jal;
  reg  [19:0] rob_uop_2_25_br_mask;
  reg  [5:0]  rob_uop_2_25_ftq_idx;
  reg         rob_uop_2_25_edge_inst;
  reg  [5:0]  rob_uop_2_25_pc_lob;
  reg  [6:0]  rob_uop_2_25_pdst;
  reg  [6:0]  rob_uop_2_25_stale_pdst;
  reg         rob_uop_2_25_is_fencei;
  reg         rob_uop_2_25_uses_ldq;
  reg         rob_uop_2_25_uses_stq;
  reg         rob_uop_2_25_is_sys_pc2epc;
  reg         rob_uop_2_25_flush_on_commit;
  reg  [5:0]  rob_uop_2_25_ldst;
  reg         rob_uop_2_25_ldst_val;
  reg  [1:0]  rob_uop_2_25_dst_rtype;
  reg         rob_uop_2_25_fp_val;
  reg  [1:0]  rob_uop_2_25_debug_fsrc;
  reg  [6:0]  rob_uop_2_26_uopc;
  reg         rob_uop_2_26_is_rvc;
  reg         rob_uop_2_26_is_br;
  reg         rob_uop_2_26_is_jalr;
  reg         rob_uop_2_26_is_jal;
  reg  [19:0] rob_uop_2_26_br_mask;
  reg  [5:0]  rob_uop_2_26_ftq_idx;
  reg         rob_uop_2_26_edge_inst;
  reg  [5:0]  rob_uop_2_26_pc_lob;
  reg  [6:0]  rob_uop_2_26_pdst;
  reg  [6:0]  rob_uop_2_26_stale_pdst;
  reg         rob_uop_2_26_is_fencei;
  reg         rob_uop_2_26_uses_ldq;
  reg         rob_uop_2_26_uses_stq;
  reg         rob_uop_2_26_is_sys_pc2epc;
  reg         rob_uop_2_26_flush_on_commit;
  reg  [5:0]  rob_uop_2_26_ldst;
  reg         rob_uop_2_26_ldst_val;
  reg  [1:0]  rob_uop_2_26_dst_rtype;
  reg         rob_uop_2_26_fp_val;
  reg  [1:0]  rob_uop_2_26_debug_fsrc;
  reg  [6:0]  rob_uop_2_27_uopc;
  reg         rob_uop_2_27_is_rvc;
  reg         rob_uop_2_27_is_br;
  reg         rob_uop_2_27_is_jalr;
  reg         rob_uop_2_27_is_jal;
  reg  [19:0] rob_uop_2_27_br_mask;
  reg  [5:0]  rob_uop_2_27_ftq_idx;
  reg         rob_uop_2_27_edge_inst;
  reg  [5:0]  rob_uop_2_27_pc_lob;
  reg  [6:0]  rob_uop_2_27_pdst;
  reg  [6:0]  rob_uop_2_27_stale_pdst;
  reg         rob_uop_2_27_is_fencei;
  reg         rob_uop_2_27_uses_ldq;
  reg         rob_uop_2_27_uses_stq;
  reg         rob_uop_2_27_is_sys_pc2epc;
  reg         rob_uop_2_27_flush_on_commit;
  reg  [5:0]  rob_uop_2_27_ldst;
  reg         rob_uop_2_27_ldst_val;
  reg  [1:0]  rob_uop_2_27_dst_rtype;
  reg         rob_uop_2_27_fp_val;
  reg  [1:0]  rob_uop_2_27_debug_fsrc;
  reg  [6:0]  rob_uop_2_28_uopc;
  reg         rob_uop_2_28_is_rvc;
  reg         rob_uop_2_28_is_br;
  reg         rob_uop_2_28_is_jalr;
  reg         rob_uop_2_28_is_jal;
  reg  [19:0] rob_uop_2_28_br_mask;
  reg  [5:0]  rob_uop_2_28_ftq_idx;
  reg         rob_uop_2_28_edge_inst;
  reg  [5:0]  rob_uop_2_28_pc_lob;
  reg  [6:0]  rob_uop_2_28_pdst;
  reg  [6:0]  rob_uop_2_28_stale_pdst;
  reg         rob_uop_2_28_is_fencei;
  reg         rob_uop_2_28_uses_ldq;
  reg         rob_uop_2_28_uses_stq;
  reg         rob_uop_2_28_is_sys_pc2epc;
  reg         rob_uop_2_28_flush_on_commit;
  reg  [5:0]  rob_uop_2_28_ldst;
  reg         rob_uop_2_28_ldst_val;
  reg  [1:0]  rob_uop_2_28_dst_rtype;
  reg         rob_uop_2_28_fp_val;
  reg  [1:0]  rob_uop_2_28_debug_fsrc;
  reg  [6:0]  rob_uop_2_29_uopc;
  reg         rob_uop_2_29_is_rvc;
  reg         rob_uop_2_29_is_br;
  reg         rob_uop_2_29_is_jalr;
  reg         rob_uop_2_29_is_jal;
  reg  [19:0] rob_uop_2_29_br_mask;
  reg  [5:0]  rob_uop_2_29_ftq_idx;
  reg         rob_uop_2_29_edge_inst;
  reg  [5:0]  rob_uop_2_29_pc_lob;
  reg  [6:0]  rob_uop_2_29_pdst;
  reg  [6:0]  rob_uop_2_29_stale_pdst;
  reg         rob_uop_2_29_is_fencei;
  reg         rob_uop_2_29_uses_ldq;
  reg         rob_uop_2_29_uses_stq;
  reg         rob_uop_2_29_is_sys_pc2epc;
  reg         rob_uop_2_29_flush_on_commit;
  reg  [5:0]  rob_uop_2_29_ldst;
  reg         rob_uop_2_29_ldst_val;
  reg  [1:0]  rob_uop_2_29_dst_rtype;
  reg         rob_uop_2_29_fp_val;
  reg  [1:0]  rob_uop_2_29_debug_fsrc;
  reg  [6:0]  rob_uop_2_30_uopc;
  reg         rob_uop_2_30_is_rvc;
  reg         rob_uop_2_30_is_br;
  reg         rob_uop_2_30_is_jalr;
  reg         rob_uop_2_30_is_jal;
  reg  [19:0] rob_uop_2_30_br_mask;
  reg  [5:0]  rob_uop_2_30_ftq_idx;
  reg         rob_uop_2_30_edge_inst;
  reg  [5:0]  rob_uop_2_30_pc_lob;
  reg  [6:0]  rob_uop_2_30_pdst;
  reg  [6:0]  rob_uop_2_30_stale_pdst;
  reg         rob_uop_2_30_is_fencei;
  reg         rob_uop_2_30_uses_ldq;
  reg         rob_uop_2_30_uses_stq;
  reg         rob_uop_2_30_is_sys_pc2epc;
  reg         rob_uop_2_30_flush_on_commit;
  reg  [5:0]  rob_uop_2_30_ldst;
  reg         rob_uop_2_30_ldst_val;
  reg  [1:0]  rob_uop_2_30_dst_rtype;
  reg         rob_uop_2_30_fp_val;
  reg  [1:0]  rob_uop_2_30_debug_fsrc;
  reg  [6:0]  rob_uop_2_31_uopc;
  reg         rob_uop_2_31_is_rvc;
  reg         rob_uop_2_31_is_br;
  reg         rob_uop_2_31_is_jalr;
  reg         rob_uop_2_31_is_jal;
  reg  [19:0] rob_uop_2_31_br_mask;
  reg  [5:0]  rob_uop_2_31_ftq_idx;
  reg         rob_uop_2_31_edge_inst;
  reg  [5:0]  rob_uop_2_31_pc_lob;
  reg  [6:0]  rob_uop_2_31_pdst;
  reg  [6:0]  rob_uop_2_31_stale_pdst;
  reg         rob_uop_2_31_is_fencei;
  reg         rob_uop_2_31_uses_ldq;
  reg         rob_uop_2_31_uses_stq;
  reg         rob_uop_2_31_is_sys_pc2epc;
  reg         rob_uop_2_31_flush_on_commit;
  reg  [5:0]  rob_uop_2_31_ldst;
  reg         rob_uop_2_31_ldst_val;
  reg  [1:0]  rob_uop_2_31_dst_rtype;
  reg         rob_uop_2_31_fp_val;
  reg  [1:0]  rob_uop_2_31_debug_fsrc;
  reg         rob_exception_2_0;
  reg         rob_exception_2_1;
  reg         rob_exception_2_2;
  reg         rob_exception_2_3;
  reg         rob_exception_2_4;
  reg         rob_exception_2_5;
  reg         rob_exception_2_6;
  reg         rob_exception_2_7;
  reg         rob_exception_2_8;
  reg         rob_exception_2_9;
  reg         rob_exception_2_10;
  reg         rob_exception_2_11;
  reg         rob_exception_2_12;
  reg         rob_exception_2_13;
  reg         rob_exception_2_14;
  reg         rob_exception_2_15;
  reg         rob_exception_2_16;
  reg         rob_exception_2_17;
  reg         rob_exception_2_18;
  reg         rob_exception_2_19;
  reg         rob_exception_2_20;
  reg         rob_exception_2_21;
  reg         rob_exception_2_22;
  reg         rob_exception_2_23;
  reg         rob_exception_2_24;
  reg         rob_exception_2_25;
  reg         rob_exception_2_26;
  reg         rob_exception_2_27;
  reg         rob_exception_2_28;
  reg         rob_exception_2_29;
  reg         rob_exception_2_30;
  reg         rob_exception_2_31;
  reg         rob_predicated_2_0;
  reg         rob_predicated_2_1;
  reg         rob_predicated_2_2;
  reg         rob_predicated_2_3;
  reg         rob_predicated_2_4;
  reg         rob_predicated_2_5;
  reg         rob_predicated_2_6;
  reg         rob_predicated_2_7;
  reg         rob_predicated_2_8;
  reg         rob_predicated_2_9;
  reg         rob_predicated_2_10;
  reg         rob_predicated_2_11;
  reg         rob_predicated_2_12;
  reg         rob_predicated_2_13;
  reg         rob_predicated_2_14;
  reg         rob_predicated_2_15;
  reg         rob_predicated_2_16;
  reg         rob_predicated_2_17;
  reg         rob_predicated_2_18;
  reg         rob_predicated_2_19;
  reg         rob_predicated_2_20;
  reg         rob_predicated_2_21;
  reg         rob_predicated_2_22;
  reg         rob_predicated_2_23;
  reg         rob_predicated_2_24;
  reg         rob_predicated_2_25;
  reg         rob_predicated_2_26;
  reg         rob_predicated_2_27;
  reg         rob_predicated_2_28;
  reg         rob_predicated_2_29;
  reg         rob_predicated_2_30;
  reg         rob_predicated_2_31;
  reg         casez_tmp_155;
  always @(*) begin
    casez (rob_tail)
      5'b00000:
        casez_tmp_155 = rob_val_2_0;
      5'b00001:
        casez_tmp_155 = rob_val_2_1;
      5'b00010:
        casez_tmp_155 = rob_val_2_2;
      5'b00011:
        casez_tmp_155 = rob_val_2_3;
      5'b00100:
        casez_tmp_155 = rob_val_2_4;
      5'b00101:
        casez_tmp_155 = rob_val_2_5;
      5'b00110:
        casez_tmp_155 = rob_val_2_6;
      5'b00111:
        casez_tmp_155 = rob_val_2_7;
      5'b01000:
        casez_tmp_155 = rob_val_2_8;
      5'b01001:
        casez_tmp_155 = rob_val_2_9;
      5'b01010:
        casez_tmp_155 = rob_val_2_10;
      5'b01011:
        casez_tmp_155 = rob_val_2_11;
      5'b01100:
        casez_tmp_155 = rob_val_2_12;
      5'b01101:
        casez_tmp_155 = rob_val_2_13;
      5'b01110:
        casez_tmp_155 = rob_val_2_14;
      5'b01111:
        casez_tmp_155 = rob_val_2_15;
      5'b10000:
        casez_tmp_155 = rob_val_2_16;
      5'b10001:
        casez_tmp_155 = rob_val_2_17;
      5'b10010:
        casez_tmp_155 = rob_val_2_18;
      5'b10011:
        casez_tmp_155 = rob_val_2_19;
      5'b10100:
        casez_tmp_155 = rob_val_2_20;
      5'b10101:
        casez_tmp_155 = rob_val_2_21;
      5'b10110:
        casez_tmp_155 = rob_val_2_22;
      5'b10111:
        casez_tmp_155 = rob_val_2_23;
      5'b11000:
        casez_tmp_155 = rob_val_2_24;
      5'b11001:
        casez_tmp_155 = rob_val_2_25;
      5'b11010:
        casez_tmp_155 = rob_val_2_26;
      5'b11011:
        casez_tmp_155 = rob_val_2_27;
      5'b11100:
        casez_tmp_155 = rob_val_2_28;
      5'b11101:
        casez_tmp_155 = rob_val_2_29;
      5'b11110:
        casez_tmp_155 = rob_val_2_30;
      default:
        casez_tmp_155 = rob_val_2_31;
    endcase
  end // always @(*)
  wire        _GEN_33 = io_wb_resps_0_valid & io_wb_resps_0_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_34 = io_wb_resps_1_valid & io_wb_resps_1_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_35 = io_wb_resps_2_valid & io_wb_resps_2_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_36 = io_wb_resps_3_valid & io_wb_resps_3_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_37 = io_wb_resps_4_valid & io_wb_resps_4_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_38 = io_wb_resps_5_valid & io_wb_resps_5_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_39 = io_wb_resps_6_valid & io_wb_resps_6_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_40 = io_wb_resps_7_valid & io_wb_resps_7_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_41 = io_wb_resps_8_valid & io_wb_resps_8_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_42 = io_wb_resps_9_valid & io_wb_resps_9_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_43 = io_lsu_clr_bsy_0_valid & io_lsu_clr_bsy_0_bits[1:0] == 2'h2;
  reg         casez_tmp_156;
  always @(*) begin
    casez (io_lsu_clr_bsy_0_bits[6:2])
      5'b00000:
        casez_tmp_156 = rob_val_2_0;
      5'b00001:
        casez_tmp_156 = rob_val_2_1;
      5'b00010:
        casez_tmp_156 = rob_val_2_2;
      5'b00011:
        casez_tmp_156 = rob_val_2_3;
      5'b00100:
        casez_tmp_156 = rob_val_2_4;
      5'b00101:
        casez_tmp_156 = rob_val_2_5;
      5'b00110:
        casez_tmp_156 = rob_val_2_6;
      5'b00111:
        casez_tmp_156 = rob_val_2_7;
      5'b01000:
        casez_tmp_156 = rob_val_2_8;
      5'b01001:
        casez_tmp_156 = rob_val_2_9;
      5'b01010:
        casez_tmp_156 = rob_val_2_10;
      5'b01011:
        casez_tmp_156 = rob_val_2_11;
      5'b01100:
        casez_tmp_156 = rob_val_2_12;
      5'b01101:
        casez_tmp_156 = rob_val_2_13;
      5'b01110:
        casez_tmp_156 = rob_val_2_14;
      5'b01111:
        casez_tmp_156 = rob_val_2_15;
      5'b10000:
        casez_tmp_156 = rob_val_2_16;
      5'b10001:
        casez_tmp_156 = rob_val_2_17;
      5'b10010:
        casez_tmp_156 = rob_val_2_18;
      5'b10011:
        casez_tmp_156 = rob_val_2_19;
      5'b10100:
        casez_tmp_156 = rob_val_2_20;
      5'b10101:
        casez_tmp_156 = rob_val_2_21;
      5'b10110:
        casez_tmp_156 = rob_val_2_22;
      5'b10111:
        casez_tmp_156 = rob_val_2_23;
      5'b11000:
        casez_tmp_156 = rob_val_2_24;
      5'b11001:
        casez_tmp_156 = rob_val_2_25;
      5'b11010:
        casez_tmp_156 = rob_val_2_26;
      5'b11011:
        casez_tmp_156 = rob_val_2_27;
      5'b11100:
        casez_tmp_156 = rob_val_2_28;
      5'b11101:
        casez_tmp_156 = rob_val_2_29;
      5'b11110:
        casez_tmp_156 = rob_val_2_30;
      default:
        casez_tmp_156 = rob_val_2_31;
    endcase
  end // always @(*)
  reg         casez_tmp_157;
  always @(*) begin
    casez (io_lsu_clr_bsy_0_bits[6:2])
      5'b00000:
        casez_tmp_157 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_157 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_157 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_157 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_157 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_157 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_157 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_157 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_157 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_157 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_157 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_157 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_157 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_157 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_157 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_157 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_157 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_157 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_157 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_157 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_157 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_157 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_157 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_157 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_157 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_157 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_157 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_157 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_157 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_157 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_157 = rob_bsy_2_30;
      default:
        casez_tmp_157 = rob_bsy_2_31;
    endcase
  end // always @(*)
  wire        _GEN_44 = io_lsu_clr_bsy_1_valid & io_lsu_clr_bsy_1_bits[1:0] == 2'h2;
  reg         casez_tmp_158;
  always @(*) begin
    casez (io_lsu_clr_bsy_1_bits[6:2])
      5'b00000:
        casez_tmp_158 = rob_val_2_0;
      5'b00001:
        casez_tmp_158 = rob_val_2_1;
      5'b00010:
        casez_tmp_158 = rob_val_2_2;
      5'b00011:
        casez_tmp_158 = rob_val_2_3;
      5'b00100:
        casez_tmp_158 = rob_val_2_4;
      5'b00101:
        casez_tmp_158 = rob_val_2_5;
      5'b00110:
        casez_tmp_158 = rob_val_2_6;
      5'b00111:
        casez_tmp_158 = rob_val_2_7;
      5'b01000:
        casez_tmp_158 = rob_val_2_8;
      5'b01001:
        casez_tmp_158 = rob_val_2_9;
      5'b01010:
        casez_tmp_158 = rob_val_2_10;
      5'b01011:
        casez_tmp_158 = rob_val_2_11;
      5'b01100:
        casez_tmp_158 = rob_val_2_12;
      5'b01101:
        casez_tmp_158 = rob_val_2_13;
      5'b01110:
        casez_tmp_158 = rob_val_2_14;
      5'b01111:
        casez_tmp_158 = rob_val_2_15;
      5'b10000:
        casez_tmp_158 = rob_val_2_16;
      5'b10001:
        casez_tmp_158 = rob_val_2_17;
      5'b10010:
        casez_tmp_158 = rob_val_2_18;
      5'b10011:
        casez_tmp_158 = rob_val_2_19;
      5'b10100:
        casez_tmp_158 = rob_val_2_20;
      5'b10101:
        casez_tmp_158 = rob_val_2_21;
      5'b10110:
        casez_tmp_158 = rob_val_2_22;
      5'b10111:
        casez_tmp_158 = rob_val_2_23;
      5'b11000:
        casez_tmp_158 = rob_val_2_24;
      5'b11001:
        casez_tmp_158 = rob_val_2_25;
      5'b11010:
        casez_tmp_158 = rob_val_2_26;
      5'b11011:
        casez_tmp_158 = rob_val_2_27;
      5'b11100:
        casez_tmp_158 = rob_val_2_28;
      5'b11101:
        casez_tmp_158 = rob_val_2_29;
      5'b11110:
        casez_tmp_158 = rob_val_2_30;
      default:
        casez_tmp_158 = rob_val_2_31;
    endcase
  end // always @(*)
  reg         casez_tmp_159;
  always @(*) begin
    casez (io_lsu_clr_bsy_1_bits[6:2])
      5'b00000:
        casez_tmp_159 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_159 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_159 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_159 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_159 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_159 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_159 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_159 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_159 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_159 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_159 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_159 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_159 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_159 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_159 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_159 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_159 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_159 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_159 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_159 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_159 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_159 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_159 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_159 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_159 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_159 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_159 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_159 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_159 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_159 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_159 = rob_bsy_2_30;
      default:
        casez_tmp_159 = rob_bsy_2_31;
    endcase
  end // always @(*)
  wire        _GEN_45 = io_lsu_clr_bsy_2_valid & io_lsu_clr_bsy_2_bits[1:0] == 2'h2;
  reg         casez_tmp_160;
  always @(*) begin
    casez (io_lsu_clr_bsy_2_bits[6:2])
      5'b00000:
        casez_tmp_160 = rob_val_2_0;
      5'b00001:
        casez_tmp_160 = rob_val_2_1;
      5'b00010:
        casez_tmp_160 = rob_val_2_2;
      5'b00011:
        casez_tmp_160 = rob_val_2_3;
      5'b00100:
        casez_tmp_160 = rob_val_2_4;
      5'b00101:
        casez_tmp_160 = rob_val_2_5;
      5'b00110:
        casez_tmp_160 = rob_val_2_6;
      5'b00111:
        casez_tmp_160 = rob_val_2_7;
      5'b01000:
        casez_tmp_160 = rob_val_2_8;
      5'b01001:
        casez_tmp_160 = rob_val_2_9;
      5'b01010:
        casez_tmp_160 = rob_val_2_10;
      5'b01011:
        casez_tmp_160 = rob_val_2_11;
      5'b01100:
        casez_tmp_160 = rob_val_2_12;
      5'b01101:
        casez_tmp_160 = rob_val_2_13;
      5'b01110:
        casez_tmp_160 = rob_val_2_14;
      5'b01111:
        casez_tmp_160 = rob_val_2_15;
      5'b10000:
        casez_tmp_160 = rob_val_2_16;
      5'b10001:
        casez_tmp_160 = rob_val_2_17;
      5'b10010:
        casez_tmp_160 = rob_val_2_18;
      5'b10011:
        casez_tmp_160 = rob_val_2_19;
      5'b10100:
        casez_tmp_160 = rob_val_2_20;
      5'b10101:
        casez_tmp_160 = rob_val_2_21;
      5'b10110:
        casez_tmp_160 = rob_val_2_22;
      5'b10111:
        casez_tmp_160 = rob_val_2_23;
      5'b11000:
        casez_tmp_160 = rob_val_2_24;
      5'b11001:
        casez_tmp_160 = rob_val_2_25;
      5'b11010:
        casez_tmp_160 = rob_val_2_26;
      5'b11011:
        casez_tmp_160 = rob_val_2_27;
      5'b11100:
        casez_tmp_160 = rob_val_2_28;
      5'b11101:
        casez_tmp_160 = rob_val_2_29;
      5'b11110:
        casez_tmp_160 = rob_val_2_30;
      default:
        casez_tmp_160 = rob_val_2_31;
    endcase
  end // always @(*)
  reg         casez_tmp_161;
  always @(*) begin
    casez (io_lsu_clr_bsy_2_bits[6:2])
      5'b00000:
        casez_tmp_161 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_161 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_161 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_161 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_161 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_161 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_161 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_161 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_161 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_161 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_161 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_161 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_161 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_161 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_161 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_161 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_161 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_161 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_161 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_161 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_161 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_161 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_161 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_161 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_161 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_161 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_161 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_161 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_161 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_161 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_161 = rob_bsy_2_30;
      default:
        casez_tmp_161 = rob_bsy_2_31;
    endcase
  end // always @(*)
  wire        _GEN_46 = io_lxcpt_valid & io_lxcpt_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_47 = _GEN_46 & _GEN_13 & ~reset;
  reg         casez_tmp_162;
  always @(*) begin
    casez (io_lxcpt_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_162 = rob_unsafe_2_0;
      5'b00001:
        casez_tmp_162 = rob_unsafe_2_1;
      5'b00010:
        casez_tmp_162 = rob_unsafe_2_2;
      5'b00011:
        casez_tmp_162 = rob_unsafe_2_3;
      5'b00100:
        casez_tmp_162 = rob_unsafe_2_4;
      5'b00101:
        casez_tmp_162 = rob_unsafe_2_5;
      5'b00110:
        casez_tmp_162 = rob_unsafe_2_6;
      5'b00111:
        casez_tmp_162 = rob_unsafe_2_7;
      5'b01000:
        casez_tmp_162 = rob_unsafe_2_8;
      5'b01001:
        casez_tmp_162 = rob_unsafe_2_9;
      5'b01010:
        casez_tmp_162 = rob_unsafe_2_10;
      5'b01011:
        casez_tmp_162 = rob_unsafe_2_11;
      5'b01100:
        casez_tmp_162 = rob_unsafe_2_12;
      5'b01101:
        casez_tmp_162 = rob_unsafe_2_13;
      5'b01110:
        casez_tmp_162 = rob_unsafe_2_14;
      5'b01111:
        casez_tmp_162 = rob_unsafe_2_15;
      5'b10000:
        casez_tmp_162 = rob_unsafe_2_16;
      5'b10001:
        casez_tmp_162 = rob_unsafe_2_17;
      5'b10010:
        casez_tmp_162 = rob_unsafe_2_18;
      5'b10011:
        casez_tmp_162 = rob_unsafe_2_19;
      5'b10100:
        casez_tmp_162 = rob_unsafe_2_20;
      5'b10101:
        casez_tmp_162 = rob_unsafe_2_21;
      5'b10110:
        casez_tmp_162 = rob_unsafe_2_22;
      5'b10111:
        casez_tmp_162 = rob_unsafe_2_23;
      5'b11000:
        casez_tmp_162 = rob_unsafe_2_24;
      5'b11001:
        casez_tmp_162 = rob_unsafe_2_25;
      5'b11010:
        casez_tmp_162 = rob_unsafe_2_26;
      5'b11011:
        casez_tmp_162 = rob_unsafe_2_27;
      5'b11100:
        casez_tmp_162 = rob_unsafe_2_28;
      5'b11101:
        casez_tmp_162 = rob_unsafe_2_29;
      5'b11110:
        casez_tmp_162 = rob_unsafe_2_30;
      default:
        casez_tmp_162 = rob_unsafe_2_31;
    endcase
  end // always @(*)
  reg         casez_tmp_163;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_163 = rob_val_2_0;
      5'b00001:
        casez_tmp_163 = rob_val_2_1;
      5'b00010:
        casez_tmp_163 = rob_val_2_2;
      5'b00011:
        casez_tmp_163 = rob_val_2_3;
      5'b00100:
        casez_tmp_163 = rob_val_2_4;
      5'b00101:
        casez_tmp_163 = rob_val_2_5;
      5'b00110:
        casez_tmp_163 = rob_val_2_6;
      5'b00111:
        casez_tmp_163 = rob_val_2_7;
      5'b01000:
        casez_tmp_163 = rob_val_2_8;
      5'b01001:
        casez_tmp_163 = rob_val_2_9;
      5'b01010:
        casez_tmp_163 = rob_val_2_10;
      5'b01011:
        casez_tmp_163 = rob_val_2_11;
      5'b01100:
        casez_tmp_163 = rob_val_2_12;
      5'b01101:
        casez_tmp_163 = rob_val_2_13;
      5'b01110:
        casez_tmp_163 = rob_val_2_14;
      5'b01111:
        casez_tmp_163 = rob_val_2_15;
      5'b10000:
        casez_tmp_163 = rob_val_2_16;
      5'b10001:
        casez_tmp_163 = rob_val_2_17;
      5'b10010:
        casez_tmp_163 = rob_val_2_18;
      5'b10011:
        casez_tmp_163 = rob_val_2_19;
      5'b10100:
        casez_tmp_163 = rob_val_2_20;
      5'b10101:
        casez_tmp_163 = rob_val_2_21;
      5'b10110:
        casez_tmp_163 = rob_val_2_22;
      5'b10111:
        casez_tmp_163 = rob_val_2_23;
      5'b11000:
        casez_tmp_163 = rob_val_2_24;
      5'b11001:
        casez_tmp_163 = rob_val_2_25;
      5'b11010:
        casez_tmp_163 = rob_val_2_26;
      5'b11011:
        casez_tmp_163 = rob_val_2_27;
      5'b11100:
        casez_tmp_163 = rob_val_2_28;
      5'b11101:
        casez_tmp_163 = rob_val_2_29;
      5'b11110:
        casez_tmp_163 = rob_val_2_30;
      default:
        casez_tmp_163 = rob_val_2_31;
    endcase
  end // always @(*)
  reg         casez_tmp_164;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_164 = rob_exception_2_0;
      5'b00001:
        casez_tmp_164 = rob_exception_2_1;
      5'b00010:
        casez_tmp_164 = rob_exception_2_2;
      5'b00011:
        casez_tmp_164 = rob_exception_2_3;
      5'b00100:
        casez_tmp_164 = rob_exception_2_4;
      5'b00101:
        casez_tmp_164 = rob_exception_2_5;
      5'b00110:
        casez_tmp_164 = rob_exception_2_6;
      5'b00111:
        casez_tmp_164 = rob_exception_2_7;
      5'b01000:
        casez_tmp_164 = rob_exception_2_8;
      5'b01001:
        casez_tmp_164 = rob_exception_2_9;
      5'b01010:
        casez_tmp_164 = rob_exception_2_10;
      5'b01011:
        casez_tmp_164 = rob_exception_2_11;
      5'b01100:
        casez_tmp_164 = rob_exception_2_12;
      5'b01101:
        casez_tmp_164 = rob_exception_2_13;
      5'b01110:
        casez_tmp_164 = rob_exception_2_14;
      5'b01111:
        casez_tmp_164 = rob_exception_2_15;
      5'b10000:
        casez_tmp_164 = rob_exception_2_16;
      5'b10001:
        casez_tmp_164 = rob_exception_2_17;
      5'b10010:
        casez_tmp_164 = rob_exception_2_18;
      5'b10011:
        casez_tmp_164 = rob_exception_2_19;
      5'b10100:
        casez_tmp_164 = rob_exception_2_20;
      5'b10101:
        casez_tmp_164 = rob_exception_2_21;
      5'b10110:
        casez_tmp_164 = rob_exception_2_22;
      5'b10111:
        casez_tmp_164 = rob_exception_2_23;
      5'b11000:
        casez_tmp_164 = rob_exception_2_24;
      5'b11001:
        casez_tmp_164 = rob_exception_2_25;
      5'b11010:
        casez_tmp_164 = rob_exception_2_26;
      5'b11011:
        casez_tmp_164 = rob_exception_2_27;
      5'b11100:
        casez_tmp_164 = rob_exception_2_28;
      5'b11101:
        casez_tmp_164 = rob_exception_2_29;
      5'b11110:
        casez_tmp_164 = rob_exception_2_30;
      default:
        casez_tmp_164 = rob_exception_2_31;
    endcase
  end // always @(*)
  wire        can_throw_exception_2 = casez_tmp_163 & casez_tmp_164;
  reg         casez_tmp_165;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_165 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_165 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_165 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_165 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_165 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_165 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_165 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_165 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_165 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_165 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_165 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_165 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_165 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_165 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_165 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_165 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_165 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_165 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_165 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_165 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_165 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_165 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_165 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_165 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_165 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_165 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_165 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_165 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_165 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_165 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_165 = rob_bsy_2_30;
      default:
        casez_tmp_165 = rob_bsy_2_31;
    endcase
  end // always @(*)
  wire        can_commit_2 = casez_tmp_163 & ~casez_tmp_165 & ~io_csr_stall;
  reg         casez_tmp_166;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_166 = rob_predicated_2_0;
      5'b00001:
        casez_tmp_166 = rob_predicated_2_1;
      5'b00010:
        casez_tmp_166 = rob_predicated_2_2;
      5'b00011:
        casez_tmp_166 = rob_predicated_2_3;
      5'b00100:
        casez_tmp_166 = rob_predicated_2_4;
      5'b00101:
        casez_tmp_166 = rob_predicated_2_5;
      5'b00110:
        casez_tmp_166 = rob_predicated_2_6;
      5'b00111:
        casez_tmp_166 = rob_predicated_2_7;
      5'b01000:
        casez_tmp_166 = rob_predicated_2_8;
      5'b01001:
        casez_tmp_166 = rob_predicated_2_9;
      5'b01010:
        casez_tmp_166 = rob_predicated_2_10;
      5'b01011:
        casez_tmp_166 = rob_predicated_2_11;
      5'b01100:
        casez_tmp_166 = rob_predicated_2_12;
      5'b01101:
        casez_tmp_166 = rob_predicated_2_13;
      5'b01110:
        casez_tmp_166 = rob_predicated_2_14;
      5'b01111:
        casez_tmp_166 = rob_predicated_2_15;
      5'b10000:
        casez_tmp_166 = rob_predicated_2_16;
      5'b10001:
        casez_tmp_166 = rob_predicated_2_17;
      5'b10010:
        casez_tmp_166 = rob_predicated_2_18;
      5'b10011:
        casez_tmp_166 = rob_predicated_2_19;
      5'b10100:
        casez_tmp_166 = rob_predicated_2_20;
      5'b10101:
        casez_tmp_166 = rob_predicated_2_21;
      5'b10110:
        casez_tmp_166 = rob_predicated_2_22;
      5'b10111:
        casez_tmp_166 = rob_predicated_2_23;
      5'b11000:
        casez_tmp_166 = rob_predicated_2_24;
      5'b11001:
        casez_tmp_166 = rob_predicated_2_25;
      5'b11010:
        casez_tmp_166 = rob_predicated_2_26;
      5'b11011:
        casez_tmp_166 = rob_predicated_2_27;
      5'b11100:
        casez_tmp_166 = rob_predicated_2_28;
      5'b11101:
        casez_tmp_166 = rob_predicated_2_29;
      5'b11110:
        casez_tmp_166 = rob_predicated_2_30;
      default:
        casez_tmp_166 = rob_predicated_2_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_167;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_167 = rob_uop_2_0_uopc;
      5'b00001:
        casez_tmp_167 = rob_uop_2_1_uopc;
      5'b00010:
        casez_tmp_167 = rob_uop_2_2_uopc;
      5'b00011:
        casez_tmp_167 = rob_uop_2_3_uopc;
      5'b00100:
        casez_tmp_167 = rob_uop_2_4_uopc;
      5'b00101:
        casez_tmp_167 = rob_uop_2_5_uopc;
      5'b00110:
        casez_tmp_167 = rob_uop_2_6_uopc;
      5'b00111:
        casez_tmp_167 = rob_uop_2_7_uopc;
      5'b01000:
        casez_tmp_167 = rob_uop_2_8_uopc;
      5'b01001:
        casez_tmp_167 = rob_uop_2_9_uopc;
      5'b01010:
        casez_tmp_167 = rob_uop_2_10_uopc;
      5'b01011:
        casez_tmp_167 = rob_uop_2_11_uopc;
      5'b01100:
        casez_tmp_167 = rob_uop_2_12_uopc;
      5'b01101:
        casez_tmp_167 = rob_uop_2_13_uopc;
      5'b01110:
        casez_tmp_167 = rob_uop_2_14_uopc;
      5'b01111:
        casez_tmp_167 = rob_uop_2_15_uopc;
      5'b10000:
        casez_tmp_167 = rob_uop_2_16_uopc;
      5'b10001:
        casez_tmp_167 = rob_uop_2_17_uopc;
      5'b10010:
        casez_tmp_167 = rob_uop_2_18_uopc;
      5'b10011:
        casez_tmp_167 = rob_uop_2_19_uopc;
      5'b10100:
        casez_tmp_167 = rob_uop_2_20_uopc;
      5'b10101:
        casez_tmp_167 = rob_uop_2_21_uopc;
      5'b10110:
        casez_tmp_167 = rob_uop_2_22_uopc;
      5'b10111:
        casez_tmp_167 = rob_uop_2_23_uopc;
      5'b11000:
        casez_tmp_167 = rob_uop_2_24_uopc;
      5'b11001:
        casez_tmp_167 = rob_uop_2_25_uopc;
      5'b11010:
        casez_tmp_167 = rob_uop_2_26_uopc;
      5'b11011:
        casez_tmp_167 = rob_uop_2_27_uopc;
      5'b11100:
        casez_tmp_167 = rob_uop_2_28_uopc;
      5'b11101:
        casez_tmp_167 = rob_uop_2_29_uopc;
      5'b11110:
        casez_tmp_167 = rob_uop_2_30_uopc;
      default:
        casez_tmp_167 = rob_uop_2_31_uopc;
    endcase
  end // always @(*)
  reg         casez_tmp_168;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_168 = rob_uop_2_0_is_rvc;
      5'b00001:
        casez_tmp_168 = rob_uop_2_1_is_rvc;
      5'b00010:
        casez_tmp_168 = rob_uop_2_2_is_rvc;
      5'b00011:
        casez_tmp_168 = rob_uop_2_3_is_rvc;
      5'b00100:
        casez_tmp_168 = rob_uop_2_4_is_rvc;
      5'b00101:
        casez_tmp_168 = rob_uop_2_5_is_rvc;
      5'b00110:
        casez_tmp_168 = rob_uop_2_6_is_rvc;
      5'b00111:
        casez_tmp_168 = rob_uop_2_7_is_rvc;
      5'b01000:
        casez_tmp_168 = rob_uop_2_8_is_rvc;
      5'b01001:
        casez_tmp_168 = rob_uop_2_9_is_rvc;
      5'b01010:
        casez_tmp_168 = rob_uop_2_10_is_rvc;
      5'b01011:
        casez_tmp_168 = rob_uop_2_11_is_rvc;
      5'b01100:
        casez_tmp_168 = rob_uop_2_12_is_rvc;
      5'b01101:
        casez_tmp_168 = rob_uop_2_13_is_rvc;
      5'b01110:
        casez_tmp_168 = rob_uop_2_14_is_rvc;
      5'b01111:
        casez_tmp_168 = rob_uop_2_15_is_rvc;
      5'b10000:
        casez_tmp_168 = rob_uop_2_16_is_rvc;
      5'b10001:
        casez_tmp_168 = rob_uop_2_17_is_rvc;
      5'b10010:
        casez_tmp_168 = rob_uop_2_18_is_rvc;
      5'b10011:
        casez_tmp_168 = rob_uop_2_19_is_rvc;
      5'b10100:
        casez_tmp_168 = rob_uop_2_20_is_rvc;
      5'b10101:
        casez_tmp_168 = rob_uop_2_21_is_rvc;
      5'b10110:
        casez_tmp_168 = rob_uop_2_22_is_rvc;
      5'b10111:
        casez_tmp_168 = rob_uop_2_23_is_rvc;
      5'b11000:
        casez_tmp_168 = rob_uop_2_24_is_rvc;
      5'b11001:
        casez_tmp_168 = rob_uop_2_25_is_rvc;
      5'b11010:
        casez_tmp_168 = rob_uop_2_26_is_rvc;
      5'b11011:
        casez_tmp_168 = rob_uop_2_27_is_rvc;
      5'b11100:
        casez_tmp_168 = rob_uop_2_28_is_rvc;
      5'b11101:
        casez_tmp_168 = rob_uop_2_29_is_rvc;
      5'b11110:
        casez_tmp_168 = rob_uop_2_30_is_rvc;
      default:
        casez_tmp_168 = rob_uop_2_31_is_rvc;
    endcase
  end // always @(*)
  reg         casez_tmp_169;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_169 = rob_uop_2_0_is_br;
      5'b00001:
        casez_tmp_169 = rob_uop_2_1_is_br;
      5'b00010:
        casez_tmp_169 = rob_uop_2_2_is_br;
      5'b00011:
        casez_tmp_169 = rob_uop_2_3_is_br;
      5'b00100:
        casez_tmp_169 = rob_uop_2_4_is_br;
      5'b00101:
        casez_tmp_169 = rob_uop_2_5_is_br;
      5'b00110:
        casez_tmp_169 = rob_uop_2_6_is_br;
      5'b00111:
        casez_tmp_169 = rob_uop_2_7_is_br;
      5'b01000:
        casez_tmp_169 = rob_uop_2_8_is_br;
      5'b01001:
        casez_tmp_169 = rob_uop_2_9_is_br;
      5'b01010:
        casez_tmp_169 = rob_uop_2_10_is_br;
      5'b01011:
        casez_tmp_169 = rob_uop_2_11_is_br;
      5'b01100:
        casez_tmp_169 = rob_uop_2_12_is_br;
      5'b01101:
        casez_tmp_169 = rob_uop_2_13_is_br;
      5'b01110:
        casez_tmp_169 = rob_uop_2_14_is_br;
      5'b01111:
        casez_tmp_169 = rob_uop_2_15_is_br;
      5'b10000:
        casez_tmp_169 = rob_uop_2_16_is_br;
      5'b10001:
        casez_tmp_169 = rob_uop_2_17_is_br;
      5'b10010:
        casez_tmp_169 = rob_uop_2_18_is_br;
      5'b10011:
        casez_tmp_169 = rob_uop_2_19_is_br;
      5'b10100:
        casez_tmp_169 = rob_uop_2_20_is_br;
      5'b10101:
        casez_tmp_169 = rob_uop_2_21_is_br;
      5'b10110:
        casez_tmp_169 = rob_uop_2_22_is_br;
      5'b10111:
        casez_tmp_169 = rob_uop_2_23_is_br;
      5'b11000:
        casez_tmp_169 = rob_uop_2_24_is_br;
      5'b11001:
        casez_tmp_169 = rob_uop_2_25_is_br;
      5'b11010:
        casez_tmp_169 = rob_uop_2_26_is_br;
      5'b11011:
        casez_tmp_169 = rob_uop_2_27_is_br;
      5'b11100:
        casez_tmp_169 = rob_uop_2_28_is_br;
      5'b11101:
        casez_tmp_169 = rob_uop_2_29_is_br;
      5'b11110:
        casez_tmp_169 = rob_uop_2_30_is_br;
      default:
        casez_tmp_169 = rob_uop_2_31_is_br;
    endcase
  end // always @(*)
  reg         casez_tmp_170;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_170 = rob_uop_2_0_is_jalr;
      5'b00001:
        casez_tmp_170 = rob_uop_2_1_is_jalr;
      5'b00010:
        casez_tmp_170 = rob_uop_2_2_is_jalr;
      5'b00011:
        casez_tmp_170 = rob_uop_2_3_is_jalr;
      5'b00100:
        casez_tmp_170 = rob_uop_2_4_is_jalr;
      5'b00101:
        casez_tmp_170 = rob_uop_2_5_is_jalr;
      5'b00110:
        casez_tmp_170 = rob_uop_2_6_is_jalr;
      5'b00111:
        casez_tmp_170 = rob_uop_2_7_is_jalr;
      5'b01000:
        casez_tmp_170 = rob_uop_2_8_is_jalr;
      5'b01001:
        casez_tmp_170 = rob_uop_2_9_is_jalr;
      5'b01010:
        casez_tmp_170 = rob_uop_2_10_is_jalr;
      5'b01011:
        casez_tmp_170 = rob_uop_2_11_is_jalr;
      5'b01100:
        casez_tmp_170 = rob_uop_2_12_is_jalr;
      5'b01101:
        casez_tmp_170 = rob_uop_2_13_is_jalr;
      5'b01110:
        casez_tmp_170 = rob_uop_2_14_is_jalr;
      5'b01111:
        casez_tmp_170 = rob_uop_2_15_is_jalr;
      5'b10000:
        casez_tmp_170 = rob_uop_2_16_is_jalr;
      5'b10001:
        casez_tmp_170 = rob_uop_2_17_is_jalr;
      5'b10010:
        casez_tmp_170 = rob_uop_2_18_is_jalr;
      5'b10011:
        casez_tmp_170 = rob_uop_2_19_is_jalr;
      5'b10100:
        casez_tmp_170 = rob_uop_2_20_is_jalr;
      5'b10101:
        casez_tmp_170 = rob_uop_2_21_is_jalr;
      5'b10110:
        casez_tmp_170 = rob_uop_2_22_is_jalr;
      5'b10111:
        casez_tmp_170 = rob_uop_2_23_is_jalr;
      5'b11000:
        casez_tmp_170 = rob_uop_2_24_is_jalr;
      5'b11001:
        casez_tmp_170 = rob_uop_2_25_is_jalr;
      5'b11010:
        casez_tmp_170 = rob_uop_2_26_is_jalr;
      5'b11011:
        casez_tmp_170 = rob_uop_2_27_is_jalr;
      5'b11100:
        casez_tmp_170 = rob_uop_2_28_is_jalr;
      5'b11101:
        casez_tmp_170 = rob_uop_2_29_is_jalr;
      5'b11110:
        casez_tmp_170 = rob_uop_2_30_is_jalr;
      default:
        casez_tmp_170 = rob_uop_2_31_is_jalr;
    endcase
  end // always @(*)
  reg         casez_tmp_171;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_171 = rob_uop_2_0_is_jal;
      5'b00001:
        casez_tmp_171 = rob_uop_2_1_is_jal;
      5'b00010:
        casez_tmp_171 = rob_uop_2_2_is_jal;
      5'b00011:
        casez_tmp_171 = rob_uop_2_3_is_jal;
      5'b00100:
        casez_tmp_171 = rob_uop_2_4_is_jal;
      5'b00101:
        casez_tmp_171 = rob_uop_2_5_is_jal;
      5'b00110:
        casez_tmp_171 = rob_uop_2_6_is_jal;
      5'b00111:
        casez_tmp_171 = rob_uop_2_7_is_jal;
      5'b01000:
        casez_tmp_171 = rob_uop_2_8_is_jal;
      5'b01001:
        casez_tmp_171 = rob_uop_2_9_is_jal;
      5'b01010:
        casez_tmp_171 = rob_uop_2_10_is_jal;
      5'b01011:
        casez_tmp_171 = rob_uop_2_11_is_jal;
      5'b01100:
        casez_tmp_171 = rob_uop_2_12_is_jal;
      5'b01101:
        casez_tmp_171 = rob_uop_2_13_is_jal;
      5'b01110:
        casez_tmp_171 = rob_uop_2_14_is_jal;
      5'b01111:
        casez_tmp_171 = rob_uop_2_15_is_jal;
      5'b10000:
        casez_tmp_171 = rob_uop_2_16_is_jal;
      5'b10001:
        casez_tmp_171 = rob_uop_2_17_is_jal;
      5'b10010:
        casez_tmp_171 = rob_uop_2_18_is_jal;
      5'b10011:
        casez_tmp_171 = rob_uop_2_19_is_jal;
      5'b10100:
        casez_tmp_171 = rob_uop_2_20_is_jal;
      5'b10101:
        casez_tmp_171 = rob_uop_2_21_is_jal;
      5'b10110:
        casez_tmp_171 = rob_uop_2_22_is_jal;
      5'b10111:
        casez_tmp_171 = rob_uop_2_23_is_jal;
      5'b11000:
        casez_tmp_171 = rob_uop_2_24_is_jal;
      5'b11001:
        casez_tmp_171 = rob_uop_2_25_is_jal;
      5'b11010:
        casez_tmp_171 = rob_uop_2_26_is_jal;
      5'b11011:
        casez_tmp_171 = rob_uop_2_27_is_jal;
      5'b11100:
        casez_tmp_171 = rob_uop_2_28_is_jal;
      5'b11101:
        casez_tmp_171 = rob_uop_2_29_is_jal;
      5'b11110:
        casez_tmp_171 = rob_uop_2_30_is_jal;
      default:
        casez_tmp_171 = rob_uop_2_31_is_jal;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_172;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_172 = rob_uop_2_0_ftq_idx;
      5'b00001:
        casez_tmp_172 = rob_uop_2_1_ftq_idx;
      5'b00010:
        casez_tmp_172 = rob_uop_2_2_ftq_idx;
      5'b00011:
        casez_tmp_172 = rob_uop_2_3_ftq_idx;
      5'b00100:
        casez_tmp_172 = rob_uop_2_4_ftq_idx;
      5'b00101:
        casez_tmp_172 = rob_uop_2_5_ftq_idx;
      5'b00110:
        casez_tmp_172 = rob_uop_2_6_ftq_idx;
      5'b00111:
        casez_tmp_172 = rob_uop_2_7_ftq_idx;
      5'b01000:
        casez_tmp_172 = rob_uop_2_8_ftq_idx;
      5'b01001:
        casez_tmp_172 = rob_uop_2_9_ftq_idx;
      5'b01010:
        casez_tmp_172 = rob_uop_2_10_ftq_idx;
      5'b01011:
        casez_tmp_172 = rob_uop_2_11_ftq_idx;
      5'b01100:
        casez_tmp_172 = rob_uop_2_12_ftq_idx;
      5'b01101:
        casez_tmp_172 = rob_uop_2_13_ftq_idx;
      5'b01110:
        casez_tmp_172 = rob_uop_2_14_ftq_idx;
      5'b01111:
        casez_tmp_172 = rob_uop_2_15_ftq_idx;
      5'b10000:
        casez_tmp_172 = rob_uop_2_16_ftq_idx;
      5'b10001:
        casez_tmp_172 = rob_uop_2_17_ftq_idx;
      5'b10010:
        casez_tmp_172 = rob_uop_2_18_ftq_idx;
      5'b10011:
        casez_tmp_172 = rob_uop_2_19_ftq_idx;
      5'b10100:
        casez_tmp_172 = rob_uop_2_20_ftq_idx;
      5'b10101:
        casez_tmp_172 = rob_uop_2_21_ftq_idx;
      5'b10110:
        casez_tmp_172 = rob_uop_2_22_ftq_idx;
      5'b10111:
        casez_tmp_172 = rob_uop_2_23_ftq_idx;
      5'b11000:
        casez_tmp_172 = rob_uop_2_24_ftq_idx;
      5'b11001:
        casez_tmp_172 = rob_uop_2_25_ftq_idx;
      5'b11010:
        casez_tmp_172 = rob_uop_2_26_ftq_idx;
      5'b11011:
        casez_tmp_172 = rob_uop_2_27_ftq_idx;
      5'b11100:
        casez_tmp_172 = rob_uop_2_28_ftq_idx;
      5'b11101:
        casez_tmp_172 = rob_uop_2_29_ftq_idx;
      5'b11110:
        casez_tmp_172 = rob_uop_2_30_ftq_idx;
      default:
        casez_tmp_172 = rob_uop_2_31_ftq_idx;
    endcase
  end // always @(*)
  reg         casez_tmp_173;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_173 = rob_uop_2_0_edge_inst;
      5'b00001:
        casez_tmp_173 = rob_uop_2_1_edge_inst;
      5'b00010:
        casez_tmp_173 = rob_uop_2_2_edge_inst;
      5'b00011:
        casez_tmp_173 = rob_uop_2_3_edge_inst;
      5'b00100:
        casez_tmp_173 = rob_uop_2_4_edge_inst;
      5'b00101:
        casez_tmp_173 = rob_uop_2_5_edge_inst;
      5'b00110:
        casez_tmp_173 = rob_uop_2_6_edge_inst;
      5'b00111:
        casez_tmp_173 = rob_uop_2_7_edge_inst;
      5'b01000:
        casez_tmp_173 = rob_uop_2_8_edge_inst;
      5'b01001:
        casez_tmp_173 = rob_uop_2_9_edge_inst;
      5'b01010:
        casez_tmp_173 = rob_uop_2_10_edge_inst;
      5'b01011:
        casez_tmp_173 = rob_uop_2_11_edge_inst;
      5'b01100:
        casez_tmp_173 = rob_uop_2_12_edge_inst;
      5'b01101:
        casez_tmp_173 = rob_uop_2_13_edge_inst;
      5'b01110:
        casez_tmp_173 = rob_uop_2_14_edge_inst;
      5'b01111:
        casez_tmp_173 = rob_uop_2_15_edge_inst;
      5'b10000:
        casez_tmp_173 = rob_uop_2_16_edge_inst;
      5'b10001:
        casez_tmp_173 = rob_uop_2_17_edge_inst;
      5'b10010:
        casez_tmp_173 = rob_uop_2_18_edge_inst;
      5'b10011:
        casez_tmp_173 = rob_uop_2_19_edge_inst;
      5'b10100:
        casez_tmp_173 = rob_uop_2_20_edge_inst;
      5'b10101:
        casez_tmp_173 = rob_uop_2_21_edge_inst;
      5'b10110:
        casez_tmp_173 = rob_uop_2_22_edge_inst;
      5'b10111:
        casez_tmp_173 = rob_uop_2_23_edge_inst;
      5'b11000:
        casez_tmp_173 = rob_uop_2_24_edge_inst;
      5'b11001:
        casez_tmp_173 = rob_uop_2_25_edge_inst;
      5'b11010:
        casez_tmp_173 = rob_uop_2_26_edge_inst;
      5'b11011:
        casez_tmp_173 = rob_uop_2_27_edge_inst;
      5'b11100:
        casez_tmp_173 = rob_uop_2_28_edge_inst;
      5'b11101:
        casez_tmp_173 = rob_uop_2_29_edge_inst;
      5'b11110:
        casez_tmp_173 = rob_uop_2_30_edge_inst;
      default:
        casez_tmp_173 = rob_uop_2_31_edge_inst;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_174;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_174 = rob_uop_2_0_pc_lob;
      5'b00001:
        casez_tmp_174 = rob_uop_2_1_pc_lob;
      5'b00010:
        casez_tmp_174 = rob_uop_2_2_pc_lob;
      5'b00011:
        casez_tmp_174 = rob_uop_2_3_pc_lob;
      5'b00100:
        casez_tmp_174 = rob_uop_2_4_pc_lob;
      5'b00101:
        casez_tmp_174 = rob_uop_2_5_pc_lob;
      5'b00110:
        casez_tmp_174 = rob_uop_2_6_pc_lob;
      5'b00111:
        casez_tmp_174 = rob_uop_2_7_pc_lob;
      5'b01000:
        casez_tmp_174 = rob_uop_2_8_pc_lob;
      5'b01001:
        casez_tmp_174 = rob_uop_2_9_pc_lob;
      5'b01010:
        casez_tmp_174 = rob_uop_2_10_pc_lob;
      5'b01011:
        casez_tmp_174 = rob_uop_2_11_pc_lob;
      5'b01100:
        casez_tmp_174 = rob_uop_2_12_pc_lob;
      5'b01101:
        casez_tmp_174 = rob_uop_2_13_pc_lob;
      5'b01110:
        casez_tmp_174 = rob_uop_2_14_pc_lob;
      5'b01111:
        casez_tmp_174 = rob_uop_2_15_pc_lob;
      5'b10000:
        casez_tmp_174 = rob_uop_2_16_pc_lob;
      5'b10001:
        casez_tmp_174 = rob_uop_2_17_pc_lob;
      5'b10010:
        casez_tmp_174 = rob_uop_2_18_pc_lob;
      5'b10011:
        casez_tmp_174 = rob_uop_2_19_pc_lob;
      5'b10100:
        casez_tmp_174 = rob_uop_2_20_pc_lob;
      5'b10101:
        casez_tmp_174 = rob_uop_2_21_pc_lob;
      5'b10110:
        casez_tmp_174 = rob_uop_2_22_pc_lob;
      5'b10111:
        casez_tmp_174 = rob_uop_2_23_pc_lob;
      5'b11000:
        casez_tmp_174 = rob_uop_2_24_pc_lob;
      5'b11001:
        casez_tmp_174 = rob_uop_2_25_pc_lob;
      5'b11010:
        casez_tmp_174 = rob_uop_2_26_pc_lob;
      5'b11011:
        casez_tmp_174 = rob_uop_2_27_pc_lob;
      5'b11100:
        casez_tmp_174 = rob_uop_2_28_pc_lob;
      5'b11101:
        casez_tmp_174 = rob_uop_2_29_pc_lob;
      5'b11110:
        casez_tmp_174 = rob_uop_2_30_pc_lob;
      default:
        casez_tmp_174 = rob_uop_2_31_pc_lob;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_175;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_175 = rob_uop_2_0_pdst;
      5'b00001:
        casez_tmp_175 = rob_uop_2_1_pdst;
      5'b00010:
        casez_tmp_175 = rob_uop_2_2_pdst;
      5'b00011:
        casez_tmp_175 = rob_uop_2_3_pdst;
      5'b00100:
        casez_tmp_175 = rob_uop_2_4_pdst;
      5'b00101:
        casez_tmp_175 = rob_uop_2_5_pdst;
      5'b00110:
        casez_tmp_175 = rob_uop_2_6_pdst;
      5'b00111:
        casez_tmp_175 = rob_uop_2_7_pdst;
      5'b01000:
        casez_tmp_175 = rob_uop_2_8_pdst;
      5'b01001:
        casez_tmp_175 = rob_uop_2_9_pdst;
      5'b01010:
        casez_tmp_175 = rob_uop_2_10_pdst;
      5'b01011:
        casez_tmp_175 = rob_uop_2_11_pdst;
      5'b01100:
        casez_tmp_175 = rob_uop_2_12_pdst;
      5'b01101:
        casez_tmp_175 = rob_uop_2_13_pdst;
      5'b01110:
        casez_tmp_175 = rob_uop_2_14_pdst;
      5'b01111:
        casez_tmp_175 = rob_uop_2_15_pdst;
      5'b10000:
        casez_tmp_175 = rob_uop_2_16_pdst;
      5'b10001:
        casez_tmp_175 = rob_uop_2_17_pdst;
      5'b10010:
        casez_tmp_175 = rob_uop_2_18_pdst;
      5'b10011:
        casez_tmp_175 = rob_uop_2_19_pdst;
      5'b10100:
        casez_tmp_175 = rob_uop_2_20_pdst;
      5'b10101:
        casez_tmp_175 = rob_uop_2_21_pdst;
      5'b10110:
        casez_tmp_175 = rob_uop_2_22_pdst;
      5'b10111:
        casez_tmp_175 = rob_uop_2_23_pdst;
      5'b11000:
        casez_tmp_175 = rob_uop_2_24_pdst;
      5'b11001:
        casez_tmp_175 = rob_uop_2_25_pdst;
      5'b11010:
        casez_tmp_175 = rob_uop_2_26_pdst;
      5'b11011:
        casez_tmp_175 = rob_uop_2_27_pdst;
      5'b11100:
        casez_tmp_175 = rob_uop_2_28_pdst;
      5'b11101:
        casez_tmp_175 = rob_uop_2_29_pdst;
      5'b11110:
        casez_tmp_175 = rob_uop_2_30_pdst;
      default:
        casez_tmp_175 = rob_uop_2_31_pdst;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_176;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_176 = rob_uop_2_0_stale_pdst;
      5'b00001:
        casez_tmp_176 = rob_uop_2_1_stale_pdst;
      5'b00010:
        casez_tmp_176 = rob_uop_2_2_stale_pdst;
      5'b00011:
        casez_tmp_176 = rob_uop_2_3_stale_pdst;
      5'b00100:
        casez_tmp_176 = rob_uop_2_4_stale_pdst;
      5'b00101:
        casez_tmp_176 = rob_uop_2_5_stale_pdst;
      5'b00110:
        casez_tmp_176 = rob_uop_2_6_stale_pdst;
      5'b00111:
        casez_tmp_176 = rob_uop_2_7_stale_pdst;
      5'b01000:
        casez_tmp_176 = rob_uop_2_8_stale_pdst;
      5'b01001:
        casez_tmp_176 = rob_uop_2_9_stale_pdst;
      5'b01010:
        casez_tmp_176 = rob_uop_2_10_stale_pdst;
      5'b01011:
        casez_tmp_176 = rob_uop_2_11_stale_pdst;
      5'b01100:
        casez_tmp_176 = rob_uop_2_12_stale_pdst;
      5'b01101:
        casez_tmp_176 = rob_uop_2_13_stale_pdst;
      5'b01110:
        casez_tmp_176 = rob_uop_2_14_stale_pdst;
      5'b01111:
        casez_tmp_176 = rob_uop_2_15_stale_pdst;
      5'b10000:
        casez_tmp_176 = rob_uop_2_16_stale_pdst;
      5'b10001:
        casez_tmp_176 = rob_uop_2_17_stale_pdst;
      5'b10010:
        casez_tmp_176 = rob_uop_2_18_stale_pdst;
      5'b10011:
        casez_tmp_176 = rob_uop_2_19_stale_pdst;
      5'b10100:
        casez_tmp_176 = rob_uop_2_20_stale_pdst;
      5'b10101:
        casez_tmp_176 = rob_uop_2_21_stale_pdst;
      5'b10110:
        casez_tmp_176 = rob_uop_2_22_stale_pdst;
      5'b10111:
        casez_tmp_176 = rob_uop_2_23_stale_pdst;
      5'b11000:
        casez_tmp_176 = rob_uop_2_24_stale_pdst;
      5'b11001:
        casez_tmp_176 = rob_uop_2_25_stale_pdst;
      5'b11010:
        casez_tmp_176 = rob_uop_2_26_stale_pdst;
      5'b11011:
        casez_tmp_176 = rob_uop_2_27_stale_pdst;
      5'b11100:
        casez_tmp_176 = rob_uop_2_28_stale_pdst;
      5'b11101:
        casez_tmp_176 = rob_uop_2_29_stale_pdst;
      5'b11110:
        casez_tmp_176 = rob_uop_2_30_stale_pdst;
      default:
        casez_tmp_176 = rob_uop_2_31_stale_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_177;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_177 = rob_uop_2_0_is_fencei;
      5'b00001:
        casez_tmp_177 = rob_uop_2_1_is_fencei;
      5'b00010:
        casez_tmp_177 = rob_uop_2_2_is_fencei;
      5'b00011:
        casez_tmp_177 = rob_uop_2_3_is_fencei;
      5'b00100:
        casez_tmp_177 = rob_uop_2_4_is_fencei;
      5'b00101:
        casez_tmp_177 = rob_uop_2_5_is_fencei;
      5'b00110:
        casez_tmp_177 = rob_uop_2_6_is_fencei;
      5'b00111:
        casez_tmp_177 = rob_uop_2_7_is_fencei;
      5'b01000:
        casez_tmp_177 = rob_uop_2_8_is_fencei;
      5'b01001:
        casez_tmp_177 = rob_uop_2_9_is_fencei;
      5'b01010:
        casez_tmp_177 = rob_uop_2_10_is_fencei;
      5'b01011:
        casez_tmp_177 = rob_uop_2_11_is_fencei;
      5'b01100:
        casez_tmp_177 = rob_uop_2_12_is_fencei;
      5'b01101:
        casez_tmp_177 = rob_uop_2_13_is_fencei;
      5'b01110:
        casez_tmp_177 = rob_uop_2_14_is_fencei;
      5'b01111:
        casez_tmp_177 = rob_uop_2_15_is_fencei;
      5'b10000:
        casez_tmp_177 = rob_uop_2_16_is_fencei;
      5'b10001:
        casez_tmp_177 = rob_uop_2_17_is_fencei;
      5'b10010:
        casez_tmp_177 = rob_uop_2_18_is_fencei;
      5'b10011:
        casez_tmp_177 = rob_uop_2_19_is_fencei;
      5'b10100:
        casez_tmp_177 = rob_uop_2_20_is_fencei;
      5'b10101:
        casez_tmp_177 = rob_uop_2_21_is_fencei;
      5'b10110:
        casez_tmp_177 = rob_uop_2_22_is_fencei;
      5'b10111:
        casez_tmp_177 = rob_uop_2_23_is_fencei;
      5'b11000:
        casez_tmp_177 = rob_uop_2_24_is_fencei;
      5'b11001:
        casez_tmp_177 = rob_uop_2_25_is_fencei;
      5'b11010:
        casez_tmp_177 = rob_uop_2_26_is_fencei;
      5'b11011:
        casez_tmp_177 = rob_uop_2_27_is_fencei;
      5'b11100:
        casez_tmp_177 = rob_uop_2_28_is_fencei;
      5'b11101:
        casez_tmp_177 = rob_uop_2_29_is_fencei;
      5'b11110:
        casez_tmp_177 = rob_uop_2_30_is_fencei;
      default:
        casez_tmp_177 = rob_uop_2_31_is_fencei;
    endcase
  end // always @(*)
  reg         casez_tmp_178;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_178 = rob_uop_2_0_uses_ldq;
      5'b00001:
        casez_tmp_178 = rob_uop_2_1_uses_ldq;
      5'b00010:
        casez_tmp_178 = rob_uop_2_2_uses_ldq;
      5'b00011:
        casez_tmp_178 = rob_uop_2_3_uses_ldq;
      5'b00100:
        casez_tmp_178 = rob_uop_2_4_uses_ldq;
      5'b00101:
        casez_tmp_178 = rob_uop_2_5_uses_ldq;
      5'b00110:
        casez_tmp_178 = rob_uop_2_6_uses_ldq;
      5'b00111:
        casez_tmp_178 = rob_uop_2_7_uses_ldq;
      5'b01000:
        casez_tmp_178 = rob_uop_2_8_uses_ldq;
      5'b01001:
        casez_tmp_178 = rob_uop_2_9_uses_ldq;
      5'b01010:
        casez_tmp_178 = rob_uop_2_10_uses_ldq;
      5'b01011:
        casez_tmp_178 = rob_uop_2_11_uses_ldq;
      5'b01100:
        casez_tmp_178 = rob_uop_2_12_uses_ldq;
      5'b01101:
        casez_tmp_178 = rob_uop_2_13_uses_ldq;
      5'b01110:
        casez_tmp_178 = rob_uop_2_14_uses_ldq;
      5'b01111:
        casez_tmp_178 = rob_uop_2_15_uses_ldq;
      5'b10000:
        casez_tmp_178 = rob_uop_2_16_uses_ldq;
      5'b10001:
        casez_tmp_178 = rob_uop_2_17_uses_ldq;
      5'b10010:
        casez_tmp_178 = rob_uop_2_18_uses_ldq;
      5'b10011:
        casez_tmp_178 = rob_uop_2_19_uses_ldq;
      5'b10100:
        casez_tmp_178 = rob_uop_2_20_uses_ldq;
      5'b10101:
        casez_tmp_178 = rob_uop_2_21_uses_ldq;
      5'b10110:
        casez_tmp_178 = rob_uop_2_22_uses_ldq;
      5'b10111:
        casez_tmp_178 = rob_uop_2_23_uses_ldq;
      5'b11000:
        casez_tmp_178 = rob_uop_2_24_uses_ldq;
      5'b11001:
        casez_tmp_178 = rob_uop_2_25_uses_ldq;
      5'b11010:
        casez_tmp_178 = rob_uop_2_26_uses_ldq;
      5'b11011:
        casez_tmp_178 = rob_uop_2_27_uses_ldq;
      5'b11100:
        casez_tmp_178 = rob_uop_2_28_uses_ldq;
      5'b11101:
        casez_tmp_178 = rob_uop_2_29_uses_ldq;
      5'b11110:
        casez_tmp_178 = rob_uop_2_30_uses_ldq;
      default:
        casez_tmp_178 = rob_uop_2_31_uses_ldq;
    endcase
  end // always @(*)
  reg         casez_tmp_179;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_179 = rob_uop_2_0_uses_stq;
      5'b00001:
        casez_tmp_179 = rob_uop_2_1_uses_stq;
      5'b00010:
        casez_tmp_179 = rob_uop_2_2_uses_stq;
      5'b00011:
        casez_tmp_179 = rob_uop_2_3_uses_stq;
      5'b00100:
        casez_tmp_179 = rob_uop_2_4_uses_stq;
      5'b00101:
        casez_tmp_179 = rob_uop_2_5_uses_stq;
      5'b00110:
        casez_tmp_179 = rob_uop_2_6_uses_stq;
      5'b00111:
        casez_tmp_179 = rob_uop_2_7_uses_stq;
      5'b01000:
        casez_tmp_179 = rob_uop_2_8_uses_stq;
      5'b01001:
        casez_tmp_179 = rob_uop_2_9_uses_stq;
      5'b01010:
        casez_tmp_179 = rob_uop_2_10_uses_stq;
      5'b01011:
        casez_tmp_179 = rob_uop_2_11_uses_stq;
      5'b01100:
        casez_tmp_179 = rob_uop_2_12_uses_stq;
      5'b01101:
        casez_tmp_179 = rob_uop_2_13_uses_stq;
      5'b01110:
        casez_tmp_179 = rob_uop_2_14_uses_stq;
      5'b01111:
        casez_tmp_179 = rob_uop_2_15_uses_stq;
      5'b10000:
        casez_tmp_179 = rob_uop_2_16_uses_stq;
      5'b10001:
        casez_tmp_179 = rob_uop_2_17_uses_stq;
      5'b10010:
        casez_tmp_179 = rob_uop_2_18_uses_stq;
      5'b10011:
        casez_tmp_179 = rob_uop_2_19_uses_stq;
      5'b10100:
        casez_tmp_179 = rob_uop_2_20_uses_stq;
      5'b10101:
        casez_tmp_179 = rob_uop_2_21_uses_stq;
      5'b10110:
        casez_tmp_179 = rob_uop_2_22_uses_stq;
      5'b10111:
        casez_tmp_179 = rob_uop_2_23_uses_stq;
      5'b11000:
        casez_tmp_179 = rob_uop_2_24_uses_stq;
      5'b11001:
        casez_tmp_179 = rob_uop_2_25_uses_stq;
      5'b11010:
        casez_tmp_179 = rob_uop_2_26_uses_stq;
      5'b11011:
        casez_tmp_179 = rob_uop_2_27_uses_stq;
      5'b11100:
        casez_tmp_179 = rob_uop_2_28_uses_stq;
      5'b11101:
        casez_tmp_179 = rob_uop_2_29_uses_stq;
      5'b11110:
        casez_tmp_179 = rob_uop_2_30_uses_stq;
      default:
        casez_tmp_179 = rob_uop_2_31_uses_stq;
    endcase
  end // always @(*)
  reg         casez_tmp_180;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_180 = rob_uop_2_0_is_sys_pc2epc;
      5'b00001:
        casez_tmp_180 = rob_uop_2_1_is_sys_pc2epc;
      5'b00010:
        casez_tmp_180 = rob_uop_2_2_is_sys_pc2epc;
      5'b00011:
        casez_tmp_180 = rob_uop_2_3_is_sys_pc2epc;
      5'b00100:
        casez_tmp_180 = rob_uop_2_4_is_sys_pc2epc;
      5'b00101:
        casez_tmp_180 = rob_uop_2_5_is_sys_pc2epc;
      5'b00110:
        casez_tmp_180 = rob_uop_2_6_is_sys_pc2epc;
      5'b00111:
        casez_tmp_180 = rob_uop_2_7_is_sys_pc2epc;
      5'b01000:
        casez_tmp_180 = rob_uop_2_8_is_sys_pc2epc;
      5'b01001:
        casez_tmp_180 = rob_uop_2_9_is_sys_pc2epc;
      5'b01010:
        casez_tmp_180 = rob_uop_2_10_is_sys_pc2epc;
      5'b01011:
        casez_tmp_180 = rob_uop_2_11_is_sys_pc2epc;
      5'b01100:
        casez_tmp_180 = rob_uop_2_12_is_sys_pc2epc;
      5'b01101:
        casez_tmp_180 = rob_uop_2_13_is_sys_pc2epc;
      5'b01110:
        casez_tmp_180 = rob_uop_2_14_is_sys_pc2epc;
      5'b01111:
        casez_tmp_180 = rob_uop_2_15_is_sys_pc2epc;
      5'b10000:
        casez_tmp_180 = rob_uop_2_16_is_sys_pc2epc;
      5'b10001:
        casez_tmp_180 = rob_uop_2_17_is_sys_pc2epc;
      5'b10010:
        casez_tmp_180 = rob_uop_2_18_is_sys_pc2epc;
      5'b10011:
        casez_tmp_180 = rob_uop_2_19_is_sys_pc2epc;
      5'b10100:
        casez_tmp_180 = rob_uop_2_20_is_sys_pc2epc;
      5'b10101:
        casez_tmp_180 = rob_uop_2_21_is_sys_pc2epc;
      5'b10110:
        casez_tmp_180 = rob_uop_2_22_is_sys_pc2epc;
      5'b10111:
        casez_tmp_180 = rob_uop_2_23_is_sys_pc2epc;
      5'b11000:
        casez_tmp_180 = rob_uop_2_24_is_sys_pc2epc;
      5'b11001:
        casez_tmp_180 = rob_uop_2_25_is_sys_pc2epc;
      5'b11010:
        casez_tmp_180 = rob_uop_2_26_is_sys_pc2epc;
      5'b11011:
        casez_tmp_180 = rob_uop_2_27_is_sys_pc2epc;
      5'b11100:
        casez_tmp_180 = rob_uop_2_28_is_sys_pc2epc;
      5'b11101:
        casez_tmp_180 = rob_uop_2_29_is_sys_pc2epc;
      5'b11110:
        casez_tmp_180 = rob_uop_2_30_is_sys_pc2epc;
      default:
        casez_tmp_180 = rob_uop_2_31_is_sys_pc2epc;
    endcase
  end // always @(*)
  reg         casez_tmp_181;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_181 = rob_uop_2_0_flush_on_commit;
      5'b00001:
        casez_tmp_181 = rob_uop_2_1_flush_on_commit;
      5'b00010:
        casez_tmp_181 = rob_uop_2_2_flush_on_commit;
      5'b00011:
        casez_tmp_181 = rob_uop_2_3_flush_on_commit;
      5'b00100:
        casez_tmp_181 = rob_uop_2_4_flush_on_commit;
      5'b00101:
        casez_tmp_181 = rob_uop_2_5_flush_on_commit;
      5'b00110:
        casez_tmp_181 = rob_uop_2_6_flush_on_commit;
      5'b00111:
        casez_tmp_181 = rob_uop_2_7_flush_on_commit;
      5'b01000:
        casez_tmp_181 = rob_uop_2_8_flush_on_commit;
      5'b01001:
        casez_tmp_181 = rob_uop_2_9_flush_on_commit;
      5'b01010:
        casez_tmp_181 = rob_uop_2_10_flush_on_commit;
      5'b01011:
        casez_tmp_181 = rob_uop_2_11_flush_on_commit;
      5'b01100:
        casez_tmp_181 = rob_uop_2_12_flush_on_commit;
      5'b01101:
        casez_tmp_181 = rob_uop_2_13_flush_on_commit;
      5'b01110:
        casez_tmp_181 = rob_uop_2_14_flush_on_commit;
      5'b01111:
        casez_tmp_181 = rob_uop_2_15_flush_on_commit;
      5'b10000:
        casez_tmp_181 = rob_uop_2_16_flush_on_commit;
      5'b10001:
        casez_tmp_181 = rob_uop_2_17_flush_on_commit;
      5'b10010:
        casez_tmp_181 = rob_uop_2_18_flush_on_commit;
      5'b10011:
        casez_tmp_181 = rob_uop_2_19_flush_on_commit;
      5'b10100:
        casez_tmp_181 = rob_uop_2_20_flush_on_commit;
      5'b10101:
        casez_tmp_181 = rob_uop_2_21_flush_on_commit;
      5'b10110:
        casez_tmp_181 = rob_uop_2_22_flush_on_commit;
      5'b10111:
        casez_tmp_181 = rob_uop_2_23_flush_on_commit;
      5'b11000:
        casez_tmp_181 = rob_uop_2_24_flush_on_commit;
      5'b11001:
        casez_tmp_181 = rob_uop_2_25_flush_on_commit;
      5'b11010:
        casez_tmp_181 = rob_uop_2_26_flush_on_commit;
      5'b11011:
        casez_tmp_181 = rob_uop_2_27_flush_on_commit;
      5'b11100:
        casez_tmp_181 = rob_uop_2_28_flush_on_commit;
      5'b11101:
        casez_tmp_181 = rob_uop_2_29_flush_on_commit;
      5'b11110:
        casez_tmp_181 = rob_uop_2_30_flush_on_commit;
      default:
        casez_tmp_181 = rob_uop_2_31_flush_on_commit;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_182;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_182 = rob_uop_2_0_ldst;
      5'b00001:
        casez_tmp_182 = rob_uop_2_1_ldst;
      5'b00010:
        casez_tmp_182 = rob_uop_2_2_ldst;
      5'b00011:
        casez_tmp_182 = rob_uop_2_3_ldst;
      5'b00100:
        casez_tmp_182 = rob_uop_2_4_ldst;
      5'b00101:
        casez_tmp_182 = rob_uop_2_5_ldst;
      5'b00110:
        casez_tmp_182 = rob_uop_2_6_ldst;
      5'b00111:
        casez_tmp_182 = rob_uop_2_7_ldst;
      5'b01000:
        casez_tmp_182 = rob_uop_2_8_ldst;
      5'b01001:
        casez_tmp_182 = rob_uop_2_9_ldst;
      5'b01010:
        casez_tmp_182 = rob_uop_2_10_ldst;
      5'b01011:
        casez_tmp_182 = rob_uop_2_11_ldst;
      5'b01100:
        casez_tmp_182 = rob_uop_2_12_ldst;
      5'b01101:
        casez_tmp_182 = rob_uop_2_13_ldst;
      5'b01110:
        casez_tmp_182 = rob_uop_2_14_ldst;
      5'b01111:
        casez_tmp_182 = rob_uop_2_15_ldst;
      5'b10000:
        casez_tmp_182 = rob_uop_2_16_ldst;
      5'b10001:
        casez_tmp_182 = rob_uop_2_17_ldst;
      5'b10010:
        casez_tmp_182 = rob_uop_2_18_ldst;
      5'b10011:
        casez_tmp_182 = rob_uop_2_19_ldst;
      5'b10100:
        casez_tmp_182 = rob_uop_2_20_ldst;
      5'b10101:
        casez_tmp_182 = rob_uop_2_21_ldst;
      5'b10110:
        casez_tmp_182 = rob_uop_2_22_ldst;
      5'b10111:
        casez_tmp_182 = rob_uop_2_23_ldst;
      5'b11000:
        casez_tmp_182 = rob_uop_2_24_ldst;
      5'b11001:
        casez_tmp_182 = rob_uop_2_25_ldst;
      5'b11010:
        casez_tmp_182 = rob_uop_2_26_ldst;
      5'b11011:
        casez_tmp_182 = rob_uop_2_27_ldst;
      5'b11100:
        casez_tmp_182 = rob_uop_2_28_ldst;
      5'b11101:
        casez_tmp_182 = rob_uop_2_29_ldst;
      5'b11110:
        casez_tmp_182 = rob_uop_2_30_ldst;
      default:
        casez_tmp_182 = rob_uop_2_31_ldst;
    endcase
  end // always @(*)
  reg         casez_tmp_183;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_183 = rob_uop_2_0_ldst_val;
      5'b00001:
        casez_tmp_183 = rob_uop_2_1_ldst_val;
      5'b00010:
        casez_tmp_183 = rob_uop_2_2_ldst_val;
      5'b00011:
        casez_tmp_183 = rob_uop_2_3_ldst_val;
      5'b00100:
        casez_tmp_183 = rob_uop_2_4_ldst_val;
      5'b00101:
        casez_tmp_183 = rob_uop_2_5_ldst_val;
      5'b00110:
        casez_tmp_183 = rob_uop_2_6_ldst_val;
      5'b00111:
        casez_tmp_183 = rob_uop_2_7_ldst_val;
      5'b01000:
        casez_tmp_183 = rob_uop_2_8_ldst_val;
      5'b01001:
        casez_tmp_183 = rob_uop_2_9_ldst_val;
      5'b01010:
        casez_tmp_183 = rob_uop_2_10_ldst_val;
      5'b01011:
        casez_tmp_183 = rob_uop_2_11_ldst_val;
      5'b01100:
        casez_tmp_183 = rob_uop_2_12_ldst_val;
      5'b01101:
        casez_tmp_183 = rob_uop_2_13_ldst_val;
      5'b01110:
        casez_tmp_183 = rob_uop_2_14_ldst_val;
      5'b01111:
        casez_tmp_183 = rob_uop_2_15_ldst_val;
      5'b10000:
        casez_tmp_183 = rob_uop_2_16_ldst_val;
      5'b10001:
        casez_tmp_183 = rob_uop_2_17_ldst_val;
      5'b10010:
        casez_tmp_183 = rob_uop_2_18_ldst_val;
      5'b10011:
        casez_tmp_183 = rob_uop_2_19_ldst_val;
      5'b10100:
        casez_tmp_183 = rob_uop_2_20_ldst_val;
      5'b10101:
        casez_tmp_183 = rob_uop_2_21_ldst_val;
      5'b10110:
        casez_tmp_183 = rob_uop_2_22_ldst_val;
      5'b10111:
        casez_tmp_183 = rob_uop_2_23_ldst_val;
      5'b11000:
        casez_tmp_183 = rob_uop_2_24_ldst_val;
      5'b11001:
        casez_tmp_183 = rob_uop_2_25_ldst_val;
      5'b11010:
        casez_tmp_183 = rob_uop_2_26_ldst_val;
      5'b11011:
        casez_tmp_183 = rob_uop_2_27_ldst_val;
      5'b11100:
        casez_tmp_183 = rob_uop_2_28_ldst_val;
      5'b11101:
        casez_tmp_183 = rob_uop_2_29_ldst_val;
      5'b11110:
        casez_tmp_183 = rob_uop_2_30_ldst_val;
      default:
        casez_tmp_183 = rob_uop_2_31_ldst_val;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_184;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_184 = rob_uop_2_0_dst_rtype;
      5'b00001:
        casez_tmp_184 = rob_uop_2_1_dst_rtype;
      5'b00010:
        casez_tmp_184 = rob_uop_2_2_dst_rtype;
      5'b00011:
        casez_tmp_184 = rob_uop_2_3_dst_rtype;
      5'b00100:
        casez_tmp_184 = rob_uop_2_4_dst_rtype;
      5'b00101:
        casez_tmp_184 = rob_uop_2_5_dst_rtype;
      5'b00110:
        casez_tmp_184 = rob_uop_2_6_dst_rtype;
      5'b00111:
        casez_tmp_184 = rob_uop_2_7_dst_rtype;
      5'b01000:
        casez_tmp_184 = rob_uop_2_8_dst_rtype;
      5'b01001:
        casez_tmp_184 = rob_uop_2_9_dst_rtype;
      5'b01010:
        casez_tmp_184 = rob_uop_2_10_dst_rtype;
      5'b01011:
        casez_tmp_184 = rob_uop_2_11_dst_rtype;
      5'b01100:
        casez_tmp_184 = rob_uop_2_12_dst_rtype;
      5'b01101:
        casez_tmp_184 = rob_uop_2_13_dst_rtype;
      5'b01110:
        casez_tmp_184 = rob_uop_2_14_dst_rtype;
      5'b01111:
        casez_tmp_184 = rob_uop_2_15_dst_rtype;
      5'b10000:
        casez_tmp_184 = rob_uop_2_16_dst_rtype;
      5'b10001:
        casez_tmp_184 = rob_uop_2_17_dst_rtype;
      5'b10010:
        casez_tmp_184 = rob_uop_2_18_dst_rtype;
      5'b10011:
        casez_tmp_184 = rob_uop_2_19_dst_rtype;
      5'b10100:
        casez_tmp_184 = rob_uop_2_20_dst_rtype;
      5'b10101:
        casez_tmp_184 = rob_uop_2_21_dst_rtype;
      5'b10110:
        casez_tmp_184 = rob_uop_2_22_dst_rtype;
      5'b10111:
        casez_tmp_184 = rob_uop_2_23_dst_rtype;
      5'b11000:
        casez_tmp_184 = rob_uop_2_24_dst_rtype;
      5'b11001:
        casez_tmp_184 = rob_uop_2_25_dst_rtype;
      5'b11010:
        casez_tmp_184 = rob_uop_2_26_dst_rtype;
      5'b11011:
        casez_tmp_184 = rob_uop_2_27_dst_rtype;
      5'b11100:
        casez_tmp_184 = rob_uop_2_28_dst_rtype;
      5'b11101:
        casez_tmp_184 = rob_uop_2_29_dst_rtype;
      5'b11110:
        casez_tmp_184 = rob_uop_2_30_dst_rtype;
      default:
        casez_tmp_184 = rob_uop_2_31_dst_rtype;
    endcase
  end // always @(*)
  reg         casez_tmp_185;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_185 = rob_uop_2_0_fp_val;
      5'b00001:
        casez_tmp_185 = rob_uop_2_1_fp_val;
      5'b00010:
        casez_tmp_185 = rob_uop_2_2_fp_val;
      5'b00011:
        casez_tmp_185 = rob_uop_2_3_fp_val;
      5'b00100:
        casez_tmp_185 = rob_uop_2_4_fp_val;
      5'b00101:
        casez_tmp_185 = rob_uop_2_5_fp_val;
      5'b00110:
        casez_tmp_185 = rob_uop_2_6_fp_val;
      5'b00111:
        casez_tmp_185 = rob_uop_2_7_fp_val;
      5'b01000:
        casez_tmp_185 = rob_uop_2_8_fp_val;
      5'b01001:
        casez_tmp_185 = rob_uop_2_9_fp_val;
      5'b01010:
        casez_tmp_185 = rob_uop_2_10_fp_val;
      5'b01011:
        casez_tmp_185 = rob_uop_2_11_fp_val;
      5'b01100:
        casez_tmp_185 = rob_uop_2_12_fp_val;
      5'b01101:
        casez_tmp_185 = rob_uop_2_13_fp_val;
      5'b01110:
        casez_tmp_185 = rob_uop_2_14_fp_val;
      5'b01111:
        casez_tmp_185 = rob_uop_2_15_fp_val;
      5'b10000:
        casez_tmp_185 = rob_uop_2_16_fp_val;
      5'b10001:
        casez_tmp_185 = rob_uop_2_17_fp_val;
      5'b10010:
        casez_tmp_185 = rob_uop_2_18_fp_val;
      5'b10011:
        casez_tmp_185 = rob_uop_2_19_fp_val;
      5'b10100:
        casez_tmp_185 = rob_uop_2_20_fp_val;
      5'b10101:
        casez_tmp_185 = rob_uop_2_21_fp_val;
      5'b10110:
        casez_tmp_185 = rob_uop_2_22_fp_val;
      5'b10111:
        casez_tmp_185 = rob_uop_2_23_fp_val;
      5'b11000:
        casez_tmp_185 = rob_uop_2_24_fp_val;
      5'b11001:
        casez_tmp_185 = rob_uop_2_25_fp_val;
      5'b11010:
        casez_tmp_185 = rob_uop_2_26_fp_val;
      5'b11011:
        casez_tmp_185 = rob_uop_2_27_fp_val;
      5'b11100:
        casez_tmp_185 = rob_uop_2_28_fp_val;
      5'b11101:
        casez_tmp_185 = rob_uop_2_29_fp_val;
      5'b11110:
        casez_tmp_185 = rob_uop_2_30_fp_val;
      default:
        casez_tmp_185 = rob_uop_2_31_fp_val;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_186;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_186 = rob_uop_2_0_debug_fsrc;
      5'b00001:
        casez_tmp_186 = rob_uop_2_1_debug_fsrc;
      5'b00010:
        casez_tmp_186 = rob_uop_2_2_debug_fsrc;
      5'b00011:
        casez_tmp_186 = rob_uop_2_3_debug_fsrc;
      5'b00100:
        casez_tmp_186 = rob_uop_2_4_debug_fsrc;
      5'b00101:
        casez_tmp_186 = rob_uop_2_5_debug_fsrc;
      5'b00110:
        casez_tmp_186 = rob_uop_2_6_debug_fsrc;
      5'b00111:
        casez_tmp_186 = rob_uop_2_7_debug_fsrc;
      5'b01000:
        casez_tmp_186 = rob_uop_2_8_debug_fsrc;
      5'b01001:
        casez_tmp_186 = rob_uop_2_9_debug_fsrc;
      5'b01010:
        casez_tmp_186 = rob_uop_2_10_debug_fsrc;
      5'b01011:
        casez_tmp_186 = rob_uop_2_11_debug_fsrc;
      5'b01100:
        casez_tmp_186 = rob_uop_2_12_debug_fsrc;
      5'b01101:
        casez_tmp_186 = rob_uop_2_13_debug_fsrc;
      5'b01110:
        casez_tmp_186 = rob_uop_2_14_debug_fsrc;
      5'b01111:
        casez_tmp_186 = rob_uop_2_15_debug_fsrc;
      5'b10000:
        casez_tmp_186 = rob_uop_2_16_debug_fsrc;
      5'b10001:
        casez_tmp_186 = rob_uop_2_17_debug_fsrc;
      5'b10010:
        casez_tmp_186 = rob_uop_2_18_debug_fsrc;
      5'b10011:
        casez_tmp_186 = rob_uop_2_19_debug_fsrc;
      5'b10100:
        casez_tmp_186 = rob_uop_2_20_debug_fsrc;
      5'b10101:
        casez_tmp_186 = rob_uop_2_21_debug_fsrc;
      5'b10110:
        casez_tmp_186 = rob_uop_2_22_debug_fsrc;
      5'b10111:
        casez_tmp_186 = rob_uop_2_23_debug_fsrc;
      5'b11000:
        casez_tmp_186 = rob_uop_2_24_debug_fsrc;
      5'b11001:
        casez_tmp_186 = rob_uop_2_25_debug_fsrc;
      5'b11010:
        casez_tmp_186 = rob_uop_2_26_debug_fsrc;
      5'b11011:
        casez_tmp_186 = rob_uop_2_27_debug_fsrc;
      5'b11100:
        casez_tmp_186 = rob_uop_2_28_debug_fsrc;
      5'b11101:
        casez_tmp_186 = rob_uop_2_29_debug_fsrc;
      5'b11110:
        casez_tmp_186 = rob_uop_2_30_debug_fsrc;
      default:
        casez_tmp_186 = rob_uop_2_31_debug_fsrc;
    endcase
  end // always @(*)
  wire        _GEN_48 = io_brupdate_b2_mispredict & io_brupdate_b2_uop_rob_idx[1:0] == 2'h2;
  wire        rbk_row_2 = _io_commit_rollback_T_3 & ~full;
  reg         casez_tmp_187;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_187 = rob_val_2_0;
      5'b00001:
        casez_tmp_187 = rob_val_2_1;
      5'b00010:
        casez_tmp_187 = rob_val_2_2;
      5'b00011:
        casez_tmp_187 = rob_val_2_3;
      5'b00100:
        casez_tmp_187 = rob_val_2_4;
      5'b00101:
        casez_tmp_187 = rob_val_2_5;
      5'b00110:
        casez_tmp_187 = rob_val_2_6;
      5'b00111:
        casez_tmp_187 = rob_val_2_7;
      5'b01000:
        casez_tmp_187 = rob_val_2_8;
      5'b01001:
        casez_tmp_187 = rob_val_2_9;
      5'b01010:
        casez_tmp_187 = rob_val_2_10;
      5'b01011:
        casez_tmp_187 = rob_val_2_11;
      5'b01100:
        casez_tmp_187 = rob_val_2_12;
      5'b01101:
        casez_tmp_187 = rob_val_2_13;
      5'b01110:
        casez_tmp_187 = rob_val_2_14;
      5'b01111:
        casez_tmp_187 = rob_val_2_15;
      5'b10000:
        casez_tmp_187 = rob_val_2_16;
      5'b10001:
        casez_tmp_187 = rob_val_2_17;
      5'b10010:
        casez_tmp_187 = rob_val_2_18;
      5'b10011:
        casez_tmp_187 = rob_val_2_19;
      5'b10100:
        casez_tmp_187 = rob_val_2_20;
      5'b10101:
        casez_tmp_187 = rob_val_2_21;
      5'b10110:
        casez_tmp_187 = rob_val_2_22;
      5'b10111:
        casez_tmp_187 = rob_val_2_23;
      5'b11000:
        casez_tmp_187 = rob_val_2_24;
      5'b11001:
        casez_tmp_187 = rob_val_2_25;
      5'b11010:
        casez_tmp_187 = rob_val_2_26;
      5'b11011:
        casez_tmp_187 = rob_val_2_27;
      5'b11100:
        casez_tmp_187 = rob_val_2_28;
      5'b11101:
        casez_tmp_187 = rob_val_2_29;
      5'b11110:
        casez_tmp_187 = rob_val_2_30;
      default:
        casez_tmp_187 = rob_val_2_31;
    endcase
  end // always @(*)
  wire        _io_commit_rbk_valids_2_output = rbk_row_2 & casez_tmp_187;
  reg  [4:0]  casez_tmp_188;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_188 = rob_fflags_2_0;
      5'b00001:
        casez_tmp_188 = rob_fflags_2_1;
      5'b00010:
        casez_tmp_188 = rob_fflags_2_2;
      5'b00011:
        casez_tmp_188 = rob_fflags_2_3;
      5'b00100:
        casez_tmp_188 = rob_fflags_2_4;
      5'b00101:
        casez_tmp_188 = rob_fflags_2_5;
      5'b00110:
        casez_tmp_188 = rob_fflags_2_6;
      5'b00111:
        casez_tmp_188 = rob_fflags_2_7;
      5'b01000:
        casez_tmp_188 = rob_fflags_2_8;
      5'b01001:
        casez_tmp_188 = rob_fflags_2_9;
      5'b01010:
        casez_tmp_188 = rob_fflags_2_10;
      5'b01011:
        casez_tmp_188 = rob_fflags_2_11;
      5'b01100:
        casez_tmp_188 = rob_fflags_2_12;
      5'b01101:
        casez_tmp_188 = rob_fflags_2_13;
      5'b01110:
        casez_tmp_188 = rob_fflags_2_14;
      5'b01111:
        casez_tmp_188 = rob_fflags_2_15;
      5'b10000:
        casez_tmp_188 = rob_fflags_2_16;
      5'b10001:
        casez_tmp_188 = rob_fflags_2_17;
      5'b10010:
        casez_tmp_188 = rob_fflags_2_18;
      5'b10011:
        casez_tmp_188 = rob_fflags_2_19;
      5'b10100:
        casez_tmp_188 = rob_fflags_2_20;
      5'b10101:
        casez_tmp_188 = rob_fflags_2_21;
      5'b10110:
        casez_tmp_188 = rob_fflags_2_22;
      5'b10111:
        casez_tmp_188 = rob_fflags_2_23;
      5'b11000:
        casez_tmp_188 = rob_fflags_2_24;
      5'b11001:
        casez_tmp_188 = rob_fflags_2_25;
      5'b11010:
        casez_tmp_188 = rob_fflags_2_26;
      5'b11011:
        casez_tmp_188 = rob_fflags_2_27;
      5'b11100:
        casez_tmp_188 = rob_fflags_2_28;
      5'b11101:
        casez_tmp_188 = rob_fflags_2_29;
      5'b11110:
        casez_tmp_188 = rob_fflags_2_30;
      default:
        casez_tmp_188 = rob_fflags_2_31;
    endcase
  end // always @(*)
  reg         casez_tmp_189;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_189 = rob_uop_2_0_uses_ldq;
      5'b00001:
        casez_tmp_189 = rob_uop_2_1_uses_ldq;
      5'b00010:
        casez_tmp_189 = rob_uop_2_2_uses_ldq;
      5'b00011:
        casez_tmp_189 = rob_uop_2_3_uses_ldq;
      5'b00100:
        casez_tmp_189 = rob_uop_2_4_uses_ldq;
      5'b00101:
        casez_tmp_189 = rob_uop_2_5_uses_ldq;
      5'b00110:
        casez_tmp_189 = rob_uop_2_6_uses_ldq;
      5'b00111:
        casez_tmp_189 = rob_uop_2_7_uses_ldq;
      5'b01000:
        casez_tmp_189 = rob_uop_2_8_uses_ldq;
      5'b01001:
        casez_tmp_189 = rob_uop_2_9_uses_ldq;
      5'b01010:
        casez_tmp_189 = rob_uop_2_10_uses_ldq;
      5'b01011:
        casez_tmp_189 = rob_uop_2_11_uses_ldq;
      5'b01100:
        casez_tmp_189 = rob_uop_2_12_uses_ldq;
      5'b01101:
        casez_tmp_189 = rob_uop_2_13_uses_ldq;
      5'b01110:
        casez_tmp_189 = rob_uop_2_14_uses_ldq;
      5'b01111:
        casez_tmp_189 = rob_uop_2_15_uses_ldq;
      5'b10000:
        casez_tmp_189 = rob_uop_2_16_uses_ldq;
      5'b10001:
        casez_tmp_189 = rob_uop_2_17_uses_ldq;
      5'b10010:
        casez_tmp_189 = rob_uop_2_18_uses_ldq;
      5'b10011:
        casez_tmp_189 = rob_uop_2_19_uses_ldq;
      5'b10100:
        casez_tmp_189 = rob_uop_2_20_uses_ldq;
      5'b10101:
        casez_tmp_189 = rob_uop_2_21_uses_ldq;
      5'b10110:
        casez_tmp_189 = rob_uop_2_22_uses_ldq;
      5'b10111:
        casez_tmp_189 = rob_uop_2_23_uses_ldq;
      5'b11000:
        casez_tmp_189 = rob_uop_2_24_uses_ldq;
      5'b11001:
        casez_tmp_189 = rob_uop_2_25_uses_ldq;
      5'b11010:
        casez_tmp_189 = rob_uop_2_26_uses_ldq;
      5'b11011:
        casez_tmp_189 = rob_uop_2_27_uses_ldq;
      5'b11100:
        casez_tmp_189 = rob_uop_2_28_uses_ldq;
      5'b11101:
        casez_tmp_189 = rob_uop_2_29_uses_ldq;
      5'b11110:
        casez_tmp_189 = rob_uop_2_30_uses_ldq;
      default:
        casez_tmp_189 = rob_uop_2_31_uses_ldq;
    endcase
  end // always @(*)
  reg         casez_tmp_190;
  always @(*) begin
    casez (rob_pnr)
      5'b00000:
        casez_tmp_190 = rob_unsafe_2_0;
      5'b00001:
        casez_tmp_190 = rob_unsafe_2_1;
      5'b00010:
        casez_tmp_190 = rob_unsafe_2_2;
      5'b00011:
        casez_tmp_190 = rob_unsafe_2_3;
      5'b00100:
        casez_tmp_190 = rob_unsafe_2_4;
      5'b00101:
        casez_tmp_190 = rob_unsafe_2_5;
      5'b00110:
        casez_tmp_190 = rob_unsafe_2_6;
      5'b00111:
        casez_tmp_190 = rob_unsafe_2_7;
      5'b01000:
        casez_tmp_190 = rob_unsafe_2_8;
      5'b01001:
        casez_tmp_190 = rob_unsafe_2_9;
      5'b01010:
        casez_tmp_190 = rob_unsafe_2_10;
      5'b01011:
        casez_tmp_190 = rob_unsafe_2_11;
      5'b01100:
        casez_tmp_190 = rob_unsafe_2_12;
      5'b01101:
        casez_tmp_190 = rob_unsafe_2_13;
      5'b01110:
        casez_tmp_190 = rob_unsafe_2_14;
      5'b01111:
        casez_tmp_190 = rob_unsafe_2_15;
      5'b10000:
        casez_tmp_190 = rob_unsafe_2_16;
      5'b10001:
        casez_tmp_190 = rob_unsafe_2_17;
      5'b10010:
        casez_tmp_190 = rob_unsafe_2_18;
      5'b10011:
        casez_tmp_190 = rob_unsafe_2_19;
      5'b10100:
        casez_tmp_190 = rob_unsafe_2_20;
      5'b10101:
        casez_tmp_190 = rob_unsafe_2_21;
      5'b10110:
        casez_tmp_190 = rob_unsafe_2_22;
      5'b10111:
        casez_tmp_190 = rob_unsafe_2_23;
      5'b11000:
        casez_tmp_190 = rob_unsafe_2_24;
      5'b11001:
        casez_tmp_190 = rob_unsafe_2_25;
      5'b11010:
        casez_tmp_190 = rob_unsafe_2_26;
      5'b11011:
        casez_tmp_190 = rob_unsafe_2_27;
      5'b11100:
        casez_tmp_190 = rob_unsafe_2_28;
      5'b11101:
        casez_tmp_190 = rob_unsafe_2_29;
      5'b11110:
        casez_tmp_190 = rob_unsafe_2_30;
      default:
        casez_tmp_190 = rob_unsafe_2_31;
    endcase
  end // always @(*)
  reg         casez_tmp_191;
  always @(*) begin
    casez (rob_pnr)
      5'b00000:
        casez_tmp_191 = rob_exception_2_0;
      5'b00001:
        casez_tmp_191 = rob_exception_2_1;
      5'b00010:
        casez_tmp_191 = rob_exception_2_2;
      5'b00011:
        casez_tmp_191 = rob_exception_2_3;
      5'b00100:
        casez_tmp_191 = rob_exception_2_4;
      5'b00101:
        casez_tmp_191 = rob_exception_2_5;
      5'b00110:
        casez_tmp_191 = rob_exception_2_6;
      5'b00111:
        casez_tmp_191 = rob_exception_2_7;
      5'b01000:
        casez_tmp_191 = rob_exception_2_8;
      5'b01001:
        casez_tmp_191 = rob_exception_2_9;
      5'b01010:
        casez_tmp_191 = rob_exception_2_10;
      5'b01011:
        casez_tmp_191 = rob_exception_2_11;
      5'b01100:
        casez_tmp_191 = rob_exception_2_12;
      5'b01101:
        casez_tmp_191 = rob_exception_2_13;
      5'b01110:
        casez_tmp_191 = rob_exception_2_14;
      5'b01111:
        casez_tmp_191 = rob_exception_2_15;
      5'b10000:
        casez_tmp_191 = rob_exception_2_16;
      5'b10001:
        casez_tmp_191 = rob_exception_2_17;
      5'b10010:
        casez_tmp_191 = rob_exception_2_18;
      5'b10011:
        casez_tmp_191 = rob_exception_2_19;
      5'b10100:
        casez_tmp_191 = rob_exception_2_20;
      5'b10101:
        casez_tmp_191 = rob_exception_2_21;
      5'b10110:
        casez_tmp_191 = rob_exception_2_22;
      5'b10111:
        casez_tmp_191 = rob_exception_2_23;
      5'b11000:
        casez_tmp_191 = rob_exception_2_24;
      5'b11001:
        casez_tmp_191 = rob_exception_2_25;
      5'b11010:
        casez_tmp_191 = rob_exception_2_26;
      5'b11011:
        casez_tmp_191 = rob_exception_2_27;
      5'b11100:
        casez_tmp_191 = rob_exception_2_28;
      5'b11101:
        casez_tmp_191 = rob_exception_2_29;
      5'b11110:
        casez_tmp_191 = rob_exception_2_30;
      default:
        casez_tmp_191 = rob_exception_2_31;
    endcase
  end // always @(*)
  reg         casez_tmp_192;
  always @(*) begin
    casez (rob_pnr)
      5'b00000:
        casez_tmp_192 = rob_val_2_0;
      5'b00001:
        casez_tmp_192 = rob_val_2_1;
      5'b00010:
        casez_tmp_192 = rob_val_2_2;
      5'b00011:
        casez_tmp_192 = rob_val_2_3;
      5'b00100:
        casez_tmp_192 = rob_val_2_4;
      5'b00101:
        casez_tmp_192 = rob_val_2_5;
      5'b00110:
        casez_tmp_192 = rob_val_2_6;
      5'b00111:
        casez_tmp_192 = rob_val_2_7;
      5'b01000:
        casez_tmp_192 = rob_val_2_8;
      5'b01001:
        casez_tmp_192 = rob_val_2_9;
      5'b01010:
        casez_tmp_192 = rob_val_2_10;
      5'b01011:
        casez_tmp_192 = rob_val_2_11;
      5'b01100:
        casez_tmp_192 = rob_val_2_12;
      5'b01101:
        casez_tmp_192 = rob_val_2_13;
      5'b01110:
        casez_tmp_192 = rob_val_2_14;
      5'b01111:
        casez_tmp_192 = rob_val_2_15;
      5'b10000:
        casez_tmp_192 = rob_val_2_16;
      5'b10001:
        casez_tmp_192 = rob_val_2_17;
      5'b10010:
        casez_tmp_192 = rob_val_2_18;
      5'b10011:
        casez_tmp_192 = rob_val_2_19;
      5'b10100:
        casez_tmp_192 = rob_val_2_20;
      5'b10101:
        casez_tmp_192 = rob_val_2_21;
      5'b10110:
        casez_tmp_192 = rob_val_2_22;
      5'b10111:
        casez_tmp_192 = rob_val_2_23;
      5'b11000:
        casez_tmp_192 = rob_val_2_24;
      5'b11001:
        casez_tmp_192 = rob_val_2_25;
      5'b11010:
        casez_tmp_192 = rob_val_2_26;
      5'b11011:
        casez_tmp_192 = rob_val_2_27;
      5'b11100:
        casez_tmp_192 = rob_val_2_28;
      5'b11101:
        casez_tmp_192 = rob_val_2_29;
      5'b11110:
        casez_tmp_192 = rob_val_2_30;
      default:
        casez_tmp_192 = rob_val_2_31;
    endcase
  end // always @(*)
  reg         casez_tmp_193;
  always @(*) begin
    casez (io_wb_resps_0_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_193 = rob_val_2_0;
      5'b00001:
        casez_tmp_193 = rob_val_2_1;
      5'b00010:
        casez_tmp_193 = rob_val_2_2;
      5'b00011:
        casez_tmp_193 = rob_val_2_3;
      5'b00100:
        casez_tmp_193 = rob_val_2_4;
      5'b00101:
        casez_tmp_193 = rob_val_2_5;
      5'b00110:
        casez_tmp_193 = rob_val_2_6;
      5'b00111:
        casez_tmp_193 = rob_val_2_7;
      5'b01000:
        casez_tmp_193 = rob_val_2_8;
      5'b01001:
        casez_tmp_193 = rob_val_2_9;
      5'b01010:
        casez_tmp_193 = rob_val_2_10;
      5'b01011:
        casez_tmp_193 = rob_val_2_11;
      5'b01100:
        casez_tmp_193 = rob_val_2_12;
      5'b01101:
        casez_tmp_193 = rob_val_2_13;
      5'b01110:
        casez_tmp_193 = rob_val_2_14;
      5'b01111:
        casez_tmp_193 = rob_val_2_15;
      5'b10000:
        casez_tmp_193 = rob_val_2_16;
      5'b10001:
        casez_tmp_193 = rob_val_2_17;
      5'b10010:
        casez_tmp_193 = rob_val_2_18;
      5'b10011:
        casez_tmp_193 = rob_val_2_19;
      5'b10100:
        casez_tmp_193 = rob_val_2_20;
      5'b10101:
        casez_tmp_193 = rob_val_2_21;
      5'b10110:
        casez_tmp_193 = rob_val_2_22;
      5'b10111:
        casez_tmp_193 = rob_val_2_23;
      5'b11000:
        casez_tmp_193 = rob_val_2_24;
      5'b11001:
        casez_tmp_193 = rob_val_2_25;
      5'b11010:
        casez_tmp_193 = rob_val_2_26;
      5'b11011:
        casez_tmp_193 = rob_val_2_27;
      5'b11100:
        casez_tmp_193 = rob_val_2_28;
      5'b11101:
        casez_tmp_193 = rob_val_2_29;
      5'b11110:
        casez_tmp_193 = rob_val_2_30;
      default:
        casez_tmp_193 = rob_val_2_31;
    endcase
  end // always @(*)
  reg         casez_tmp_194;
  always @(*) begin
    casez (io_wb_resps_0_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_194 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_194 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_194 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_194 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_194 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_194 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_194 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_194 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_194 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_194 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_194 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_194 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_194 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_194 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_194 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_194 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_194 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_194 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_194 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_194 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_194 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_194 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_194 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_194 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_194 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_194 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_194 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_194 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_194 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_194 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_194 = rob_bsy_2_30;
      default:
        casez_tmp_194 = rob_bsy_2_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_195;
  always @(*) begin
    casez (io_wb_resps_0_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_195 = rob_uop_2_0_pdst;
      5'b00001:
        casez_tmp_195 = rob_uop_2_1_pdst;
      5'b00010:
        casez_tmp_195 = rob_uop_2_2_pdst;
      5'b00011:
        casez_tmp_195 = rob_uop_2_3_pdst;
      5'b00100:
        casez_tmp_195 = rob_uop_2_4_pdst;
      5'b00101:
        casez_tmp_195 = rob_uop_2_5_pdst;
      5'b00110:
        casez_tmp_195 = rob_uop_2_6_pdst;
      5'b00111:
        casez_tmp_195 = rob_uop_2_7_pdst;
      5'b01000:
        casez_tmp_195 = rob_uop_2_8_pdst;
      5'b01001:
        casez_tmp_195 = rob_uop_2_9_pdst;
      5'b01010:
        casez_tmp_195 = rob_uop_2_10_pdst;
      5'b01011:
        casez_tmp_195 = rob_uop_2_11_pdst;
      5'b01100:
        casez_tmp_195 = rob_uop_2_12_pdst;
      5'b01101:
        casez_tmp_195 = rob_uop_2_13_pdst;
      5'b01110:
        casez_tmp_195 = rob_uop_2_14_pdst;
      5'b01111:
        casez_tmp_195 = rob_uop_2_15_pdst;
      5'b10000:
        casez_tmp_195 = rob_uop_2_16_pdst;
      5'b10001:
        casez_tmp_195 = rob_uop_2_17_pdst;
      5'b10010:
        casez_tmp_195 = rob_uop_2_18_pdst;
      5'b10011:
        casez_tmp_195 = rob_uop_2_19_pdst;
      5'b10100:
        casez_tmp_195 = rob_uop_2_20_pdst;
      5'b10101:
        casez_tmp_195 = rob_uop_2_21_pdst;
      5'b10110:
        casez_tmp_195 = rob_uop_2_22_pdst;
      5'b10111:
        casez_tmp_195 = rob_uop_2_23_pdst;
      5'b11000:
        casez_tmp_195 = rob_uop_2_24_pdst;
      5'b11001:
        casez_tmp_195 = rob_uop_2_25_pdst;
      5'b11010:
        casez_tmp_195 = rob_uop_2_26_pdst;
      5'b11011:
        casez_tmp_195 = rob_uop_2_27_pdst;
      5'b11100:
        casez_tmp_195 = rob_uop_2_28_pdst;
      5'b11101:
        casez_tmp_195 = rob_uop_2_29_pdst;
      5'b11110:
        casez_tmp_195 = rob_uop_2_30_pdst;
      default:
        casez_tmp_195 = rob_uop_2_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_196;
  always @(*) begin
    casez (io_wb_resps_0_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_196 = rob_uop_2_0_ldst_val;
      5'b00001:
        casez_tmp_196 = rob_uop_2_1_ldst_val;
      5'b00010:
        casez_tmp_196 = rob_uop_2_2_ldst_val;
      5'b00011:
        casez_tmp_196 = rob_uop_2_3_ldst_val;
      5'b00100:
        casez_tmp_196 = rob_uop_2_4_ldst_val;
      5'b00101:
        casez_tmp_196 = rob_uop_2_5_ldst_val;
      5'b00110:
        casez_tmp_196 = rob_uop_2_6_ldst_val;
      5'b00111:
        casez_tmp_196 = rob_uop_2_7_ldst_val;
      5'b01000:
        casez_tmp_196 = rob_uop_2_8_ldst_val;
      5'b01001:
        casez_tmp_196 = rob_uop_2_9_ldst_val;
      5'b01010:
        casez_tmp_196 = rob_uop_2_10_ldst_val;
      5'b01011:
        casez_tmp_196 = rob_uop_2_11_ldst_val;
      5'b01100:
        casez_tmp_196 = rob_uop_2_12_ldst_val;
      5'b01101:
        casez_tmp_196 = rob_uop_2_13_ldst_val;
      5'b01110:
        casez_tmp_196 = rob_uop_2_14_ldst_val;
      5'b01111:
        casez_tmp_196 = rob_uop_2_15_ldst_val;
      5'b10000:
        casez_tmp_196 = rob_uop_2_16_ldst_val;
      5'b10001:
        casez_tmp_196 = rob_uop_2_17_ldst_val;
      5'b10010:
        casez_tmp_196 = rob_uop_2_18_ldst_val;
      5'b10011:
        casez_tmp_196 = rob_uop_2_19_ldst_val;
      5'b10100:
        casez_tmp_196 = rob_uop_2_20_ldst_val;
      5'b10101:
        casez_tmp_196 = rob_uop_2_21_ldst_val;
      5'b10110:
        casez_tmp_196 = rob_uop_2_22_ldst_val;
      5'b10111:
        casez_tmp_196 = rob_uop_2_23_ldst_val;
      5'b11000:
        casez_tmp_196 = rob_uop_2_24_ldst_val;
      5'b11001:
        casez_tmp_196 = rob_uop_2_25_ldst_val;
      5'b11010:
        casez_tmp_196 = rob_uop_2_26_ldst_val;
      5'b11011:
        casez_tmp_196 = rob_uop_2_27_ldst_val;
      5'b11100:
        casez_tmp_196 = rob_uop_2_28_ldst_val;
      5'b11101:
        casez_tmp_196 = rob_uop_2_29_ldst_val;
      5'b11110:
        casez_tmp_196 = rob_uop_2_30_ldst_val;
      default:
        casez_tmp_196 = rob_uop_2_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_197;
  always @(*) begin
    casez (io_wb_resps_1_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_197 = rob_val_2_0;
      5'b00001:
        casez_tmp_197 = rob_val_2_1;
      5'b00010:
        casez_tmp_197 = rob_val_2_2;
      5'b00011:
        casez_tmp_197 = rob_val_2_3;
      5'b00100:
        casez_tmp_197 = rob_val_2_4;
      5'b00101:
        casez_tmp_197 = rob_val_2_5;
      5'b00110:
        casez_tmp_197 = rob_val_2_6;
      5'b00111:
        casez_tmp_197 = rob_val_2_7;
      5'b01000:
        casez_tmp_197 = rob_val_2_8;
      5'b01001:
        casez_tmp_197 = rob_val_2_9;
      5'b01010:
        casez_tmp_197 = rob_val_2_10;
      5'b01011:
        casez_tmp_197 = rob_val_2_11;
      5'b01100:
        casez_tmp_197 = rob_val_2_12;
      5'b01101:
        casez_tmp_197 = rob_val_2_13;
      5'b01110:
        casez_tmp_197 = rob_val_2_14;
      5'b01111:
        casez_tmp_197 = rob_val_2_15;
      5'b10000:
        casez_tmp_197 = rob_val_2_16;
      5'b10001:
        casez_tmp_197 = rob_val_2_17;
      5'b10010:
        casez_tmp_197 = rob_val_2_18;
      5'b10011:
        casez_tmp_197 = rob_val_2_19;
      5'b10100:
        casez_tmp_197 = rob_val_2_20;
      5'b10101:
        casez_tmp_197 = rob_val_2_21;
      5'b10110:
        casez_tmp_197 = rob_val_2_22;
      5'b10111:
        casez_tmp_197 = rob_val_2_23;
      5'b11000:
        casez_tmp_197 = rob_val_2_24;
      5'b11001:
        casez_tmp_197 = rob_val_2_25;
      5'b11010:
        casez_tmp_197 = rob_val_2_26;
      5'b11011:
        casez_tmp_197 = rob_val_2_27;
      5'b11100:
        casez_tmp_197 = rob_val_2_28;
      5'b11101:
        casez_tmp_197 = rob_val_2_29;
      5'b11110:
        casez_tmp_197 = rob_val_2_30;
      default:
        casez_tmp_197 = rob_val_2_31;
    endcase
  end // always @(*)
  reg         casez_tmp_198;
  always @(*) begin
    casez (io_wb_resps_1_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_198 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_198 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_198 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_198 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_198 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_198 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_198 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_198 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_198 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_198 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_198 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_198 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_198 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_198 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_198 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_198 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_198 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_198 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_198 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_198 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_198 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_198 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_198 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_198 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_198 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_198 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_198 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_198 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_198 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_198 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_198 = rob_bsy_2_30;
      default:
        casez_tmp_198 = rob_bsy_2_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_199;
  always @(*) begin
    casez (io_wb_resps_1_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_199 = rob_uop_2_0_pdst;
      5'b00001:
        casez_tmp_199 = rob_uop_2_1_pdst;
      5'b00010:
        casez_tmp_199 = rob_uop_2_2_pdst;
      5'b00011:
        casez_tmp_199 = rob_uop_2_3_pdst;
      5'b00100:
        casez_tmp_199 = rob_uop_2_4_pdst;
      5'b00101:
        casez_tmp_199 = rob_uop_2_5_pdst;
      5'b00110:
        casez_tmp_199 = rob_uop_2_6_pdst;
      5'b00111:
        casez_tmp_199 = rob_uop_2_7_pdst;
      5'b01000:
        casez_tmp_199 = rob_uop_2_8_pdst;
      5'b01001:
        casez_tmp_199 = rob_uop_2_9_pdst;
      5'b01010:
        casez_tmp_199 = rob_uop_2_10_pdst;
      5'b01011:
        casez_tmp_199 = rob_uop_2_11_pdst;
      5'b01100:
        casez_tmp_199 = rob_uop_2_12_pdst;
      5'b01101:
        casez_tmp_199 = rob_uop_2_13_pdst;
      5'b01110:
        casez_tmp_199 = rob_uop_2_14_pdst;
      5'b01111:
        casez_tmp_199 = rob_uop_2_15_pdst;
      5'b10000:
        casez_tmp_199 = rob_uop_2_16_pdst;
      5'b10001:
        casez_tmp_199 = rob_uop_2_17_pdst;
      5'b10010:
        casez_tmp_199 = rob_uop_2_18_pdst;
      5'b10011:
        casez_tmp_199 = rob_uop_2_19_pdst;
      5'b10100:
        casez_tmp_199 = rob_uop_2_20_pdst;
      5'b10101:
        casez_tmp_199 = rob_uop_2_21_pdst;
      5'b10110:
        casez_tmp_199 = rob_uop_2_22_pdst;
      5'b10111:
        casez_tmp_199 = rob_uop_2_23_pdst;
      5'b11000:
        casez_tmp_199 = rob_uop_2_24_pdst;
      5'b11001:
        casez_tmp_199 = rob_uop_2_25_pdst;
      5'b11010:
        casez_tmp_199 = rob_uop_2_26_pdst;
      5'b11011:
        casez_tmp_199 = rob_uop_2_27_pdst;
      5'b11100:
        casez_tmp_199 = rob_uop_2_28_pdst;
      5'b11101:
        casez_tmp_199 = rob_uop_2_29_pdst;
      5'b11110:
        casez_tmp_199 = rob_uop_2_30_pdst;
      default:
        casez_tmp_199 = rob_uop_2_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_200;
  always @(*) begin
    casez (io_wb_resps_1_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_200 = rob_uop_2_0_ldst_val;
      5'b00001:
        casez_tmp_200 = rob_uop_2_1_ldst_val;
      5'b00010:
        casez_tmp_200 = rob_uop_2_2_ldst_val;
      5'b00011:
        casez_tmp_200 = rob_uop_2_3_ldst_val;
      5'b00100:
        casez_tmp_200 = rob_uop_2_4_ldst_val;
      5'b00101:
        casez_tmp_200 = rob_uop_2_5_ldst_val;
      5'b00110:
        casez_tmp_200 = rob_uop_2_6_ldst_val;
      5'b00111:
        casez_tmp_200 = rob_uop_2_7_ldst_val;
      5'b01000:
        casez_tmp_200 = rob_uop_2_8_ldst_val;
      5'b01001:
        casez_tmp_200 = rob_uop_2_9_ldst_val;
      5'b01010:
        casez_tmp_200 = rob_uop_2_10_ldst_val;
      5'b01011:
        casez_tmp_200 = rob_uop_2_11_ldst_val;
      5'b01100:
        casez_tmp_200 = rob_uop_2_12_ldst_val;
      5'b01101:
        casez_tmp_200 = rob_uop_2_13_ldst_val;
      5'b01110:
        casez_tmp_200 = rob_uop_2_14_ldst_val;
      5'b01111:
        casez_tmp_200 = rob_uop_2_15_ldst_val;
      5'b10000:
        casez_tmp_200 = rob_uop_2_16_ldst_val;
      5'b10001:
        casez_tmp_200 = rob_uop_2_17_ldst_val;
      5'b10010:
        casez_tmp_200 = rob_uop_2_18_ldst_val;
      5'b10011:
        casez_tmp_200 = rob_uop_2_19_ldst_val;
      5'b10100:
        casez_tmp_200 = rob_uop_2_20_ldst_val;
      5'b10101:
        casez_tmp_200 = rob_uop_2_21_ldst_val;
      5'b10110:
        casez_tmp_200 = rob_uop_2_22_ldst_val;
      5'b10111:
        casez_tmp_200 = rob_uop_2_23_ldst_val;
      5'b11000:
        casez_tmp_200 = rob_uop_2_24_ldst_val;
      5'b11001:
        casez_tmp_200 = rob_uop_2_25_ldst_val;
      5'b11010:
        casez_tmp_200 = rob_uop_2_26_ldst_val;
      5'b11011:
        casez_tmp_200 = rob_uop_2_27_ldst_val;
      5'b11100:
        casez_tmp_200 = rob_uop_2_28_ldst_val;
      5'b11101:
        casez_tmp_200 = rob_uop_2_29_ldst_val;
      5'b11110:
        casez_tmp_200 = rob_uop_2_30_ldst_val;
      default:
        casez_tmp_200 = rob_uop_2_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_201;
  always @(*) begin
    casez (io_wb_resps_2_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_201 = rob_val_2_0;
      5'b00001:
        casez_tmp_201 = rob_val_2_1;
      5'b00010:
        casez_tmp_201 = rob_val_2_2;
      5'b00011:
        casez_tmp_201 = rob_val_2_3;
      5'b00100:
        casez_tmp_201 = rob_val_2_4;
      5'b00101:
        casez_tmp_201 = rob_val_2_5;
      5'b00110:
        casez_tmp_201 = rob_val_2_6;
      5'b00111:
        casez_tmp_201 = rob_val_2_7;
      5'b01000:
        casez_tmp_201 = rob_val_2_8;
      5'b01001:
        casez_tmp_201 = rob_val_2_9;
      5'b01010:
        casez_tmp_201 = rob_val_2_10;
      5'b01011:
        casez_tmp_201 = rob_val_2_11;
      5'b01100:
        casez_tmp_201 = rob_val_2_12;
      5'b01101:
        casez_tmp_201 = rob_val_2_13;
      5'b01110:
        casez_tmp_201 = rob_val_2_14;
      5'b01111:
        casez_tmp_201 = rob_val_2_15;
      5'b10000:
        casez_tmp_201 = rob_val_2_16;
      5'b10001:
        casez_tmp_201 = rob_val_2_17;
      5'b10010:
        casez_tmp_201 = rob_val_2_18;
      5'b10011:
        casez_tmp_201 = rob_val_2_19;
      5'b10100:
        casez_tmp_201 = rob_val_2_20;
      5'b10101:
        casez_tmp_201 = rob_val_2_21;
      5'b10110:
        casez_tmp_201 = rob_val_2_22;
      5'b10111:
        casez_tmp_201 = rob_val_2_23;
      5'b11000:
        casez_tmp_201 = rob_val_2_24;
      5'b11001:
        casez_tmp_201 = rob_val_2_25;
      5'b11010:
        casez_tmp_201 = rob_val_2_26;
      5'b11011:
        casez_tmp_201 = rob_val_2_27;
      5'b11100:
        casez_tmp_201 = rob_val_2_28;
      5'b11101:
        casez_tmp_201 = rob_val_2_29;
      5'b11110:
        casez_tmp_201 = rob_val_2_30;
      default:
        casez_tmp_201 = rob_val_2_31;
    endcase
  end // always @(*)
  reg         casez_tmp_202;
  always @(*) begin
    casez (io_wb_resps_2_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_202 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_202 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_202 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_202 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_202 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_202 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_202 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_202 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_202 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_202 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_202 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_202 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_202 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_202 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_202 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_202 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_202 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_202 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_202 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_202 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_202 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_202 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_202 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_202 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_202 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_202 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_202 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_202 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_202 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_202 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_202 = rob_bsy_2_30;
      default:
        casez_tmp_202 = rob_bsy_2_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_203;
  always @(*) begin
    casez (io_wb_resps_2_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_203 = rob_uop_2_0_pdst;
      5'b00001:
        casez_tmp_203 = rob_uop_2_1_pdst;
      5'b00010:
        casez_tmp_203 = rob_uop_2_2_pdst;
      5'b00011:
        casez_tmp_203 = rob_uop_2_3_pdst;
      5'b00100:
        casez_tmp_203 = rob_uop_2_4_pdst;
      5'b00101:
        casez_tmp_203 = rob_uop_2_5_pdst;
      5'b00110:
        casez_tmp_203 = rob_uop_2_6_pdst;
      5'b00111:
        casez_tmp_203 = rob_uop_2_7_pdst;
      5'b01000:
        casez_tmp_203 = rob_uop_2_8_pdst;
      5'b01001:
        casez_tmp_203 = rob_uop_2_9_pdst;
      5'b01010:
        casez_tmp_203 = rob_uop_2_10_pdst;
      5'b01011:
        casez_tmp_203 = rob_uop_2_11_pdst;
      5'b01100:
        casez_tmp_203 = rob_uop_2_12_pdst;
      5'b01101:
        casez_tmp_203 = rob_uop_2_13_pdst;
      5'b01110:
        casez_tmp_203 = rob_uop_2_14_pdst;
      5'b01111:
        casez_tmp_203 = rob_uop_2_15_pdst;
      5'b10000:
        casez_tmp_203 = rob_uop_2_16_pdst;
      5'b10001:
        casez_tmp_203 = rob_uop_2_17_pdst;
      5'b10010:
        casez_tmp_203 = rob_uop_2_18_pdst;
      5'b10011:
        casez_tmp_203 = rob_uop_2_19_pdst;
      5'b10100:
        casez_tmp_203 = rob_uop_2_20_pdst;
      5'b10101:
        casez_tmp_203 = rob_uop_2_21_pdst;
      5'b10110:
        casez_tmp_203 = rob_uop_2_22_pdst;
      5'b10111:
        casez_tmp_203 = rob_uop_2_23_pdst;
      5'b11000:
        casez_tmp_203 = rob_uop_2_24_pdst;
      5'b11001:
        casez_tmp_203 = rob_uop_2_25_pdst;
      5'b11010:
        casez_tmp_203 = rob_uop_2_26_pdst;
      5'b11011:
        casez_tmp_203 = rob_uop_2_27_pdst;
      5'b11100:
        casez_tmp_203 = rob_uop_2_28_pdst;
      5'b11101:
        casez_tmp_203 = rob_uop_2_29_pdst;
      5'b11110:
        casez_tmp_203 = rob_uop_2_30_pdst;
      default:
        casez_tmp_203 = rob_uop_2_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_204;
  always @(*) begin
    casez (io_wb_resps_2_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_204 = rob_uop_2_0_ldst_val;
      5'b00001:
        casez_tmp_204 = rob_uop_2_1_ldst_val;
      5'b00010:
        casez_tmp_204 = rob_uop_2_2_ldst_val;
      5'b00011:
        casez_tmp_204 = rob_uop_2_3_ldst_val;
      5'b00100:
        casez_tmp_204 = rob_uop_2_4_ldst_val;
      5'b00101:
        casez_tmp_204 = rob_uop_2_5_ldst_val;
      5'b00110:
        casez_tmp_204 = rob_uop_2_6_ldst_val;
      5'b00111:
        casez_tmp_204 = rob_uop_2_7_ldst_val;
      5'b01000:
        casez_tmp_204 = rob_uop_2_8_ldst_val;
      5'b01001:
        casez_tmp_204 = rob_uop_2_9_ldst_val;
      5'b01010:
        casez_tmp_204 = rob_uop_2_10_ldst_val;
      5'b01011:
        casez_tmp_204 = rob_uop_2_11_ldst_val;
      5'b01100:
        casez_tmp_204 = rob_uop_2_12_ldst_val;
      5'b01101:
        casez_tmp_204 = rob_uop_2_13_ldst_val;
      5'b01110:
        casez_tmp_204 = rob_uop_2_14_ldst_val;
      5'b01111:
        casez_tmp_204 = rob_uop_2_15_ldst_val;
      5'b10000:
        casez_tmp_204 = rob_uop_2_16_ldst_val;
      5'b10001:
        casez_tmp_204 = rob_uop_2_17_ldst_val;
      5'b10010:
        casez_tmp_204 = rob_uop_2_18_ldst_val;
      5'b10011:
        casez_tmp_204 = rob_uop_2_19_ldst_val;
      5'b10100:
        casez_tmp_204 = rob_uop_2_20_ldst_val;
      5'b10101:
        casez_tmp_204 = rob_uop_2_21_ldst_val;
      5'b10110:
        casez_tmp_204 = rob_uop_2_22_ldst_val;
      5'b10111:
        casez_tmp_204 = rob_uop_2_23_ldst_val;
      5'b11000:
        casez_tmp_204 = rob_uop_2_24_ldst_val;
      5'b11001:
        casez_tmp_204 = rob_uop_2_25_ldst_val;
      5'b11010:
        casez_tmp_204 = rob_uop_2_26_ldst_val;
      5'b11011:
        casez_tmp_204 = rob_uop_2_27_ldst_val;
      5'b11100:
        casez_tmp_204 = rob_uop_2_28_ldst_val;
      5'b11101:
        casez_tmp_204 = rob_uop_2_29_ldst_val;
      5'b11110:
        casez_tmp_204 = rob_uop_2_30_ldst_val;
      default:
        casez_tmp_204 = rob_uop_2_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_205;
  always @(*) begin
    casez (io_wb_resps_3_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_205 = rob_val_2_0;
      5'b00001:
        casez_tmp_205 = rob_val_2_1;
      5'b00010:
        casez_tmp_205 = rob_val_2_2;
      5'b00011:
        casez_tmp_205 = rob_val_2_3;
      5'b00100:
        casez_tmp_205 = rob_val_2_4;
      5'b00101:
        casez_tmp_205 = rob_val_2_5;
      5'b00110:
        casez_tmp_205 = rob_val_2_6;
      5'b00111:
        casez_tmp_205 = rob_val_2_7;
      5'b01000:
        casez_tmp_205 = rob_val_2_8;
      5'b01001:
        casez_tmp_205 = rob_val_2_9;
      5'b01010:
        casez_tmp_205 = rob_val_2_10;
      5'b01011:
        casez_tmp_205 = rob_val_2_11;
      5'b01100:
        casez_tmp_205 = rob_val_2_12;
      5'b01101:
        casez_tmp_205 = rob_val_2_13;
      5'b01110:
        casez_tmp_205 = rob_val_2_14;
      5'b01111:
        casez_tmp_205 = rob_val_2_15;
      5'b10000:
        casez_tmp_205 = rob_val_2_16;
      5'b10001:
        casez_tmp_205 = rob_val_2_17;
      5'b10010:
        casez_tmp_205 = rob_val_2_18;
      5'b10011:
        casez_tmp_205 = rob_val_2_19;
      5'b10100:
        casez_tmp_205 = rob_val_2_20;
      5'b10101:
        casez_tmp_205 = rob_val_2_21;
      5'b10110:
        casez_tmp_205 = rob_val_2_22;
      5'b10111:
        casez_tmp_205 = rob_val_2_23;
      5'b11000:
        casez_tmp_205 = rob_val_2_24;
      5'b11001:
        casez_tmp_205 = rob_val_2_25;
      5'b11010:
        casez_tmp_205 = rob_val_2_26;
      5'b11011:
        casez_tmp_205 = rob_val_2_27;
      5'b11100:
        casez_tmp_205 = rob_val_2_28;
      5'b11101:
        casez_tmp_205 = rob_val_2_29;
      5'b11110:
        casez_tmp_205 = rob_val_2_30;
      default:
        casez_tmp_205 = rob_val_2_31;
    endcase
  end // always @(*)
  reg         casez_tmp_206;
  always @(*) begin
    casez (io_wb_resps_3_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_206 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_206 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_206 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_206 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_206 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_206 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_206 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_206 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_206 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_206 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_206 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_206 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_206 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_206 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_206 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_206 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_206 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_206 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_206 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_206 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_206 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_206 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_206 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_206 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_206 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_206 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_206 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_206 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_206 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_206 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_206 = rob_bsy_2_30;
      default:
        casez_tmp_206 = rob_bsy_2_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_207;
  always @(*) begin
    casez (io_wb_resps_3_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_207 = rob_uop_2_0_pdst;
      5'b00001:
        casez_tmp_207 = rob_uop_2_1_pdst;
      5'b00010:
        casez_tmp_207 = rob_uop_2_2_pdst;
      5'b00011:
        casez_tmp_207 = rob_uop_2_3_pdst;
      5'b00100:
        casez_tmp_207 = rob_uop_2_4_pdst;
      5'b00101:
        casez_tmp_207 = rob_uop_2_5_pdst;
      5'b00110:
        casez_tmp_207 = rob_uop_2_6_pdst;
      5'b00111:
        casez_tmp_207 = rob_uop_2_7_pdst;
      5'b01000:
        casez_tmp_207 = rob_uop_2_8_pdst;
      5'b01001:
        casez_tmp_207 = rob_uop_2_9_pdst;
      5'b01010:
        casez_tmp_207 = rob_uop_2_10_pdst;
      5'b01011:
        casez_tmp_207 = rob_uop_2_11_pdst;
      5'b01100:
        casez_tmp_207 = rob_uop_2_12_pdst;
      5'b01101:
        casez_tmp_207 = rob_uop_2_13_pdst;
      5'b01110:
        casez_tmp_207 = rob_uop_2_14_pdst;
      5'b01111:
        casez_tmp_207 = rob_uop_2_15_pdst;
      5'b10000:
        casez_tmp_207 = rob_uop_2_16_pdst;
      5'b10001:
        casez_tmp_207 = rob_uop_2_17_pdst;
      5'b10010:
        casez_tmp_207 = rob_uop_2_18_pdst;
      5'b10011:
        casez_tmp_207 = rob_uop_2_19_pdst;
      5'b10100:
        casez_tmp_207 = rob_uop_2_20_pdst;
      5'b10101:
        casez_tmp_207 = rob_uop_2_21_pdst;
      5'b10110:
        casez_tmp_207 = rob_uop_2_22_pdst;
      5'b10111:
        casez_tmp_207 = rob_uop_2_23_pdst;
      5'b11000:
        casez_tmp_207 = rob_uop_2_24_pdst;
      5'b11001:
        casez_tmp_207 = rob_uop_2_25_pdst;
      5'b11010:
        casez_tmp_207 = rob_uop_2_26_pdst;
      5'b11011:
        casez_tmp_207 = rob_uop_2_27_pdst;
      5'b11100:
        casez_tmp_207 = rob_uop_2_28_pdst;
      5'b11101:
        casez_tmp_207 = rob_uop_2_29_pdst;
      5'b11110:
        casez_tmp_207 = rob_uop_2_30_pdst;
      default:
        casez_tmp_207 = rob_uop_2_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_208;
  always @(*) begin
    casez (io_wb_resps_3_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_208 = rob_uop_2_0_ldst_val;
      5'b00001:
        casez_tmp_208 = rob_uop_2_1_ldst_val;
      5'b00010:
        casez_tmp_208 = rob_uop_2_2_ldst_val;
      5'b00011:
        casez_tmp_208 = rob_uop_2_3_ldst_val;
      5'b00100:
        casez_tmp_208 = rob_uop_2_4_ldst_val;
      5'b00101:
        casez_tmp_208 = rob_uop_2_5_ldst_val;
      5'b00110:
        casez_tmp_208 = rob_uop_2_6_ldst_val;
      5'b00111:
        casez_tmp_208 = rob_uop_2_7_ldst_val;
      5'b01000:
        casez_tmp_208 = rob_uop_2_8_ldst_val;
      5'b01001:
        casez_tmp_208 = rob_uop_2_9_ldst_val;
      5'b01010:
        casez_tmp_208 = rob_uop_2_10_ldst_val;
      5'b01011:
        casez_tmp_208 = rob_uop_2_11_ldst_val;
      5'b01100:
        casez_tmp_208 = rob_uop_2_12_ldst_val;
      5'b01101:
        casez_tmp_208 = rob_uop_2_13_ldst_val;
      5'b01110:
        casez_tmp_208 = rob_uop_2_14_ldst_val;
      5'b01111:
        casez_tmp_208 = rob_uop_2_15_ldst_val;
      5'b10000:
        casez_tmp_208 = rob_uop_2_16_ldst_val;
      5'b10001:
        casez_tmp_208 = rob_uop_2_17_ldst_val;
      5'b10010:
        casez_tmp_208 = rob_uop_2_18_ldst_val;
      5'b10011:
        casez_tmp_208 = rob_uop_2_19_ldst_val;
      5'b10100:
        casez_tmp_208 = rob_uop_2_20_ldst_val;
      5'b10101:
        casez_tmp_208 = rob_uop_2_21_ldst_val;
      5'b10110:
        casez_tmp_208 = rob_uop_2_22_ldst_val;
      5'b10111:
        casez_tmp_208 = rob_uop_2_23_ldst_val;
      5'b11000:
        casez_tmp_208 = rob_uop_2_24_ldst_val;
      5'b11001:
        casez_tmp_208 = rob_uop_2_25_ldst_val;
      5'b11010:
        casez_tmp_208 = rob_uop_2_26_ldst_val;
      5'b11011:
        casez_tmp_208 = rob_uop_2_27_ldst_val;
      5'b11100:
        casez_tmp_208 = rob_uop_2_28_ldst_val;
      5'b11101:
        casez_tmp_208 = rob_uop_2_29_ldst_val;
      5'b11110:
        casez_tmp_208 = rob_uop_2_30_ldst_val;
      default:
        casez_tmp_208 = rob_uop_2_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_209;
  always @(*) begin
    casez (io_wb_resps_4_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_209 = rob_val_2_0;
      5'b00001:
        casez_tmp_209 = rob_val_2_1;
      5'b00010:
        casez_tmp_209 = rob_val_2_2;
      5'b00011:
        casez_tmp_209 = rob_val_2_3;
      5'b00100:
        casez_tmp_209 = rob_val_2_4;
      5'b00101:
        casez_tmp_209 = rob_val_2_5;
      5'b00110:
        casez_tmp_209 = rob_val_2_6;
      5'b00111:
        casez_tmp_209 = rob_val_2_7;
      5'b01000:
        casez_tmp_209 = rob_val_2_8;
      5'b01001:
        casez_tmp_209 = rob_val_2_9;
      5'b01010:
        casez_tmp_209 = rob_val_2_10;
      5'b01011:
        casez_tmp_209 = rob_val_2_11;
      5'b01100:
        casez_tmp_209 = rob_val_2_12;
      5'b01101:
        casez_tmp_209 = rob_val_2_13;
      5'b01110:
        casez_tmp_209 = rob_val_2_14;
      5'b01111:
        casez_tmp_209 = rob_val_2_15;
      5'b10000:
        casez_tmp_209 = rob_val_2_16;
      5'b10001:
        casez_tmp_209 = rob_val_2_17;
      5'b10010:
        casez_tmp_209 = rob_val_2_18;
      5'b10011:
        casez_tmp_209 = rob_val_2_19;
      5'b10100:
        casez_tmp_209 = rob_val_2_20;
      5'b10101:
        casez_tmp_209 = rob_val_2_21;
      5'b10110:
        casez_tmp_209 = rob_val_2_22;
      5'b10111:
        casez_tmp_209 = rob_val_2_23;
      5'b11000:
        casez_tmp_209 = rob_val_2_24;
      5'b11001:
        casez_tmp_209 = rob_val_2_25;
      5'b11010:
        casez_tmp_209 = rob_val_2_26;
      5'b11011:
        casez_tmp_209 = rob_val_2_27;
      5'b11100:
        casez_tmp_209 = rob_val_2_28;
      5'b11101:
        casez_tmp_209 = rob_val_2_29;
      5'b11110:
        casez_tmp_209 = rob_val_2_30;
      default:
        casez_tmp_209 = rob_val_2_31;
    endcase
  end // always @(*)
  reg         casez_tmp_210;
  always @(*) begin
    casez (io_wb_resps_4_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_210 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_210 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_210 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_210 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_210 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_210 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_210 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_210 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_210 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_210 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_210 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_210 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_210 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_210 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_210 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_210 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_210 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_210 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_210 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_210 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_210 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_210 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_210 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_210 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_210 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_210 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_210 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_210 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_210 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_210 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_210 = rob_bsy_2_30;
      default:
        casez_tmp_210 = rob_bsy_2_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_211;
  always @(*) begin
    casez (io_wb_resps_4_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_211 = rob_uop_2_0_pdst;
      5'b00001:
        casez_tmp_211 = rob_uop_2_1_pdst;
      5'b00010:
        casez_tmp_211 = rob_uop_2_2_pdst;
      5'b00011:
        casez_tmp_211 = rob_uop_2_3_pdst;
      5'b00100:
        casez_tmp_211 = rob_uop_2_4_pdst;
      5'b00101:
        casez_tmp_211 = rob_uop_2_5_pdst;
      5'b00110:
        casez_tmp_211 = rob_uop_2_6_pdst;
      5'b00111:
        casez_tmp_211 = rob_uop_2_7_pdst;
      5'b01000:
        casez_tmp_211 = rob_uop_2_8_pdst;
      5'b01001:
        casez_tmp_211 = rob_uop_2_9_pdst;
      5'b01010:
        casez_tmp_211 = rob_uop_2_10_pdst;
      5'b01011:
        casez_tmp_211 = rob_uop_2_11_pdst;
      5'b01100:
        casez_tmp_211 = rob_uop_2_12_pdst;
      5'b01101:
        casez_tmp_211 = rob_uop_2_13_pdst;
      5'b01110:
        casez_tmp_211 = rob_uop_2_14_pdst;
      5'b01111:
        casez_tmp_211 = rob_uop_2_15_pdst;
      5'b10000:
        casez_tmp_211 = rob_uop_2_16_pdst;
      5'b10001:
        casez_tmp_211 = rob_uop_2_17_pdst;
      5'b10010:
        casez_tmp_211 = rob_uop_2_18_pdst;
      5'b10011:
        casez_tmp_211 = rob_uop_2_19_pdst;
      5'b10100:
        casez_tmp_211 = rob_uop_2_20_pdst;
      5'b10101:
        casez_tmp_211 = rob_uop_2_21_pdst;
      5'b10110:
        casez_tmp_211 = rob_uop_2_22_pdst;
      5'b10111:
        casez_tmp_211 = rob_uop_2_23_pdst;
      5'b11000:
        casez_tmp_211 = rob_uop_2_24_pdst;
      5'b11001:
        casez_tmp_211 = rob_uop_2_25_pdst;
      5'b11010:
        casez_tmp_211 = rob_uop_2_26_pdst;
      5'b11011:
        casez_tmp_211 = rob_uop_2_27_pdst;
      5'b11100:
        casez_tmp_211 = rob_uop_2_28_pdst;
      5'b11101:
        casez_tmp_211 = rob_uop_2_29_pdst;
      5'b11110:
        casez_tmp_211 = rob_uop_2_30_pdst;
      default:
        casez_tmp_211 = rob_uop_2_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_212;
  always @(*) begin
    casez (io_wb_resps_4_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_212 = rob_uop_2_0_ldst_val;
      5'b00001:
        casez_tmp_212 = rob_uop_2_1_ldst_val;
      5'b00010:
        casez_tmp_212 = rob_uop_2_2_ldst_val;
      5'b00011:
        casez_tmp_212 = rob_uop_2_3_ldst_val;
      5'b00100:
        casez_tmp_212 = rob_uop_2_4_ldst_val;
      5'b00101:
        casez_tmp_212 = rob_uop_2_5_ldst_val;
      5'b00110:
        casez_tmp_212 = rob_uop_2_6_ldst_val;
      5'b00111:
        casez_tmp_212 = rob_uop_2_7_ldst_val;
      5'b01000:
        casez_tmp_212 = rob_uop_2_8_ldst_val;
      5'b01001:
        casez_tmp_212 = rob_uop_2_9_ldst_val;
      5'b01010:
        casez_tmp_212 = rob_uop_2_10_ldst_val;
      5'b01011:
        casez_tmp_212 = rob_uop_2_11_ldst_val;
      5'b01100:
        casez_tmp_212 = rob_uop_2_12_ldst_val;
      5'b01101:
        casez_tmp_212 = rob_uop_2_13_ldst_val;
      5'b01110:
        casez_tmp_212 = rob_uop_2_14_ldst_val;
      5'b01111:
        casez_tmp_212 = rob_uop_2_15_ldst_val;
      5'b10000:
        casez_tmp_212 = rob_uop_2_16_ldst_val;
      5'b10001:
        casez_tmp_212 = rob_uop_2_17_ldst_val;
      5'b10010:
        casez_tmp_212 = rob_uop_2_18_ldst_val;
      5'b10011:
        casez_tmp_212 = rob_uop_2_19_ldst_val;
      5'b10100:
        casez_tmp_212 = rob_uop_2_20_ldst_val;
      5'b10101:
        casez_tmp_212 = rob_uop_2_21_ldst_val;
      5'b10110:
        casez_tmp_212 = rob_uop_2_22_ldst_val;
      5'b10111:
        casez_tmp_212 = rob_uop_2_23_ldst_val;
      5'b11000:
        casez_tmp_212 = rob_uop_2_24_ldst_val;
      5'b11001:
        casez_tmp_212 = rob_uop_2_25_ldst_val;
      5'b11010:
        casez_tmp_212 = rob_uop_2_26_ldst_val;
      5'b11011:
        casez_tmp_212 = rob_uop_2_27_ldst_val;
      5'b11100:
        casez_tmp_212 = rob_uop_2_28_ldst_val;
      5'b11101:
        casez_tmp_212 = rob_uop_2_29_ldst_val;
      5'b11110:
        casez_tmp_212 = rob_uop_2_30_ldst_val;
      default:
        casez_tmp_212 = rob_uop_2_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_213;
  always @(*) begin
    casez (io_wb_resps_5_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_213 = rob_val_2_0;
      5'b00001:
        casez_tmp_213 = rob_val_2_1;
      5'b00010:
        casez_tmp_213 = rob_val_2_2;
      5'b00011:
        casez_tmp_213 = rob_val_2_3;
      5'b00100:
        casez_tmp_213 = rob_val_2_4;
      5'b00101:
        casez_tmp_213 = rob_val_2_5;
      5'b00110:
        casez_tmp_213 = rob_val_2_6;
      5'b00111:
        casez_tmp_213 = rob_val_2_7;
      5'b01000:
        casez_tmp_213 = rob_val_2_8;
      5'b01001:
        casez_tmp_213 = rob_val_2_9;
      5'b01010:
        casez_tmp_213 = rob_val_2_10;
      5'b01011:
        casez_tmp_213 = rob_val_2_11;
      5'b01100:
        casez_tmp_213 = rob_val_2_12;
      5'b01101:
        casez_tmp_213 = rob_val_2_13;
      5'b01110:
        casez_tmp_213 = rob_val_2_14;
      5'b01111:
        casez_tmp_213 = rob_val_2_15;
      5'b10000:
        casez_tmp_213 = rob_val_2_16;
      5'b10001:
        casez_tmp_213 = rob_val_2_17;
      5'b10010:
        casez_tmp_213 = rob_val_2_18;
      5'b10011:
        casez_tmp_213 = rob_val_2_19;
      5'b10100:
        casez_tmp_213 = rob_val_2_20;
      5'b10101:
        casez_tmp_213 = rob_val_2_21;
      5'b10110:
        casez_tmp_213 = rob_val_2_22;
      5'b10111:
        casez_tmp_213 = rob_val_2_23;
      5'b11000:
        casez_tmp_213 = rob_val_2_24;
      5'b11001:
        casez_tmp_213 = rob_val_2_25;
      5'b11010:
        casez_tmp_213 = rob_val_2_26;
      5'b11011:
        casez_tmp_213 = rob_val_2_27;
      5'b11100:
        casez_tmp_213 = rob_val_2_28;
      5'b11101:
        casez_tmp_213 = rob_val_2_29;
      5'b11110:
        casez_tmp_213 = rob_val_2_30;
      default:
        casez_tmp_213 = rob_val_2_31;
    endcase
  end // always @(*)
  reg         casez_tmp_214;
  always @(*) begin
    casez (io_wb_resps_5_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_214 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_214 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_214 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_214 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_214 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_214 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_214 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_214 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_214 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_214 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_214 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_214 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_214 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_214 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_214 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_214 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_214 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_214 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_214 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_214 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_214 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_214 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_214 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_214 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_214 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_214 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_214 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_214 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_214 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_214 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_214 = rob_bsy_2_30;
      default:
        casez_tmp_214 = rob_bsy_2_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_215;
  always @(*) begin
    casez (io_wb_resps_5_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_215 = rob_uop_2_0_pdst;
      5'b00001:
        casez_tmp_215 = rob_uop_2_1_pdst;
      5'b00010:
        casez_tmp_215 = rob_uop_2_2_pdst;
      5'b00011:
        casez_tmp_215 = rob_uop_2_3_pdst;
      5'b00100:
        casez_tmp_215 = rob_uop_2_4_pdst;
      5'b00101:
        casez_tmp_215 = rob_uop_2_5_pdst;
      5'b00110:
        casez_tmp_215 = rob_uop_2_6_pdst;
      5'b00111:
        casez_tmp_215 = rob_uop_2_7_pdst;
      5'b01000:
        casez_tmp_215 = rob_uop_2_8_pdst;
      5'b01001:
        casez_tmp_215 = rob_uop_2_9_pdst;
      5'b01010:
        casez_tmp_215 = rob_uop_2_10_pdst;
      5'b01011:
        casez_tmp_215 = rob_uop_2_11_pdst;
      5'b01100:
        casez_tmp_215 = rob_uop_2_12_pdst;
      5'b01101:
        casez_tmp_215 = rob_uop_2_13_pdst;
      5'b01110:
        casez_tmp_215 = rob_uop_2_14_pdst;
      5'b01111:
        casez_tmp_215 = rob_uop_2_15_pdst;
      5'b10000:
        casez_tmp_215 = rob_uop_2_16_pdst;
      5'b10001:
        casez_tmp_215 = rob_uop_2_17_pdst;
      5'b10010:
        casez_tmp_215 = rob_uop_2_18_pdst;
      5'b10011:
        casez_tmp_215 = rob_uop_2_19_pdst;
      5'b10100:
        casez_tmp_215 = rob_uop_2_20_pdst;
      5'b10101:
        casez_tmp_215 = rob_uop_2_21_pdst;
      5'b10110:
        casez_tmp_215 = rob_uop_2_22_pdst;
      5'b10111:
        casez_tmp_215 = rob_uop_2_23_pdst;
      5'b11000:
        casez_tmp_215 = rob_uop_2_24_pdst;
      5'b11001:
        casez_tmp_215 = rob_uop_2_25_pdst;
      5'b11010:
        casez_tmp_215 = rob_uop_2_26_pdst;
      5'b11011:
        casez_tmp_215 = rob_uop_2_27_pdst;
      5'b11100:
        casez_tmp_215 = rob_uop_2_28_pdst;
      5'b11101:
        casez_tmp_215 = rob_uop_2_29_pdst;
      5'b11110:
        casez_tmp_215 = rob_uop_2_30_pdst;
      default:
        casez_tmp_215 = rob_uop_2_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_216;
  always @(*) begin
    casez (io_wb_resps_5_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_216 = rob_uop_2_0_ldst_val;
      5'b00001:
        casez_tmp_216 = rob_uop_2_1_ldst_val;
      5'b00010:
        casez_tmp_216 = rob_uop_2_2_ldst_val;
      5'b00011:
        casez_tmp_216 = rob_uop_2_3_ldst_val;
      5'b00100:
        casez_tmp_216 = rob_uop_2_4_ldst_val;
      5'b00101:
        casez_tmp_216 = rob_uop_2_5_ldst_val;
      5'b00110:
        casez_tmp_216 = rob_uop_2_6_ldst_val;
      5'b00111:
        casez_tmp_216 = rob_uop_2_7_ldst_val;
      5'b01000:
        casez_tmp_216 = rob_uop_2_8_ldst_val;
      5'b01001:
        casez_tmp_216 = rob_uop_2_9_ldst_val;
      5'b01010:
        casez_tmp_216 = rob_uop_2_10_ldst_val;
      5'b01011:
        casez_tmp_216 = rob_uop_2_11_ldst_val;
      5'b01100:
        casez_tmp_216 = rob_uop_2_12_ldst_val;
      5'b01101:
        casez_tmp_216 = rob_uop_2_13_ldst_val;
      5'b01110:
        casez_tmp_216 = rob_uop_2_14_ldst_val;
      5'b01111:
        casez_tmp_216 = rob_uop_2_15_ldst_val;
      5'b10000:
        casez_tmp_216 = rob_uop_2_16_ldst_val;
      5'b10001:
        casez_tmp_216 = rob_uop_2_17_ldst_val;
      5'b10010:
        casez_tmp_216 = rob_uop_2_18_ldst_val;
      5'b10011:
        casez_tmp_216 = rob_uop_2_19_ldst_val;
      5'b10100:
        casez_tmp_216 = rob_uop_2_20_ldst_val;
      5'b10101:
        casez_tmp_216 = rob_uop_2_21_ldst_val;
      5'b10110:
        casez_tmp_216 = rob_uop_2_22_ldst_val;
      5'b10111:
        casez_tmp_216 = rob_uop_2_23_ldst_val;
      5'b11000:
        casez_tmp_216 = rob_uop_2_24_ldst_val;
      5'b11001:
        casez_tmp_216 = rob_uop_2_25_ldst_val;
      5'b11010:
        casez_tmp_216 = rob_uop_2_26_ldst_val;
      5'b11011:
        casez_tmp_216 = rob_uop_2_27_ldst_val;
      5'b11100:
        casez_tmp_216 = rob_uop_2_28_ldst_val;
      5'b11101:
        casez_tmp_216 = rob_uop_2_29_ldst_val;
      5'b11110:
        casez_tmp_216 = rob_uop_2_30_ldst_val;
      default:
        casez_tmp_216 = rob_uop_2_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_217;
  always @(*) begin
    casez (io_wb_resps_6_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_217 = rob_val_2_0;
      5'b00001:
        casez_tmp_217 = rob_val_2_1;
      5'b00010:
        casez_tmp_217 = rob_val_2_2;
      5'b00011:
        casez_tmp_217 = rob_val_2_3;
      5'b00100:
        casez_tmp_217 = rob_val_2_4;
      5'b00101:
        casez_tmp_217 = rob_val_2_5;
      5'b00110:
        casez_tmp_217 = rob_val_2_6;
      5'b00111:
        casez_tmp_217 = rob_val_2_7;
      5'b01000:
        casez_tmp_217 = rob_val_2_8;
      5'b01001:
        casez_tmp_217 = rob_val_2_9;
      5'b01010:
        casez_tmp_217 = rob_val_2_10;
      5'b01011:
        casez_tmp_217 = rob_val_2_11;
      5'b01100:
        casez_tmp_217 = rob_val_2_12;
      5'b01101:
        casez_tmp_217 = rob_val_2_13;
      5'b01110:
        casez_tmp_217 = rob_val_2_14;
      5'b01111:
        casez_tmp_217 = rob_val_2_15;
      5'b10000:
        casez_tmp_217 = rob_val_2_16;
      5'b10001:
        casez_tmp_217 = rob_val_2_17;
      5'b10010:
        casez_tmp_217 = rob_val_2_18;
      5'b10011:
        casez_tmp_217 = rob_val_2_19;
      5'b10100:
        casez_tmp_217 = rob_val_2_20;
      5'b10101:
        casez_tmp_217 = rob_val_2_21;
      5'b10110:
        casez_tmp_217 = rob_val_2_22;
      5'b10111:
        casez_tmp_217 = rob_val_2_23;
      5'b11000:
        casez_tmp_217 = rob_val_2_24;
      5'b11001:
        casez_tmp_217 = rob_val_2_25;
      5'b11010:
        casez_tmp_217 = rob_val_2_26;
      5'b11011:
        casez_tmp_217 = rob_val_2_27;
      5'b11100:
        casez_tmp_217 = rob_val_2_28;
      5'b11101:
        casez_tmp_217 = rob_val_2_29;
      5'b11110:
        casez_tmp_217 = rob_val_2_30;
      default:
        casez_tmp_217 = rob_val_2_31;
    endcase
  end // always @(*)
  reg         casez_tmp_218;
  always @(*) begin
    casez (io_wb_resps_6_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_218 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_218 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_218 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_218 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_218 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_218 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_218 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_218 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_218 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_218 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_218 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_218 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_218 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_218 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_218 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_218 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_218 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_218 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_218 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_218 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_218 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_218 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_218 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_218 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_218 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_218 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_218 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_218 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_218 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_218 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_218 = rob_bsy_2_30;
      default:
        casez_tmp_218 = rob_bsy_2_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_219;
  always @(*) begin
    casez (io_wb_resps_6_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_219 = rob_uop_2_0_pdst;
      5'b00001:
        casez_tmp_219 = rob_uop_2_1_pdst;
      5'b00010:
        casez_tmp_219 = rob_uop_2_2_pdst;
      5'b00011:
        casez_tmp_219 = rob_uop_2_3_pdst;
      5'b00100:
        casez_tmp_219 = rob_uop_2_4_pdst;
      5'b00101:
        casez_tmp_219 = rob_uop_2_5_pdst;
      5'b00110:
        casez_tmp_219 = rob_uop_2_6_pdst;
      5'b00111:
        casez_tmp_219 = rob_uop_2_7_pdst;
      5'b01000:
        casez_tmp_219 = rob_uop_2_8_pdst;
      5'b01001:
        casez_tmp_219 = rob_uop_2_9_pdst;
      5'b01010:
        casez_tmp_219 = rob_uop_2_10_pdst;
      5'b01011:
        casez_tmp_219 = rob_uop_2_11_pdst;
      5'b01100:
        casez_tmp_219 = rob_uop_2_12_pdst;
      5'b01101:
        casez_tmp_219 = rob_uop_2_13_pdst;
      5'b01110:
        casez_tmp_219 = rob_uop_2_14_pdst;
      5'b01111:
        casez_tmp_219 = rob_uop_2_15_pdst;
      5'b10000:
        casez_tmp_219 = rob_uop_2_16_pdst;
      5'b10001:
        casez_tmp_219 = rob_uop_2_17_pdst;
      5'b10010:
        casez_tmp_219 = rob_uop_2_18_pdst;
      5'b10011:
        casez_tmp_219 = rob_uop_2_19_pdst;
      5'b10100:
        casez_tmp_219 = rob_uop_2_20_pdst;
      5'b10101:
        casez_tmp_219 = rob_uop_2_21_pdst;
      5'b10110:
        casez_tmp_219 = rob_uop_2_22_pdst;
      5'b10111:
        casez_tmp_219 = rob_uop_2_23_pdst;
      5'b11000:
        casez_tmp_219 = rob_uop_2_24_pdst;
      5'b11001:
        casez_tmp_219 = rob_uop_2_25_pdst;
      5'b11010:
        casez_tmp_219 = rob_uop_2_26_pdst;
      5'b11011:
        casez_tmp_219 = rob_uop_2_27_pdst;
      5'b11100:
        casez_tmp_219 = rob_uop_2_28_pdst;
      5'b11101:
        casez_tmp_219 = rob_uop_2_29_pdst;
      5'b11110:
        casez_tmp_219 = rob_uop_2_30_pdst;
      default:
        casez_tmp_219 = rob_uop_2_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_220;
  always @(*) begin
    casez (io_wb_resps_6_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_220 = rob_uop_2_0_ldst_val;
      5'b00001:
        casez_tmp_220 = rob_uop_2_1_ldst_val;
      5'b00010:
        casez_tmp_220 = rob_uop_2_2_ldst_val;
      5'b00011:
        casez_tmp_220 = rob_uop_2_3_ldst_val;
      5'b00100:
        casez_tmp_220 = rob_uop_2_4_ldst_val;
      5'b00101:
        casez_tmp_220 = rob_uop_2_5_ldst_val;
      5'b00110:
        casez_tmp_220 = rob_uop_2_6_ldst_val;
      5'b00111:
        casez_tmp_220 = rob_uop_2_7_ldst_val;
      5'b01000:
        casez_tmp_220 = rob_uop_2_8_ldst_val;
      5'b01001:
        casez_tmp_220 = rob_uop_2_9_ldst_val;
      5'b01010:
        casez_tmp_220 = rob_uop_2_10_ldst_val;
      5'b01011:
        casez_tmp_220 = rob_uop_2_11_ldst_val;
      5'b01100:
        casez_tmp_220 = rob_uop_2_12_ldst_val;
      5'b01101:
        casez_tmp_220 = rob_uop_2_13_ldst_val;
      5'b01110:
        casez_tmp_220 = rob_uop_2_14_ldst_val;
      5'b01111:
        casez_tmp_220 = rob_uop_2_15_ldst_val;
      5'b10000:
        casez_tmp_220 = rob_uop_2_16_ldst_val;
      5'b10001:
        casez_tmp_220 = rob_uop_2_17_ldst_val;
      5'b10010:
        casez_tmp_220 = rob_uop_2_18_ldst_val;
      5'b10011:
        casez_tmp_220 = rob_uop_2_19_ldst_val;
      5'b10100:
        casez_tmp_220 = rob_uop_2_20_ldst_val;
      5'b10101:
        casez_tmp_220 = rob_uop_2_21_ldst_val;
      5'b10110:
        casez_tmp_220 = rob_uop_2_22_ldst_val;
      5'b10111:
        casez_tmp_220 = rob_uop_2_23_ldst_val;
      5'b11000:
        casez_tmp_220 = rob_uop_2_24_ldst_val;
      5'b11001:
        casez_tmp_220 = rob_uop_2_25_ldst_val;
      5'b11010:
        casez_tmp_220 = rob_uop_2_26_ldst_val;
      5'b11011:
        casez_tmp_220 = rob_uop_2_27_ldst_val;
      5'b11100:
        casez_tmp_220 = rob_uop_2_28_ldst_val;
      5'b11101:
        casez_tmp_220 = rob_uop_2_29_ldst_val;
      5'b11110:
        casez_tmp_220 = rob_uop_2_30_ldst_val;
      default:
        casez_tmp_220 = rob_uop_2_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_221;
  always @(*) begin
    casez (io_wb_resps_7_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_221 = rob_val_2_0;
      5'b00001:
        casez_tmp_221 = rob_val_2_1;
      5'b00010:
        casez_tmp_221 = rob_val_2_2;
      5'b00011:
        casez_tmp_221 = rob_val_2_3;
      5'b00100:
        casez_tmp_221 = rob_val_2_4;
      5'b00101:
        casez_tmp_221 = rob_val_2_5;
      5'b00110:
        casez_tmp_221 = rob_val_2_6;
      5'b00111:
        casez_tmp_221 = rob_val_2_7;
      5'b01000:
        casez_tmp_221 = rob_val_2_8;
      5'b01001:
        casez_tmp_221 = rob_val_2_9;
      5'b01010:
        casez_tmp_221 = rob_val_2_10;
      5'b01011:
        casez_tmp_221 = rob_val_2_11;
      5'b01100:
        casez_tmp_221 = rob_val_2_12;
      5'b01101:
        casez_tmp_221 = rob_val_2_13;
      5'b01110:
        casez_tmp_221 = rob_val_2_14;
      5'b01111:
        casez_tmp_221 = rob_val_2_15;
      5'b10000:
        casez_tmp_221 = rob_val_2_16;
      5'b10001:
        casez_tmp_221 = rob_val_2_17;
      5'b10010:
        casez_tmp_221 = rob_val_2_18;
      5'b10011:
        casez_tmp_221 = rob_val_2_19;
      5'b10100:
        casez_tmp_221 = rob_val_2_20;
      5'b10101:
        casez_tmp_221 = rob_val_2_21;
      5'b10110:
        casez_tmp_221 = rob_val_2_22;
      5'b10111:
        casez_tmp_221 = rob_val_2_23;
      5'b11000:
        casez_tmp_221 = rob_val_2_24;
      5'b11001:
        casez_tmp_221 = rob_val_2_25;
      5'b11010:
        casez_tmp_221 = rob_val_2_26;
      5'b11011:
        casez_tmp_221 = rob_val_2_27;
      5'b11100:
        casez_tmp_221 = rob_val_2_28;
      5'b11101:
        casez_tmp_221 = rob_val_2_29;
      5'b11110:
        casez_tmp_221 = rob_val_2_30;
      default:
        casez_tmp_221 = rob_val_2_31;
    endcase
  end // always @(*)
  reg         casez_tmp_222;
  always @(*) begin
    casez (io_wb_resps_7_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_222 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_222 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_222 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_222 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_222 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_222 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_222 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_222 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_222 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_222 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_222 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_222 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_222 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_222 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_222 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_222 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_222 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_222 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_222 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_222 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_222 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_222 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_222 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_222 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_222 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_222 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_222 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_222 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_222 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_222 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_222 = rob_bsy_2_30;
      default:
        casez_tmp_222 = rob_bsy_2_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_223;
  always @(*) begin
    casez (io_wb_resps_7_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_223 = rob_uop_2_0_pdst;
      5'b00001:
        casez_tmp_223 = rob_uop_2_1_pdst;
      5'b00010:
        casez_tmp_223 = rob_uop_2_2_pdst;
      5'b00011:
        casez_tmp_223 = rob_uop_2_3_pdst;
      5'b00100:
        casez_tmp_223 = rob_uop_2_4_pdst;
      5'b00101:
        casez_tmp_223 = rob_uop_2_5_pdst;
      5'b00110:
        casez_tmp_223 = rob_uop_2_6_pdst;
      5'b00111:
        casez_tmp_223 = rob_uop_2_7_pdst;
      5'b01000:
        casez_tmp_223 = rob_uop_2_8_pdst;
      5'b01001:
        casez_tmp_223 = rob_uop_2_9_pdst;
      5'b01010:
        casez_tmp_223 = rob_uop_2_10_pdst;
      5'b01011:
        casez_tmp_223 = rob_uop_2_11_pdst;
      5'b01100:
        casez_tmp_223 = rob_uop_2_12_pdst;
      5'b01101:
        casez_tmp_223 = rob_uop_2_13_pdst;
      5'b01110:
        casez_tmp_223 = rob_uop_2_14_pdst;
      5'b01111:
        casez_tmp_223 = rob_uop_2_15_pdst;
      5'b10000:
        casez_tmp_223 = rob_uop_2_16_pdst;
      5'b10001:
        casez_tmp_223 = rob_uop_2_17_pdst;
      5'b10010:
        casez_tmp_223 = rob_uop_2_18_pdst;
      5'b10011:
        casez_tmp_223 = rob_uop_2_19_pdst;
      5'b10100:
        casez_tmp_223 = rob_uop_2_20_pdst;
      5'b10101:
        casez_tmp_223 = rob_uop_2_21_pdst;
      5'b10110:
        casez_tmp_223 = rob_uop_2_22_pdst;
      5'b10111:
        casez_tmp_223 = rob_uop_2_23_pdst;
      5'b11000:
        casez_tmp_223 = rob_uop_2_24_pdst;
      5'b11001:
        casez_tmp_223 = rob_uop_2_25_pdst;
      5'b11010:
        casez_tmp_223 = rob_uop_2_26_pdst;
      5'b11011:
        casez_tmp_223 = rob_uop_2_27_pdst;
      5'b11100:
        casez_tmp_223 = rob_uop_2_28_pdst;
      5'b11101:
        casez_tmp_223 = rob_uop_2_29_pdst;
      5'b11110:
        casez_tmp_223 = rob_uop_2_30_pdst;
      default:
        casez_tmp_223 = rob_uop_2_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_224;
  always @(*) begin
    casez (io_wb_resps_7_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_224 = rob_uop_2_0_ldst_val;
      5'b00001:
        casez_tmp_224 = rob_uop_2_1_ldst_val;
      5'b00010:
        casez_tmp_224 = rob_uop_2_2_ldst_val;
      5'b00011:
        casez_tmp_224 = rob_uop_2_3_ldst_val;
      5'b00100:
        casez_tmp_224 = rob_uop_2_4_ldst_val;
      5'b00101:
        casez_tmp_224 = rob_uop_2_5_ldst_val;
      5'b00110:
        casez_tmp_224 = rob_uop_2_6_ldst_val;
      5'b00111:
        casez_tmp_224 = rob_uop_2_7_ldst_val;
      5'b01000:
        casez_tmp_224 = rob_uop_2_8_ldst_val;
      5'b01001:
        casez_tmp_224 = rob_uop_2_9_ldst_val;
      5'b01010:
        casez_tmp_224 = rob_uop_2_10_ldst_val;
      5'b01011:
        casez_tmp_224 = rob_uop_2_11_ldst_val;
      5'b01100:
        casez_tmp_224 = rob_uop_2_12_ldst_val;
      5'b01101:
        casez_tmp_224 = rob_uop_2_13_ldst_val;
      5'b01110:
        casez_tmp_224 = rob_uop_2_14_ldst_val;
      5'b01111:
        casez_tmp_224 = rob_uop_2_15_ldst_val;
      5'b10000:
        casez_tmp_224 = rob_uop_2_16_ldst_val;
      5'b10001:
        casez_tmp_224 = rob_uop_2_17_ldst_val;
      5'b10010:
        casez_tmp_224 = rob_uop_2_18_ldst_val;
      5'b10011:
        casez_tmp_224 = rob_uop_2_19_ldst_val;
      5'b10100:
        casez_tmp_224 = rob_uop_2_20_ldst_val;
      5'b10101:
        casez_tmp_224 = rob_uop_2_21_ldst_val;
      5'b10110:
        casez_tmp_224 = rob_uop_2_22_ldst_val;
      5'b10111:
        casez_tmp_224 = rob_uop_2_23_ldst_val;
      5'b11000:
        casez_tmp_224 = rob_uop_2_24_ldst_val;
      5'b11001:
        casez_tmp_224 = rob_uop_2_25_ldst_val;
      5'b11010:
        casez_tmp_224 = rob_uop_2_26_ldst_val;
      5'b11011:
        casez_tmp_224 = rob_uop_2_27_ldst_val;
      5'b11100:
        casez_tmp_224 = rob_uop_2_28_ldst_val;
      5'b11101:
        casez_tmp_224 = rob_uop_2_29_ldst_val;
      5'b11110:
        casez_tmp_224 = rob_uop_2_30_ldst_val;
      default:
        casez_tmp_224 = rob_uop_2_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_225;
  always @(*) begin
    casez (io_wb_resps_8_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_225 = rob_val_2_0;
      5'b00001:
        casez_tmp_225 = rob_val_2_1;
      5'b00010:
        casez_tmp_225 = rob_val_2_2;
      5'b00011:
        casez_tmp_225 = rob_val_2_3;
      5'b00100:
        casez_tmp_225 = rob_val_2_4;
      5'b00101:
        casez_tmp_225 = rob_val_2_5;
      5'b00110:
        casez_tmp_225 = rob_val_2_6;
      5'b00111:
        casez_tmp_225 = rob_val_2_7;
      5'b01000:
        casez_tmp_225 = rob_val_2_8;
      5'b01001:
        casez_tmp_225 = rob_val_2_9;
      5'b01010:
        casez_tmp_225 = rob_val_2_10;
      5'b01011:
        casez_tmp_225 = rob_val_2_11;
      5'b01100:
        casez_tmp_225 = rob_val_2_12;
      5'b01101:
        casez_tmp_225 = rob_val_2_13;
      5'b01110:
        casez_tmp_225 = rob_val_2_14;
      5'b01111:
        casez_tmp_225 = rob_val_2_15;
      5'b10000:
        casez_tmp_225 = rob_val_2_16;
      5'b10001:
        casez_tmp_225 = rob_val_2_17;
      5'b10010:
        casez_tmp_225 = rob_val_2_18;
      5'b10011:
        casez_tmp_225 = rob_val_2_19;
      5'b10100:
        casez_tmp_225 = rob_val_2_20;
      5'b10101:
        casez_tmp_225 = rob_val_2_21;
      5'b10110:
        casez_tmp_225 = rob_val_2_22;
      5'b10111:
        casez_tmp_225 = rob_val_2_23;
      5'b11000:
        casez_tmp_225 = rob_val_2_24;
      5'b11001:
        casez_tmp_225 = rob_val_2_25;
      5'b11010:
        casez_tmp_225 = rob_val_2_26;
      5'b11011:
        casez_tmp_225 = rob_val_2_27;
      5'b11100:
        casez_tmp_225 = rob_val_2_28;
      5'b11101:
        casez_tmp_225 = rob_val_2_29;
      5'b11110:
        casez_tmp_225 = rob_val_2_30;
      default:
        casez_tmp_225 = rob_val_2_31;
    endcase
  end // always @(*)
  reg         casez_tmp_226;
  always @(*) begin
    casez (io_wb_resps_8_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_226 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_226 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_226 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_226 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_226 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_226 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_226 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_226 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_226 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_226 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_226 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_226 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_226 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_226 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_226 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_226 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_226 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_226 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_226 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_226 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_226 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_226 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_226 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_226 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_226 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_226 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_226 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_226 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_226 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_226 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_226 = rob_bsy_2_30;
      default:
        casez_tmp_226 = rob_bsy_2_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_227;
  always @(*) begin
    casez (io_wb_resps_8_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_227 = rob_uop_2_0_pdst;
      5'b00001:
        casez_tmp_227 = rob_uop_2_1_pdst;
      5'b00010:
        casez_tmp_227 = rob_uop_2_2_pdst;
      5'b00011:
        casez_tmp_227 = rob_uop_2_3_pdst;
      5'b00100:
        casez_tmp_227 = rob_uop_2_4_pdst;
      5'b00101:
        casez_tmp_227 = rob_uop_2_5_pdst;
      5'b00110:
        casez_tmp_227 = rob_uop_2_6_pdst;
      5'b00111:
        casez_tmp_227 = rob_uop_2_7_pdst;
      5'b01000:
        casez_tmp_227 = rob_uop_2_8_pdst;
      5'b01001:
        casez_tmp_227 = rob_uop_2_9_pdst;
      5'b01010:
        casez_tmp_227 = rob_uop_2_10_pdst;
      5'b01011:
        casez_tmp_227 = rob_uop_2_11_pdst;
      5'b01100:
        casez_tmp_227 = rob_uop_2_12_pdst;
      5'b01101:
        casez_tmp_227 = rob_uop_2_13_pdst;
      5'b01110:
        casez_tmp_227 = rob_uop_2_14_pdst;
      5'b01111:
        casez_tmp_227 = rob_uop_2_15_pdst;
      5'b10000:
        casez_tmp_227 = rob_uop_2_16_pdst;
      5'b10001:
        casez_tmp_227 = rob_uop_2_17_pdst;
      5'b10010:
        casez_tmp_227 = rob_uop_2_18_pdst;
      5'b10011:
        casez_tmp_227 = rob_uop_2_19_pdst;
      5'b10100:
        casez_tmp_227 = rob_uop_2_20_pdst;
      5'b10101:
        casez_tmp_227 = rob_uop_2_21_pdst;
      5'b10110:
        casez_tmp_227 = rob_uop_2_22_pdst;
      5'b10111:
        casez_tmp_227 = rob_uop_2_23_pdst;
      5'b11000:
        casez_tmp_227 = rob_uop_2_24_pdst;
      5'b11001:
        casez_tmp_227 = rob_uop_2_25_pdst;
      5'b11010:
        casez_tmp_227 = rob_uop_2_26_pdst;
      5'b11011:
        casez_tmp_227 = rob_uop_2_27_pdst;
      5'b11100:
        casez_tmp_227 = rob_uop_2_28_pdst;
      5'b11101:
        casez_tmp_227 = rob_uop_2_29_pdst;
      5'b11110:
        casez_tmp_227 = rob_uop_2_30_pdst;
      default:
        casez_tmp_227 = rob_uop_2_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_228;
  always @(*) begin
    casez (io_wb_resps_8_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_228 = rob_uop_2_0_ldst_val;
      5'b00001:
        casez_tmp_228 = rob_uop_2_1_ldst_val;
      5'b00010:
        casez_tmp_228 = rob_uop_2_2_ldst_val;
      5'b00011:
        casez_tmp_228 = rob_uop_2_3_ldst_val;
      5'b00100:
        casez_tmp_228 = rob_uop_2_4_ldst_val;
      5'b00101:
        casez_tmp_228 = rob_uop_2_5_ldst_val;
      5'b00110:
        casez_tmp_228 = rob_uop_2_6_ldst_val;
      5'b00111:
        casez_tmp_228 = rob_uop_2_7_ldst_val;
      5'b01000:
        casez_tmp_228 = rob_uop_2_8_ldst_val;
      5'b01001:
        casez_tmp_228 = rob_uop_2_9_ldst_val;
      5'b01010:
        casez_tmp_228 = rob_uop_2_10_ldst_val;
      5'b01011:
        casez_tmp_228 = rob_uop_2_11_ldst_val;
      5'b01100:
        casez_tmp_228 = rob_uop_2_12_ldst_val;
      5'b01101:
        casez_tmp_228 = rob_uop_2_13_ldst_val;
      5'b01110:
        casez_tmp_228 = rob_uop_2_14_ldst_val;
      5'b01111:
        casez_tmp_228 = rob_uop_2_15_ldst_val;
      5'b10000:
        casez_tmp_228 = rob_uop_2_16_ldst_val;
      5'b10001:
        casez_tmp_228 = rob_uop_2_17_ldst_val;
      5'b10010:
        casez_tmp_228 = rob_uop_2_18_ldst_val;
      5'b10011:
        casez_tmp_228 = rob_uop_2_19_ldst_val;
      5'b10100:
        casez_tmp_228 = rob_uop_2_20_ldst_val;
      5'b10101:
        casez_tmp_228 = rob_uop_2_21_ldst_val;
      5'b10110:
        casez_tmp_228 = rob_uop_2_22_ldst_val;
      5'b10111:
        casez_tmp_228 = rob_uop_2_23_ldst_val;
      5'b11000:
        casez_tmp_228 = rob_uop_2_24_ldst_val;
      5'b11001:
        casez_tmp_228 = rob_uop_2_25_ldst_val;
      5'b11010:
        casez_tmp_228 = rob_uop_2_26_ldst_val;
      5'b11011:
        casez_tmp_228 = rob_uop_2_27_ldst_val;
      5'b11100:
        casez_tmp_228 = rob_uop_2_28_ldst_val;
      5'b11101:
        casez_tmp_228 = rob_uop_2_29_ldst_val;
      5'b11110:
        casez_tmp_228 = rob_uop_2_30_ldst_val;
      default:
        casez_tmp_228 = rob_uop_2_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_229;
  always @(*) begin
    casez (io_wb_resps_9_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_229 = rob_val_2_0;
      5'b00001:
        casez_tmp_229 = rob_val_2_1;
      5'b00010:
        casez_tmp_229 = rob_val_2_2;
      5'b00011:
        casez_tmp_229 = rob_val_2_3;
      5'b00100:
        casez_tmp_229 = rob_val_2_4;
      5'b00101:
        casez_tmp_229 = rob_val_2_5;
      5'b00110:
        casez_tmp_229 = rob_val_2_6;
      5'b00111:
        casez_tmp_229 = rob_val_2_7;
      5'b01000:
        casez_tmp_229 = rob_val_2_8;
      5'b01001:
        casez_tmp_229 = rob_val_2_9;
      5'b01010:
        casez_tmp_229 = rob_val_2_10;
      5'b01011:
        casez_tmp_229 = rob_val_2_11;
      5'b01100:
        casez_tmp_229 = rob_val_2_12;
      5'b01101:
        casez_tmp_229 = rob_val_2_13;
      5'b01110:
        casez_tmp_229 = rob_val_2_14;
      5'b01111:
        casez_tmp_229 = rob_val_2_15;
      5'b10000:
        casez_tmp_229 = rob_val_2_16;
      5'b10001:
        casez_tmp_229 = rob_val_2_17;
      5'b10010:
        casez_tmp_229 = rob_val_2_18;
      5'b10011:
        casez_tmp_229 = rob_val_2_19;
      5'b10100:
        casez_tmp_229 = rob_val_2_20;
      5'b10101:
        casez_tmp_229 = rob_val_2_21;
      5'b10110:
        casez_tmp_229 = rob_val_2_22;
      5'b10111:
        casez_tmp_229 = rob_val_2_23;
      5'b11000:
        casez_tmp_229 = rob_val_2_24;
      5'b11001:
        casez_tmp_229 = rob_val_2_25;
      5'b11010:
        casez_tmp_229 = rob_val_2_26;
      5'b11011:
        casez_tmp_229 = rob_val_2_27;
      5'b11100:
        casez_tmp_229 = rob_val_2_28;
      5'b11101:
        casez_tmp_229 = rob_val_2_29;
      5'b11110:
        casez_tmp_229 = rob_val_2_30;
      default:
        casez_tmp_229 = rob_val_2_31;
    endcase
  end // always @(*)
  reg         casez_tmp_230;
  always @(*) begin
    casez (io_wb_resps_9_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_230 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_230 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_230 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_230 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_230 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_230 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_230 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_230 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_230 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_230 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_230 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_230 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_230 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_230 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_230 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_230 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_230 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_230 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_230 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_230 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_230 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_230 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_230 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_230 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_230 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_230 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_230 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_230 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_230 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_230 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_230 = rob_bsy_2_30;
      default:
        casez_tmp_230 = rob_bsy_2_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_231;
  always @(*) begin
    casez (io_wb_resps_9_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_231 = rob_uop_2_0_pdst;
      5'b00001:
        casez_tmp_231 = rob_uop_2_1_pdst;
      5'b00010:
        casez_tmp_231 = rob_uop_2_2_pdst;
      5'b00011:
        casez_tmp_231 = rob_uop_2_3_pdst;
      5'b00100:
        casez_tmp_231 = rob_uop_2_4_pdst;
      5'b00101:
        casez_tmp_231 = rob_uop_2_5_pdst;
      5'b00110:
        casez_tmp_231 = rob_uop_2_6_pdst;
      5'b00111:
        casez_tmp_231 = rob_uop_2_7_pdst;
      5'b01000:
        casez_tmp_231 = rob_uop_2_8_pdst;
      5'b01001:
        casez_tmp_231 = rob_uop_2_9_pdst;
      5'b01010:
        casez_tmp_231 = rob_uop_2_10_pdst;
      5'b01011:
        casez_tmp_231 = rob_uop_2_11_pdst;
      5'b01100:
        casez_tmp_231 = rob_uop_2_12_pdst;
      5'b01101:
        casez_tmp_231 = rob_uop_2_13_pdst;
      5'b01110:
        casez_tmp_231 = rob_uop_2_14_pdst;
      5'b01111:
        casez_tmp_231 = rob_uop_2_15_pdst;
      5'b10000:
        casez_tmp_231 = rob_uop_2_16_pdst;
      5'b10001:
        casez_tmp_231 = rob_uop_2_17_pdst;
      5'b10010:
        casez_tmp_231 = rob_uop_2_18_pdst;
      5'b10011:
        casez_tmp_231 = rob_uop_2_19_pdst;
      5'b10100:
        casez_tmp_231 = rob_uop_2_20_pdst;
      5'b10101:
        casez_tmp_231 = rob_uop_2_21_pdst;
      5'b10110:
        casez_tmp_231 = rob_uop_2_22_pdst;
      5'b10111:
        casez_tmp_231 = rob_uop_2_23_pdst;
      5'b11000:
        casez_tmp_231 = rob_uop_2_24_pdst;
      5'b11001:
        casez_tmp_231 = rob_uop_2_25_pdst;
      5'b11010:
        casez_tmp_231 = rob_uop_2_26_pdst;
      5'b11011:
        casez_tmp_231 = rob_uop_2_27_pdst;
      5'b11100:
        casez_tmp_231 = rob_uop_2_28_pdst;
      5'b11101:
        casez_tmp_231 = rob_uop_2_29_pdst;
      5'b11110:
        casez_tmp_231 = rob_uop_2_30_pdst;
      default:
        casez_tmp_231 = rob_uop_2_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_232;
  always @(*) begin
    casez (io_wb_resps_9_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_232 = rob_uop_2_0_ldst_val;
      5'b00001:
        casez_tmp_232 = rob_uop_2_1_ldst_val;
      5'b00010:
        casez_tmp_232 = rob_uop_2_2_ldst_val;
      5'b00011:
        casez_tmp_232 = rob_uop_2_3_ldst_val;
      5'b00100:
        casez_tmp_232 = rob_uop_2_4_ldst_val;
      5'b00101:
        casez_tmp_232 = rob_uop_2_5_ldst_val;
      5'b00110:
        casez_tmp_232 = rob_uop_2_6_ldst_val;
      5'b00111:
        casez_tmp_232 = rob_uop_2_7_ldst_val;
      5'b01000:
        casez_tmp_232 = rob_uop_2_8_ldst_val;
      5'b01001:
        casez_tmp_232 = rob_uop_2_9_ldst_val;
      5'b01010:
        casez_tmp_232 = rob_uop_2_10_ldst_val;
      5'b01011:
        casez_tmp_232 = rob_uop_2_11_ldst_val;
      5'b01100:
        casez_tmp_232 = rob_uop_2_12_ldst_val;
      5'b01101:
        casez_tmp_232 = rob_uop_2_13_ldst_val;
      5'b01110:
        casez_tmp_232 = rob_uop_2_14_ldst_val;
      5'b01111:
        casez_tmp_232 = rob_uop_2_15_ldst_val;
      5'b10000:
        casez_tmp_232 = rob_uop_2_16_ldst_val;
      5'b10001:
        casez_tmp_232 = rob_uop_2_17_ldst_val;
      5'b10010:
        casez_tmp_232 = rob_uop_2_18_ldst_val;
      5'b10011:
        casez_tmp_232 = rob_uop_2_19_ldst_val;
      5'b10100:
        casez_tmp_232 = rob_uop_2_20_ldst_val;
      5'b10101:
        casez_tmp_232 = rob_uop_2_21_ldst_val;
      5'b10110:
        casez_tmp_232 = rob_uop_2_22_ldst_val;
      5'b10111:
        casez_tmp_232 = rob_uop_2_23_ldst_val;
      5'b11000:
        casez_tmp_232 = rob_uop_2_24_ldst_val;
      5'b11001:
        casez_tmp_232 = rob_uop_2_25_ldst_val;
      5'b11010:
        casez_tmp_232 = rob_uop_2_26_ldst_val;
      5'b11011:
        casez_tmp_232 = rob_uop_2_27_ldst_val;
      5'b11100:
        casez_tmp_232 = rob_uop_2_28_ldst_val;
      5'b11101:
        casez_tmp_232 = rob_uop_2_29_ldst_val;
      5'b11110:
        casez_tmp_232 = rob_uop_2_30_ldst_val;
      default:
        casez_tmp_232 = rob_uop_2_31_ldst_val;
    endcase
  end // always @(*)
  reg         rob_val_3_0;
  reg         rob_val_3_1;
  reg         rob_val_3_2;
  reg         rob_val_3_3;
  reg         rob_val_3_4;
  reg         rob_val_3_5;
  reg         rob_val_3_6;
  reg         rob_val_3_7;
  reg         rob_val_3_8;
  reg         rob_val_3_9;
  reg         rob_val_3_10;
  reg         rob_val_3_11;
  reg         rob_val_3_12;
  reg         rob_val_3_13;
  reg         rob_val_3_14;
  reg         rob_val_3_15;
  reg         rob_val_3_16;
  reg         rob_val_3_17;
  reg         rob_val_3_18;
  reg         rob_val_3_19;
  reg         rob_val_3_20;
  reg         rob_val_3_21;
  reg         rob_val_3_22;
  reg         rob_val_3_23;
  reg         rob_val_3_24;
  reg         rob_val_3_25;
  reg         rob_val_3_26;
  reg         rob_val_3_27;
  reg         rob_val_3_28;
  reg         rob_val_3_29;
  reg         rob_val_3_30;
  reg         rob_val_3_31;
  reg         rob_bsy_3_0;
  reg         rob_bsy_3_1;
  reg         rob_bsy_3_2;
  reg         rob_bsy_3_3;
  reg         rob_bsy_3_4;
  reg         rob_bsy_3_5;
  reg         rob_bsy_3_6;
  reg         rob_bsy_3_7;
  reg         rob_bsy_3_8;
  reg         rob_bsy_3_9;
  reg         rob_bsy_3_10;
  reg         rob_bsy_3_11;
  reg         rob_bsy_3_12;
  reg         rob_bsy_3_13;
  reg         rob_bsy_3_14;
  reg         rob_bsy_3_15;
  reg         rob_bsy_3_16;
  reg         rob_bsy_3_17;
  reg         rob_bsy_3_18;
  reg         rob_bsy_3_19;
  reg         rob_bsy_3_20;
  reg         rob_bsy_3_21;
  reg         rob_bsy_3_22;
  reg         rob_bsy_3_23;
  reg         rob_bsy_3_24;
  reg         rob_bsy_3_25;
  reg         rob_bsy_3_26;
  reg         rob_bsy_3_27;
  reg         rob_bsy_3_28;
  reg         rob_bsy_3_29;
  reg         rob_bsy_3_30;
  reg         rob_bsy_3_31;
  reg         rob_unsafe_3_0;
  reg         rob_unsafe_3_1;
  reg         rob_unsafe_3_2;
  reg         rob_unsafe_3_3;
  reg         rob_unsafe_3_4;
  reg         rob_unsafe_3_5;
  reg         rob_unsafe_3_6;
  reg         rob_unsafe_3_7;
  reg         rob_unsafe_3_8;
  reg         rob_unsafe_3_9;
  reg         rob_unsafe_3_10;
  reg         rob_unsafe_3_11;
  reg         rob_unsafe_3_12;
  reg         rob_unsafe_3_13;
  reg         rob_unsafe_3_14;
  reg         rob_unsafe_3_15;
  reg         rob_unsafe_3_16;
  reg         rob_unsafe_3_17;
  reg         rob_unsafe_3_18;
  reg         rob_unsafe_3_19;
  reg         rob_unsafe_3_20;
  reg         rob_unsafe_3_21;
  reg         rob_unsafe_3_22;
  reg         rob_unsafe_3_23;
  reg         rob_unsafe_3_24;
  reg         rob_unsafe_3_25;
  reg         rob_unsafe_3_26;
  reg         rob_unsafe_3_27;
  reg         rob_unsafe_3_28;
  reg         rob_unsafe_3_29;
  reg         rob_unsafe_3_30;
  reg         rob_unsafe_3_31;
  reg  [6:0]  rob_uop_3_0_uopc;
  reg         rob_uop_3_0_is_rvc;
  reg         rob_uop_3_0_is_br;
  reg         rob_uop_3_0_is_jalr;
  reg         rob_uop_3_0_is_jal;
  reg  [19:0] rob_uop_3_0_br_mask;
  reg  [5:0]  rob_uop_3_0_ftq_idx;
  reg         rob_uop_3_0_edge_inst;
  reg  [5:0]  rob_uop_3_0_pc_lob;
  reg  [6:0]  rob_uop_3_0_pdst;
  reg  [6:0]  rob_uop_3_0_stale_pdst;
  reg         rob_uop_3_0_is_fencei;
  reg         rob_uop_3_0_uses_ldq;
  reg         rob_uop_3_0_uses_stq;
  reg         rob_uop_3_0_is_sys_pc2epc;
  reg         rob_uop_3_0_flush_on_commit;
  reg  [5:0]  rob_uop_3_0_ldst;
  reg         rob_uop_3_0_ldst_val;
  reg  [1:0]  rob_uop_3_0_dst_rtype;
  reg         rob_uop_3_0_fp_val;
  reg  [1:0]  rob_uop_3_0_debug_fsrc;
  reg  [6:0]  rob_uop_3_1_uopc;
  reg         rob_uop_3_1_is_rvc;
  reg         rob_uop_3_1_is_br;
  reg         rob_uop_3_1_is_jalr;
  reg         rob_uop_3_1_is_jal;
  reg  [19:0] rob_uop_3_1_br_mask;
  reg  [5:0]  rob_uop_3_1_ftq_idx;
  reg         rob_uop_3_1_edge_inst;
  reg  [5:0]  rob_uop_3_1_pc_lob;
  reg  [6:0]  rob_uop_3_1_pdst;
  reg  [6:0]  rob_uop_3_1_stale_pdst;
  reg         rob_uop_3_1_is_fencei;
  reg         rob_uop_3_1_uses_ldq;
  reg         rob_uop_3_1_uses_stq;
  reg         rob_uop_3_1_is_sys_pc2epc;
  reg         rob_uop_3_1_flush_on_commit;
  reg  [5:0]  rob_uop_3_1_ldst;
  reg         rob_uop_3_1_ldst_val;
  reg  [1:0]  rob_uop_3_1_dst_rtype;
  reg         rob_uop_3_1_fp_val;
  reg  [1:0]  rob_uop_3_1_debug_fsrc;
  reg  [6:0]  rob_uop_3_2_uopc;
  reg         rob_uop_3_2_is_rvc;
  reg         rob_uop_3_2_is_br;
  reg         rob_uop_3_2_is_jalr;
  reg         rob_uop_3_2_is_jal;
  reg  [19:0] rob_uop_3_2_br_mask;
  reg  [5:0]  rob_uop_3_2_ftq_idx;
  reg         rob_uop_3_2_edge_inst;
  reg  [5:0]  rob_uop_3_2_pc_lob;
  reg  [6:0]  rob_uop_3_2_pdst;
  reg  [6:0]  rob_uop_3_2_stale_pdst;
  reg         rob_uop_3_2_is_fencei;
  reg         rob_uop_3_2_uses_ldq;
  reg         rob_uop_3_2_uses_stq;
  reg         rob_uop_3_2_is_sys_pc2epc;
  reg         rob_uop_3_2_flush_on_commit;
  reg  [5:0]  rob_uop_3_2_ldst;
  reg         rob_uop_3_2_ldst_val;
  reg  [1:0]  rob_uop_3_2_dst_rtype;
  reg         rob_uop_3_2_fp_val;
  reg  [1:0]  rob_uop_3_2_debug_fsrc;
  reg  [6:0]  rob_uop_3_3_uopc;
  reg         rob_uop_3_3_is_rvc;
  reg         rob_uop_3_3_is_br;
  reg         rob_uop_3_3_is_jalr;
  reg         rob_uop_3_3_is_jal;
  reg  [19:0] rob_uop_3_3_br_mask;
  reg  [5:0]  rob_uop_3_3_ftq_idx;
  reg         rob_uop_3_3_edge_inst;
  reg  [5:0]  rob_uop_3_3_pc_lob;
  reg  [6:0]  rob_uop_3_3_pdst;
  reg  [6:0]  rob_uop_3_3_stale_pdst;
  reg         rob_uop_3_3_is_fencei;
  reg         rob_uop_3_3_uses_ldq;
  reg         rob_uop_3_3_uses_stq;
  reg         rob_uop_3_3_is_sys_pc2epc;
  reg         rob_uop_3_3_flush_on_commit;
  reg  [5:0]  rob_uop_3_3_ldst;
  reg         rob_uop_3_3_ldst_val;
  reg  [1:0]  rob_uop_3_3_dst_rtype;
  reg         rob_uop_3_3_fp_val;
  reg  [1:0]  rob_uop_3_3_debug_fsrc;
  reg  [6:0]  rob_uop_3_4_uopc;
  reg         rob_uop_3_4_is_rvc;
  reg         rob_uop_3_4_is_br;
  reg         rob_uop_3_4_is_jalr;
  reg         rob_uop_3_4_is_jal;
  reg  [19:0] rob_uop_3_4_br_mask;
  reg  [5:0]  rob_uop_3_4_ftq_idx;
  reg         rob_uop_3_4_edge_inst;
  reg  [5:0]  rob_uop_3_4_pc_lob;
  reg  [6:0]  rob_uop_3_4_pdst;
  reg  [6:0]  rob_uop_3_4_stale_pdst;
  reg         rob_uop_3_4_is_fencei;
  reg         rob_uop_3_4_uses_ldq;
  reg         rob_uop_3_4_uses_stq;
  reg         rob_uop_3_4_is_sys_pc2epc;
  reg         rob_uop_3_4_flush_on_commit;
  reg  [5:0]  rob_uop_3_4_ldst;
  reg         rob_uop_3_4_ldst_val;
  reg  [1:0]  rob_uop_3_4_dst_rtype;
  reg         rob_uop_3_4_fp_val;
  reg  [1:0]  rob_uop_3_4_debug_fsrc;
  reg  [6:0]  rob_uop_3_5_uopc;
  reg         rob_uop_3_5_is_rvc;
  reg         rob_uop_3_5_is_br;
  reg         rob_uop_3_5_is_jalr;
  reg         rob_uop_3_5_is_jal;
  reg  [19:0] rob_uop_3_5_br_mask;
  reg  [5:0]  rob_uop_3_5_ftq_idx;
  reg         rob_uop_3_5_edge_inst;
  reg  [5:0]  rob_uop_3_5_pc_lob;
  reg  [6:0]  rob_uop_3_5_pdst;
  reg  [6:0]  rob_uop_3_5_stale_pdst;
  reg         rob_uop_3_5_is_fencei;
  reg         rob_uop_3_5_uses_ldq;
  reg         rob_uop_3_5_uses_stq;
  reg         rob_uop_3_5_is_sys_pc2epc;
  reg         rob_uop_3_5_flush_on_commit;
  reg  [5:0]  rob_uop_3_5_ldst;
  reg         rob_uop_3_5_ldst_val;
  reg  [1:0]  rob_uop_3_5_dst_rtype;
  reg         rob_uop_3_5_fp_val;
  reg  [1:0]  rob_uop_3_5_debug_fsrc;
  reg  [6:0]  rob_uop_3_6_uopc;
  reg         rob_uop_3_6_is_rvc;
  reg         rob_uop_3_6_is_br;
  reg         rob_uop_3_6_is_jalr;
  reg         rob_uop_3_6_is_jal;
  reg  [19:0] rob_uop_3_6_br_mask;
  reg  [5:0]  rob_uop_3_6_ftq_idx;
  reg         rob_uop_3_6_edge_inst;
  reg  [5:0]  rob_uop_3_6_pc_lob;
  reg  [6:0]  rob_uop_3_6_pdst;
  reg  [6:0]  rob_uop_3_6_stale_pdst;
  reg         rob_uop_3_6_is_fencei;
  reg         rob_uop_3_6_uses_ldq;
  reg         rob_uop_3_6_uses_stq;
  reg         rob_uop_3_6_is_sys_pc2epc;
  reg         rob_uop_3_6_flush_on_commit;
  reg  [5:0]  rob_uop_3_6_ldst;
  reg         rob_uop_3_6_ldst_val;
  reg  [1:0]  rob_uop_3_6_dst_rtype;
  reg         rob_uop_3_6_fp_val;
  reg  [1:0]  rob_uop_3_6_debug_fsrc;
  reg  [6:0]  rob_uop_3_7_uopc;
  reg         rob_uop_3_7_is_rvc;
  reg         rob_uop_3_7_is_br;
  reg         rob_uop_3_7_is_jalr;
  reg         rob_uop_3_7_is_jal;
  reg  [19:0] rob_uop_3_7_br_mask;
  reg  [5:0]  rob_uop_3_7_ftq_idx;
  reg         rob_uop_3_7_edge_inst;
  reg  [5:0]  rob_uop_3_7_pc_lob;
  reg  [6:0]  rob_uop_3_7_pdst;
  reg  [6:0]  rob_uop_3_7_stale_pdst;
  reg         rob_uop_3_7_is_fencei;
  reg         rob_uop_3_7_uses_ldq;
  reg         rob_uop_3_7_uses_stq;
  reg         rob_uop_3_7_is_sys_pc2epc;
  reg         rob_uop_3_7_flush_on_commit;
  reg  [5:0]  rob_uop_3_7_ldst;
  reg         rob_uop_3_7_ldst_val;
  reg  [1:0]  rob_uop_3_7_dst_rtype;
  reg         rob_uop_3_7_fp_val;
  reg  [1:0]  rob_uop_3_7_debug_fsrc;
  reg  [6:0]  rob_uop_3_8_uopc;
  reg         rob_uop_3_8_is_rvc;
  reg         rob_uop_3_8_is_br;
  reg         rob_uop_3_8_is_jalr;
  reg         rob_uop_3_8_is_jal;
  reg  [19:0] rob_uop_3_8_br_mask;
  reg  [5:0]  rob_uop_3_8_ftq_idx;
  reg         rob_uop_3_8_edge_inst;
  reg  [5:0]  rob_uop_3_8_pc_lob;
  reg  [6:0]  rob_uop_3_8_pdst;
  reg  [6:0]  rob_uop_3_8_stale_pdst;
  reg         rob_uop_3_8_is_fencei;
  reg         rob_uop_3_8_uses_ldq;
  reg         rob_uop_3_8_uses_stq;
  reg         rob_uop_3_8_is_sys_pc2epc;
  reg         rob_uop_3_8_flush_on_commit;
  reg  [5:0]  rob_uop_3_8_ldst;
  reg         rob_uop_3_8_ldst_val;
  reg  [1:0]  rob_uop_3_8_dst_rtype;
  reg         rob_uop_3_8_fp_val;
  reg  [1:0]  rob_uop_3_8_debug_fsrc;
  reg  [6:0]  rob_uop_3_9_uopc;
  reg         rob_uop_3_9_is_rvc;
  reg         rob_uop_3_9_is_br;
  reg         rob_uop_3_9_is_jalr;
  reg         rob_uop_3_9_is_jal;
  reg  [19:0] rob_uop_3_9_br_mask;
  reg  [5:0]  rob_uop_3_9_ftq_idx;
  reg         rob_uop_3_9_edge_inst;
  reg  [5:0]  rob_uop_3_9_pc_lob;
  reg  [6:0]  rob_uop_3_9_pdst;
  reg  [6:0]  rob_uop_3_9_stale_pdst;
  reg         rob_uop_3_9_is_fencei;
  reg         rob_uop_3_9_uses_ldq;
  reg         rob_uop_3_9_uses_stq;
  reg         rob_uop_3_9_is_sys_pc2epc;
  reg         rob_uop_3_9_flush_on_commit;
  reg  [5:0]  rob_uop_3_9_ldst;
  reg         rob_uop_3_9_ldst_val;
  reg  [1:0]  rob_uop_3_9_dst_rtype;
  reg         rob_uop_3_9_fp_val;
  reg  [1:0]  rob_uop_3_9_debug_fsrc;
  reg  [6:0]  rob_uop_3_10_uopc;
  reg         rob_uop_3_10_is_rvc;
  reg         rob_uop_3_10_is_br;
  reg         rob_uop_3_10_is_jalr;
  reg         rob_uop_3_10_is_jal;
  reg  [19:0] rob_uop_3_10_br_mask;
  reg  [5:0]  rob_uop_3_10_ftq_idx;
  reg         rob_uop_3_10_edge_inst;
  reg  [5:0]  rob_uop_3_10_pc_lob;
  reg  [6:0]  rob_uop_3_10_pdst;
  reg  [6:0]  rob_uop_3_10_stale_pdst;
  reg         rob_uop_3_10_is_fencei;
  reg         rob_uop_3_10_uses_ldq;
  reg         rob_uop_3_10_uses_stq;
  reg         rob_uop_3_10_is_sys_pc2epc;
  reg         rob_uop_3_10_flush_on_commit;
  reg  [5:0]  rob_uop_3_10_ldst;
  reg         rob_uop_3_10_ldst_val;
  reg  [1:0]  rob_uop_3_10_dst_rtype;
  reg         rob_uop_3_10_fp_val;
  reg  [1:0]  rob_uop_3_10_debug_fsrc;
  reg  [6:0]  rob_uop_3_11_uopc;
  reg         rob_uop_3_11_is_rvc;
  reg         rob_uop_3_11_is_br;
  reg         rob_uop_3_11_is_jalr;
  reg         rob_uop_3_11_is_jal;
  reg  [19:0] rob_uop_3_11_br_mask;
  reg  [5:0]  rob_uop_3_11_ftq_idx;
  reg         rob_uop_3_11_edge_inst;
  reg  [5:0]  rob_uop_3_11_pc_lob;
  reg  [6:0]  rob_uop_3_11_pdst;
  reg  [6:0]  rob_uop_3_11_stale_pdst;
  reg         rob_uop_3_11_is_fencei;
  reg         rob_uop_3_11_uses_ldq;
  reg         rob_uop_3_11_uses_stq;
  reg         rob_uop_3_11_is_sys_pc2epc;
  reg         rob_uop_3_11_flush_on_commit;
  reg  [5:0]  rob_uop_3_11_ldst;
  reg         rob_uop_3_11_ldst_val;
  reg  [1:0]  rob_uop_3_11_dst_rtype;
  reg         rob_uop_3_11_fp_val;
  reg  [1:0]  rob_uop_3_11_debug_fsrc;
  reg  [6:0]  rob_uop_3_12_uopc;
  reg         rob_uop_3_12_is_rvc;
  reg         rob_uop_3_12_is_br;
  reg         rob_uop_3_12_is_jalr;
  reg         rob_uop_3_12_is_jal;
  reg  [19:0] rob_uop_3_12_br_mask;
  reg  [5:0]  rob_uop_3_12_ftq_idx;
  reg         rob_uop_3_12_edge_inst;
  reg  [5:0]  rob_uop_3_12_pc_lob;
  reg  [6:0]  rob_uop_3_12_pdst;
  reg  [6:0]  rob_uop_3_12_stale_pdst;
  reg         rob_uop_3_12_is_fencei;
  reg         rob_uop_3_12_uses_ldq;
  reg         rob_uop_3_12_uses_stq;
  reg         rob_uop_3_12_is_sys_pc2epc;
  reg         rob_uop_3_12_flush_on_commit;
  reg  [5:0]  rob_uop_3_12_ldst;
  reg         rob_uop_3_12_ldst_val;
  reg  [1:0]  rob_uop_3_12_dst_rtype;
  reg         rob_uop_3_12_fp_val;
  reg  [1:0]  rob_uop_3_12_debug_fsrc;
  reg  [6:0]  rob_uop_3_13_uopc;
  reg         rob_uop_3_13_is_rvc;
  reg         rob_uop_3_13_is_br;
  reg         rob_uop_3_13_is_jalr;
  reg         rob_uop_3_13_is_jal;
  reg  [19:0] rob_uop_3_13_br_mask;
  reg  [5:0]  rob_uop_3_13_ftq_idx;
  reg         rob_uop_3_13_edge_inst;
  reg  [5:0]  rob_uop_3_13_pc_lob;
  reg  [6:0]  rob_uop_3_13_pdst;
  reg  [6:0]  rob_uop_3_13_stale_pdst;
  reg         rob_uop_3_13_is_fencei;
  reg         rob_uop_3_13_uses_ldq;
  reg         rob_uop_3_13_uses_stq;
  reg         rob_uop_3_13_is_sys_pc2epc;
  reg         rob_uop_3_13_flush_on_commit;
  reg  [5:0]  rob_uop_3_13_ldst;
  reg         rob_uop_3_13_ldst_val;
  reg  [1:0]  rob_uop_3_13_dst_rtype;
  reg         rob_uop_3_13_fp_val;
  reg  [1:0]  rob_uop_3_13_debug_fsrc;
  reg  [6:0]  rob_uop_3_14_uopc;
  reg         rob_uop_3_14_is_rvc;
  reg         rob_uop_3_14_is_br;
  reg         rob_uop_3_14_is_jalr;
  reg         rob_uop_3_14_is_jal;
  reg  [19:0] rob_uop_3_14_br_mask;
  reg  [5:0]  rob_uop_3_14_ftq_idx;
  reg         rob_uop_3_14_edge_inst;
  reg  [5:0]  rob_uop_3_14_pc_lob;
  reg  [6:0]  rob_uop_3_14_pdst;
  reg  [6:0]  rob_uop_3_14_stale_pdst;
  reg         rob_uop_3_14_is_fencei;
  reg         rob_uop_3_14_uses_ldq;
  reg         rob_uop_3_14_uses_stq;
  reg         rob_uop_3_14_is_sys_pc2epc;
  reg         rob_uop_3_14_flush_on_commit;
  reg  [5:0]  rob_uop_3_14_ldst;
  reg         rob_uop_3_14_ldst_val;
  reg  [1:0]  rob_uop_3_14_dst_rtype;
  reg         rob_uop_3_14_fp_val;
  reg  [1:0]  rob_uop_3_14_debug_fsrc;
  reg  [6:0]  rob_uop_3_15_uopc;
  reg         rob_uop_3_15_is_rvc;
  reg         rob_uop_3_15_is_br;
  reg         rob_uop_3_15_is_jalr;
  reg         rob_uop_3_15_is_jal;
  reg  [19:0] rob_uop_3_15_br_mask;
  reg  [5:0]  rob_uop_3_15_ftq_idx;
  reg         rob_uop_3_15_edge_inst;
  reg  [5:0]  rob_uop_3_15_pc_lob;
  reg  [6:0]  rob_uop_3_15_pdst;
  reg  [6:0]  rob_uop_3_15_stale_pdst;
  reg         rob_uop_3_15_is_fencei;
  reg         rob_uop_3_15_uses_ldq;
  reg         rob_uop_3_15_uses_stq;
  reg         rob_uop_3_15_is_sys_pc2epc;
  reg         rob_uop_3_15_flush_on_commit;
  reg  [5:0]  rob_uop_3_15_ldst;
  reg         rob_uop_3_15_ldst_val;
  reg  [1:0]  rob_uop_3_15_dst_rtype;
  reg         rob_uop_3_15_fp_val;
  reg  [1:0]  rob_uop_3_15_debug_fsrc;
  reg  [6:0]  rob_uop_3_16_uopc;
  reg         rob_uop_3_16_is_rvc;
  reg         rob_uop_3_16_is_br;
  reg         rob_uop_3_16_is_jalr;
  reg         rob_uop_3_16_is_jal;
  reg  [19:0] rob_uop_3_16_br_mask;
  reg  [5:0]  rob_uop_3_16_ftq_idx;
  reg         rob_uop_3_16_edge_inst;
  reg  [5:0]  rob_uop_3_16_pc_lob;
  reg  [6:0]  rob_uop_3_16_pdst;
  reg  [6:0]  rob_uop_3_16_stale_pdst;
  reg         rob_uop_3_16_is_fencei;
  reg         rob_uop_3_16_uses_ldq;
  reg         rob_uop_3_16_uses_stq;
  reg         rob_uop_3_16_is_sys_pc2epc;
  reg         rob_uop_3_16_flush_on_commit;
  reg  [5:0]  rob_uop_3_16_ldst;
  reg         rob_uop_3_16_ldst_val;
  reg  [1:0]  rob_uop_3_16_dst_rtype;
  reg         rob_uop_3_16_fp_val;
  reg  [1:0]  rob_uop_3_16_debug_fsrc;
  reg  [6:0]  rob_uop_3_17_uopc;
  reg         rob_uop_3_17_is_rvc;
  reg         rob_uop_3_17_is_br;
  reg         rob_uop_3_17_is_jalr;
  reg         rob_uop_3_17_is_jal;
  reg  [19:0] rob_uop_3_17_br_mask;
  reg  [5:0]  rob_uop_3_17_ftq_idx;
  reg         rob_uop_3_17_edge_inst;
  reg  [5:0]  rob_uop_3_17_pc_lob;
  reg  [6:0]  rob_uop_3_17_pdst;
  reg  [6:0]  rob_uop_3_17_stale_pdst;
  reg         rob_uop_3_17_is_fencei;
  reg         rob_uop_3_17_uses_ldq;
  reg         rob_uop_3_17_uses_stq;
  reg         rob_uop_3_17_is_sys_pc2epc;
  reg         rob_uop_3_17_flush_on_commit;
  reg  [5:0]  rob_uop_3_17_ldst;
  reg         rob_uop_3_17_ldst_val;
  reg  [1:0]  rob_uop_3_17_dst_rtype;
  reg         rob_uop_3_17_fp_val;
  reg  [1:0]  rob_uop_3_17_debug_fsrc;
  reg  [6:0]  rob_uop_3_18_uopc;
  reg         rob_uop_3_18_is_rvc;
  reg         rob_uop_3_18_is_br;
  reg         rob_uop_3_18_is_jalr;
  reg         rob_uop_3_18_is_jal;
  reg  [19:0] rob_uop_3_18_br_mask;
  reg  [5:0]  rob_uop_3_18_ftq_idx;
  reg         rob_uop_3_18_edge_inst;
  reg  [5:0]  rob_uop_3_18_pc_lob;
  reg  [6:0]  rob_uop_3_18_pdst;
  reg  [6:0]  rob_uop_3_18_stale_pdst;
  reg         rob_uop_3_18_is_fencei;
  reg         rob_uop_3_18_uses_ldq;
  reg         rob_uop_3_18_uses_stq;
  reg         rob_uop_3_18_is_sys_pc2epc;
  reg         rob_uop_3_18_flush_on_commit;
  reg  [5:0]  rob_uop_3_18_ldst;
  reg         rob_uop_3_18_ldst_val;
  reg  [1:0]  rob_uop_3_18_dst_rtype;
  reg         rob_uop_3_18_fp_val;
  reg  [1:0]  rob_uop_3_18_debug_fsrc;
  reg  [6:0]  rob_uop_3_19_uopc;
  reg         rob_uop_3_19_is_rvc;
  reg         rob_uop_3_19_is_br;
  reg         rob_uop_3_19_is_jalr;
  reg         rob_uop_3_19_is_jal;
  reg  [19:0] rob_uop_3_19_br_mask;
  reg  [5:0]  rob_uop_3_19_ftq_idx;
  reg         rob_uop_3_19_edge_inst;
  reg  [5:0]  rob_uop_3_19_pc_lob;
  reg  [6:0]  rob_uop_3_19_pdst;
  reg  [6:0]  rob_uop_3_19_stale_pdst;
  reg         rob_uop_3_19_is_fencei;
  reg         rob_uop_3_19_uses_ldq;
  reg         rob_uop_3_19_uses_stq;
  reg         rob_uop_3_19_is_sys_pc2epc;
  reg         rob_uop_3_19_flush_on_commit;
  reg  [5:0]  rob_uop_3_19_ldst;
  reg         rob_uop_3_19_ldst_val;
  reg  [1:0]  rob_uop_3_19_dst_rtype;
  reg         rob_uop_3_19_fp_val;
  reg  [1:0]  rob_uop_3_19_debug_fsrc;
  reg  [6:0]  rob_uop_3_20_uopc;
  reg         rob_uop_3_20_is_rvc;
  reg         rob_uop_3_20_is_br;
  reg         rob_uop_3_20_is_jalr;
  reg         rob_uop_3_20_is_jal;
  reg  [19:0] rob_uop_3_20_br_mask;
  reg  [5:0]  rob_uop_3_20_ftq_idx;
  reg         rob_uop_3_20_edge_inst;
  reg  [5:0]  rob_uop_3_20_pc_lob;
  reg  [6:0]  rob_uop_3_20_pdst;
  reg  [6:0]  rob_uop_3_20_stale_pdst;
  reg         rob_uop_3_20_is_fencei;
  reg         rob_uop_3_20_uses_ldq;
  reg         rob_uop_3_20_uses_stq;
  reg         rob_uop_3_20_is_sys_pc2epc;
  reg         rob_uop_3_20_flush_on_commit;
  reg  [5:0]  rob_uop_3_20_ldst;
  reg         rob_uop_3_20_ldst_val;
  reg  [1:0]  rob_uop_3_20_dst_rtype;
  reg         rob_uop_3_20_fp_val;
  reg  [1:0]  rob_uop_3_20_debug_fsrc;
  reg  [6:0]  rob_uop_3_21_uopc;
  reg         rob_uop_3_21_is_rvc;
  reg         rob_uop_3_21_is_br;
  reg         rob_uop_3_21_is_jalr;
  reg         rob_uop_3_21_is_jal;
  reg  [19:0] rob_uop_3_21_br_mask;
  reg  [5:0]  rob_uop_3_21_ftq_idx;
  reg         rob_uop_3_21_edge_inst;
  reg  [5:0]  rob_uop_3_21_pc_lob;
  reg  [6:0]  rob_uop_3_21_pdst;
  reg  [6:0]  rob_uop_3_21_stale_pdst;
  reg         rob_uop_3_21_is_fencei;
  reg         rob_uop_3_21_uses_ldq;
  reg         rob_uop_3_21_uses_stq;
  reg         rob_uop_3_21_is_sys_pc2epc;
  reg         rob_uop_3_21_flush_on_commit;
  reg  [5:0]  rob_uop_3_21_ldst;
  reg         rob_uop_3_21_ldst_val;
  reg  [1:0]  rob_uop_3_21_dst_rtype;
  reg         rob_uop_3_21_fp_val;
  reg  [1:0]  rob_uop_3_21_debug_fsrc;
  reg  [6:0]  rob_uop_3_22_uopc;
  reg         rob_uop_3_22_is_rvc;
  reg         rob_uop_3_22_is_br;
  reg         rob_uop_3_22_is_jalr;
  reg         rob_uop_3_22_is_jal;
  reg  [19:0] rob_uop_3_22_br_mask;
  reg  [5:0]  rob_uop_3_22_ftq_idx;
  reg         rob_uop_3_22_edge_inst;
  reg  [5:0]  rob_uop_3_22_pc_lob;
  reg  [6:0]  rob_uop_3_22_pdst;
  reg  [6:0]  rob_uop_3_22_stale_pdst;
  reg         rob_uop_3_22_is_fencei;
  reg         rob_uop_3_22_uses_ldq;
  reg         rob_uop_3_22_uses_stq;
  reg         rob_uop_3_22_is_sys_pc2epc;
  reg         rob_uop_3_22_flush_on_commit;
  reg  [5:0]  rob_uop_3_22_ldst;
  reg         rob_uop_3_22_ldst_val;
  reg  [1:0]  rob_uop_3_22_dst_rtype;
  reg         rob_uop_3_22_fp_val;
  reg  [1:0]  rob_uop_3_22_debug_fsrc;
  reg  [6:0]  rob_uop_3_23_uopc;
  reg         rob_uop_3_23_is_rvc;
  reg         rob_uop_3_23_is_br;
  reg         rob_uop_3_23_is_jalr;
  reg         rob_uop_3_23_is_jal;
  reg  [19:0] rob_uop_3_23_br_mask;
  reg  [5:0]  rob_uop_3_23_ftq_idx;
  reg         rob_uop_3_23_edge_inst;
  reg  [5:0]  rob_uop_3_23_pc_lob;
  reg  [6:0]  rob_uop_3_23_pdst;
  reg  [6:0]  rob_uop_3_23_stale_pdst;
  reg         rob_uop_3_23_is_fencei;
  reg         rob_uop_3_23_uses_ldq;
  reg         rob_uop_3_23_uses_stq;
  reg         rob_uop_3_23_is_sys_pc2epc;
  reg         rob_uop_3_23_flush_on_commit;
  reg  [5:0]  rob_uop_3_23_ldst;
  reg         rob_uop_3_23_ldst_val;
  reg  [1:0]  rob_uop_3_23_dst_rtype;
  reg         rob_uop_3_23_fp_val;
  reg  [1:0]  rob_uop_3_23_debug_fsrc;
  reg  [6:0]  rob_uop_3_24_uopc;
  reg         rob_uop_3_24_is_rvc;
  reg         rob_uop_3_24_is_br;
  reg         rob_uop_3_24_is_jalr;
  reg         rob_uop_3_24_is_jal;
  reg  [19:0] rob_uop_3_24_br_mask;
  reg  [5:0]  rob_uop_3_24_ftq_idx;
  reg         rob_uop_3_24_edge_inst;
  reg  [5:0]  rob_uop_3_24_pc_lob;
  reg  [6:0]  rob_uop_3_24_pdst;
  reg  [6:0]  rob_uop_3_24_stale_pdst;
  reg         rob_uop_3_24_is_fencei;
  reg         rob_uop_3_24_uses_ldq;
  reg         rob_uop_3_24_uses_stq;
  reg         rob_uop_3_24_is_sys_pc2epc;
  reg         rob_uop_3_24_flush_on_commit;
  reg  [5:0]  rob_uop_3_24_ldst;
  reg         rob_uop_3_24_ldst_val;
  reg  [1:0]  rob_uop_3_24_dst_rtype;
  reg         rob_uop_3_24_fp_val;
  reg  [1:0]  rob_uop_3_24_debug_fsrc;
  reg  [6:0]  rob_uop_3_25_uopc;
  reg         rob_uop_3_25_is_rvc;
  reg         rob_uop_3_25_is_br;
  reg         rob_uop_3_25_is_jalr;
  reg         rob_uop_3_25_is_jal;
  reg  [19:0] rob_uop_3_25_br_mask;
  reg  [5:0]  rob_uop_3_25_ftq_idx;
  reg         rob_uop_3_25_edge_inst;
  reg  [5:0]  rob_uop_3_25_pc_lob;
  reg  [6:0]  rob_uop_3_25_pdst;
  reg  [6:0]  rob_uop_3_25_stale_pdst;
  reg         rob_uop_3_25_is_fencei;
  reg         rob_uop_3_25_uses_ldq;
  reg         rob_uop_3_25_uses_stq;
  reg         rob_uop_3_25_is_sys_pc2epc;
  reg         rob_uop_3_25_flush_on_commit;
  reg  [5:0]  rob_uop_3_25_ldst;
  reg         rob_uop_3_25_ldst_val;
  reg  [1:0]  rob_uop_3_25_dst_rtype;
  reg         rob_uop_3_25_fp_val;
  reg  [1:0]  rob_uop_3_25_debug_fsrc;
  reg  [6:0]  rob_uop_3_26_uopc;
  reg         rob_uop_3_26_is_rvc;
  reg         rob_uop_3_26_is_br;
  reg         rob_uop_3_26_is_jalr;
  reg         rob_uop_3_26_is_jal;
  reg  [19:0] rob_uop_3_26_br_mask;
  reg  [5:0]  rob_uop_3_26_ftq_idx;
  reg         rob_uop_3_26_edge_inst;
  reg  [5:0]  rob_uop_3_26_pc_lob;
  reg  [6:0]  rob_uop_3_26_pdst;
  reg  [6:0]  rob_uop_3_26_stale_pdst;
  reg         rob_uop_3_26_is_fencei;
  reg         rob_uop_3_26_uses_ldq;
  reg         rob_uop_3_26_uses_stq;
  reg         rob_uop_3_26_is_sys_pc2epc;
  reg         rob_uop_3_26_flush_on_commit;
  reg  [5:0]  rob_uop_3_26_ldst;
  reg         rob_uop_3_26_ldst_val;
  reg  [1:0]  rob_uop_3_26_dst_rtype;
  reg         rob_uop_3_26_fp_val;
  reg  [1:0]  rob_uop_3_26_debug_fsrc;
  reg  [6:0]  rob_uop_3_27_uopc;
  reg         rob_uop_3_27_is_rvc;
  reg         rob_uop_3_27_is_br;
  reg         rob_uop_3_27_is_jalr;
  reg         rob_uop_3_27_is_jal;
  reg  [19:0] rob_uop_3_27_br_mask;
  reg  [5:0]  rob_uop_3_27_ftq_idx;
  reg         rob_uop_3_27_edge_inst;
  reg  [5:0]  rob_uop_3_27_pc_lob;
  reg  [6:0]  rob_uop_3_27_pdst;
  reg  [6:0]  rob_uop_3_27_stale_pdst;
  reg         rob_uop_3_27_is_fencei;
  reg         rob_uop_3_27_uses_ldq;
  reg         rob_uop_3_27_uses_stq;
  reg         rob_uop_3_27_is_sys_pc2epc;
  reg         rob_uop_3_27_flush_on_commit;
  reg  [5:0]  rob_uop_3_27_ldst;
  reg         rob_uop_3_27_ldst_val;
  reg  [1:0]  rob_uop_3_27_dst_rtype;
  reg         rob_uop_3_27_fp_val;
  reg  [1:0]  rob_uop_3_27_debug_fsrc;
  reg  [6:0]  rob_uop_3_28_uopc;
  reg         rob_uop_3_28_is_rvc;
  reg         rob_uop_3_28_is_br;
  reg         rob_uop_3_28_is_jalr;
  reg         rob_uop_3_28_is_jal;
  reg  [19:0] rob_uop_3_28_br_mask;
  reg  [5:0]  rob_uop_3_28_ftq_idx;
  reg         rob_uop_3_28_edge_inst;
  reg  [5:0]  rob_uop_3_28_pc_lob;
  reg  [6:0]  rob_uop_3_28_pdst;
  reg  [6:0]  rob_uop_3_28_stale_pdst;
  reg         rob_uop_3_28_is_fencei;
  reg         rob_uop_3_28_uses_ldq;
  reg         rob_uop_3_28_uses_stq;
  reg         rob_uop_3_28_is_sys_pc2epc;
  reg         rob_uop_3_28_flush_on_commit;
  reg  [5:0]  rob_uop_3_28_ldst;
  reg         rob_uop_3_28_ldst_val;
  reg  [1:0]  rob_uop_3_28_dst_rtype;
  reg         rob_uop_3_28_fp_val;
  reg  [1:0]  rob_uop_3_28_debug_fsrc;
  reg  [6:0]  rob_uop_3_29_uopc;
  reg         rob_uop_3_29_is_rvc;
  reg         rob_uop_3_29_is_br;
  reg         rob_uop_3_29_is_jalr;
  reg         rob_uop_3_29_is_jal;
  reg  [19:0] rob_uop_3_29_br_mask;
  reg  [5:0]  rob_uop_3_29_ftq_idx;
  reg         rob_uop_3_29_edge_inst;
  reg  [5:0]  rob_uop_3_29_pc_lob;
  reg  [6:0]  rob_uop_3_29_pdst;
  reg  [6:0]  rob_uop_3_29_stale_pdst;
  reg         rob_uop_3_29_is_fencei;
  reg         rob_uop_3_29_uses_ldq;
  reg         rob_uop_3_29_uses_stq;
  reg         rob_uop_3_29_is_sys_pc2epc;
  reg         rob_uop_3_29_flush_on_commit;
  reg  [5:0]  rob_uop_3_29_ldst;
  reg         rob_uop_3_29_ldst_val;
  reg  [1:0]  rob_uop_3_29_dst_rtype;
  reg         rob_uop_3_29_fp_val;
  reg  [1:0]  rob_uop_3_29_debug_fsrc;
  reg  [6:0]  rob_uop_3_30_uopc;
  reg         rob_uop_3_30_is_rvc;
  reg         rob_uop_3_30_is_br;
  reg         rob_uop_3_30_is_jalr;
  reg         rob_uop_3_30_is_jal;
  reg  [19:0] rob_uop_3_30_br_mask;
  reg  [5:0]  rob_uop_3_30_ftq_idx;
  reg         rob_uop_3_30_edge_inst;
  reg  [5:0]  rob_uop_3_30_pc_lob;
  reg  [6:0]  rob_uop_3_30_pdst;
  reg  [6:0]  rob_uop_3_30_stale_pdst;
  reg         rob_uop_3_30_is_fencei;
  reg         rob_uop_3_30_uses_ldq;
  reg         rob_uop_3_30_uses_stq;
  reg         rob_uop_3_30_is_sys_pc2epc;
  reg         rob_uop_3_30_flush_on_commit;
  reg  [5:0]  rob_uop_3_30_ldst;
  reg         rob_uop_3_30_ldst_val;
  reg  [1:0]  rob_uop_3_30_dst_rtype;
  reg         rob_uop_3_30_fp_val;
  reg  [1:0]  rob_uop_3_30_debug_fsrc;
  reg  [6:0]  rob_uop_3_31_uopc;
  reg         rob_uop_3_31_is_rvc;
  reg         rob_uop_3_31_is_br;
  reg         rob_uop_3_31_is_jalr;
  reg         rob_uop_3_31_is_jal;
  reg  [19:0] rob_uop_3_31_br_mask;
  reg  [5:0]  rob_uop_3_31_ftq_idx;
  reg         rob_uop_3_31_edge_inst;
  reg  [5:0]  rob_uop_3_31_pc_lob;
  reg  [6:0]  rob_uop_3_31_pdst;
  reg  [6:0]  rob_uop_3_31_stale_pdst;
  reg         rob_uop_3_31_is_fencei;
  reg         rob_uop_3_31_uses_ldq;
  reg         rob_uop_3_31_uses_stq;
  reg         rob_uop_3_31_is_sys_pc2epc;
  reg         rob_uop_3_31_flush_on_commit;
  reg  [5:0]  rob_uop_3_31_ldst;
  reg         rob_uop_3_31_ldst_val;
  reg  [1:0]  rob_uop_3_31_dst_rtype;
  reg         rob_uop_3_31_fp_val;
  reg  [1:0]  rob_uop_3_31_debug_fsrc;
  reg         rob_exception_3_0;
  reg         rob_exception_3_1;
  reg         rob_exception_3_2;
  reg         rob_exception_3_3;
  reg         rob_exception_3_4;
  reg         rob_exception_3_5;
  reg         rob_exception_3_6;
  reg         rob_exception_3_7;
  reg         rob_exception_3_8;
  reg         rob_exception_3_9;
  reg         rob_exception_3_10;
  reg         rob_exception_3_11;
  reg         rob_exception_3_12;
  reg         rob_exception_3_13;
  reg         rob_exception_3_14;
  reg         rob_exception_3_15;
  reg         rob_exception_3_16;
  reg         rob_exception_3_17;
  reg         rob_exception_3_18;
  reg         rob_exception_3_19;
  reg         rob_exception_3_20;
  reg         rob_exception_3_21;
  reg         rob_exception_3_22;
  reg         rob_exception_3_23;
  reg         rob_exception_3_24;
  reg         rob_exception_3_25;
  reg         rob_exception_3_26;
  reg         rob_exception_3_27;
  reg         rob_exception_3_28;
  reg         rob_exception_3_29;
  reg         rob_exception_3_30;
  reg         rob_exception_3_31;
  reg         rob_predicated_3_0;
  reg         rob_predicated_3_1;
  reg         rob_predicated_3_2;
  reg         rob_predicated_3_3;
  reg         rob_predicated_3_4;
  reg         rob_predicated_3_5;
  reg         rob_predicated_3_6;
  reg         rob_predicated_3_7;
  reg         rob_predicated_3_8;
  reg         rob_predicated_3_9;
  reg         rob_predicated_3_10;
  reg         rob_predicated_3_11;
  reg         rob_predicated_3_12;
  reg         rob_predicated_3_13;
  reg         rob_predicated_3_14;
  reg         rob_predicated_3_15;
  reg         rob_predicated_3_16;
  reg         rob_predicated_3_17;
  reg         rob_predicated_3_18;
  reg         rob_predicated_3_19;
  reg         rob_predicated_3_20;
  reg         rob_predicated_3_21;
  reg         rob_predicated_3_22;
  reg         rob_predicated_3_23;
  reg         rob_predicated_3_24;
  reg         rob_predicated_3_25;
  reg         rob_predicated_3_26;
  reg         rob_predicated_3_27;
  reg         rob_predicated_3_28;
  reg         rob_predicated_3_29;
  reg         rob_predicated_3_30;
  reg         rob_predicated_3_31;
  reg         casez_tmp_233;
  always @(*) begin
    casez (rob_tail)
      5'b00000:
        casez_tmp_233 = rob_val_3_0;
      5'b00001:
        casez_tmp_233 = rob_val_3_1;
      5'b00010:
        casez_tmp_233 = rob_val_3_2;
      5'b00011:
        casez_tmp_233 = rob_val_3_3;
      5'b00100:
        casez_tmp_233 = rob_val_3_4;
      5'b00101:
        casez_tmp_233 = rob_val_3_5;
      5'b00110:
        casez_tmp_233 = rob_val_3_6;
      5'b00111:
        casez_tmp_233 = rob_val_3_7;
      5'b01000:
        casez_tmp_233 = rob_val_3_8;
      5'b01001:
        casez_tmp_233 = rob_val_3_9;
      5'b01010:
        casez_tmp_233 = rob_val_3_10;
      5'b01011:
        casez_tmp_233 = rob_val_3_11;
      5'b01100:
        casez_tmp_233 = rob_val_3_12;
      5'b01101:
        casez_tmp_233 = rob_val_3_13;
      5'b01110:
        casez_tmp_233 = rob_val_3_14;
      5'b01111:
        casez_tmp_233 = rob_val_3_15;
      5'b10000:
        casez_tmp_233 = rob_val_3_16;
      5'b10001:
        casez_tmp_233 = rob_val_3_17;
      5'b10010:
        casez_tmp_233 = rob_val_3_18;
      5'b10011:
        casez_tmp_233 = rob_val_3_19;
      5'b10100:
        casez_tmp_233 = rob_val_3_20;
      5'b10101:
        casez_tmp_233 = rob_val_3_21;
      5'b10110:
        casez_tmp_233 = rob_val_3_22;
      5'b10111:
        casez_tmp_233 = rob_val_3_23;
      5'b11000:
        casez_tmp_233 = rob_val_3_24;
      5'b11001:
        casez_tmp_233 = rob_val_3_25;
      5'b11010:
        casez_tmp_233 = rob_val_3_26;
      5'b11011:
        casez_tmp_233 = rob_val_3_27;
      5'b11100:
        casez_tmp_233 = rob_val_3_28;
      5'b11101:
        casez_tmp_233 = rob_val_3_29;
      5'b11110:
        casez_tmp_233 = rob_val_3_30;
      default:
        casez_tmp_233 = rob_val_3_31;
    endcase
  end // always @(*)
  wire        _GEN_49 = io_wb_resps_0_valid & (&(io_wb_resps_0_bits_uop_rob_idx[1:0]));
  wire        _GEN_50 = io_wb_resps_1_valid & (&(io_wb_resps_1_bits_uop_rob_idx[1:0]));
  wire        _GEN_51 = io_wb_resps_2_valid & (&(io_wb_resps_2_bits_uop_rob_idx[1:0]));
  wire        _GEN_52 = io_wb_resps_3_valid & (&(io_wb_resps_3_bits_uop_rob_idx[1:0]));
  wire        _GEN_53 = io_wb_resps_4_valid & (&(io_wb_resps_4_bits_uop_rob_idx[1:0]));
  wire        _GEN_54 = io_wb_resps_5_valid & (&(io_wb_resps_5_bits_uop_rob_idx[1:0]));
  wire        _GEN_55 = io_wb_resps_6_valid & (&(io_wb_resps_6_bits_uop_rob_idx[1:0]));
  wire        _GEN_56 = io_wb_resps_7_valid & (&(io_wb_resps_7_bits_uop_rob_idx[1:0]));
  wire        _GEN_57 = io_wb_resps_8_valid & (&(io_wb_resps_8_bits_uop_rob_idx[1:0]));
  wire        _GEN_58 = io_wb_resps_9_valid & (&(io_wb_resps_9_bits_uop_rob_idx[1:0]));
  wire        _GEN_59 = io_lsu_clr_bsy_0_valid & (&(io_lsu_clr_bsy_0_bits[1:0]));
  reg         casez_tmp_234;
  always @(*) begin
    casez (io_lsu_clr_bsy_0_bits[6:2])
      5'b00000:
        casez_tmp_234 = rob_val_3_0;
      5'b00001:
        casez_tmp_234 = rob_val_3_1;
      5'b00010:
        casez_tmp_234 = rob_val_3_2;
      5'b00011:
        casez_tmp_234 = rob_val_3_3;
      5'b00100:
        casez_tmp_234 = rob_val_3_4;
      5'b00101:
        casez_tmp_234 = rob_val_3_5;
      5'b00110:
        casez_tmp_234 = rob_val_3_6;
      5'b00111:
        casez_tmp_234 = rob_val_3_7;
      5'b01000:
        casez_tmp_234 = rob_val_3_8;
      5'b01001:
        casez_tmp_234 = rob_val_3_9;
      5'b01010:
        casez_tmp_234 = rob_val_3_10;
      5'b01011:
        casez_tmp_234 = rob_val_3_11;
      5'b01100:
        casez_tmp_234 = rob_val_3_12;
      5'b01101:
        casez_tmp_234 = rob_val_3_13;
      5'b01110:
        casez_tmp_234 = rob_val_3_14;
      5'b01111:
        casez_tmp_234 = rob_val_3_15;
      5'b10000:
        casez_tmp_234 = rob_val_3_16;
      5'b10001:
        casez_tmp_234 = rob_val_3_17;
      5'b10010:
        casez_tmp_234 = rob_val_3_18;
      5'b10011:
        casez_tmp_234 = rob_val_3_19;
      5'b10100:
        casez_tmp_234 = rob_val_3_20;
      5'b10101:
        casez_tmp_234 = rob_val_3_21;
      5'b10110:
        casez_tmp_234 = rob_val_3_22;
      5'b10111:
        casez_tmp_234 = rob_val_3_23;
      5'b11000:
        casez_tmp_234 = rob_val_3_24;
      5'b11001:
        casez_tmp_234 = rob_val_3_25;
      5'b11010:
        casez_tmp_234 = rob_val_3_26;
      5'b11011:
        casez_tmp_234 = rob_val_3_27;
      5'b11100:
        casez_tmp_234 = rob_val_3_28;
      5'b11101:
        casez_tmp_234 = rob_val_3_29;
      5'b11110:
        casez_tmp_234 = rob_val_3_30;
      default:
        casez_tmp_234 = rob_val_3_31;
    endcase
  end // always @(*)
  reg         casez_tmp_235;
  always @(*) begin
    casez (io_lsu_clr_bsy_0_bits[6:2])
      5'b00000:
        casez_tmp_235 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_235 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_235 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_235 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_235 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_235 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_235 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_235 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_235 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_235 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_235 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_235 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_235 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_235 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_235 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_235 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_235 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_235 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_235 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_235 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_235 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_235 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_235 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_235 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_235 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_235 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_235 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_235 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_235 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_235 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_235 = rob_bsy_3_30;
      default:
        casez_tmp_235 = rob_bsy_3_31;
    endcase
  end // always @(*)
  wire        _GEN_60 = io_lsu_clr_bsy_1_valid & (&(io_lsu_clr_bsy_1_bits[1:0]));
  reg         casez_tmp_236;
  always @(*) begin
    casez (io_lsu_clr_bsy_1_bits[6:2])
      5'b00000:
        casez_tmp_236 = rob_val_3_0;
      5'b00001:
        casez_tmp_236 = rob_val_3_1;
      5'b00010:
        casez_tmp_236 = rob_val_3_2;
      5'b00011:
        casez_tmp_236 = rob_val_3_3;
      5'b00100:
        casez_tmp_236 = rob_val_3_4;
      5'b00101:
        casez_tmp_236 = rob_val_3_5;
      5'b00110:
        casez_tmp_236 = rob_val_3_6;
      5'b00111:
        casez_tmp_236 = rob_val_3_7;
      5'b01000:
        casez_tmp_236 = rob_val_3_8;
      5'b01001:
        casez_tmp_236 = rob_val_3_9;
      5'b01010:
        casez_tmp_236 = rob_val_3_10;
      5'b01011:
        casez_tmp_236 = rob_val_3_11;
      5'b01100:
        casez_tmp_236 = rob_val_3_12;
      5'b01101:
        casez_tmp_236 = rob_val_3_13;
      5'b01110:
        casez_tmp_236 = rob_val_3_14;
      5'b01111:
        casez_tmp_236 = rob_val_3_15;
      5'b10000:
        casez_tmp_236 = rob_val_3_16;
      5'b10001:
        casez_tmp_236 = rob_val_3_17;
      5'b10010:
        casez_tmp_236 = rob_val_3_18;
      5'b10011:
        casez_tmp_236 = rob_val_3_19;
      5'b10100:
        casez_tmp_236 = rob_val_3_20;
      5'b10101:
        casez_tmp_236 = rob_val_3_21;
      5'b10110:
        casez_tmp_236 = rob_val_3_22;
      5'b10111:
        casez_tmp_236 = rob_val_3_23;
      5'b11000:
        casez_tmp_236 = rob_val_3_24;
      5'b11001:
        casez_tmp_236 = rob_val_3_25;
      5'b11010:
        casez_tmp_236 = rob_val_3_26;
      5'b11011:
        casez_tmp_236 = rob_val_3_27;
      5'b11100:
        casez_tmp_236 = rob_val_3_28;
      5'b11101:
        casez_tmp_236 = rob_val_3_29;
      5'b11110:
        casez_tmp_236 = rob_val_3_30;
      default:
        casez_tmp_236 = rob_val_3_31;
    endcase
  end // always @(*)
  reg         casez_tmp_237;
  always @(*) begin
    casez (io_lsu_clr_bsy_1_bits[6:2])
      5'b00000:
        casez_tmp_237 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_237 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_237 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_237 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_237 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_237 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_237 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_237 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_237 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_237 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_237 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_237 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_237 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_237 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_237 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_237 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_237 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_237 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_237 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_237 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_237 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_237 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_237 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_237 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_237 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_237 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_237 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_237 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_237 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_237 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_237 = rob_bsy_3_30;
      default:
        casez_tmp_237 = rob_bsy_3_31;
    endcase
  end // always @(*)
  wire        _GEN_61 = io_lsu_clr_bsy_2_valid & (&(io_lsu_clr_bsy_2_bits[1:0]));
  reg         casez_tmp_238;
  always @(*) begin
    casez (io_lsu_clr_bsy_2_bits[6:2])
      5'b00000:
        casez_tmp_238 = rob_val_3_0;
      5'b00001:
        casez_tmp_238 = rob_val_3_1;
      5'b00010:
        casez_tmp_238 = rob_val_3_2;
      5'b00011:
        casez_tmp_238 = rob_val_3_3;
      5'b00100:
        casez_tmp_238 = rob_val_3_4;
      5'b00101:
        casez_tmp_238 = rob_val_3_5;
      5'b00110:
        casez_tmp_238 = rob_val_3_6;
      5'b00111:
        casez_tmp_238 = rob_val_3_7;
      5'b01000:
        casez_tmp_238 = rob_val_3_8;
      5'b01001:
        casez_tmp_238 = rob_val_3_9;
      5'b01010:
        casez_tmp_238 = rob_val_3_10;
      5'b01011:
        casez_tmp_238 = rob_val_3_11;
      5'b01100:
        casez_tmp_238 = rob_val_3_12;
      5'b01101:
        casez_tmp_238 = rob_val_3_13;
      5'b01110:
        casez_tmp_238 = rob_val_3_14;
      5'b01111:
        casez_tmp_238 = rob_val_3_15;
      5'b10000:
        casez_tmp_238 = rob_val_3_16;
      5'b10001:
        casez_tmp_238 = rob_val_3_17;
      5'b10010:
        casez_tmp_238 = rob_val_3_18;
      5'b10011:
        casez_tmp_238 = rob_val_3_19;
      5'b10100:
        casez_tmp_238 = rob_val_3_20;
      5'b10101:
        casez_tmp_238 = rob_val_3_21;
      5'b10110:
        casez_tmp_238 = rob_val_3_22;
      5'b10111:
        casez_tmp_238 = rob_val_3_23;
      5'b11000:
        casez_tmp_238 = rob_val_3_24;
      5'b11001:
        casez_tmp_238 = rob_val_3_25;
      5'b11010:
        casez_tmp_238 = rob_val_3_26;
      5'b11011:
        casez_tmp_238 = rob_val_3_27;
      5'b11100:
        casez_tmp_238 = rob_val_3_28;
      5'b11101:
        casez_tmp_238 = rob_val_3_29;
      5'b11110:
        casez_tmp_238 = rob_val_3_30;
      default:
        casez_tmp_238 = rob_val_3_31;
    endcase
  end // always @(*)
  reg         casez_tmp_239;
  always @(*) begin
    casez (io_lsu_clr_bsy_2_bits[6:2])
      5'b00000:
        casez_tmp_239 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_239 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_239 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_239 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_239 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_239 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_239 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_239 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_239 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_239 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_239 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_239 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_239 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_239 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_239 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_239 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_239 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_239 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_239 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_239 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_239 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_239 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_239 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_239 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_239 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_239 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_239 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_239 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_239 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_239 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_239 = rob_bsy_3_30;
      default:
        casez_tmp_239 = rob_bsy_3_31;
    endcase
  end // always @(*)
  wire        _GEN_62 = io_lxcpt_valid & (&(io_lxcpt_bits_uop_rob_idx[1:0]));
  wire        _GEN_63 = _GEN_62 & _GEN_13 & ~reset;
  reg         casez_tmp_240;
  always @(*) begin
    casez (io_lxcpt_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_240 = rob_unsafe_3_0;
      5'b00001:
        casez_tmp_240 = rob_unsafe_3_1;
      5'b00010:
        casez_tmp_240 = rob_unsafe_3_2;
      5'b00011:
        casez_tmp_240 = rob_unsafe_3_3;
      5'b00100:
        casez_tmp_240 = rob_unsafe_3_4;
      5'b00101:
        casez_tmp_240 = rob_unsafe_3_5;
      5'b00110:
        casez_tmp_240 = rob_unsafe_3_6;
      5'b00111:
        casez_tmp_240 = rob_unsafe_3_7;
      5'b01000:
        casez_tmp_240 = rob_unsafe_3_8;
      5'b01001:
        casez_tmp_240 = rob_unsafe_3_9;
      5'b01010:
        casez_tmp_240 = rob_unsafe_3_10;
      5'b01011:
        casez_tmp_240 = rob_unsafe_3_11;
      5'b01100:
        casez_tmp_240 = rob_unsafe_3_12;
      5'b01101:
        casez_tmp_240 = rob_unsafe_3_13;
      5'b01110:
        casez_tmp_240 = rob_unsafe_3_14;
      5'b01111:
        casez_tmp_240 = rob_unsafe_3_15;
      5'b10000:
        casez_tmp_240 = rob_unsafe_3_16;
      5'b10001:
        casez_tmp_240 = rob_unsafe_3_17;
      5'b10010:
        casez_tmp_240 = rob_unsafe_3_18;
      5'b10011:
        casez_tmp_240 = rob_unsafe_3_19;
      5'b10100:
        casez_tmp_240 = rob_unsafe_3_20;
      5'b10101:
        casez_tmp_240 = rob_unsafe_3_21;
      5'b10110:
        casez_tmp_240 = rob_unsafe_3_22;
      5'b10111:
        casez_tmp_240 = rob_unsafe_3_23;
      5'b11000:
        casez_tmp_240 = rob_unsafe_3_24;
      5'b11001:
        casez_tmp_240 = rob_unsafe_3_25;
      5'b11010:
        casez_tmp_240 = rob_unsafe_3_26;
      5'b11011:
        casez_tmp_240 = rob_unsafe_3_27;
      5'b11100:
        casez_tmp_240 = rob_unsafe_3_28;
      5'b11101:
        casez_tmp_240 = rob_unsafe_3_29;
      5'b11110:
        casez_tmp_240 = rob_unsafe_3_30;
      default:
        casez_tmp_240 = rob_unsafe_3_31;
    endcase
  end // always @(*)
  reg         casez_tmp_241;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_241 = rob_val_3_0;
      5'b00001:
        casez_tmp_241 = rob_val_3_1;
      5'b00010:
        casez_tmp_241 = rob_val_3_2;
      5'b00011:
        casez_tmp_241 = rob_val_3_3;
      5'b00100:
        casez_tmp_241 = rob_val_3_4;
      5'b00101:
        casez_tmp_241 = rob_val_3_5;
      5'b00110:
        casez_tmp_241 = rob_val_3_6;
      5'b00111:
        casez_tmp_241 = rob_val_3_7;
      5'b01000:
        casez_tmp_241 = rob_val_3_8;
      5'b01001:
        casez_tmp_241 = rob_val_3_9;
      5'b01010:
        casez_tmp_241 = rob_val_3_10;
      5'b01011:
        casez_tmp_241 = rob_val_3_11;
      5'b01100:
        casez_tmp_241 = rob_val_3_12;
      5'b01101:
        casez_tmp_241 = rob_val_3_13;
      5'b01110:
        casez_tmp_241 = rob_val_3_14;
      5'b01111:
        casez_tmp_241 = rob_val_3_15;
      5'b10000:
        casez_tmp_241 = rob_val_3_16;
      5'b10001:
        casez_tmp_241 = rob_val_3_17;
      5'b10010:
        casez_tmp_241 = rob_val_3_18;
      5'b10011:
        casez_tmp_241 = rob_val_3_19;
      5'b10100:
        casez_tmp_241 = rob_val_3_20;
      5'b10101:
        casez_tmp_241 = rob_val_3_21;
      5'b10110:
        casez_tmp_241 = rob_val_3_22;
      5'b10111:
        casez_tmp_241 = rob_val_3_23;
      5'b11000:
        casez_tmp_241 = rob_val_3_24;
      5'b11001:
        casez_tmp_241 = rob_val_3_25;
      5'b11010:
        casez_tmp_241 = rob_val_3_26;
      5'b11011:
        casez_tmp_241 = rob_val_3_27;
      5'b11100:
        casez_tmp_241 = rob_val_3_28;
      5'b11101:
        casez_tmp_241 = rob_val_3_29;
      5'b11110:
        casez_tmp_241 = rob_val_3_30;
      default:
        casez_tmp_241 = rob_val_3_31;
    endcase
  end // always @(*)
  reg         casez_tmp_242;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_242 = rob_exception_3_0;
      5'b00001:
        casez_tmp_242 = rob_exception_3_1;
      5'b00010:
        casez_tmp_242 = rob_exception_3_2;
      5'b00011:
        casez_tmp_242 = rob_exception_3_3;
      5'b00100:
        casez_tmp_242 = rob_exception_3_4;
      5'b00101:
        casez_tmp_242 = rob_exception_3_5;
      5'b00110:
        casez_tmp_242 = rob_exception_3_6;
      5'b00111:
        casez_tmp_242 = rob_exception_3_7;
      5'b01000:
        casez_tmp_242 = rob_exception_3_8;
      5'b01001:
        casez_tmp_242 = rob_exception_3_9;
      5'b01010:
        casez_tmp_242 = rob_exception_3_10;
      5'b01011:
        casez_tmp_242 = rob_exception_3_11;
      5'b01100:
        casez_tmp_242 = rob_exception_3_12;
      5'b01101:
        casez_tmp_242 = rob_exception_3_13;
      5'b01110:
        casez_tmp_242 = rob_exception_3_14;
      5'b01111:
        casez_tmp_242 = rob_exception_3_15;
      5'b10000:
        casez_tmp_242 = rob_exception_3_16;
      5'b10001:
        casez_tmp_242 = rob_exception_3_17;
      5'b10010:
        casez_tmp_242 = rob_exception_3_18;
      5'b10011:
        casez_tmp_242 = rob_exception_3_19;
      5'b10100:
        casez_tmp_242 = rob_exception_3_20;
      5'b10101:
        casez_tmp_242 = rob_exception_3_21;
      5'b10110:
        casez_tmp_242 = rob_exception_3_22;
      5'b10111:
        casez_tmp_242 = rob_exception_3_23;
      5'b11000:
        casez_tmp_242 = rob_exception_3_24;
      5'b11001:
        casez_tmp_242 = rob_exception_3_25;
      5'b11010:
        casez_tmp_242 = rob_exception_3_26;
      5'b11011:
        casez_tmp_242 = rob_exception_3_27;
      5'b11100:
        casez_tmp_242 = rob_exception_3_28;
      5'b11101:
        casez_tmp_242 = rob_exception_3_29;
      5'b11110:
        casez_tmp_242 = rob_exception_3_30;
      default:
        casez_tmp_242 = rob_exception_3_31;
    endcase
  end // always @(*)
  wire        can_throw_exception_3 = casez_tmp_241 & casez_tmp_242;
  reg         casez_tmp_243;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_243 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_243 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_243 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_243 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_243 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_243 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_243 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_243 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_243 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_243 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_243 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_243 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_243 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_243 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_243 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_243 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_243 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_243 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_243 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_243 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_243 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_243 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_243 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_243 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_243 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_243 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_243 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_243 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_243 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_243 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_243 = rob_bsy_3_30;
      default:
        casez_tmp_243 = rob_bsy_3_31;
    endcase
  end // always @(*)
  reg         casez_tmp_244;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_244 = rob_predicated_3_0;
      5'b00001:
        casez_tmp_244 = rob_predicated_3_1;
      5'b00010:
        casez_tmp_244 = rob_predicated_3_2;
      5'b00011:
        casez_tmp_244 = rob_predicated_3_3;
      5'b00100:
        casez_tmp_244 = rob_predicated_3_4;
      5'b00101:
        casez_tmp_244 = rob_predicated_3_5;
      5'b00110:
        casez_tmp_244 = rob_predicated_3_6;
      5'b00111:
        casez_tmp_244 = rob_predicated_3_7;
      5'b01000:
        casez_tmp_244 = rob_predicated_3_8;
      5'b01001:
        casez_tmp_244 = rob_predicated_3_9;
      5'b01010:
        casez_tmp_244 = rob_predicated_3_10;
      5'b01011:
        casez_tmp_244 = rob_predicated_3_11;
      5'b01100:
        casez_tmp_244 = rob_predicated_3_12;
      5'b01101:
        casez_tmp_244 = rob_predicated_3_13;
      5'b01110:
        casez_tmp_244 = rob_predicated_3_14;
      5'b01111:
        casez_tmp_244 = rob_predicated_3_15;
      5'b10000:
        casez_tmp_244 = rob_predicated_3_16;
      5'b10001:
        casez_tmp_244 = rob_predicated_3_17;
      5'b10010:
        casez_tmp_244 = rob_predicated_3_18;
      5'b10011:
        casez_tmp_244 = rob_predicated_3_19;
      5'b10100:
        casez_tmp_244 = rob_predicated_3_20;
      5'b10101:
        casez_tmp_244 = rob_predicated_3_21;
      5'b10110:
        casez_tmp_244 = rob_predicated_3_22;
      5'b10111:
        casez_tmp_244 = rob_predicated_3_23;
      5'b11000:
        casez_tmp_244 = rob_predicated_3_24;
      5'b11001:
        casez_tmp_244 = rob_predicated_3_25;
      5'b11010:
        casez_tmp_244 = rob_predicated_3_26;
      5'b11011:
        casez_tmp_244 = rob_predicated_3_27;
      5'b11100:
        casez_tmp_244 = rob_predicated_3_28;
      5'b11101:
        casez_tmp_244 = rob_predicated_3_29;
      5'b11110:
        casez_tmp_244 = rob_predicated_3_30;
      default:
        casez_tmp_244 = rob_predicated_3_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_245;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_245 = rob_uop_3_0_uopc;
      5'b00001:
        casez_tmp_245 = rob_uop_3_1_uopc;
      5'b00010:
        casez_tmp_245 = rob_uop_3_2_uopc;
      5'b00011:
        casez_tmp_245 = rob_uop_3_3_uopc;
      5'b00100:
        casez_tmp_245 = rob_uop_3_4_uopc;
      5'b00101:
        casez_tmp_245 = rob_uop_3_5_uopc;
      5'b00110:
        casez_tmp_245 = rob_uop_3_6_uopc;
      5'b00111:
        casez_tmp_245 = rob_uop_3_7_uopc;
      5'b01000:
        casez_tmp_245 = rob_uop_3_8_uopc;
      5'b01001:
        casez_tmp_245 = rob_uop_3_9_uopc;
      5'b01010:
        casez_tmp_245 = rob_uop_3_10_uopc;
      5'b01011:
        casez_tmp_245 = rob_uop_3_11_uopc;
      5'b01100:
        casez_tmp_245 = rob_uop_3_12_uopc;
      5'b01101:
        casez_tmp_245 = rob_uop_3_13_uopc;
      5'b01110:
        casez_tmp_245 = rob_uop_3_14_uopc;
      5'b01111:
        casez_tmp_245 = rob_uop_3_15_uopc;
      5'b10000:
        casez_tmp_245 = rob_uop_3_16_uopc;
      5'b10001:
        casez_tmp_245 = rob_uop_3_17_uopc;
      5'b10010:
        casez_tmp_245 = rob_uop_3_18_uopc;
      5'b10011:
        casez_tmp_245 = rob_uop_3_19_uopc;
      5'b10100:
        casez_tmp_245 = rob_uop_3_20_uopc;
      5'b10101:
        casez_tmp_245 = rob_uop_3_21_uopc;
      5'b10110:
        casez_tmp_245 = rob_uop_3_22_uopc;
      5'b10111:
        casez_tmp_245 = rob_uop_3_23_uopc;
      5'b11000:
        casez_tmp_245 = rob_uop_3_24_uopc;
      5'b11001:
        casez_tmp_245 = rob_uop_3_25_uopc;
      5'b11010:
        casez_tmp_245 = rob_uop_3_26_uopc;
      5'b11011:
        casez_tmp_245 = rob_uop_3_27_uopc;
      5'b11100:
        casez_tmp_245 = rob_uop_3_28_uopc;
      5'b11101:
        casez_tmp_245 = rob_uop_3_29_uopc;
      5'b11110:
        casez_tmp_245 = rob_uop_3_30_uopc;
      default:
        casez_tmp_245 = rob_uop_3_31_uopc;
    endcase
  end // always @(*)
  reg         casez_tmp_246;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_246 = rob_uop_3_0_is_rvc;
      5'b00001:
        casez_tmp_246 = rob_uop_3_1_is_rvc;
      5'b00010:
        casez_tmp_246 = rob_uop_3_2_is_rvc;
      5'b00011:
        casez_tmp_246 = rob_uop_3_3_is_rvc;
      5'b00100:
        casez_tmp_246 = rob_uop_3_4_is_rvc;
      5'b00101:
        casez_tmp_246 = rob_uop_3_5_is_rvc;
      5'b00110:
        casez_tmp_246 = rob_uop_3_6_is_rvc;
      5'b00111:
        casez_tmp_246 = rob_uop_3_7_is_rvc;
      5'b01000:
        casez_tmp_246 = rob_uop_3_8_is_rvc;
      5'b01001:
        casez_tmp_246 = rob_uop_3_9_is_rvc;
      5'b01010:
        casez_tmp_246 = rob_uop_3_10_is_rvc;
      5'b01011:
        casez_tmp_246 = rob_uop_3_11_is_rvc;
      5'b01100:
        casez_tmp_246 = rob_uop_3_12_is_rvc;
      5'b01101:
        casez_tmp_246 = rob_uop_3_13_is_rvc;
      5'b01110:
        casez_tmp_246 = rob_uop_3_14_is_rvc;
      5'b01111:
        casez_tmp_246 = rob_uop_3_15_is_rvc;
      5'b10000:
        casez_tmp_246 = rob_uop_3_16_is_rvc;
      5'b10001:
        casez_tmp_246 = rob_uop_3_17_is_rvc;
      5'b10010:
        casez_tmp_246 = rob_uop_3_18_is_rvc;
      5'b10011:
        casez_tmp_246 = rob_uop_3_19_is_rvc;
      5'b10100:
        casez_tmp_246 = rob_uop_3_20_is_rvc;
      5'b10101:
        casez_tmp_246 = rob_uop_3_21_is_rvc;
      5'b10110:
        casez_tmp_246 = rob_uop_3_22_is_rvc;
      5'b10111:
        casez_tmp_246 = rob_uop_3_23_is_rvc;
      5'b11000:
        casez_tmp_246 = rob_uop_3_24_is_rvc;
      5'b11001:
        casez_tmp_246 = rob_uop_3_25_is_rvc;
      5'b11010:
        casez_tmp_246 = rob_uop_3_26_is_rvc;
      5'b11011:
        casez_tmp_246 = rob_uop_3_27_is_rvc;
      5'b11100:
        casez_tmp_246 = rob_uop_3_28_is_rvc;
      5'b11101:
        casez_tmp_246 = rob_uop_3_29_is_rvc;
      5'b11110:
        casez_tmp_246 = rob_uop_3_30_is_rvc;
      default:
        casez_tmp_246 = rob_uop_3_31_is_rvc;
    endcase
  end // always @(*)
  reg         casez_tmp_247;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_247 = rob_uop_3_0_is_br;
      5'b00001:
        casez_tmp_247 = rob_uop_3_1_is_br;
      5'b00010:
        casez_tmp_247 = rob_uop_3_2_is_br;
      5'b00011:
        casez_tmp_247 = rob_uop_3_3_is_br;
      5'b00100:
        casez_tmp_247 = rob_uop_3_4_is_br;
      5'b00101:
        casez_tmp_247 = rob_uop_3_5_is_br;
      5'b00110:
        casez_tmp_247 = rob_uop_3_6_is_br;
      5'b00111:
        casez_tmp_247 = rob_uop_3_7_is_br;
      5'b01000:
        casez_tmp_247 = rob_uop_3_8_is_br;
      5'b01001:
        casez_tmp_247 = rob_uop_3_9_is_br;
      5'b01010:
        casez_tmp_247 = rob_uop_3_10_is_br;
      5'b01011:
        casez_tmp_247 = rob_uop_3_11_is_br;
      5'b01100:
        casez_tmp_247 = rob_uop_3_12_is_br;
      5'b01101:
        casez_tmp_247 = rob_uop_3_13_is_br;
      5'b01110:
        casez_tmp_247 = rob_uop_3_14_is_br;
      5'b01111:
        casez_tmp_247 = rob_uop_3_15_is_br;
      5'b10000:
        casez_tmp_247 = rob_uop_3_16_is_br;
      5'b10001:
        casez_tmp_247 = rob_uop_3_17_is_br;
      5'b10010:
        casez_tmp_247 = rob_uop_3_18_is_br;
      5'b10011:
        casez_tmp_247 = rob_uop_3_19_is_br;
      5'b10100:
        casez_tmp_247 = rob_uop_3_20_is_br;
      5'b10101:
        casez_tmp_247 = rob_uop_3_21_is_br;
      5'b10110:
        casez_tmp_247 = rob_uop_3_22_is_br;
      5'b10111:
        casez_tmp_247 = rob_uop_3_23_is_br;
      5'b11000:
        casez_tmp_247 = rob_uop_3_24_is_br;
      5'b11001:
        casez_tmp_247 = rob_uop_3_25_is_br;
      5'b11010:
        casez_tmp_247 = rob_uop_3_26_is_br;
      5'b11011:
        casez_tmp_247 = rob_uop_3_27_is_br;
      5'b11100:
        casez_tmp_247 = rob_uop_3_28_is_br;
      5'b11101:
        casez_tmp_247 = rob_uop_3_29_is_br;
      5'b11110:
        casez_tmp_247 = rob_uop_3_30_is_br;
      default:
        casez_tmp_247 = rob_uop_3_31_is_br;
    endcase
  end // always @(*)
  reg         casez_tmp_248;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_248 = rob_uop_3_0_is_jalr;
      5'b00001:
        casez_tmp_248 = rob_uop_3_1_is_jalr;
      5'b00010:
        casez_tmp_248 = rob_uop_3_2_is_jalr;
      5'b00011:
        casez_tmp_248 = rob_uop_3_3_is_jalr;
      5'b00100:
        casez_tmp_248 = rob_uop_3_4_is_jalr;
      5'b00101:
        casez_tmp_248 = rob_uop_3_5_is_jalr;
      5'b00110:
        casez_tmp_248 = rob_uop_3_6_is_jalr;
      5'b00111:
        casez_tmp_248 = rob_uop_3_7_is_jalr;
      5'b01000:
        casez_tmp_248 = rob_uop_3_8_is_jalr;
      5'b01001:
        casez_tmp_248 = rob_uop_3_9_is_jalr;
      5'b01010:
        casez_tmp_248 = rob_uop_3_10_is_jalr;
      5'b01011:
        casez_tmp_248 = rob_uop_3_11_is_jalr;
      5'b01100:
        casez_tmp_248 = rob_uop_3_12_is_jalr;
      5'b01101:
        casez_tmp_248 = rob_uop_3_13_is_jalr;
      5'b01110:
        casez_tmp_248 = rob_uop_3_14_is_jalr;
      5'b01111:
        casez_tmp_248 = rob_uop_3_15_is_jalr;
      5'b10000:
        casez_tmp_248 = rob_uop_3_16_is_jalr;
      5'b10001:
        casez_tmp_248 = rob_uop_3_17_is_jalr;
      5'b10010:
        casez_tmp_248 = rob_uop_3_18_is_jalr;
      5'b10011:
        casez_tmp_248 = rob_uop_3_19_is_jalr;
      5'b10100:
        casez_tmp_248 = rob_uop_3_20_is_jalr;
      5'b10101:
        casez_tmp_248 = rob_uop_3_21_is_jalr;
      5'b10110:
        casez_tmp_248 = rob_uop_3_22_is_jalr;
      5'b10111:
        casez_tmp_248 = rob_uop_3_23_is_jalr;
      5'b11000:
        casez_tmp_248 = rob_uop_3_24_is_jalr;
      5'b11001:
        casez_tmp_248 = rob_uop_3_25_is_jalr;
      5'b11010:
        casez_tmp_248 = rob_uop_3_26_is_jalr;
      5'b11011:
        casez_tmp_248 = rob_uop_3_27_is_jalr;
      5'b11100:
        casez_tmp_248 = rob_uop_3_28_is_jalr;
      5'b11101:
        casez_tmp_248 = rob_uop_3_29_is_jalr;
      5'b11110:
        casez_tmp_248 = rob_uop_3_30_is_jalr;
      default:
        casez_tmp_248 = rob_uop_3_31_is_jalr;
    endcase
  end // always @(*)
  reg         casez_tmp_249;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_249 = rob_uop_3_0_is_jal;
      5'b00001:
        casez_tmp_249 = rob_uop_3_1_is_jal;
      5'b00010:
        casez_tmp_249 = rob_uop_3_2_is_jal;
      5'b00011:
        casez_tmp_249 = rob_uop_3_3_is_jal;
      5'b00100:
        casez_tmp_249 = rob_uop_3_4_is_jal;
      5'b00101:
        casez_tmp_249 = rob_uop_3_5_is_jal;
      5'b00110:
        casez_tmp_249 = rob_uop_3_6_is_jal;
      5'b00111:
        casez_tmp_249 = rob_uop_3_7_is_jal;
      5'b01000:
        casez_tmp_249 = rob_uop_3_8_is_jal;
      5'b01001:
        casez_tmp_249 = rob_uop_3_9_is_jal;
      5'b01010:
        casez_tmp_249 = rob_uop_3_10_is_jal;
      5'b01011:
        casez_tmp_249 = rob_uop_3_11_is_jal;
      5'b01100:
        casez_tmp_249 = rob_uop_3_12_is_jal;
      5'b01101:
        casez_tmp_249 = rob_uop_3_13_is_jal;
      5'b01110:
        casez_tmp_249 = rob_uop_3_14_is_jal;
      5'b01111:
        casez_tmp_249 = rob_uop_3_15_is_jal;
      5'b10000:
        casez_tmp_249 = rob_uop_3_16_is_jal;
      5'b10001:
        casez_tmp_249 = rob_uop_3_17_is_jal;
      5'b10010:
        casez_tmp_249 = rob_uop_3_18_is_jal;
      5'b10011:
        casez_tmp_249 = rob_uop_3_19_is_jal;
      5'b10100:
        casez_tmp_249 = rob_uop_3_20_is_jal;
      5'b10101:
        casez_tmp_249 = rob_uop_3_21_is_jal;
      5'b10110:
        casez_tmp_249 = rob_uop_3_22_is_jal;
      5'b10111:
        casez_tmp_249 = rob_uop_3_23_is_jal;
      5'b11000:
        casez_tmp_249 = rob_uop_3_24_is_jal;
      5'b11001:
        casez_tmp_249 = rob_uop_3_25_is_jal;
      5'b11010:
        casez_tmp_249 = rob_uop_3_26_is_jal;
      5'b11011:
        casez_tmp_249 = rob_uop_3_27_is_jal;
      5'b11100:
        casez_tmp_249 = rob_uop_3_28_is_jal;
      5'b11101:
        casez_tmp_249 = rob_uop_3_29_is_jal;
      5'b11110:
        casez_tmp_249 = rob_uop_3_30_is_jal;
      default:
        casez_tmp_249 = rob_uop_3_31_is_jal;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_250;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_250 = rob_uop_3_0_ftq_idx;
      5'b00001:
        casez_tmp_250 = rob_uop_3_1_ftq_idx;
      5'b00010:
        casez_tmp_250 = rob_uop_3_2_ftq_idx;
      5'b00011:
        casez_tmp_250 = rob_uop_3_3_ftq_idx;
      5'b00100:
        casez_tmp_250 = rob_uop_3_4_ftq_idx;
      5'b00101:
        casez_tmp_250 = rob_uop_3_5_ftq_idx;
      5'b00110:
        casez_tmp_250 = rob_uop_3_6_ftq_idx;
      5'b00111:
        casez_tmp_250 = rob_uop_3_7_ftq_idx;
      5'b01000:
        casez_tmp_250 = rob_uop_3_8_ftq_idx;
      5'b01001:
        casez_tmp_250 = rob_uop_3_9_ftq_idx;
      5'b01010:
        casez_tmp_250 = rob_uop_3_10_ftq_idx;
      5'b01011:
        casez_tmp_250 = rob_uop_3_11_ftq_idx;
      5'b01100:
        casez_tmp_250 = rob_uop_3_12_ftq_idx;
      5'b01101:
        casez_tmp_250 = rob_uop_3_13_ftq_idx;
      5'b01110:
        casez_tmp_250 = rob_uop_3_14_ftq_idx;
      5'b01111:
        casez_tmp_250 = rob_uop_3_15_ftq_idx;
      5'b10000:
        casez_tmp_250 = rob_uop_3_16_ftq_idx;
      5'b10001:
        casez_tmp_250 = rob_uop_3_17_ftq_idx;
      5'b10010:
        casez_tmp_250 = rob_uop_3_18_ftq_idx;
      5'b10011:
        casez_tmp_250 = rob_uop_3_19_ftq_idx;
      5'b10100:
        casez_tmp_250 = rob_uop_3_20_ftq_idx;
      5'b10101:
        casez_tmp_250 = rob_uop_3_21_ftq_idx;
      5'b10110:
        casez_tmp_250 = rob_uop_3_22_ftq_idx;
      5'b10111:
        casez_tmp_250 = rob_uop_3_23_ftq_idx;
      5'b11000:
        casez_tmp_250 = rob_uop_3_24_ftq_idx;
      5'b11001:
        casez_tmp_250 = rob_uop_3_25_ftq_idx;
      5'b11010:
        casez_tmp_250 = rob_uop_3_26_ftq_idx;
      5'b11011:
        casez_tmp_250 = rob_uop_3_27_ftq_idx;
      5'b11100:
        casez_tmp_250 = rob_uop_3_28_ftq_idx;
      5'b11101:
        casez_tmp_250 = rob_uop_3_29_ftq_idx;
      5'b11110:
        casez_tmp_250 = rob_uop_3_30_ftq_idx;
      default:
        casez_tmp_250 = rob_uop_3_31_ftq_idx;
    endcase
  end // always @(*)
  reg         casez_tmp_251;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_251 = rob_uop_3_0_edge_inst;
      5'b00001:
        casez_tmp_251 = rob_uop_3_1_edge_inst;
      5'b00010:
        casez_tmp_251 = rob_uop_3_2_edge_inst;
      5'b00011:
        casez_tmp_251 = rob_uop_3_3_edge_inst;
      5'b00100:
        casez_tmp_251 = rob_uop_3_4_edge_inst;
      5'b00101:
        casez_tmp_251 = rob_uop_3_5_edge_inst;
      5'b00110:
        casez_tmp_251 = rob_uop_3_6_edge_inst;
      5'b00111:
        casez_tmp_251 = rob_uop_3_7_edge_inst;
      5'b01000:
        casez_tmp_251 = rob_uop_3_8_edge_inst;
      5'b01001:
        casez_tmp_251 = rob_uop_3_9_edge_inst;
      5'b01010:
        casez_tmp_251 = rob_uop_3_10_edge_inst;
      5'b01011:
        casez_tmp_251 = rob_uop_3_11_edge_inst;
      5'b01100:
        casez_tmp_251 = rob_uop_3_12_edge_inst;
      5'b01101:
        casez_tmp_251 = rob_uop_3_13_edge_inst;
      5'b01110:
        casez_tmp_251 = rob_uop_3_14_edge_inst;
      5'b01111:
        casez_tmp_251 = rob_uop_3_15_edge_inst;
      5'b10000:
        casez_tmp_251 = rob_uop_3_16_edge_inst;
      5'b10001:
        casez_tmp_251 = rob_uop_3_17_edge_inst;
      5'b10010:
        casez_tmp_251 = rob_uop_3_18_edge_inst;
      5'b10011:
        casez_tmp_251 = rob_uop_3_19_edge_inst;
      5'b10100:
        casez_tmp_251 = rob_uop_3_20_edge_inst;
      5'b10101:
        casez_tmp_251 = rob_uop_3_21_edge_inst;
      5'b10110:
        casez_tmp_251 = rob_uop_3_22_edge_inst;
      5'b10111:
        casez_tmp_251 = rob_uop_3_23_edge_inst;
      5'b11000:
        casez_tmp_251 = rob_uop_3_24_edge_inst;
      5'b11001:
        casez_tmp_251 = rob_uop_3_25_edge_inst;
      5'b11010:
        casez_tmp_251 = rob_uop_3_26_edge_inst;
      5'b11011:
        casez_tmp_251 = rob_uop_3_27_edge_inst;
      5'b11100:
        casez_tmp_251 = rob_uop_3_28_edge_inst;
      5'b11101:
        casez_tmp_251 = rob_uop_3_29_edge_inst;
      5'b11110:
        casez_tmp_251 = rob_uop_3_30_edge_inst;
      default:
        casez_tmp_251 = rob_uop_3_31_edge_inst;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_252;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_252 = rob_uop_3_0_pc_lob;
      5'b00001:
        casez_tmp_252 = rob_uop_3_1_pc_lob;
      5'b00010:
        casez_tmp_252 = rob_uop_3_2_pc_lob;
      5'b00011:
        casez_tmp_252 = rob_uop_3_3_pc_lob;
      5'b00100:
        casez_tmp_252 = rob_uop_3_4_pc_lob;
      5'b00101:
        casez_tmp_252 = rob_uop_3_5_pc_lob;
      5'b00110:
        casez_tmp_252 = rob_uop_3_6_pc_lob;
      5'b00111:
        casez_tmp_252 = rob_uop_3_7_pc_lob;
      5'b01000:
        casez_tmp_252 = rob_uop_3_8_pc_lob;
      5'b01001:
        casez_tmp_252 = rob_uop_3_9_pc_lob;
      5'b01010:
        casez_tmp_252 = rob_uop_3_10_pc_lob;
      5'b01011:
        casez_tmp_252 = rob_uop_3_11_pc_lob;
      5'b01100:
        casez_tmp_252 = rob_uop_3_12_pc_lob;
      5'b01101:
        casez_tmp_252 = rob_uop_3_13_pc_lob;
      5'b01110:
        casez_tmp_252 = rob_uop_3_14_pc_lob;
      5'b01111:
        casez_tmp_252 = rob_uop_3_15_pc_lob;
      5'b10000:
        casez_tmp_252 = rob_uop_3_16_pc_lob;
      5'b10001:
        casez_tmp_252 = rob_uop_3_17_pc_lob;
      5'b10010:
        casez_tmp_252 = rob_uop_3_18_pc_lob;
      5'b10011:
        casez_tmp_252 = rob_uop_3_19_pc_lob;
      5'b10100:
        casez_tmp_252 = rob_uop_3_20_pc_lob;
      5'b10101:
        casez_tmp_252 = rob_uop_3_21_pc_lob;
      5'b10110:
        casez_tmp_252 = rob_uop_3_22_pc_lob;
      5'b10111:
        casez_tmp_252 = rob_uop_3_23_pc_lob;
      5'b11000:
        casez_tmp_252 = rob_uop_3_24_pc_lob;
      5'b11001:
        casez_tmp_252 = rob_uop_3_25_pc_lob;
      5'b11010:
        casez_tmp_252 = rob_uop_3_26_pc_lob;
      5'b11011:
        casez_tmp_252 = rob_uop_3_27_pc_lob;
      5'b11100:
        casez_tmp_252 = rob_uop_3_28_pc_lob;
      5'b11101:
        casez_tmp_252 = rob_uop_3_29_pc_lob;
      5'b11110:
        casez_tmp_252 = rob_uop_3_30_pc_lob;
      default:
        casez_tmp_252 = rob_uop_3_31_pc_lob;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_253;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_253 = rob_uop_3_0_pdst;
      5'b00001:
        casez_tmp_253 = rob_uop_3_1_pdst;
      5'b00010:
        casez_tmp_253 = rob_uop_3_2_pdst;
      5'b00011:
        casez_tmp_253 = rob_uop_3_3_pdst;
      5'b00100:
        casez_tmp_253 = rob_uop_3_4_pdst;
      5'b00101:
        casez_tmp_253 = rob_uop_3_5_pdst;
      5'b00110:
        casez_tmp_253 = rob_uop_3_6_pdst;
      5'b00111:
        casez_tmp_253 = rob_uop_3_7_pdst;
      5'b01000:
        casez_tmp_253 = rob_uop_3_8_pdst;
      5'b01001:
        casez_tmp_253 = rob_uop_3_9_pdst;
      5'b01010:
        casez_tmp_253 = rob_uop_3_10_pdst;
      5'b01011:
        casez_tmp_253 = rob_uop_3_11_pdst;
      5'b01100:
        casez_tmp_253 = rob_uop_3_12_pdst;
      5'b01101:
        casez_tmp_253 = rob_uop_3_13_pdst;
      5'b01110:
        casez_tmp_253 = rob_uop_3_14_pdst;
      5'b01111:
        casez_tmp_253 = rob_uop_3_15_pdst;
      5'b10000:
        casez_tmp_253 = rob_uop_3_16_pdst;
      5'b10001:
        casez_tmp_253 = rob_uop_3_17_pdst;
      5'b10010:
        casez_tmp_253 = rob_uop_3_18_pdst;
      5'b10011:
        casez_tmp_253 = rob_uop_3_19_pdst;
      5'b10100:
        casez_tmp_253 = rob_uop_3_20_pdst;
      5'b10101:
        casez_tmp_253 = rob_uop_3_21_pdst;
      5'b10110:
        casez_tmp_253 = rob_uop_3_22_pdst;
      5'b10111:
        casez_tmp_253 = rob_uop_3_23_pdst;
      5'b11000:
        casez_tmp_253 = rob_uop_3_24_pdst;
      5'b11001:
        casez_tmp_253 = rob_uop_3_25_pdst;
      5'b11010:
        casez_tmp_253 = rob_uop_3_26_pdst;
      5'b11011:
        casez_tmp_253 = rob_uop_3_27_pdst;
      5'b11100:
        casez_tmp_253 = rob_uop_3_28_pdst;
      5'b11101:
        casez_tmp_253 = rob_uop_3_29_pdst;
      5'b11110:
        casez_tmp_253 = rob_uop_3_30_pdst;
      default:
        casez_tmp_253 = rob_uop_3_31_pdst;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_254;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_254 = rob_uop_3_0_stale_pdst;
      5'b00001:
        casez_tmp_254 = rob_uop_3_1_stale_pdst;
      5'b00010:
        casez_tmp_254 = rob_uop_3_2_stale_pdst;
      5'b00011:
        casez_tmp_254 = rob_uop_3_3_stale_pdst;
      5'b00100:
        casez_tmp_254 = rob_uop_3_4_stale_pdst;
      5'b00101:
        casez_tmp_254 = rob_uop_3_5_stale_pdst;
      5'b00110:
        casez_tmp_254 = rob_uop_3_6_stale_pdst;
      5'b00111:
        casez_tmp_254 = rob_uop_3_7_stale_pdst;
      5'b01000:
        casez_tmp_254 = rob_uop_3_8_stale_pdst;
      5'b01001:
        casez_tmp_254 = rob_uop_3_9_stale_pdst;
      5'b01010:
        casez_tmp_254 = rob_uop_3_10_stale_pdst;
      5'b01011:
        casez_tmp_254 = rob_uop_3_11_stale_pdst;
      5'b01100:
        casez_tmp_254 = rob_uop_3_12_stale_pdst;
      5'b01101:
        casez_tmp_254 = rob_uop_3_13_stale_pdst;
      5'b01110:
        casez_tmp_254 = rob_uop_3_14_stale_pdst;
      5'b01111:
        casez_tmp_254 = rob_uop_3_15_stale_pdst;
      5'b10000:
        casez_tmp_254 = rob_uop_3_16_stale_pdst;
      5'b10001:
        casez_tmp_254 = rob_uop_3_17_stale_pdst;
      5'b10010:
        casez_tmp_254 = rob_uop_3_18_stale_pdst;
      5'b10011:
        casez_tmp_254 = rob_uop_3_19_stale_pdst;
      5'b10100:
        casez_tmp_254 = rob_uop_3_20_stale_pdst;
      5'b10101:
        casez_tmp_254 = rob_uop_3_21_stale_pdst;
      5'b10110:
        casez_tmp_254 = rob_uop_3_22_stale_pdst;
      5'b10111:
        casez_tmp_254 = rob_uop_3_23_stale_pdst;
      5'b11000:
        casez_tmp_254 = rob_uop_3_24_stale_pdst;
      5'b11001:
        casez_tmp_254 = rob_uop_3_25_stale_pdst;
      5'b11010:
        casez_tmp_254 = rob_uop_3_26_stale_pdst;
      5'b11011:
        casez_tmp_254 = rob_uop_3_27_stale_pdst;
      5'b11100:
        casez_tmp_254 = rob_uop_3_28_stale_pdst;
      5'b11101:
        casez_tmp_254 = rob_uop_3_29_stale_pdst;
      5'b11110:
        casez_tmp_254 = rob_uop_3_30_stale_pdst;
      default:
        casez_tmp_254 = rob_uop_3_31_stale_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_255;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_255 = rob_uop_3_0_is_fencei;
      5'b00001:
        casez_tmp_255 = rob_uop_3_1_is_fencei;
      5'b00010:
        casez_tmp_255 = rob_uop_3_2_is_fencei;
      5'b00011:
        casez_tmp_255 = rob_uop_3_3_is_fencei;
      5'b00100:
        casez_tmp_255 = rob_uop_3_4_is_fencei;
      5'b00101:
        casez_tmp_255 = rob_uop_3_5_is_fencei;
      5'b00110:
        casez_tmp_255 = rob_uop_3_6_is_fencei;
      5'b00111:
        casez_tmp_255 = rob_uop_3_7_is_fencei;
      5'b01000:
        casez_tmp_255 = rob_uop_3_8_is_fencei;
      5'b01001:
        casez_tmp_255 = rob_uop_3_9_is_fencei;
      5'b01010:
        casez_tmp_255 = rob_uop_3_10_is_fencei;
      5'b01011:
        casez_tmp_255 = rob_uop_3_11_is_fencei;
      5'b01100:
        casez_tmp_255 = rob_uop_3_12_is_fencei;
      5'b01101:
        casez_tmp_255 = rob_uop_3_13_is_fencei;
      5'b01110:
        casez_tmp_255 = rob_uop_3_14_is_fencei;
      5'b01111:
        casez_tmp_255 = rob_uop_3_15_is_fencei;
      5'b10000:
        casez_tmp_255 = rob_uop_3_16_is_fencei;
      5'b10001:
        casez_tmp_255 = rob_uop_3_17_is_fencei;
      5'b10010:
        casez_tmp_255 = rob_uop_3_18_is_fencei;
      5'b10011:
        casez_tmp_255 = rob_uop_3_19_is_fencei;
      5'b10100:
        casez_tmp_255 = rob_uop_3_20_is_fencei;
      5'b10101:
        casez_tmp_255 = rob_uop_3_21_is_fencei;
      5'b10110:
        casez_tmp_255 = rob_uop_3_22_is_fencei;
      5'b10111:
        casez_tmp_255 = rob_uop_3_23_is_fencei;
      5'b11000:
        casez_tmp_255 = rob_uop_3_24_is_fencei;
      5'b11001:
        casez_tmp_255 = rob_uop_3_25_is_fencei;
      5'b11010:
        casez_tmp_255 = rob_uop_3_26_is_fencei;
      5'b11011:
        casez_tmp_255 = rob_uop_3_27_is_fencei;
      5'b11100:
        casez_tmp_255 = rob_uop_3_28_is_fencei;
      5'b11101:
        casez_tmp_255 = rob_uop_3_29_is_fencei;
      5'b11110:
        casez_tmp_255 = rob_uop_3_30_is_fencei;
      default:
        casez_tmp_255 = rob_uop_3_31_is_fencei;
    endcase
  end // always @(*)
  reg         casez_tmp_256;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_256 = rob_uop_3_0_uses_ldq;
      5'b00001:
        casez_tmp_256 = rob_uop_3_1_uses_ldq;
      5'b00010:
        casez_tmp_256 = rob_uop_3_2_uses_ldq;
      5'b00011:
        casez_tmp_256 = rob_uop_3_3_uses_ldq;
      5'b00100:
        casez_tmp_256 = rob_uop_3_4_uses_ldq;
      5'b00101:
        casez_tmp_256 = rob_uop_3_5_uses_ldq;
      5'b00110:
        casez_tmp_256 = rob_uop_3_6_uses_ldq;
      5'b00111:
        casez_tmp_256 = rob_uop_3_7_uses_ldq;
      5'b01000:
        casez_tmp_256 = rob_uop_3_8_uses_ldq;
      5'b01001:
        casez_tmp_256 = rob_uop_3_9_uses_ldq;
      5'b01010:
        casez_tmp_256 = rob_uop_3_10_uses_ldq;
      5'b01011:
        casez_tmp_256 = rob_uop_3_11_uses_ldq;
      5'b01100:
        casez_tmp_256 = rob_uop_3_12_uses_ldq;
      5'b01101:
        casez_tmp_256 = rob_uop_3_13_uses_ldq;
      5'b01110:
        casez_tmp_256 = rob_uop_3_14_uses_ldq;
      5'b01111:
        casez_tmp_256 = rob_uop_3_15_uses_ldq;
      5'b10000:
        casez_tmp_256 = rob_uop_3_16_uses_ldq;
      5'b10001:
        casez_tmp_256 = rob_uop_3_17_uses_ldq;
      5'b10010:
        casez_tmp_256 = rob_uop_3_18_uses_ldq;
      5'b10011:
        casez_tmp_256 = rob_uop_3_19_uses_ldq;
      5'b10100:
        casez_tmp_256 = rob_uop_3_20_uses_ldq;
      5'b10101:
        casez_tmp_256 = rob_uop_3_21_uses_ldq;
      5'b10110:
        casez_tmp_256 = rob_uop_3_22_uses_ldq;
      5'b10111:
        casez_tmp_256 = rob_uop_3_23_uses_ldq;
      5'b11000:
        casez_tmp_256 = rob_uop_3_24_uses_ldq;
      5'b11001:
        casez_tmp_256 = rob_uop_3_25_uses_ldq;
      5'b11010:
        casez_tmp_256 = rob_uop_3_26_uses_ldq;
      5'b11011:
        casez_tmp_256 = rob_uop_3_27_uses_ldq;
      5'b11100:
        casez_tmp_256 = rob_uop_3_28_uses_ldq;
      5'b11101:
        casez_tmp_256 = rob_uop_3_29_uses_ldq;
      5'b11110:
        casez_tmp_256 = rob_uop_3_30_uses_ldq;
      default:
        casez_tmp_256 = rob_uop_3_31_uses_ldq;
    endcase
  end // always @(*)
  reg         casez_tmp_257;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_257 = rob_uop_3_0_uses_stq;
      5'b00001:
        casez_tmp_257 = rob_uop_3_1_uses_stq;
      5'b00010:
        casez_tmp_257 = rob_uop_3_2_uses_stq;
      5'b00011:
        casez_tmp_257 = rob_uop_3_3_uses_stq;
      5'b00100:
        casez_tmp_257 = rob_uop_3_4_uses_stq;
      5'b00101:
        casez_tmp_257 = rob_uop_3_5_uses_stq;
      5'b00110:
        casez_tmp_257 = rob_uop_3_6_uses_stq;
      5'b00111:
        casez_tmp_257 = rob_uop_3_7_uses_stq;
      5'b01000:
        casez_tmp_257 = rob_uop_3_8_uses_stq;
      5'b01001:
        casez_tmp_257 = rob_uop_3_9_uses_stq;
      5'b01010:
        casez_tmp_257 = rob_uop_3_10_uses_stq;
      5'b01011:
        casez_tmp_257 = rob_uop_3_11_uses_stq;
      5'b01100:
        casez_tmp_257 = rob_uop_3_12_uses_stq;
      5'b01101:
        casez_tmp_257 = rob_uop_3_13_uses_stq;
      5'b01110:
        casez_tmp_257 = rob_uop_3_14_uses_stq;
      5'b01111:
        casez_tmp_257 = rob_uop_3_15_uses_stq;
      5'b10000:
        casez_tmp_257 = rob_uop_3_16_uses_stq;
      5'b10001:
        casez_tmp_257 = rob_uop_3_17_uses_stq;
      5'b10010:
        casez_tmp_257 = rob_uop_3_18_uses_stq;
      5'b10011:
        casez_tmp_257 = rob_uop_3_19_uses_stq;
      5'b10100:
        casez_tmp_257 = rob_uop_3_20_uses_stq;
      5'b10101:
        casez_tmp_257 = rob_uop_3_21_uses_stq;
      5'b10110:
        casez_tmp_257 = rob_uop_3_22_uses_stq;
      5'b10111:
        casez_tmp_257 = rob_uop_3_23_uses_stq;
      5'b11000:
        casez_tmp_257 = rob_uop_3_24_uses_stq;
      5'b11001:
        casez_tmp_257 = rob_uop_3_25_uses_stq;
      5'b11010:
        casez_tmp_257 = rob_uop_3_26_uses_stq;
      5'b11011:
        casez_tmp_257 = rob_uop_3_27_uses_stq;
      5'b11100:
        casez_tmp_257 = rob_uop_3_28_uses_stq;
      5'b11101:
        casez_tmp_257 = rob_uop_3_29_uses_stq;
      5'b11110:
        casez_tmp_257 = rob_uop_3_30_uses_stq;
      default:
        casez_tmp_257 = rob_uop_3_31_uses_stq;
    endcase
  end // always @(*)
  reg         casez_tmp_258;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_258 = rob_uop_3_0_is_sys_pc2epc;
      5'b00001:
        casez_tmp_258 = rob_uop_3_1_is_sys_pc2epc;
      5'b00010:
        casez_tmp_258 = rob_uop_3_2_is_sys_pc2epc;
      5'b00011:
        casez_tmp_258 = rob_uop_3_3_is_sys_pc2epc;
      5'b00100:
        casez_tmp_258 = rob_uop_3_4_is_sys_pc2epc;
      5'b00101:
        casez_tmp_258 = rob_uop_3_5_is_sys_pc2epc;
      5'b00110:
        casez_tmp_258 = rob_uop_3_6_is_sys_pc2epc;
      5'b00111:
        casez_tmp_258 = rob_uop_3_7_is_sys_pc2epc;
      5'b01000:
        casez_tmp_258 = rob_uop_3_8_is_sys_pc2epc;
      5'b01001:
        casez_tmp_258 = rob_uop_3_9_is_sys_pc2epc;
      5'b01010:
        casez_tmp_258 = rob_uop_3_10_is_sys_pc2epc;
      5'b01011:
        casez_tmp_258 = rob_uop_3_11_is_sys_pc2epc;
      5'b01100:
        casez_tmp_258 = rob_uop_3_12_is_sys_pc2epc;
      5'b01101:
        casez_tmp_258 = rob_uop_3_13_is_sys_pc2epc;
      5'b01110:
        casez_tmp_258 = rob_uop_3_14_is_sys_pc2epc;
      5'b01111:
        casez_tmp_258 = rob_uop_3_15_is_sys_pc2epc;
      5'b10000:
        casez_tmp_258 = rob_uop_3_16_is_sys_pc2epc;
      5'b10001:
        casez_tmp_258 = rob_uop_3_17_is_sys_pc2epc;
      5'b10010:
        casez_tmp_258 = rob_uop_3_18_is_sys_pc2epc;
      5'b10011:
        casez_tmp_258 = rob_uop_3_19_is_sys_pc2epc;
      5'b10100:
        casez_tmp_258 = rob_uop_3_20_is_sys_pc2epc;
      5'b10101:
        casez_tmp_258 = rob_uop_3_21_is_sys_pc2epc;
      5'b10110:
        casez_tmp_258 = rob_uop_3_22_is_sys_pc2epc;
      5'b10111:
        casez_tmp_258 = rob_uop_3_23_is_sys_pc2epc;
      5'b11000:
        casez_tmp_258 = rob_uop_3_24_is_sys_pc2epc;
      5'b11001:
        casez_tmp_258 = rob_uop_3_25_is_sys_pc2epc;
      5'b11010:
        casez_tmp_258 = rob_uop_3_26_is_sys_pc2epc;
      5'b11011:
        casez_tmp_258 = rob_uop_3_27_is_sys_pc2epc;
      5'b11100:
        casez_tmp_258 = rob_uop_3_28_is_sys_pc2epc;
      5'b11101:
        casez_tmp_258 = rob_uop_3_29_is_sys_pc2epc;
      5'b11110:
        casez_tmp_258 = rob_uop_3_30_is_sys_pc2epc;
      default:
        casez_tmp_258 = rob_uop_3_31_is_sys_pc2epc;
    endcase
  end // always @(*)
  reg         casez_tmp_259;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_259 = rob_uop_3_0_flush_on_commit;
      5'b00001:
        casez_tmp_259 = rob_uop_3_1_flush_on_commit;
      5'b00010:
        casez_tmp_259 = rob_uop_3_2_flush_on_commit;
      5'b00011:
        casez_tmp_259 = rob_uop_3_3_flush_on_commit;
      5'b00100:
        casez_tmp_259 = rob_uop_3_4_flush_on_commit;
      5'b00101:
        casez_tmp_259 = rob_uop_3_5_flush_on_commit;
      5'b00110:
        casez_tmp_259 = rob_uop_3_6_flush_on_commit;
      5'b00111:
        casez_tmp_259 = rob_uop_3_7_flush_on_commit;
      5'b01000:
        casez_tmp_259 = rob_uop_3_8_flush_on_commit;
      5'b01001:
        casez_tmp_259 = rob_uop_3_9_flush_on_commit;
      5'b01010:
        casez_tmp_259 = rob_uop_3_10_flush_on_commit;
      5'b01011:
        casez_tmp_259 = rob_uop_3_11_flush_on_commit;
      5'b01100:
        casez_tmp_259 = rob_uop_3_12_flush_on_commit;
      5'b01101:
        casez_tmp_259 = rob_uop_3_13_flush_on_commit;
      5'b01110:
        casez_tmp_259 = rob_uop_3_14_flush_on_commit;
      5'b01111:
        casez_tmp_259 = rob_uop_3_15_flush_on_commit;
      5'b10000:
        casez_tmp_259 = rob_uop_3_16_flush_on_commit;
      5'b10001:
        casez_tmp_259 = rob_uop_3_17_flush_on_commit;
      5'b10010:
        casez_tmp_259 = rob_uop_3_18_flush_on_commit;
      5'b10011:
        casez_tmp_259 = rob_uop_3_19_flush_on_commit;
      5'b10100:
        casez_tmp_259 = rob_uop_3_20_flush_on_commit;
      5'b10101:
        casez_tmp_259 = rob_uop_3_21_flush_on_commit;
      5'b10110:
        casez_tmp_259 = rob_uop_3_22_flush_on_commit;
      5'b10111:
        casez_tmp_259 = rob_uop_3_23_flush_on_commit;
      5'b11000:
        casez_tmp_259 = rob_uop_3_24_flush_on_commit;
      5'b11001:
        casez_tmp_259 = rob_uop_3_25_flush_on_commit;
      5'b11010:
        casez_tmp_259 = rob_uop_3_26_flush_on_commit;
      5'b11011:
        casez_tmp_259 = rob_uop_3_27_flush_on_commit;
      5'b11100:
        casez_tmp_259 = rob_uop_3_28_flush_on_commit;
      5'b11101:
        casez_tmp_259 = rob_uop_3_29_flush_on_commit;
      5'b11110:
        casez_tmp_259 = rob_uop_3_30_flush_on_commit;
      default:
        casez_tmp_259 = rob_uop_3_31_flush_on_commit;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_260;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_260 = rob_uop_3_0_ldst;
      5'b00001:
        casez_tmp_260 = rob_uop_3_1_ldst;
      5'b00010:
        casez_tmp_260 = rob_uop_3_2_ldst;
      5'b00011:
        casez_tmp_260 = rob_uop_3_3_ldst;
      5'b00100:
        casez_tmp_260 = rob_uop_3_4_ldst;
      5'b00101:
        casez_tmp_260 = rob_uop_3_5_ldst;
      5'b00110:
        casez_tmp_260 = rob_uop_3_6_ldst;
      5'b00111:
        casez_tmp_260 = rob_uop_3_7_ldst;
      5'b01000:
        casez_tmp_260 = rob_uop_3_8_ldst;
      5'b01001:
        casez_tmp_260 = rob_uop_3_9_ldst;
      5'b01010:
        casez_tmp_260 = rob_uop_3_10_ldst;
      5'b01011:
        casez_tmp_260 = rob_uop_3_11_ldst;
      5'b01100:
        casez_tmp_260 = rob_uop_3_12_ldst;
      5'b01101:
        casez_tmp_260 = rob_uop_3_13_ldst;
      5'b01110:
        casez_tmp_260 = rob_uop_3_14_ldst;
      5'b01111:
        casez_tmp_260 = rob_uop_3_15_ldst;
      5'b10000:
        casez_tmp_260 = rob_uop_3_16_ldst;
      5'b10001:
        casez_tmp_260 = rob_uop_3_17_ldst;
      5'b10010:
        casez_tmp_260 = rob_uop_3_18_ldst;
      5'b10011:
        casez_tmp_260 = rob_uop_3_19_ldst;
      5'b10100:
        casez_tmp_260 = rob_uop_3_20_ldst;
      5'b10101:
        casez_tmp_260 = rob_uop_3_21_ldst;
      5'b10110:
        casez_tmp_260 = rob_uop_3_22_ldst;
      5'b10111:
        casez_tmp_260 = rob_uop_3_23_ldst;
      5'b11000:
        casez_tmp_260 = rob_uop_3_24_ldst;
      5'b11001:
        casez_tmp_260 = rob_uop_3_25_ldst;
      5'b11010:
        casez_tmp_260 = rob_uop_3_26_ldst;
      5'b11011:
        casez_tmp_260 = rob_uop_3_27_ldst;
      5'b11100:
        casez_tmp_260 = rob_uop_3_28_ldst;
      5'b11101:
        casez_tmp_260 = rob_uop_3_29_ldst;
      5'b11110:
        casez_tmp_260 = rob_uop_3_30_ldst;
      default:
        casez_tmp_260 = rob_uop_3_31_ldst;
    endcase
  end // always @(*)
  reg         casez_tmp_261;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_261 = rob_uop_3_0_ldst_val;
      5'b00001:
        casez_tmp_261 = rob_uop_3_1_ldst_val;
      5'b00010:
        casez_tmp_261 = rob_uop_3_2_ldst_val;
      5'b00011:
        casez_tmp_261 = rob_uop_3_3_ldst_val;
      5'b00100:
        casez_tmp_261 = rob_uop_3_4_ldst_val;
      5'b00101:
        casez_tmp_261 = rob_uop_3_5_ldst_val;
      5'b00110:
        casez_tmp_261 = rob_uop_3_6_ldst_val;
      5'b00111:
        casez_tmp_261 = rob_uop_3_7_ldst_val;
      5'b01000:
        casez_tmp_261 = rob_uop_3_8_ldst_val;
      5'b01001:
        casez_tmp_261 = rob_uop_3_9_ldst_val;
      5'b01010:
        casez_tmp_261 = rob_uop_3_10_ldst_val;
      5'b01011:
        casez_tmp_261 = rob_uop_3_11_ldst_val;
      5'b01100:
        casez_tmp_261 = rob_uop_3_12_ldst_val;
      5'b01101:
        casez_tmp_261 = rob_uop_3_13_ldst_val;
      5'b01110:
        casez_tmp_261 = rob_uop_3_14_ldst_val;
      5'b01111:
        casez_tmp_261 = rob_uop_3_15_ldst_val;
      5'b10000:
        casez_tmp_261 = rob_uop_3_16_ldst_val;
      5'b10001:
        casez_tmp_261 = rob_uop_3_17_ldst_val;
      5'b10010:
        casez_tmp_261 = rob_uop_3_18_ldst_val;
      5'b10011:
        casez_tmp_261 = rob_uop_3_19_ldst_val;
      5'b10100:
        casez_tmp_261 = rob_uop_3_20_ldst_val;
      5'b10101:
        casez_tmp_261 = rob_uop_3_21_ldst_val;
      5'b10110:
        casez_tmp_261 = rob_uop_3_22_ldst_val;
      5'b10111:
        casez_tmp_261 = rob_uop_3_23_ldst_val;
      5'b11000:
        casez_tmp_261 = rob_uop_3_24_ldst_val;
      5'b11001:
        casez_tmp_261 = rob_uop_3_25_ldst_val;
      5'b11010:
        casez_tmp_261 = rob_uop_3_26_ldst_val;
      5'b11011:
        casez_tmp_261 = rob_uop_3_27_ldst_val;
      5'b11100:
        casez_tmp_261 = rob_uop_3_28_ldst_val;
      5'b11101:
        casez_tmp_261 = rob_uop_3_29_ldst_val;
      5'b11110:
        casez_tmp_261 = rob_uop_3_30_ldst_val;
      default:
        casez_tmp_261 = rob_uop_3_31_ldst_val;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_262;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_262 = rob_uop_3_0_dst_rtype;
      5'b00001:
        casez_tmp_262 = rob_uop_3_1_dst_rtype;
      5'b00010:
        casez_tmp_262 = rob_uop_3_2_dst_rtype;
      5'b00011:
        casez_tmp_262 = rob_uop_3_3_dst_rtype;
      5'b00100:
        casez_tmp_262 = rob_uop_3_4_dst_rtype;
      5'b00101:
        casez_tmp_262 = rob_uop_3_5_dst_rtype;
      5'b00110:
        casez_tmp_262 = rob_uop_3_6_dst_rtype;
      5'b00111:
        casez_tmp_262 = rob_uop_3_7_dst_rtype;
      5'b01000:
        casez_tmp_262 = rob_uop_3_8_dst_rtype;
      5'b01001:
        casez_tmp_262 = rob_uop_3_9_dst_rtype;
      5'b01010:
        casez_tmp_262 = rob_uop_3_10_dst_rtype;
      5'b01011:
        casez_tmp_262 = rob_uop_3_11_dst_rtype;
      5'b01100:
        casez_tmp_262 = rob_uop_3_12_dst_rtype;
      5'b01101:
        casez_tmp_262 = rob_uop_3_13_dst_rtype;
      5'b01110:
        casez_tmp_262 = rob_uop_3_14_dst_rtype;
      5'b01111:
        casez_tmp_262 = rob_uop_3_15_dst_rtype;
      5'b10000:
        casez_tmp_262 = rob_uop_3_16_dst_rtype;
      5'b10001:
        casez_tmp_262 = rob_uop_3_17_dst_rtype;
      5'b10010:
        casez_tmp_262 = rob_uop_3_18_dst_rtype;
      5'b10011:
        casez_tmp_262 = rob_uop_3_19_dst_rtype;
      5'b10100:
        casez_tmp_262 = rob_uop_3_20_dst_rtype;
      5'b10101:
        casez_tmp_262 = rob_uop_3_21_dst_rtype;
      5'b10110:
        casez_tmp_262 = rob_uop_3_22_dst_rtype;
      5'b10111:
        casez_tmp_262 = rob_uop_3_23_dst_rtype;
      5'b11000:
        casez_tmp_262 = rob_uop_3_24_dst_rtype;
      5'b11001:
        casez_tmp_262 = rob_uop_3_25_dst_rtype;
      5'b11010:
        casez_tmp_262 = rob_uop_3_26_dst_rtype;
      5'b11011:
        casez_tmp_262 = rob_uop_3_27_dst_rtype;
      5'b11100:
        casez_tmp_262 = rob_uop_3_28_dst_rtype;
      5'b11101:
        casez_tmp_262 = rob_uop_3_29_dst_rtype;
      5'b11110:
        casez_tmp_262 = rob_uop_3_30_dst_rtype;
      default:
        casez_tmp_262 = rob_uop_3_31_dst_rtype;
    endcase
  end // always @(*)
  reg         casez_tmp_263;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_263 = rob_uop_3_0_fp_val;
      5'b00001:
        casez_tmp_263 = rob_uop_3_1_fp_val;
      5'b00010:
        casez_tmp_263 = rob_uop_3_2_fp_val;
      5'b00011:
        casez_tmp_263 = rob_uop_3_3_fp_val;
      5'b00100:
        casez_tmp_263 = rob_uop_3_4_fp_val;
      5'b00101:
        casez_tmp_263 = rob_uop_3_5_fp_val;
      5'b00110:
        casez_tmp_263 = rob_uop_3_6_fp_val;
      5'b00111:
        casez_tmp_263 = rob_uop_3_7_fp_val;
      5'b01000:
        casez_tmp_263 = rob_uop_3_8_fp_val;
      5'b01001:
        casez_tmp_263 = rob_uop_3_9_fp_val;
      5'b01010:
        casez_tmp_263 = rob_uop_3_10_fp_val;
      5'b01011:
        casez_tmp_263 = rob_uop_3_11_fp_val;
      5'b01100:
        casez_tmp_263 = rob_uop_3_12_fp_val;
      5'b01101:
        casez_tmp_263 = rob_uop_3_13_fp_val;
      5'b01110:
        casez_tmp_263 = rob_uop_3_14_fp_val;
      5'b01111:
        casez_tmp_263 = rob_uop_3_15_fp_val;
      5'b10000:
        casez_tmp_263 = rob_uop_3_16_fp_val;
      5'b10001:
        casez_tmp_263 = rob_uop_3_17_fp_val;
      5'b10010:
        casez_tmp_263 = rob_uop_3_18_fp_val;
      5'b10011:
        casez_tmp_263 = rob_uop_3_19_fp_val;
      5'b10100:
        casez_tmp_263 = rob_uop_3_20_fp_val;
      5'b10101:
        casez_tmp_263 = rob_uop_3_21_fp_val;
      5'b10110:
        casez_tmp_263 = rob_uop_3_22_fp_val;
      5'b10111:
        casez_tmp_263 = rob_uop_3_23_fp_val;
      5'b11000:
        casez_tmp_263 = rob_uop_3_24_fp_val;
      5'b11001:
        casez_tmp_263 = rob_uop_3_25_fp_val;
      5'b11010:
        casez_tmp_263 = rob_uop_3_26_fp_val;
      5'b11011:
        casez_tmp_263 = rob_uop_3_27_fp_val;
      5'b11100:
        casez_tmp_263 = rob_uop_3_28_fp_val;
      5'b11101:
        casez_tmp_263 = rob_uop_3_29_fp_val;
      5'b11110:
        casez_tmp_263 = rob_uop_3_30_fp_val;
      default:
        casez_tmp_263 = rob_uop_3_31_fp_val;
    endcase
  end // always @(*)
  reg  [1:0]  casez_tmp_264;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_264 = rob_uop_3_0_debug_fsrc;
      5'b00001:
        casez_tmp_264 = rob_uop_3_1_debug_fsrc;
      5'b00010:
        casez_tmp_264 = rob_uop_3_2_debug_fsrc;
      5'b00011:
        casez_tmp_264 = rob_uop_3_3_debug_fsrc;
      5'b00100:
        casez_tmp_264 = rob_uop_3_4_debug_fsrc;
      5'b00101:
        casez_tmp_264 = rob_uop_3_5_debug_fsrc;
      5'b00110:
        casez_tmp_264 = rob_uop_3_6_debug_fsrc;
      5'b00111:
        casez_tmp_264 = rob_uop_3_7_debug_fsrc;
      5'b01000:
        casez_tmp_264 = rob_uop_3_8_debug_fsrc;
      5'b01001:
        casez_tmp_264 = rob_uop_3_9_debug_fsrc;
      5'b01010:
        casez_tmp_264 = rob_uop_3_10_debug_fsrc;
      5'b01011:
        casez_tmp_264 = rob_uop_3_11_debug_fsrc;
      5'b01100:
        casez_tmp_264 = rob_uop_3_12_debug_fsrc;
      5'b01101:
        casez_tmp_264 = rob_uop_3_13_debug_fsrc;
      5'b01110:
        casez_tmp_264 = rob_uop_3_14_debug_fsrc;
      5'b01111:
        casez_tmp_264 = rob_uop_3_15_debug_fsrc;
      5'b10000:
        casez_tmp_264 = rob_uop_3_16_debug_fsrc;
      5'b10001:
        casez_tmp_264 = rob_uop_3_17_debug_fsrc;
      5'b10010:
        casez_tmp_264 = rob_uop_3_18_debug_fsrc;
      5'b10011:
        casez_tmp_264 = rob_uop_3_19_debug_fsrc;
      5'b10100:
        casez_tmp_264 = rob_uop_3_20_debug_fsrc;
      5'b10101:
        casez_tmp_264 = rob_uop_3_21_debug_fsrc;
      5'b10110:
        casez_tmp_264 = rob_uop_3_22_debug_fsrc;
      5'b10111:
        casez_tmp_264 = rob_uop_3_23_debug_fsrc;
      5'b11000:
        casez_tmp_264 = rob_uop_3_24_debug_fsrc;
      5'b11001:
        casez_tmp_264 = rob_uop_3_25_debug_fsrc;
      5'b11010:
        casez_tmp_264 = rob_uop_3_26_debug_fsrc;
      5'b11011:
        casez_tmp_264 = rob_uop_3_27_debug_fsrc;
      5'b11100:
        casez_tmp_264 = rob_uop_3_28_debug_fsrc;
      5'b11101:
        casez_tmp_264 = rob_uop_3_29_debug_fsrc;
      5'b11110:
        casez_tmp_264 = rob_uop_3_30_debug_fsrc;
      default:
        casez_tmp_264 = rob_uop_3_31_debug_fsrc;
    endcase
  end // always @(*)
  wire        _GEN_64 = io_brupdate_b2_mispredict & (&(io_brupdate_b2_uop_rob_idx[1:0]));
  wire        rbk_row_3 = _io_commit_rollback_T_3 & ~full;
  reg         casez_tmp_265;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_265 = rob_val_3_0;
      5'b00001:
        casez_tmp_265 = rob_val_3_1;
      5'b00010:
        casez_tmp_265 = rob_val_3_2;
      5'b00011:
        casez_tmp_265 = rob_val_3_3;
      5'b00100:
        casez_tmp_265 = rob_val_3_4;
      5'b00101:
        casez_tmp_265 = rob_val_3_5;
      5'b00110:
        casez_tmp_265 = rob_val_3_6;
      5'b00111:
        casez_tmp_265 = rob_val_3_7;
      5'b01000:
        casez_tmp_265 = rob_val_3_8;
      5'b01001:
        casez_tmp_265 = rob_val_3_9;
      5'b01010:
        casez_tmp_265 = rob_val_3_10;
      5'b01011:
        casez_tmp_265 = rob_val_3_11;
      5'b01100:
        casez_tmp_265 = rob_val_3_12;
      5'b01101:
        casez_tmp_265 = rob_val_3_13;
      5'b01110:
        casez_tmp_265 = rob_val_3_14;
      5'b01111:
        casez_tmp_265 = rob_val_3_15;
      5'b10000:
        casez_tmp_265 = rob_val_3_16;
      5'b10001:
        casez_tmp_265 = rob_val_3_17;
      5'b10010:
        casez_tmp_265 = rob_val_3_18;
      5'b10011:
        casez_tmp_265 = rob_val_3_19;
      5'b10100:
        casez_tmp_265 = rob_val_3_20;
      5'b10101:
        casez_tmp_265 = rob_val_3_21;
      5'b10110:
        casez_tmp_265 = rob_val_3_22;
      5'b10111:
        casez_tmp_265 = rob_val_3_23;
      5'b11000:
        casez_tmp_265 = rob_val_3_24;
      5'b11001:
        casez_tmp_265 = rob_val_3_25;
      5'b11010:
        casez_tmp_265 = rob_val_3_26;
      5'b11011:
        casez_tmp_265 = rob_val_3_27;
      5'b11100:
        casez_tmp_265 = rob_val_3_28;
      5'b11101:
        casez_tmp_265 = rob_val_3_29;
      5'b11110:
        casez_tmp_265 = rob_val_3_30;
      default:
        casez_tmp_265 = rob_val_3_31;
    endcase
  end // always @(*)
  wire        _io_commit_rbk_valids_3_output = rbk_row_3 & casez_tmp_265;
  reg  [4:0]  casez_tmp_266;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_266 = rob_fflags_3_0;
      5'b00001:
        casez_tmp_266 = rob_fflags_3_1;
      5'b00010:
        casez_tmp_266 = rob_fflags_3_2;
      5'b00011:
        casez_tmp_266 = rob_fflags_3_3;
      5'b00100:
        casez_tmp_266 = rob_fflags_3_4;
      5'b00101:
        casez_tmp_266 = rob_fflags_3_5;
      5'b00110:
        casez_tmp_266 = rob_fflags_3_6;
      5'b00111:
        casez_tmp_266 = rob_fflags_3_7;
      5'b01000:
        casez_tmp_266 = rob_fflags_3_8;
      5'b01001:
        casez_tmp_266 = rob_fflags_3_9;
      5'b01010:
        casez_tmp_266 = rob_fflags_3_10;
      5'b01011:
        casez_tmp_266 = rob_fflags_3_11;
      5'b01100:
        casez_tmp_266 = rob_fflags_3_12;
      5'b01101:
        casez_tmp_266 = rob_fflags_3_13;
      5'b01110:
        casez_tmp_266 = rob_fflags_3_14;
      5'b01111:
        casez_tmp_266 = rob_fflags_3_15;
      5'b10000:
        casez_tmp_266 = rob_fflags_3_16;
      5'b10001:
        casez_tmp_266 = rob_fflags_3_17;
      5'b10010:
        casez_tmp_266 = rob_fflags_3_18;
      5'b10011:
        casez_tmp_266 = rob_fflags_3_19;
      5'b10100:
        casez_tmp_266 = rob_fflags_3_20;
      5'b10101:
        casez_tmp_266 = rob_fflags_3_21;
      5'b10110:
        casez_tmp_266 = rob_fflags_3_22;
      5'b10111:
        casez_tmp_266 = rob_fflags_3_23;
      5'b11000:
        casez_tmp_266 = rob_fflags_3_24;
      5'b11001:
        casez_tmp_266 = rob_fflags_3_25;
      5'b11010:
        casez_tmp_266 = rob_fflags_3_26;
      5'b11011:
        casez_tmp_266 = rob_fflags_3_27;
      5'b11100:
        casez_tmp_266 = rob_fflags_3_28;
      5'b11101:
        casez_tmp_266 = rob_fflags_3_29;
      5'b11110:
        casez_tmp_266 = rob_fflags_3_30;
      default:
        casez_tmp_266 = rob_fflags_3_31;
    endcase
  end // always @(*)
  reg         casez_tmp_267;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_267 = rob_uop_3_0_uses_ldq;
      5'b00001:
        casez_tmp_267 = rob_uop_3_1_uses_ldq;
      5'b00010:
        casez_tmp_267 = rob_uop_3_2_uses_ldq;
      5'b00011:
        casez_tmp_267 = rob_uop_3_3_uses_ldq;
      5'b00100:
        casez_tmp_267 = rob_uop_3_4_uses_ldq;
      5'b00101:
        casez_tmp_267 = rob_uop_3_5_uses_ldq;
      5'b00110:
        casez_tmp_267 = rob_uop_3_6_uses_ldq;
      5'b00111:
        casez_tmp_267 = rob_uop_3_7_uses_ldq;
      5'b01000:
        casez_tmp_267 = rob_uop_3_8_uses_ldq;
      5'b01001:
        casez_tmp_267 = rob_uop_3_9_uses_ldq;
      5'b01010:
        casez_tmp_267 = rob_uop_3_10_uses_ldq;
      5'b01011:
        casez_tmp_267 = rob_uop_3_11_uses_ldq;
      5'b01100:
        casez_tmp_267 = rob_uop_3_12_uses_ldq;
      5'b01101:
        casez_tmp_267 = rob_uop_3_13_uses_ldq;
      5'b01110:
        casez_tmp_267 = rob_uop_3_14_uses_ldq;
      5'b01111:
        casez_tmp_267 = rob_uop_3_15_uses_ldq;
      5'b10000:
        casez_tmp_267 = rob_uop_3_16_uses_ldq;
      5'b10001:
        casez_tmp_267 = rob_uop_3_17_uses_ldq;
      5'b10010:
        casez_tmp_267 = rob_uop_3_18_uses_ldq;
      5'b10011:
        casez_tmp_267 = rob_uop_3_19_uses_ldq;
      5'b10100:
        casez_tmp_267 = rob_uop_3_20_uses_ldq;
      5'b10101:
        casez_tmp_267 = rob_uop_3_21_uses_ldq;
      5'b10110:
        casez_tmp_267 = rob_uop_3_22_uses_ldq;
      5'b10111:
        casez_tmp_267 = rob_uop_3_23_uses_ldq;
      5'b11000:
        casez_tmp_267 = rob_uop_3_24_uses_ldq;
      5'b11001:
        casez_tmp_267 = rob_uop_3_25_uses_ldq;
      5'b11010:
        casez_tmp_267 = rob_uop_3_26_uses_ldq;
      5'b11011:
        casez_tmp_267 = rob_uop_3_27_uses_ldq;
      5'b11100:
        casez_tmp_267 = rob_uop_3_28_uses_ldq;
      5'b11101:
        casez_tmp_267 = rob_uop_3_29_uses_ldq;
      5'b11110:
        casez_tmp_267 = rob_uop_3_30_uses_ldq;
      default:
        casez_tmp_267 = rob_uop_3_31_uses_ldq;
    endcase
  end // always @(*)
  reg         casez_tmp_268;
  always @(*) begin
    casez (rob_pnr)
      5'b00000:
        casez_tmp_268 = rob_unsafe_3_0;
      5'b00001:
        casez_tmp_268 = rob_unsafe_3_1;
      5'b00010:
        casez_tmp_268 = rob_unsafe_3_2;
      5'b00011:
        casez_tmp_268 = rob_unsafe_3_3;
      5'b00100:
        casez_tmp_268 = rob_unsafe_3_4;
      5'b00101:
        casez_tmp_268 = rob_unsafe_3_5;
      5'b00110:
        casez_tmp_268 = rob_unsafe_3_6;
      5'b00111:
        casez_tmp_268 = rob_unsafe_3_7;
      5'b01000:
        casez_tmp_268 = rob_unsafe_3_8;
      5'b01001:
        casez_tmp_268 = rob_unsafe_3_9;
      5'b01010:
        casez_tmp_268 = rob_unsafe_3_10;
      5'b01011:
        casez_tmp_268 = rob_unsafe_3_11;
      5'b01100:
        casez_tmp_268 = rob_unsafe_3_12;
      5'b01101:
        casez_tmp_268 = rob_unsafe_3_13;
      5'b01110:
        casez_tmp_268 = rob_unsafe_3_14;
      5'b01111:
        casez_tmp_268 = rob_unsafe_3_15;
      5'b10000:
        casez_tmp_268 = rob_unsafe_3_16;
      5'b10001:
        casez_tmp_268 = rob_unsafe_3_17;
      5'b10010:
        casez_tmp_268 = rob_unsafe_3_18;
      5'b10011:
        casez_tmp_268 = rob_unsafe_3_19;
      5'b10100:
        casez_tmp_268 = rob_unsafe_3_20;
      5'b10101:
        casez_tmp_268 = rob_unsafe_3_21;
      5'b10110:
        casez_tmp_268 = rob_unsafe_3_22;
      5'b10111:
        casez_tmp_268 = rob_unsafe_3_23;
      5'b11000:
        casez_tmp_268 = rob_unsafe_3_24;
      5'b11001:
        casez_tmp_268 = rob_unsafe_3_25;
      5'b11010:
        casez_tmp_268 = rob_unsafe_3_26;
      5'b11011:
        casez_tmp_268 = rob_unsafe_3_27;
      5'b11100:
        casez_tmp_268 = rob_unsafe_3_28;
      5'b11101:
        casez_tmp_268 = rob_unsafe_3_29;
      5'b11110:
        casez_tmp_268 = rob_unsafe_3_30;
      default:
        casez_tmp_268 = rob_unsafe_3_31;
    endcase
  end // always @(*)
  reg         casez_tmp_269;
  always @(*) begin
    casez (rob_pnr)
      5'b00000:
        casez_tmp_269 = rob_exception_3_0;
      5'b00001:
        casez_tmp_269 = rob_exception_3_1;
      5'b00010:
        casez_tmp_269 = rob_exception_3_2;
      5'b00011:
        casez_tmp_269 = rob_exception_3_3;
      5'b00100:
        casez_tmp_269 = rob_exception_3_4;
      5'b00101:
        casez_tmp_269 = rob_exception_3_5;
      5'b00110:
        casez_tmp_269 = rob_exception_3_6;
      5'b00111:
        casez_tmp_269 = rob_exception_3_7;
      5'b01000:
        casez_tmp_269 = rob_exception_3_8;
      5'b01001:
        casez_tmp_269 = rob_exception_3_9;
      5'b01010:
        casez_tmp_269 = rob_exception_3_10;
      5'b01011:
        casez_tmp_269 = rob_exception_3_11;
      5'b01100:
        casez_tmp_269 = rob_exception_3_12;
      5'b01101:
        casez_tmp_269 = rob_exception_3_13;
      5'b01110:
        casez_tmp_269 = rob_exception_3_14;
      5'b01111:
        casez_tmp_269 = rob_exception_3_15;
      5'b10000:
        casez_tmp_269 = rob_exception_3_16;
      5'b10001:
        casez_tmp_269 = rob_exception_3_17;
      5'b10010:
        casez_tmp_269 = rob_exception_3_18;
      5'b10011:
        casez_tmp_269 = rob_exception_3_19;
      5'b10100:
        casez_tmp_269 = rob_exception_3_20;
      5'b10101:
        casez_tmp_269 = rob_exception_3_21;
      5'b10110:
        casez_tmp_269 = rob_exception_3_22;
      5'b10111:
        casez_tmp_269 = rob_exception_3_23;
      5'b11000:
        casez_tmp_269 = rob_exception_3_24;
      5'b11001:
        casez_tmp_269 = rob_exception_3_25;
      5'b11010:
        casez_tmp_269 = rob_exception_3_26;
      5'b11011:
        casez_tmp_269 = rob_exception_3_27;
      5'b11100:
        casez_tmp_269 = rob_exception_3_28;
      5'b11101:
        casez_tmp_269 = rob_exception_3_29;
      5'b11110:
        casez_tmp_269 = rob_exception_3_30;
      default:
        casez_tmp_269 = rob_exception_3_31;
    endcase
  end // always @(*)
  reg         casez_tmp_270;
  always @(*) begin
    casez (rob_pnr)
      5'b00000:
        casez_tmp_270 = rob_val_3_0;
      5'b00001:
        casez_tmp_270 = rob_val_3_1;
      5'b00010:
        casez_tmp_270 = rob_val_3_2;
      5'b00011:
        casez_tmp_270 = rob_val_3_3;
      5'b00100:
        casez_tmp_270 = rob_val_3_4;
      5'b00101:
        casez_tmp_270 = rob_val_3_5;
      5'b00110:
        casez_tmp_270 = rob_val_3_6;
      5'b00111:
        casez_tmp_270 = rob_val_3_7;
      5'b01000:
        casez_tmp_270 = rob_val_3_8;
      5'b01001:
        casez_tmp_270 = rob_val_3_9;
      5'b01010:
        casez_tmp_270 = rob_val_3_10;
      5'b01011:
        casez_tmp_270 = rob_val_3_11;
      5'b01100:
        casez_tmp_270 = rob_val_3_12;
      5'b01101:
        casez_tmp_270 = rob_val_3_13;
      5'b01110:
        casez_tmp_270 = rob_val_3_14;
      5'b01111:
        casez_tmp_270 = rob_val_3_15;
      5'b10000:
        casez_tmp_270 = rob_val_3_16;
      5'b10001:
        casez_tmp_270 = rob_val_3_17;
      5'b10010:
        casez_tmp_270 = rob_val_3_18;
      5'b10011:
        casez_tmp_270 = rob_val_3_19;
      5'b10100:
        casez_tmp_270 = rob_val_3_20;
      5'b10101:
        casez_tmp_270 = rob_val_3_21;
      5'b10110:
        casez_tmp_270 = rob_val_3_22;
      5'b10111:
        casez_tmp_270 = rob_val_3_23;
      5'b11000:
        casez_tmp_270 = rob_val_3_24;
      5'b11001:
        casez_tmp_270 = rob_val_3_25;
      5'b11010:
        casez_tmp_270 = rob_val_3_26;
      5'b11011:
        casez_tmp_270 = rob_val_3_27;
      5'b11100:
        casez_tmp_270 = rob_val_3_28;
      5'b11101:
        casez_tmp_270 = rob_val_3_29;
      5'b11110:
        casez_tmp_270 = rob_val_3_30;
      default:
        casez_tmp_270 = rob_val_3_31;
    endcase
  end // always @(*)
  reg         casez_tmp_271;
  always @(*) begin
    casez (io_wb_resps_0_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_271 = rob_val_3_0;
      5'b00001:
        casez_tmp_271 = rob_val_3_1;
      5'b00010:
        casez_tmp_271 = rob_val_3_2;
      5'b00011:
        casez_tmp_271 = rob_val_3_3;
      5'b00100:
        casez_tmp_271 = rob_val_3_4;
      5'b00101:
        casez_tmp_271 = rob_val_3_5;
      5'b00110:
        casez_tmp_271 = rob_val_3_6;
      5'b00111:
        casez_tmp_271 = rob_val_3_7;
      5'b01000:
        casez_tmp_271 = rob_val_3_8;
      5'b01001:
        casez_tmp_271 = rob_val_3_9;
      5'b01010:
        casez_tmp_271 = rob_val_3_10;
      5'b01011:
        casez_tmp_271 = rob_val_3_11;
      5'b01100:
        casez_tmp_271 = rob_val_3_12;
      5'b01101:
        casez_tmp_271 = rob_val_3_13;
      5'b01110:
        casez_tmp_271 = rob_val_3_14;
      5'b01111:
        casez_tmp_271 = rob_val_3_15;
      5'b10000:
        casez_tmp_271 = rob_val_3_16;
      5'b10001:
        casez_tmp_271 = rob_val_3_17;
      5'b10010:
        casez_tmp_271 = rob_val_3_18;
      5'b10011:
        casez_tmp_271 = rob_val_3_19;
      5'b10100:
        casez_tmp_271 = rob_val_3_20;
      5'b10101:
        casez_tmp_271 = rob_val_3_21;
      5'b10110:
        casez_tmp_271 = rob_val_3_22;
      5'b10111:
        casez_tmp_271 = rob_val_3_23;
      5'b11000:
        casez_tmp_271 = rob_val_3_24;
      5'b11001:
        casez_tmp_271 = rob_val_3_25;
      5'b11010:
        casez_tmp_271 = rob_val_3_26;
      5'b11011:
        casez_tmp_271 = rob_val_3_27;
      5'b11100:
        casez_tmp_271 = rob_val_3_28;
      5'b11101:
        casez_tmp_271 = rob_val_3_29;
      5'b11110:
        casez_tmp_271 = rob_val_3_30;
      default:
        casez_tmp_271 = rob_val_3_31;
    endcase
  end // always @(*)
  reg         casez_tmp_272;
  always @(*) begin
    casez (io_wb_resps_0_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_272 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_272 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_272 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_272 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_272 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_272 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_272 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_272 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_272 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_272 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_272 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_272 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_272 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_272 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_272 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_272 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_272 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_272 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_272 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_272 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_272 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_272 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_272 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_272 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_272 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_272 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_272 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_272 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_272 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_272 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_272 = rob_bsy_3_30;
      default:
        casez_tmp_272 = rob_bsy_3_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_273;
  always @(*) begin
    casez (io_wb_resps_0_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_273 = rob_uop_3_0_pdst;
      5'b00001:
        casez_tmp_273 = rob_uop_3_1_pdst;
      5'b00010:
        casez_tmp_273 = rob_uop_3_2_pdst;
      5'b00011:
        casez_tmp_273 = rob_uop_3_3_pdst;
      5'b00100:
        casez_tmp_273 = rob_uop_3_4_pdst;
      5'b00101:
        casez_tmp_273 = rob_uop_3_5_pdst;
      5'b00110:
        casez_tmp_273 = rob_uop_3_6_pdst;
      5'b00111:
        casez_tmp_273 = rob_uop_3_7_pdst;
      5'b01000:
        casez_tmp_273 = rob_uop_3_8_pdst;
      5'b01001:
        casez_tmp_273 = rob_uop_3_9_pdst;
      5'b01010:
        casez_tmp_273 = rob_uop_3_10_pdst;
      5'b01011:
        casez_tmp_273 = rob_uop_3_11_pdst;
      5'b01100:
        casez_tmp_273 = rob_uop_3_12_pdst;
      5'b01101:
        casez_tmp_273 = rob_uop_3_13_pdst;
      5'b01110:
        casez_tmp_273 = rob_uop_3_14_pdst;
      5'b01111:
        casez_tmp_273 = rob_uop_3_15_pdst;
      5'b10000:
        casez_tmp_273 = rob_uop_3_16_pdst;
      5'b10001:
        casez_tmp_273 = rob_uop_3_17_pdst;
      5'b10010:
        casez_tmp_273 = rob_uop_3_18_pdst;
      5'b10011:
        casez_tmp_273 = rob_uop_3_19_pdst;
      5'b10100:
        casez_tmp_273 = rob_uop_3_20_pdst;
      5'b10101:
        casez_tmp_273 = rob_uop_3_21_pdst;
      5'b10110:
        casez_tmp_273 = rob_uop_3_22_pdst;
      5'b10111:
        casez_tmp_273 = rob_uop_3_23_pdst;
      5'b11000:
        casez_tmp_273 = rob_uop_3_24_pdst;
      5'b11001:
        casez_tmp_273 = rob_uop_3_25_pdst;
      5'b11010:
        casez_tmp_273 = rob_uop_3_26_pdst;
      5'b11011:
        casez_tmp_273 = rob_uop_3_27_pdst;
      5'b11100:
        casez_tmp_273 = rob_uop_3_28_pdst;
      5'b11101:
        casez_tmp_273 = rob_uop_3_29_pdst;
      5'b11110:
        casez_tmp_273 = rob_uop_3_30_pdst;
      default:
        casez_tmp_273 = rob_uop_3_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_274;
  always @(*) begin
    casez (io_wb_resps_0_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_274 = rob_uop_3_0_ldst_val;
      5'b00001:
        casez_tmp_274 = rob_uop_3_1_ldst_val;
      5'b00010:
        casez_tmp_274 = rob_uop_3_2_ldst_val;
      5'b00011:
        casez_tmp_274 = rob_uop_3_3_ldst_val;
      5'b00100:
        casez_tmp_274 = rob_uop_3_4_ldst_val;
      5'b00101:
        casez_tmp_274 = rob_uop_3_5_ldst_val;
      5'b00110:
        casez_tmp_274 = rob_uop_3_6_ldst_val;
      5'b00111:
        casez_tmp_274 = rob_uop_3_7_ldst_val;
      5'b01000:
        casez_tmp_274 = rob_uop_3_8_ldst_val;
      5'b01001:
        casez_tmp_274 = rob_uop_3_9_ldst_val;
      5'b01010:
        casez_tmp_274 = rob_uop_3_10_ldst_val;
      5'b01011:
        casez_tmp_274 = rob_uop_3_11_ldst_val;
      5'b01100:
        casez_tmp_274 = rob_uop_3_12_ldst_val;
      5'b01101:
        casez_tmp_274 = rob_uop_3_13_ldst_val;
      5'b01110:
        casez_tmp_274 = rob_uop_3_14_ldst_val;
      5'b01111:
        casez_tmp_274 = rob_uop_3_15_ldst_val;
      5'b10000:
        casez_tmp_274 = rob_uop_3_16_ldst_val;
      5'b10001:
        casez_tmp_274 = rob_uop_3_17_ldst_val;
      5'b10010:
        casez_tmp_274 = rob_uop_3_18_ldst_val;
      5'b10011:
        casez_tmp_274 = rob_uop_3_19_ldst_val;
      5'b10100:
        casez_tmp_274 = rob_uop_3_20_ldst_val;
      5'b10101:
        casez_tmp_274 = rob_uop_3_21_ldst_val;
      5'b10110:
        casez_tmp_274 = rob_uop_3_22_ldst_val;
      5'b10111:
        casez_tmp_274 = rob_uop_3_23_ldst_val;
      5'b11000:
        casez_tmp_274 = rob_uop_3_24_ldst_val;
      5'b11001:
        casez_tmp_274 = rob_uop_3_25_ldst_val;
      5'b11010:
        casez_tmp_274 = rob_uop_3_26_ldst_val;
      5'b11011:
        casez_tmp_274 = rob_uop_3_27_ldst_val;
      5'b11100:
        casez_tmp_274 = rob_uop_3_28_ldst_val;
      5'b11101:
        casez_tmp_274 = rob_uop_3_29_ldst_val;
      5'b11110:
        casez_tmp_274 = rob_uop_3_30_ldst_val;
      default:
        casez_tmp_274 = rob_uop_3_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_275;
  always @(*) begin
    casez (io_wb_resps_1_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_275 = rob_val_3_0;
      5'b00001:
        casez_tmp_275 = rob_val_3_1;
      5'b00010:
        casez_tmp_275 = rob_val_3_2;
      5'b00011:
        casez_tmp_275 = rob_val_3_3;
      5'b00100:
        casez_tmp_275 = rob_val_3_4;
      5'b00101:
        casez_tmp_275 = rob_val_3_5;
      5'b00110:
        casez_tmp_275 = rob_val_3_6;
      5'b00111:
        casez_tmp_275 = rob_val_3_7;
      5'b01000:
        casez_tmp_275 = rob_val_3_8;
      5'b01001:
        casez_tmp_275 = rob_val_3_9;
      5'b01010:
        casez_tmp_275 = rob_val_3_10;
      5'b01011:
        casez_tmp_275 = rob_val_3_11;
      5'b01100:
        casez_tmp_275 = rob_val_3_12;
      5'b01101:
        casez_tmp_275 = rob_val_3_13;
      5'b01110:
        casez_tmp_275 = rob_val_3_14;
      5'b01111:
        casez_tmp_275 = rob_val_3_15;
      5'b10000:
        casez_tmp_275 = rob_val_3_16;
      5'b10001:
        casez_tmp_275 = rob_val_3_17;
      5'b10010:
        casez_tmp_275 = rob_val_3_18;
      5'b10011:
        casez_tmp_275 = rob_val_3_19;
      5'b10100:
        casez_tmp_275 = rob_val_3_20;
      5'b10101:
        casez_tmp_275 = rob_val_3_21;
      5'b10110:
        casez_tmp_275 = rob_val_3_22;
      5'b10111:
        casez_tmp_275 = rob_val_3_23;
      5'b11000:
        casez_tmp_275 = rob_val_3_24;
      5'b11001:
        casez_tmp_275 = rob_val_3_25;
      5'b11010:
        casez_tmp_275 = rob_val_3_26;
      5'b11011:
        casez_tmp_275 = rob_val_3_27;
      5'b11100:
        casez_tmp_275 = rob_val_3_28;
      5'b11101:
        casez_tmp_275 = rob_val_3_29;
      5'b11110:
        casez_tmp_275 = rob_val_3_30;
      default:
        casez_tmp_275 = rob_val_3_31;
    endcase
  end // always @(*)
  reg         casez_tmp_276;
  always @(*) begin
    casez (io_wb_resps_1_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_276 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_276 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_276 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_276 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_276 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_276 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_276 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_276 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_276 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_276 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_276 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_276 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_276 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_276 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_276 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_276 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_276 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_276 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_276 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_276 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_276 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_276 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_276 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_276 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_276 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_276 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_276 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_276 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_276 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_276 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_276 = rob_bsy_3_30;
      default:
        casez_tmp_276 = rob_bsy_3_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_277;
  always @(*) begin
    casez (io_wb_resps_1_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_277 = rob_uop_3_0_pdst;
      5'b00001:
        casez_tmp_277 = rob_uop_3_1_pdst;
      5'b00010:
        casez_tmp_277 = rob_uop_3_2_pdst;
      5'b00011:
        casez_tmp_277 = rob_uop_3_3_pdst;
      5'b00100:
        casez_tmp_277 = rob_uop_3_4_pdst;
      5'b00101:
        casez_tmp_277 = rob_uop_3_5_pdst;
      5'b00110:
        casez_tmp_277 = rob_uop_3_6_pdst;
      5'b00111:
        casez_tmp_277 = rob_uop_3_7_pdst;
      5'b01000:
        casez_tmp_277 = rob_uop_3_8_pdst;
      5'b01001:
        casez_tmp_277 = rob_uop_3_9_pdst;
      5'b01010:
        casez_tmp_277 = rob_uop_3_10_pdst;
      5'b01011:
        casez_tmp_277 = rob_uop_3_11_pdst;
      5'b01100:
        casez_tmp_277 = rob_uop_3_12_pdst;
      5'b01101:
        casez_tmp_277 = rob_uop_3_13_pdst;
      5'b01110:
        casez_tmp_277 = rob_uop_3_14_pdst;
      5'b01111:
        casez_tmp_277 = rob_uop_3_15_pdst;
      5'b10000:
        casez_tmp_277 = rob_uop_3_16_pdst;
      5'b10001:
        casez_tmp_277 = rob_uop_3_17_pdst;
      5'b10010:
        casez_tmp_277 = rob_uop_3_18_pdst;
      5'b10011:
        casez_tmp_277 = rob_uop_3_19_pdst;
      5'b10100:
        casez_tmp_277 = rob_uop_3_20_pdst;
      5'b10101:
        casez_tmp_277 = rob_uop_3_21_pdst;
      5'b10110:
        casez_tmp_277 = rob_uop_3_22_pdst;
      5'b10111:
        casez_tmp_277 = rob_uop_3_23_pdst;
      5'b11000:
        casez_tmp_277 = rob_uop_3_24_pdst;
      5'b11001:
        casez_tmp_277 = rob_uop_3_25_pdst;
      5'b11010:
        casez_tmp_277 = rob_uop_3_26_pdst;
      5'b11011:
        casez_tmp_277 = rob_uop_3_27_pdst;
      5'b11100:
        casez_tmp_277 = rob_uop_3_28_pdst;
      5'b11101:
        casez_tmp_277 = rob_uop_3_29_pdst;
      5'b11110:
        casez_tmp_277 = rob_uop_3_30_pdst;
      default:
        casez_tmp_277 = rob_uop_3_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_278;
  always @(*) begin
    casez (io_wb_resps_1_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_278 = rob_uop_3_0_ldst_val;
      5'b00001:
        casez_tmp_278 = rob_uop_3_1_ldst_val;
      5'b00010:
        casez_tmp_278 = rob_uop_3_2_ldst_val;
      5'b00011:
        casez_tmp_278 = rob_uop_3_3_ldst_val;
      5'b00100:
        casez_tmp_278 = rob_uop_3_4_ldst_val;
      5'b00101:
        casez_tmp_278 = rob_uop_3_5_ldst_val;
      5'b00110:
        casez_tmp_278 = rob_uop_3_6_ldst_val;
      5'b00111:
        casez_tmp_278 = rob_uop_3_7_ldst_val;
      5'b01000:
        casez_tmp_278 = rob_uop_3_8_ldst_val;
      5'b01001:
        casez_tmp_278 = rob_uop_3_9_ldst_val;
      5'b01010:
        casez_tmp_278 = rob_uop_3_10_ldst_val;
      5'b01011:
        casez_tmp_278 = rob_uop_3_11_ldst_val;
      5'b01100:
        casez_tmp_278 = rob_uop_3_12_ldst_val;
      5'b01101:
        casez_tmp_278 = rob_uop_3_13_ldst_val;
      5'b01110:
        casez_tmp_278 = rob_uop_3_14_ldst_val;
      5'b01111:
        casez_tmp_278 = rob_uop_3_15_ldst_val;
      5'b10000:
        casez_tmp_278 = rob_uop_3_16_ldst_val;
      5'b10001:
        casez_tmp_278 = rob_uop_3_17_ldst_val;
      5'b10010:
        casez_tmp_278 = rob_uop_3_18_ldst_val;
      5'b10011:
        casez_tmp_278 = rob_uop_3_19_ldst_val;
      5'b10100:
        casez_tmp_278 = rob_uop_3_20_ldst_val;
      5'b10101:
        casez_tmp_278 = rob_uop_3_21_ldst_val;
      5'b10110:
        casez_tmp_278 = rob_uop_3_22_ldst_val;
      5'b10111:
        casez_tmp_278 = rob_uop_3_23_ldst_val;
      5'b11000:
        casez_tmp_278 = rob_uop_3_24_ldst_val;
      5'b11001:
        casez_tmp_278 = rob_uop_3_25_ldst_val;
      5'b11010:
        casez_tmp_278 = rob_uop_3_26_ldst_val;
      5'b11011:
        casez_tmp_278 = rob_uop_3_27_ldst_val;
      5'b11100:
        casez_tmp_278 = rob_uop_3_28_ldst_val;
      5'b11101:
        casez_tmp_278 = rob_uop_3_29_ldst_val;
      5'b11110:
        casez_tmp_278 = rob_uop_3_30_ldst_val;
      default:
        casez_tmp_278 = rob_uop_3_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_279;
  always @(*) begin
    casez (io_wb_resps_2_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_279 = rob_val_3_0;
      5'b00001:
        casez_tmp_279 = rob_val_3_1;
      5'b00010:
        casez_tmp_279 = rob_val_3_2;
      5'b00011:
        casez_tmp_279 = rob_val_3_3;
      5'b00100:
        casez_tmp_279 = rob_val_3_4;
      5'b00101:
        casez_tmp_279 = rob_val_3_5;
      5'b00110:
        casez_tmp_279 = rob_val_3_6;
      5'b00111:
        casez_tmp_279 = rob_val_3_7;
      5'b01000:
        casez_tmp_279 = rob_val_3_8;
      5'b01001:
        casez_tmp_279 = rob_val_3_9;
      5'b01010:
        casez_tmp_279 = rob_val_3_10;
      5'b01011:
        casez_tmp_279 = rob_val_3_11;
      5'b01100:
        casez_tmp_279 = rob_val_3_12;
      5'b01101:
        casez_tmp_279 = rob_val_3_13;
      5'b01110:
        casez_tmp_279 = rob_val_3_14;
      5'b01111:
        casez_tmp_279 = rob_val_3_15;
      5'b10000:
        casez_tmp_279 = rob_val_3_16;
      5'b10001:
        casez_tmp_279 = rob_val_3_17;
      5'b10010:
        casez_tmp_279 = rob_val_3_18;
      5'b10011:
        casez_tmp_279 = rob_val_3_19;
      5'b10100:
        casez_tmp_279 = rob_val_3_20;
      5'b10101:
        casez_tmp_279 = rob_val_3_21;
      5'b10110:
        casez_tmp_279 = rob_val_3_22;
      5'b10111:
        casez_tmp_279 = rob_val_3_23;
      5'b11000:
        casez_tmp_279 = rob_val_3_24;
      5'b11001:
        casez_tmp_279 = rob_val_3_25;
      5'b11010:
        casez_tmp_279 = rob_val_3_26;
      5'b11011:
        casez_tmp_279 = rob_val_3_27;
      5'b11100:
        casez_tmp_279 = rob_val_3_28;
      5'b11101:
        casez_tmp_279 = rob_val_3_29;
      5'b11110:
        casez_tmp_279 = rob_val_3_30;
      default:
        casez_tmp_279 = rob_val_3_31;
    endcase
  end // always @(*)
  reg         casez_tmp_280;
  always @(*) begin
    casez (io_wb_resps_2_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_280 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_280 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_280 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_280 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_280 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_280 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_280 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_280 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_280 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_280 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_280 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_280 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_280 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_280 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_280 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_280 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_280 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_280 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_280 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_280 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_280 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_280 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_280 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_280 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_280 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_280 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_280 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_280 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_280 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_280 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_280 = rob_bsy_3_30;
      default:
        casez_tmp_280 = rob_bsy_3_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_281;
  always @(*) begin
    casez (io_wb_resps_2_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_281 = rob_uop_3_0_pdst;
      5'b00001:
        casez_tmp_281 = rob_uop_3_1_pdst;
      5'b00010:
        casez_tmp_281 = rob_uop_3_2_pdst;
      5'b00011:
        casez_tmp_281 = rob_uop_3_3_pdst;
      5'b00100:
        casez_tmp_281 = rob_uop_3_4_pdst;
      5'b00101:
        casez_tmp_281 = rob_uop_3_5_pdst;
      5'b00110:
        casez_tmp_281 = rob_uop_3_6_pdst;
      5'b00111:
        casez_tmp_281 = rob_uop_3_7_pdst;
      5'b01000:
        casez_tmp_281 = rob_uop_3_8_pdst;
      5'b01001:
        casez_tmp_281 = rob_uop_3_9_pdst;
      5'b01010:
        casez_tmp_281 = rob_uop_3_10_pdst;
      5'b01011:
        casez_tmp_281 = rob_uop_3_11_pdst;
      5'b01100:
        casez_tmp_281 = rob_uop_3_12_pdst;
      5'b01101:
        casez_tmp_281 = rob_uop_3_13_pdst;
      5'b01110:
        casez_tmp_281 = rob_uop_3_14_pdst;
      5'b01111:
        casez_tmp_281 = rob_uop_3_15_pdst;
      5'b10000:
        casez_tmp_281 = rob_uop_3_16_pdst;
      5'b10001:
        casez_tmp_281 = rob_uop_3_17_pdst;
      5'b10010:
        casez_tmp_281 = rob_uop_3_18_pdst;
      5'b10011:
        casez_tmp_281 = rob_uop_3_19_pdst;
      5'b10100:
        casez_tmp_281 = rob_uop_3_20_pdst;
      5'b10101:
        casez_tmp_281 = rob_uop_3_21_pdst;
      5'b10110:
        casez_tmp_281 = rob_uop_3_22_pdst;
      5'b10111:
        casez_tmp_281 = rob_uop_3_23_pdst;
      5'b11000:
        casez_tmp_281 = rob_uop_3_24_pdst;
      5'b11001:
        casez_tmp_281 = rob_uop_3_25_pdst;
      5'b11010:
        casez_tmp_281 = rob_uop_3_26_pdst;
      5'b11011:
        casez_tmp_281 = rob_uop_3_27_pdst;
      5'b11100:
        casez_tmp_281 = rob_uop_3_28_pdst;
      5'b11101:
        casez_tmp_281 = rob_uop_3_29_pdst;
      5'b11110:
        casez_tmp_281 = rob_uop_3_30_pdst;
      default:
        casez_tmp_281 = rob_uop_3_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_282;
  always @(*) begin
    casez (io_wb_resps_2_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_282 = rob_uop_3_0_ldst_val;
      5'b00001:
        casez_tmp_282 = rob_uop_3_1_ldst_val;
      5'b00010:
        casez_tmp_282 = rob_uop_3_2_ldst_val;
      5'b00011:
        casez_tmp_282 = rob_uop_3_3_ldst_val;
      5'b00100:
        casez_tmp_282 = rob_uop_3_4_ldst_val;
      5'b00101:
        casez_tmp_282 = rob_uop_3_5_ldst_val;
      5'b00110:
        casez_tmp_282 = rob_uop_3_6_ldst_val;
      5'b00111:
        casez_tmp_282 = rob_uop_3_7_ldst_val;
      5'b01000:
        casez_tmp_282 = rob_uop_3_8_ldst_val;
      5'b01001:
        casez_tmp_282 = rob_uop_3_9_ldst_val;
      5'b01010:
        casez_tmp_282 = rob_uop_3_10_ldst_val;
      5'b01011:
        casez_tmp_282 = rob_uop_3_11_ldst_val;
      5'b01100:
        casez_tmp_282 = rob_uop_3_12_ldst_val;
      5'b01101:
        casez_tmp_282 = rob_uop_3_13_ldst_val;
      5'b01110:
        casez_tmp_282 = rob_uop_3_14_ldst_val;
      5'b01111:
        casez_tmp_282 = rob_uop_3_15_ldst_val;
      5'b10000:
        casez_tmp_282 = rob_uop_3_16_ldst_val;
      5'b10001:
        casez_tmp_282 = rob_uop_3_17_ldst_val;
      5'b10010:
        casez_tmp_282 = rob_uop_3_18_ldst_val;
      5'b10011:
        casez_tmp_282 = rob_uop_3_19_ldst_val;
      5'b10100:
        casez_tmp_282 = rob_uop_3_20_ldst_val;
      5'b10101:
        casez_tmp_282 = rob_uop_3_21_ldst_val;
      5'b10110:
        casez_tmp_282 = rob_uop_3_22_ldst_val;
      5'b10111:
        casez_tmp_282 = rob_uop_3_23_ldst_val;
      5'b11000:
        casez_tmp_282 = rob_uop_3_24_ldst_val;
      5'b11001:
        casez_tmp_282 = rob_uop_3_25_ldst_val;
      5'b11010:
        casez_tmp_282 = rob_uop_3_26_ldst_val;
      5'b11011:
        casez_tmp_282 = rob_uop_3_27_ldst_val;
      5'b11100:
        casez_tmp_282 = rob_uop_3_28_ldst_val;
      5'b11101:
        casez_tmp_282 = rob_uop_3_29_ldst_val;
      5'b11110:
        casez_tmp_282 = rob_uop_3_30_ldst_val;
      default:
        casez_tmp_282 = rob_uop_3_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_283;
  always @(*) begin
    casez (io_wb_resps_3_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_283 = rob_val_3_0;
      5'b00001:
        casez_tmp_283 = rob_val_3_1;
      5'b00010:
        casez_tmp_283 = rob_val_3_2;
      5'b00011:
        casez_tmp_283 = rob_val_3_3;
      5'b00100:
        casez_tmp_283 = rob_val_3_4;
      5'b00101:
        casez_tmp_283 = rob_val_3_5;
      5'b00110:
        casez_tmp_283 = rob_val_3_6;
      5'b00111:
        casez_tmp_283 = rob_val_3_7;
      5'b01000:
        casez_tmp_283 = rob_val_3_8;
      5'b01001:
        casez_tmp_283 = rob_val_3_9;
      5'b01010:
        casez_tmp_283 = rob_val_3_10;
      5'b01011:
        casez_tmp_283 = rob_val_3_11;
      5'b01100:
        casez_tmp_283 = rob_val_3_12;
      5'b01101:
        casez_tmp_283 = rob_val_3_13;
      5'b01110:
        casez_tmp_283 = rob_val_3_14;
      5'b01111:
        casez_tmp_283 = rob_val_3_15;
      5'b10000:
        casez_tmp_283 = rob_val_3_16;
      5'b10001:
        casez_tmp_283 = rob_val_3_17;
      5'b10010:
        casez_tmp_283 = rob_val_3_18;
      5'b10011:
        casez_tmp_283 = rob_val_3_19;
      5'b10100:
        casez_tmp_283 = rob_val_3_20;
      5'b10101:
        casez_tmp_283 = rob_val_3_21;
      5'b10110:
        casez_tmp_283 = rob_val_3_22;
      5'b10111:
        casez_tmp_283 = rob_val_3_23;
      5'b11000:
        casez_tmp_283 = rob_val_3_24;
      5'b11001:
        casez_tmp_283 = rob_val_3_25;
      5'b11010:
        casez_tmp_283 = rob_val_3_26;
      5'b11011:
        casez_tmp_283 = rob_val_3_27;
      5'b11100:
        casez_tmp_283 = rob_val_3_28;
      5'b11101:
        casez_tmp_283 = rob_val_3_29;
      5'b11110:
        casez_tmp_283 = rob_val_3_30;
      default:
        casez_tmp_283 = rob_val_3_31;
    endcase
  end // always @(*)
  reg         casez_tmp_284;
  always @(*) begin
    casez (io_wb_resps_3_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_284 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_284 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_284 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_284 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_284 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_284 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_284 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_284 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_284 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_284 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_284 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_284 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_284 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_284 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_284 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_284 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_284 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_284 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_284 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_284 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_284 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_284 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_284 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_284 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_284 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_284 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_284 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_284 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_284 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_284 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_284 = rob_bsy_3_30;
      default:
        casez_tmp_284 = rob_bsy_3_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_285;
  always @(*) begin
    casez (io_wb_resps_3_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_285 = rob_uop_3_0_pdst;
      5'b00001:
        casez_tmp_285 = rob_uop_3_1_pdst;
      5'b00010:
        casez_tmp_285 = rob_uop_3_2_pdst;
      5'b00011:
        casez_tmp_285 = rob_uop_3_3_pdst;
      5'b00100:
        casez_tmp_285 = rob_uop_3_4_pdst;
      5'b00101:
        casez_tmp_285 = rob_uop_3_5_pdst;
      5'b00110:
        casez_tmp_285 = rob_uop_3_6_pdst;
      5'b00111:
        casez_tmp_285 = rob_uop_3_7_pdst;
      5'b01000:
        casez_tmp_285 = rob_uop_3_8_pdst;
      5'b01001:
        casez_tmp_285 = rob_uop_3_9_pdst;
      5'b01010:
        casez_tmp_285 = rob_uop_3_10_pdst;
      5'b01011:
        casez_tmp_285 = rob_uop_3_11_pdst;
      5'b01100:
        casez_tmp_285 = rob_uop_3_12_pdst;
      5'b01101:
        casez_tmp_285 = rob_uop_3_13_pdst;
      5'b01110:
        casez_tmp_285 = rob_uop_3_14_pdst;
      5'b01111:
        casez_tmp_285 = rob_uop_3_15_pdst;
      5'b10000:
        casez_tmp_285 = rob_uop_3_16_pdst;
      5'b10001:
        casez_tmp_285 = rob_uop_3_17_pdst;
      5'b10010:
        casez_tmp_285 = rob_uop_3_18_pdst;
      5'b10011:
        casez_tmp_285 = rob_uop_3_19_pdst;
      5'b10100:
        casez_tmp_285 = rob_uop_3_20_pdst;
      5'b10101:
        casez_tmp_285 = rob_uop_3_21_pdst;
      5'b10110:
        casez_tmp_285 = rob_uop_3_22_pdst;
      5'b10111:
        casez_tmp_285 = rob_uop_3_23_pdst;
      5'b11000:
        casez_tmp_285 = rob_uop_3_24_pdst;
      5'b11001:
        casez_tmp_285 = rob_uop_3_25_pdst;
      5'b11010:
        casez_tmp_285 = rob_uop_3_26_pdst;
      5'b11011:
        casez_tmp_285 = rob_uop_3_27_pdst;
      5'b11100:
        casez_tmp_285 = rob_uop_3_28_pdst;
      5'b11101:
        casez_tmp_285 = rob_uop_3_29_pdst;
      5'b11110:
        casez_tmp_285 = rob_uop_3_30_pdst;
      default:
        casez_tmp_285 = rob_uop_3_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_286;
  always @(*) begin
    casez (io_wb_resps_3_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_286 = rob_uop_3_0_ldst_val;
      5'b00001:
        casez_tmp_286 = rob_uop_3_1_ldst_val;
      5'b00010:
        casez_tmp_286 = rob_uop_3_2_ldst_val;
      5'b00011:
        casez_tmp_286 = rob_uop_3_3_ldst_val;
      5'b00100:
        casez_tmp_286 = rob_uop_3_4_ldst_val;
      5'b00101:
        casez_tmp_286 = rob_uop_3_5_ldst_val;
      5'b00110:
        casez_tmp_286 = rob_uop_3_6_ldst_val;
      5'b00111:
        casez_tmp_286 = rob_uop_3_7_ldst_val;
      5'b01000:
        casez_tmp_286 = rob_uop_3_8_ldst_val;
      5'b01001:
        casez_tmp_286 = rob_uop_3_9_ldst_val;
      5'b01010:
        casez_tmp_286 = rob_uop_3_10_ldst_val;
      5'b01011:
        casez_tmp_286 = rob_uop_3_11_ldst_val;
      5'b01100:
        casez_tmp_286 = rob_uop_3_12_ldst_val;
      5'b01101:
        casez_tmp_286 = rob_uop_3_13_ldst_val;
      5'b01110:
        casez_tmp_286 = rob_uop_3_14_ldst_val;
      5'b01111:
        casez_tmp_286 = rob_uop_3_15_ldst_val;
      5'b10000:
        casez_tmp_286 = rob_uop_3_16_ldst_val;
      5'b10001:
        casez_tmp_286 = rob_uop_3_17_ldst_val;
      5'b10010:
        casez_tmp_286 = rob_uop_3_18_ldst_val;
      5'b10011:
        casez_tmp_286 = rob_uop_3_19_ldst_val;
      5'b10100:
        casez_tmp_286 = rob_uop_3_20_ldst_val;
      5'b10101:
        casez_tmp_286 = rob_uop_3_21_ldst_val;
      5'b10110:
        casez_tmp_286 = rob_uop_3_22_ldst_val;
      5'b10111:
        casez_tmp_286 = rob_uop_3_23_ldst_val;
      5'b11000:
        casez_tmp_286 = rob_uop_3_24_ldst_val;
      5'b11001:
        casez_tmp_286 = rob_uop_3_25_ldst_val;
      5'b11010:
        casez_tmp_286 = rob_uop_3_26_ldst_val;
      5'b11011:
        casez_tmp_286 = rob_uop_3_27_ldst_val;
      5'b11100:
        casez_tmp_286 = rob_uop_3_28_ldst_val;
      5'b11101:
        casez_tmp_286 = rob_uop_3_29_ldst_val;
      5'b11110:
        casez_tmp_286 = rob_uop_3_30_ldst_val;
      default:
        casez_tmp_286 = rob_uop_3_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_287;
  always @(*) begin
    casez (io_wb_resps_4_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_287 = rob_val_3_0;
      5'b00001:
        casez_tmp_287 = rob_val_3_1;
      5'b00010:
        casez_tmp_287 = rob_val_3_2;
      5'b00011:
        casez_tmp_287 = rob_val_3_3;
      5'b00100:
        casez_tmp_287 = rob_val_3_4;
      5'b00101:
        casez_tmp_287 = rob_val_3_5;
      5'b00110:
        casez_tmp_287 = rob_val_3_6;
      5'b00111:
        casez_tmp_287 = rob_val_3_7;
      5'b01000:
        casez_tmp_287 = rob_val_3_8;
      5'b01001:
        casez_tmp_287 = rob_val_3_9;
      5'b01010:
        casez_tmp_287 = rob_val_3_10;
      5'b01011:
        casez_tmp_287 = rob_val_3_11;
      5'b01100:
        casez_tmp_287 = rob_val_3_12;
      5'b01101:
        casez_tmp_287 = rob_val_3_13;
      5'b01110:
        casez_tmp_287 = rob_val_3_14;
      5'b01111:
        casez_tmp_287 = rob_val_3_15;
      5'b10000:
        casez_tmp_287 = rob_val_3_16;
      5'b10001:
        casez_tmp_287 = rob_val_3_17;
      5'b10010:
        casez_tmp_287 = rob_val_3_18;
      5'b10011:
        casez_tmp_287 = rob_val_3_19;
      5'b10100:
        casez_tmp_287 = rob_val_3_20;
      5'b10101:
        casez_tmp_287 = rob_val_3_21;
      5'b10110:
        casez_tmp_287 = rob_val_3_22;
      5'b10111:
        casez_tmp_287 = rob_val_3_23;
      5'b11000:
        casez_tmp_287 = rob_val_3_24;
      5'b11001:
        casez_tmp_287 = rob_val_3_25;
      5'b11010:
        casez_tmp_287 = rob_val_3_26;
      5'b11011:
        casez_tmp_287 = rob_val_3_27;
      5'b11100:
        casez_tmp_287 = rob_val_3_28;
      5'b11101:
        casez_tmp_287 = rob_val_3_29;
      5'b11110:
        casez_tmp_287 = rob_val_3_30;
      default:
        casez_tmp_287 = rob_val_3_31;
    endcase
  end // always @(*)
  reg         casez_tmp_288;
  always @(*) begin
    casez (io_wb_resps_4_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_288 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_288 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_288 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_288 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_288 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_288 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_288 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_288 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_288 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_288 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_288 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_288 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_288 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_288 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_288 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_288 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_288 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_288 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_288 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_288 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_288 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_288 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_288 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_288 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_288 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_288 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_288 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_288 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_288 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_288 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_288 = rob_bsy_3_30;
      default:
        casez_tmp_288 = rob_bsy_3_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_289;
  always @(*) begin
    casez (io_wb_resps_4_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_289 = rob_uop_3_0_pdst;
      5'b00001:
        casez_tmp_289 = rob_uop_3_1_pdst;
      5'b00010:
        casez_tmp_289 = rob_uop_3_2_pdst;
      5'b00011:
        casez_tmp_289 = rob_uop_3_3_pdst;
      5'b00100:
        casez_tmp_289 = rob_uop_3_4_pdst;
      5'b00101:
        casez_tmp_289 = rob_uop_3_5_pdst;
      5'b00110:
        casez_tmp_289 = rob_uop_3_6_pdst;
      5'b00111:
        casez_tmp_289 = rob_uop_3_7_pdst;
      5'b01000:
        casez_tmp_289 = rob_uop_3_8_pdst;
      5'b01001:
        casez_tmp_289 = rob_uop_3_9_pdst;
      5'b01010:
        casez_tmp_289 = rob_uop_3_10_pdst;
      5'b01011:
        casez_tmp_289 = rob_uop_3_11_pdst;
      5'b01100:
        casez_tmp_289 = rob_uop_3_12_pdst;
      5'b01101:
        casez_tmp_289 = rob_uop_3_13_pdst;
      5'b01110:
        casez_tmp_289 = rob_uop_3_14_pdst;
      5'b01111:
        casez_tmp_289 = rob_uop_3_15_pdst;
      5'b10000:
        casez_tmp_289 = rob_uop_3_16_pdst;
      5'b10001:
        casez_tmp_289 = rob_uop_3_17_pdst;
      5'b10010:
        casez_tmp_289 = rob_uop_3_18_pdst;
      5'b10011:
        casez_tmp_289 = rob_uop_3_19_pdst;
      5'b10100:
        casez_tmp_289 = rob_uop_3_20_pdst;
      5'b10101:
        casez_tmp_289 = rob_uop_3_21_pdst;
      5'b10110:
        casez_tmp_289 = rob_uop_3_22_pdst;
      5'b10111:
        casez_tmp_289 = rob_uop_3_23_pdst;
      5'b11000:
        casez_tmp_289 = rob_uop_3_24_pdst;
      5'b11001:
        casez_tmp_289 = rob_uop_3_25_pdst;
      5'b11010:
        casez_tmp_289 = rob_uop_3_26_pdst;
      5'b11011:
        casez_tmp_289 = rob_uop_3_27_pdst;
      5'b11100:
        casez_tmp_289 = rob_uop_3_28_pdst;
      5'b11101:
        casez_tmp_289 = rob_uop_3_29_pdst;
      5'b11110:
        casez_tmp_289 = rob_uop_3_30_pdst;
      default:
        casez_tmp_289 = rob_uop_3_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_290;
  always @(*) begin
    casez (io_wb_resps_4_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_290 = rob_uop_3_0_ldst_val;
      5'b00001:
        casez_tmp_290 = rob_uop_3_1_ldst_val;
      5'b00010:
        casez_tmp_290 = rob_uop_3_2_ldst_val;
      5'b00011:
        casez_tmp_290 = rob_uop_3_3_ldst_val;
      5'b00100:
        casez_tmp_290 = rob_uop_3_4_ldst_val;
      5'b00101:
        casez_tmp_290 = rob_uop_3_5_ldst_val;
      5'b00110:
        casez_tmp_290 = rob_uop_3_6_ldst_val;
      5'b00111:
        casez_tmp_290 = rob_uop_3_7_ldst_val;
      5'b01000:
        casez_tmp_290 = rob_uop_3_8_ldst_val;
      5'b01001:
        casez_tmp_290 = rob_uop_3_9_ldst_val;
      5'b01010:
        casez_tmp_290 = rob_uop_3_10_ldst_val;
      5'b01011:
        casez_tmp_290 = rob_uop_3_11_ldst_val;
      5'b01100:
        casez_tmp_290 = rob_uop_3_12_ldst_val;
      5'b01101:
        casez_tmp_290 = rob_uop_3_13_ldst_val;
      5'b01110:
        casez_tmp_290 = rob_uop_3_14_ldst_val;
      5'b01111:
        casez_tmp_290 = rob_uop_3_15_ldst_val;
      5'b10000:
        casez_tmp_290 = rob_uop_3_16_ldst_val;
      5'b10001:
        casez_tmp_290 = rob_uop_3_17_ldst_val;
      5'b10010:
        casez_tmp_290 = rob_uop_3_18_ldst_val;
      5'b10011:
        casez_tmp_290 = rob_uop_3_19_ldst_val;
      5'b10100:
        casez_tmp_290 = rob_uop_3_20_ldst_val;
      5'b10101:
        casez_tmp_290 = rob_uop_3_21_ldst_val;
      5'b10110:
        casez_tmp_290 = rob_uop_3_22_ldst_val;
      5'b10111:
        casez_tmp_290 = rob_uop_3_23_ldst_val;
      5'b11000:
        casez_tmp_290 = rob_uop_3_24_ldst_val;
      5'b11001:
        casez_tmp_290 = rob_uop_3_25_ldst_val;
      5'b11010:
        casez_tmp_290 = rob_uop_3_26_ldst_val;
      5'b11011:
        casez_tmp_290 = rob_uop_3_27_ldst_val;
      5'b11100:
        casez_tmp_290 = rob_uop_3_28_ldst_val;
      5'b11101:
        casez_tmp_290 = rob_uop_3_29_ldst_val;
      5'b11110:
        casez_tmp_290 = rob_uop_3_30_ldst_val;
      default:
        casez_tmp_290 = rob_uop_3_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_291;
  always @(*) begin
    casez (io_wb_resps_5_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_291 = rob_val_3_0;
      5'b00001:
        casez_tmp_291 = rob_val_3_1;
      5'b00010:
        casez_tmp_291 = rob_val_3_2;
      5'b00011:
        casez_tmp_291 = rob_val_3_3;
      5'b00100:
        casez_tmp_291 = rob_val_3_4;
      5'b00101:
        casez_tmp_291 = rob_val_3_5;
      5'b00110:
        casez_tmp_291 = rob_val_3_6;
      5'b00111:
        casez_tmp_291 = rob_val_3_7;
      5'b01000:
        casez_tmp_291 = rob_val_3_8;
      5'b01001:
        casez_tmp_291 = rob_val_3_9;
      5'b01010:
        casez_tmp_291 = rob_val_3_10;
      5'b01011:
        casez_tmp_291 = rob_val_3_11;
      5'b01100:
        casez_tmp_291 = rob_val_3_12;
      5'b01101:
        casez_tmp_291 = rob_val_3_13;
      5'b01110:
        casez_tmp_291 = rob_val_3_14;
      5'b01111:
        casez_tmp_291 = rob_val_3_15;
      5'b10000:
        casez_tmp_291 = rob_val_3_16;
      5'b10001:
        casez_tmp_291 = rob_val_3_17;
      5'b10010:
        casez_tmp_291 = rob_val_3_18;
      5'b10011:
        casez_tmp_291 = rob_val_3_19;
      5'b10100:
        casez_tmp_291 = rob_val_3_20;
      5'b10101:
        casez_tmp_291 = rob_val_3_21;
      5'b10110:
        casez_tmp_291 = rob_val_3_22;
      5'b10111:
        casez_tmp_291 = rob_val_3_23;
      5'b11000:
        casez_tmp_291 = rob_val_3_24;
      5'b11001:
        casez_tmp_291 = rob_val_3_25;
      5'b11010:
        casez_tmp_291 = rob_val_3_26;
      5'b11011:
        casez_tmp_291 = rob_val_3_27;
      5'b11100:
        casez_tmp_291 = rob_val_3_28;
      5'b11101:
        casez_tmp_291 = rob_val_3_29;
      5'b11110:
        casez_tmp_291 = rob_val_3_30;
      default:
        casez_tmp_291 = rob_val_3_31;
    endcase
  end // always @(*)
  reg         casez_tmp_292;
  always @(*) begin
    casez (io_wb_resps_5_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_292 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_292 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_292 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_292 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_292 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_292 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_292 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_292 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_292 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_292 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_292 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_292 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_292 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_292 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_292 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_292 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_292 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_292 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_292 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_292 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_292 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_292 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_292 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_292 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_292 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_292 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_292 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_292 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_292 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_292 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_292 = rob_bsy_3_30;
      default:
        casez_tmp_292 = rob_bsy_3_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_293;
  always @(*) begin
    casez (io_wb_resps_5_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_293 = rob_uop_3_0_pdst;
      5'b00001:
        casez_tmp_293 = rob_uop_3_1_pdst;
      5'b00010:
        casez_tmp_293 = rob_uop_3_2_pdst;
      5'b00011:
        casez_tmp_293 = rob_uop_3_3_pdst;
      5'b00100:
        casez_tmp_293 = rob_uop_3_4_pdst;
      5'b00101:
        casez_tmp_293 = rob_uop_3_5_pdst;
      5'b00110:
        casez_tmp_293 = rob_uop_3_6_pdst;
      5'b00111:
        casez_tmp_293 = rob_uop_3_7_pdst;
      5'b01000:
        casez_tmp_293 = rob_uop_3_8_pdst;
      5'b01001:
        casez_tmp_293 = rob_uop_3_9_pdst;
      5'b01010:
        casez_tmp_293 = rob_uop_3_10_pdst;
      5'b01011:
        casez_tmp_293 = rob_uop_3_11_pdst;
      5'b01100:
        casez_tmp_293 = rob_uop_3_12_pdst;
      5'b01101:
        casez_tmp_293 = rob_uop_3_13_pdst;
      5'b01110:
        casez_tmp_293 = rob_uop_3_14_pdst;
      5'b01111:
        casez_tmp_293 = rob_uop_3_15_pdst;
      5'b10000:
        casez_tmp_293 = rob_uop_3_16_pdst;
      5'b10001:
        casez_tmp_293 = rob_uop_3_17_pdst;
      5'b10010:
        casez_tmp_293 = rob_uop_3_18_pdst;
      5'b10011:
        casez_tmp_293 = rob_uop_3_19_pdst;
      5'b10100:
        casez_tmp_293 = rob_uop_3_20_pdst;
      5'b10101:
        casez_tmp_293 = rob_uop_3_21_pdst;
      5'b10110:
        casez_tmp_293 = rob_uop_3_22_pdst;
      5'b10111:
        casez_tmp_293 = rob_uop_3_23_pdst;
      5'b11000:
        casez_tmp_293 = rob_uop_3_24_pdst;
      5'b11001:
        casez_tmp_293 = rob_uop_3_25_pdst;
      5'b11010:
        casez_tmp_293 = rob_uop_3_26_pdst;
      5'b11011:
        casez_tmp_293 = rob_uop_3_27_pdst;
      5'b11100:
        casez_tmp_293 = rob_uop_3_28_pdst;
      5'b11101:
        casez_tmp_293 = rob_uop_3_29_pdst;
      5'b11110:
        casez_tmp_293 = rob_uop_3_30_pdst;
      default:
        casez_tmp_293 = rob_uop_3_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_294;
  always @(*) begin
    casez (io_wb_resps_5_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_294 = rob_uop_3_0_ldst_val;
      5'b00001:
        casez_tmp_294 = rob_uop_3_1_ldst_val;
      5'b00010:
        casez_tmp_294 = rob_uop_3_2_ldst_val;
      5'b00011:
        casez_tmp_294 = rob_uop_3_3_ldst_val;
      5'b00100:
        casez_tmp_294 = rob_uop_3_4_ldst_val;
      5'b00101:
        casez_tmp_294 = rob_uop_3_5_ldst_val;
      5'b00110:
        casez_tmp_294 = rob_uop_3_6_ldst_val;
      5'b00111:
        casez_tmp_294 = rob_uop_3_7_ldst_val;
      5'b01000:
        casez_tmp_294 = rob_uop_3_8_ldst_val;
      5'b01001:
        casez_tmp_294 = rob_uop_3_9_ldst_val;
      5'b01010:
        casez_tmp_294 = rob_uop_3_10_ldst_val;
      5'b01011:
        casez_tmp_294 = rob_uop_3_11_ldst_val;
      5'b01100:
        casez_tmp_294 = rob_uop_3_12_ldst_val;
      5'b01101:
        casez_tmp_294 = rob_uop_3_13_ldst_val;
      5'b01110:
        casez_tmp_294 = rob_uop_3_14_ldst_val;
      5'b01111:
        casez_tmp_294 = rob_uop_3_15_ldst_val;
      5'b10000:
        casez_tmp_294 = rob_uop_3_16_ldst_val;
      5'b10001:
        casez_tmp_294 = rob_uop_3_17_ldst_val;
      5'b10010:
        casez_tmp_294 = rob_uop_3_18_ldst_val;
      5'b10011:
        casez_tmp_294 = rob_uop_3_19_ldst_val;
      5'b10100:
        casez_tmp_294 = rob_uop_3_20_ldst_val;
      5'b10101:
        casez_tmp_294 = rob_uop_3_21_ldst_val;
      5'b10110:
        casez_tmp_294 = rob_uop_3_22_ldst_val;
      5'b10111:
        casez_tmp_294 = rob_uop_3_23_ldst_val;
      5'b11000:
        casez_tmp_294 = rob_uop_3_24_ldst_val;
      5'b11001:
        casez_tmp_294 = rob_uop_3_25_ldst_val;
      5'b11010:
        casez_tmp_294 = rob_uop_3_26_ldst_val;
      5'b11011:
        casez_tmp_294 = rob_uop_3_27_ldst_val;
      5'b11100:
        casez_tmp_294 = rob_uop_3_28_ldst_val;
      5'b11101:
        casez_tmp_294 = rob_uop_3_29_ldst_val;
      5'b11110:
        casez_tmp_294 = rob_uop_3_30_ldst_val;
      default:
        casez_tmp_294 = rob_uop_3_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_295;
  always @(*) begin
    casez (io_wb_resps_6_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_295 = rob_val_3_0;
      5'b00001:
        casez_tmp_295 = rob_val_3_1;
      5'b00010:
        casez_tmp_295 = rob_val_3_2;
      5'b00011:
        casez_tmp_295 = rob_val_3_3;
      5'b00100:
        casez_tmp_295 = rob_val_3_4;
      5'b00101:
        casez_tmp_295 = rob_val_3_5;
      5'b00110:
        casez_tmp_295 = rob_val_3_6;
      5'b00111:
        casez_tmp_295 = rob_val_3_7;
      5'b01000:
        casez_tmp_295 = rob_val_3_8;
      5'b01001:
        casez_tmp_295 = rob_val_3_9;
      5'b01010:
        casez_tmp_295 = rob_val_3_10;
      5'b01011:
        casez_tmp_295 = rob_val_3_11;
      5'b01100:
        casez_tmp_295 = rob_val_3_12;
      5'b01101:
        casez_tmp_295 = rob_val_3_13;
      5'b01110:
        casez_tmp_295 = rob_val_3_14;
      5'b01111:
        casez_tmp_295 = rob_val_3_15;
      5'b10000:
        casez_tmp_295 = rob_val_3_16;
      5'b10001:
        casez_tmp_295 = rob_val_3_17;
      5'b10010:
        casez_tmp_295 = rob_val_3_18;
      5'b10011:
        casez_tmp_295 = rob_val_3_19;
      5'b10100:
        casez_tmp_295 = rob_val_3_20;
      5'b10101:
        casez_tmp_295 = rob_val_3_21;
      5'b10110:
        casez_tmp_295 = rob_val_3_22;
      5'b10111:
        casez_tmp_295 = rob_val_3_23;
      5'b11000:
        casez_tmp_295 = rob_val_3_24;
      5'b11001:
        casez_tmp_295 = rob_val_3_25;
      5'b11010:
        casez_tmp_295 = rob_val_3_26;
      5'b11011:
        casez_tmp_295 = rob_val_3_27;
      5'b11100:
        casez_tmp_295 = rob_val_3_28;
      5'b11101:
        casez_tmp_295 = rob_val_3_29;
      5'b11110:
        casez_tmp_295 = rob_val_3_30;
      default:
        casez_tmp_295 = rob_val_3_31;
    endcase
  end // always @(*)
  reg         casez_tmp_296;
  always @(*) begin
    casez (io_wb_resps_6_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_296 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_296 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_296 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_296 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_296 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_296 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_296 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_296 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_296 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_296 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_296 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_296 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_296 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_296 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_296 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_296 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_296 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_296 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_296 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_296 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_296 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_296 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_296 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_296 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_296 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_296 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_296 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_296 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_296 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_296 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_296 = rob_bsy_3_30;
      default:
        casez_tmp_296 = rob_bsy_3_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_297;
  always @(*) begin
    casez (io_wb_resps_6_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_297 = rob_uop_3_0_pdst;
      5'b00001:
        casez_tmp_297 = rob_uop_3_1_pdst;
      5'b00010:
        casez_tmp_297 = rob_uop_3_2_pdst;
      5'b00011:
        casez_tmp_297 = rob_uop_3_3_pdst;
      5'b00100:
        casez_tmp_297 = rob_uop_3_4_pdst;
      5'b00101:
        casez_tmp_297 = rob_uop_3_5_pdst;
      5'b00110:
        casez_tmp_297 = rob_uop_3_6_pdst;
      5'b00111:
        casez_tmp_297 = rob_uop_3_7_pdst;
      5'b01000:
        casez_tmp_297 = rob_uop_3_8_pdst;
      5'b01001:
        casez_tmp_297 = rob_uop_3_9_pdst;
      5'b01010:
        casez_tmp_297 = rob_uop_3_10_pdst;
      5'b01011:
        casez_tmp_297 = rob_uop_3_11_pdst;
      5'b01100:
        casez_tmp_297 = rob_uop_3_12_pdst;
      5'b01101:
        casez_tmp_297 = rob_uop_3_13_pdst;
      5'b01110:
        casez_tmp_297 = rob_uop_3_14_pdst;
      5'b01111:
        casez_tmp_297 = rob_uop_3_15_pdst;
      5'b10000:
        casez_tmp_297 = rob_uop_3_16_pdst;
      5'b10001:
        casez_tmp_297 = rob_uop_3_17_pdst;
      5'b10010:
        casez_tmp_297 = rob_uop_3_18_pdst;
      5'b10011:
        casez_tmp_297 = rob_uop_3_19_pdst;
      5'b10100:
        casez_tmp_297 = rob_uop_3_20_pdst;
      5'b10101:
        casez_tmp_297 = rob_uop_3_21_pdst;
      5'b10110:
        casez_tmp_297 = rob_uop_3_22_pdst;
      5'b10111:
        casez_tmp_297 = rob_uop_3_23_pdst;
      5'b11000:
        casez_tmp_297 = rob_uop_3_24_pdst;
      5'b11001:
        casez_tmp_297 = rob_uop_3_25_pdst;
      5'b11010:
        casez_tmp_297 = rob_uop_3_26_pdst;
      5'b11011:
        casez_tmp_297 = rob_uop_3_27_pdst;
      5'b11100:
        casez_tmp_297 = rob_uop_3_28_pdst;
      5'b11101:
        casez_tmp_297 = rob_uop_3_29_pdst;
      5'b11110:
        casez_tmp_297 = rob_uop_3_30_pdst;
      default:
        casez_tmp_297 = rob_uop_3_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_298;
  always @(*) begin
    casez (io_wb_resps_6_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_298 = rob_uop_3_0_ldst_val;
      5'b00001:
        casez_tmp_298 = rob_uop_3_1_ldst_val;
      5'b00010:
        casez_tmp_298 = rob_uop_3_2_ldst_val;
      5'b00011:
        casez_tmp_298 = rob_uop_3_3_ldst_val;
      5'b00100:
        casez_tmp_298 = rob_uop_3_4_ldst_val;
      5'b00101:
        casez_tmp_298 = rob_uop_3_5_ldst_val;
      5'b00110:
        casez_tmp_298 = rob_uop_3_6_ldst_val;
      5'b00111:
        casez_tmp_298 = rob_uop_3_7_ldst_val;
      5'b01000:
        casez_tmp_298 = rob_uop_3_8_ldst_val;
      5'b01001:
        casez_tmp_298 = rob_uop_3_9_ldst_val;
      5'b01010:
        casez_tmp_298 = rob_uop_3_10_ldst_val;
      5'b01011:
        casez_tmp_298 = rob_uop_3_11_ldst_val;
      5'b01100:
        casez_tmp_298 = rob_uop_3_12_ldst_val;
      5'b01101:
        casez_tmp_298 = rob_uop_3_13_ldst_val;
      5'b01110:
        casez_tmp_298 = rob_uop_3_14_ldst_val;
      5'b01111:
        casez_tmp_298 = rob_uop_3_15_ldst_val;
      5'b10000:
        casez_tmp_298 = rob_uop_3_16_ldst_val;
      5'b10001:
        casez_tmp_298 = rob_uop_3_17_ldst_val;
      5'b10010:
        casez_tmp_298 = rob_uop_3_18_ldst_val;
      5'b10011:
        casez_tmp_298 = rob_uop_3_19_ldst_val;
      5'b10100:
        casez_tmp_298 = rob_uop_3_20_ldst_val;
      5'b10101:
        casez_tmp_298 = rob_uop_3_21_ldst_val;
      5'b10110:
        casez_tmp_298 = rob_uop_3_22_ldst_val;
      5'b10111:
        casez_tmp_298 = rob_uop_3_23_ldst_val;
      5'b11000:
        casez_tmp_298 = rob_uop_3_24_ldst_val;
      5'b11001:
        casez_tmp_298 = rob_uop_3_25_ldst_val;
      5'b11010:
        casez_tmp_298 = rob_uop_3_26_ldst_val;
      5'b11011:
        casez_tmp_298 = rob_uop_3_27_ldst_val;
      5'b11100:
        casez_tmp_298 = rob_uop_3_28_ldst_val;
      5'b11101:
        casez_tmp_298 = rob_uop_3_29_ldst_val;
      5'b11110:
        casez_tmp_298 = rob_uop_3_30_ldst_val;
      default:
        casez_tmp_298 = rob_uop_3_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_299;
  always @(*) begin
    casez (io_wb_resps_7_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_299 = rob_val_3_0;
      5'b00001:
        casez_tmp_299 = rob_val_3_1;
      5'b00010:
        casez_tmp_299 = rob_val_3_2;
      5'b00011:
        casez_tmp_299 = rob_val_3_3;
      5'b00100:
        casez_tmp_299 = rob_val_3_4;
      5'b00101:
        casez_tmp_299 = rob_val_3_5;
      5'b00110:
        casez_tmp_299 = rob_val_3_6;
      5'b00111:
        casez_tmp_299 = rob_val_3_7;
      5'b01000:
        casez_tmp_299 = rob_val_3_8;
      5'b01001:
        casez_tmp_299 = rob_val_3_9;
      5'b01010:
        casez_tmp_299 = rob_val_3_10;
      5'b01011:
        casez_tmp_299 = rob_val_3_11;
      5'b01100:
        casez_tmp_299 = rob_val_3_12;
      5'b01101:
        casez_tmp_299 = rob_val_3_13;
      5'b01110:
        casez_tmp_299 = rob_val_3_14;
      5'b01111:
        casez_tmp_299 = rob_val_3_15;
      5'b10000:
        casez_tmp_299 = rob_val_3_16;
      5'b10001:
        casez_tmp_299 = rob_val_3_17;
      5'b10010:
        casez_tmp_299 = rob_val_3_18;
      5'b10011:
        casez_tmp_299 = rob_val_3_19;
      5'b10100:
        casez_tmp_299 = rob_val_3_20;
      5'b10101:
        casez_tmp_299 = rob_val_3_21;
      5'b10110:
        casez_tmp_299 = rob_val_3_22;
      5'b10111:
        casez_tmp_299 = rob_val_3_23;
      5'b11000:
        casez_tmp_299 = rob_val_3_24;
      5'b11001:
        casez_tmp_299 = rob_val_3_25;
      5'b11010:
        casez_tmp_299 = rob_val_3_26;
      5'b11011:
        casez_tmp_299 = rob_val_3_27;
      5'b11100:
        casez_tmp_299 = rob_val_3_28;
      5'b11101:
        casez_tmp_299 = rob_val_3_29;
      5'b11110:
        casez_tmp_299 = rob_val_3_30;
      default:
        casez_tmp_299 = rob_val_3_31;
    endcase
  end // always @(*)
  reg         casez_tmp_300;
  always @(*) begin
    casez (io_wb_resps_7_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_300 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_300 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_300 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_300 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_300 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_300 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_300 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_300 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_300 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_300 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_300 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_300 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_300 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_300 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_300 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_300 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_300 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_300 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_300 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_300 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_300 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_300 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_300 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_300 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_300 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_300 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_300 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_300 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_300 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_300 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_300 = rob_bsy_3_30;
      default:
        casez_tmp_300 = rob_bsy_3_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_301;
  always @(*) begin
    casez (io_wb_resps_7_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_301 = rob_uop_3_0_pdst;
      5'b00001:
        casez_tmp_301 = rob_uop_3_1_pdst;
      5'b00010:
        casez_tmp_301 = rob_uop_3_2_pdst;
      5'b00011:
        casez_tmp_301 = rob_uop_3_3_pdst;
      5'b00100:
        casez_tmp_301 = rob_uop_3_4_pdst;
      5'b00101:
        casez_tmp_301 = rob_uop_3_5_pdst;
      5'b00110:
        casez_tmp_301 = rob_uop_3_6_pdst;
      5'b00111:
        casez_tmp_301 = rob_uop_3_7_pdst;
      5'b01000:
        casez_tmp_301 = rob_uop_3_8_pdst;
      5'b01001:
        casez_tmp_301 = rob_uop_3_9_pdst;
      5'b01010:
        casez_tmp_301 = rob_uop_3_10_pdst;
      5'b01011:
        casez_tmp_301 = rob_uop_3_11_pdst;
      5'b01100:
        casez_tmp_301 = rob_uop_3_12_pdst;
      5'b01101:
        casez_tmp_301 = rob_uop_3_13_pdst;
      5'b01110:
        casez_tmp_301 = rob_uop_3_14_pdst;
      5'b01111:
        casez_tmp_301 = rob_uop_3_15_pdst;
      5'b10000:
        casez_tmp_301 = rob_uop_3_16_pdst;
      5'b10001:
        casez_tmp_301 = rob_uop_3_17_pdst;
      5'b10010:
        casez_tmp_301 = rob_uop_3_18_pdst;
      5'b10011:
        casez_tmp_301 = rob_uop_3_19_pdst;
      5'b10100:
        casez_tmp_301 = rob_uop_3_20_pdst;
      5'b10101:
        casez_tmp_301 = rob_uop_3_21_pdst;
      5'b10110:
        casez_tmp_301 = rob_uop_3_22_pdst;
      5'b10111:
        casez_tmp_301 = rob_uop_3_23_pdst;
      5'b11000:
        casez_tmp_301 = rob_uop_3_24_pdst;
      5'b11001:
        casez_tmp_301 = rob_uop_3_25_pdst;
      5'b11010:
        casez_tmp_301 = rob_uop_3_26_pdst;
      5'b11011:
        casez_tmp_301 = rob_uop_3_27_pdst;
      5'b11100:
        casez_tmp_301 = rob_uop_3_28_pdst;
      5'b11101:
        casez_tmp_301 = rob_uop_3_29_pdst;
      5'b11110:
        casez_tmp_301 = rob_uop_3_30_pdst;
      default:
        casez_tmp_301 = rob_uop_3_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_302;
  always @(*) begin
    casez (io_wb_resps_7_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_302 = rob_uop_3_0_ldst_val;
      5'b00001:
        casez_tmp_302 = rob_uop_3_1_ldst_val;
      5'b00010:
        casez_tmp_302 = rob_uop_3_2_ldst_val;
      5'b00011:
        casez_tmp_302 = rob_uop_3_3_ldst_val;
      5'b00100:
        casez_tmp_302 = rob_uop_3_4_ldst_val;
      5'b00101:
        casez_tmp_302 = rob_uop_3_5_ldst_val;
      5'b00110:
        casez_tmp_302 = rob_uop_3_6_ldst_val;
      5'b00111:
        casez_tmp_302 = rob_uop_3_7_ldst_val;
      5'b01000:
        casez_tmp_302 = rob_uop_3_8_ldst_val;
      5'b01001:
        casez_tmp_302 = rob_uop_3_9_ldst_val;
      5'b01010:
        casez_tmp_302 = rob_uop_3_10_ldst_val;
      5'b01011:
        casez_tmp_302 = rob_uop_3_11_ldst_val;
      5'b01100:
        casez_tmp_302 = rob_uop_3_12_ldst_val;
      5'b01101:
        casez_tmp_302 = rob_uop_3_13_ldst_val;
      5'b01110:
        casez_tmp_302 = rob_uop_3_14_ldst_val;
      5'b01111:
        casez_tmp_302 = rob_uop_3_15_ldst_val;
      5'b10000:
        casez_tmp_302 = rob_uop_3_16_ldst_val;
      5'b10001:
        casez_tmp_302 = rob_uop_3_17_ldst_val;
      5'b10010:
        casez_tmp_302 = rob_uop_3_18_ldst_val;
      5'b10011:
        casez_tmp_302 = rob_uop_3_19_ldst_val;
      5'b10100:
        casez_tmp_302 = rob_uop_3_20_ldst_val;
      5'b10101:
        casez_tmp_302 = rob_uop_3_21_ldst_val;
      5'b10110:
        casez_tmp_302 = rob_uop_3_22_ldst_val;
      5'b10111:
        casez_tmp_302 = rob_uop_3_23_ldst_val;
      5'b11000:
        casez_tmp_302 = rob_uop_3_24_ldst_val;
      5'b11001:
        casez_tmp_302 = rob_uop_3_25_ldst_val;
      5'b11010:
        casez_tmp_302 = rob_uop_3_26_ldst_val;
      5'b11011:
        casez_tmp_302 = rob_uop_3_27_ldst_val;
      5'b11100:
        casez_tmp_302 = rob_uop_3_28_ldst_val;
      5'b11101:
        casez_tmp_302 = rob_uop_3_29_ldst_val;
      5'b11110:
        casez_tmp_302 = rob_uop_3_30_ldst_val;
      default:
        casez_tmp_302 = rob_uop_3_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_303;
  always @(*) begin
    casez (io_wb_resps_8_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_303 = rob_val_3_0;
      5'b00001:
        casez_tmp_303 = rob_val_3_1;
      5'b00010:
        casez_tmp_303 = rob_val_3_2;
      5'b00011:
        casez_tmp_303 = rob_val_3_3;
      5'b00100:
        casez_tmp_303 = rob_val_3_4;
      5'b00101:
        casez_tmp_303 = rob_val_3_5;
      5'b00110:
        casez_tmp_303 = rob_val_3_6;
      5'b00111:
        casez_tmp_303 = rob_val_3_7;
      5'b01000:
        casez_tmp_303 = rob_val_3_8;
      5'b01001:
        casez_tmp_303 = rob_val_3_9;
      5'b01010:
        casez_tmp_303 = rob_val_3_10;
      5'b01011:
        casez_tmp_303 = rob_val_3_11;
      5'b01100:
        casez_tmp_303 = rob_val_3_12;
      5'b01101:
        casez_tmp_303 = rob_val_3_13;
      5'b01110:
        casez_tmp_303 = rob_val_3_14;
      5'b01111:
        casez_tmp_303 = rob_val_3_15;
      5'b10000:
        casez_tmp_303 = rob_val_3_16;
      5'b10001:
        casez_tmp_303 = rob_val_3_17;
      5'b10010:
        casez_tmp_303 = rob_val_3_18;
      5'b10011:
        casez_tmp_303 = rob_val_3_19;
      5'b10100:
        casez_tmp_303 = rob_val_3_20;
      5'b10101:
        casez_tmp_303 = rob_val_3_21;
      5'b10110:
        casez_tmp_303 = rob_val_3_22;
      5'b10111:
        casez_tmp_303 = rob_val_3_23;
      5'b11000:
        casez_tmp_303 = rob_val_3_24;
      5'b11001:
        casez_tmp_303 = rob_val_3_25;
      5'b11010:
        casez_tmp_303 = rob_val_3_26;
      5'b11011:
        casez_tmp_303 = rob_val_3_27;
      5'b11100:
        casez_tmp_303 = rob_val_3_28;
      5'b11101:
        casez_tmp_303 = rob_val_3_29;
      5'b11110:
        casez_tmp_303 = rob_val_3_30;
      default:
        casez_tmp_303 = rob_val_3_31;
    endcase
  end // always @(*)
  reg         casez_tmp_304;
  always @(*) begin
    casez (io_wb_resps_8_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_304 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_304 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_304 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_304 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_304 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_304 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_304 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_304 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_304 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_304 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_304 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_304 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_304 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_304 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_304 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_304 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_304 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_304 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_304 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_304 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_304 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_304 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_304 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_304 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_304 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_304 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_304 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_304 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_304 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_304 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_304 = rob_bsy_3_30;
      default:
        casez_tmp_304 = rob_bsy_3_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_305;
  always @(*) begin
    casez (io_wb_resps_8_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_305 = rob_uop_3_0_pdst;
      5'b00001:
        casez_tmp_305 = rob_uop_3_1_pdst;
      5'b00010:
        casez_tmp_305 = rob_uop_3_2_pdst;
      5'b00011:
        casez_tmp_305 = rob_uop_3_3_pdst;
      5'b00100:
        casez_tmp_305 = rob_uop_3_4_pdst;
      5'b00101:
        casez_tmp_305 = rob_uop_3_5_pdst;
      5'b00110:
        casez_tmp_305 = rob_uop_3_6_pdst;
      5'b00111:
        casez_tmp_305 = rob_uop_3_7_pdst;
      5'b01000:
        casez_tmp_305 = rob_uop_3_8_pdst;
      5'b01001:
        casez_tmp_305 = rob_uop_3_9_pdst;
      5'b01010:
        casez_tmp_305 = rob_uop_3_10_pdst;
      5'b01011:
        casez_tmp_305 = rob_uop_3_11_pdst;
      5'b01100:
        casez_tmp_305 = rob_uop_3_12_pdst;
      5'b01101:
        casez_tmp_305 = rob_uop_3_13_pdst;
      5'b01110:
        casez_tmp_305 = rob_uop_3_14_pdst;
      5'b01111:
        casez_tmp_305 = rob_uop_3_15_pdst;
      5'b10000:
        casez_tmp_305 = rob_uop_3_16_pdst;
      5'b10001:
        casez_tmp_305 = rob_uop_3_17_pdst;
      5'b10010:
        casez_tmp_305 = rob_uop_3_18_pdst;
      5'b10011:
        casez_tmp_305 = rob_uop_3_19_pdst;
      5'b10100:
        casez_tmp_305 = rob_uop_3_20_pdst;
      5'b10101:
        casez_tmp_305 = rob_uop_3_21_pdst;
      5'b10110:
        casez_tmp_305 = rob_uop_3_22_pdst;
      5'b10111:
        casez_tmp_305 = rob_uop_3_23_pdst;
      5'b11000:
        casez_tmp_305 = rob_uop_3_24_pdst;
      5'b11001:
        casez_tmp_305 = rob_uop_3_25_pdst;
      5'b11010:
        casez_tmp_305 = rob_uop_3_26_pdst;
      5'b11011:
        casez_tmp_305 = rob_uop_3_27_pdst;
      5'b11100:
        casez_tmp_305 = rob_uop_3_28_pdst;
      5'b11101:
        casez_tmp_305 = rob_uop_3_29_pdst;
      5'b11110:
        casez_tmp_305 = rob_uop_3_30_pdst;
      default:
        casez_tmp_305 = rob_uop_3_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_306;
  always @(*) begin
    casez (io_wb_resps_8_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_306 = rob_uop_3_0_ldst_val;
      5'b00001:
        casez_tmp_306 = rob_uop_3_1_ldst_val;
      5'b00010:
        casez_tmp_306 = rob_uop_3_2_ldst_val;
      5'b00011:
        casez_tmp_306 = rob_uop_3_3_ldst_val;
      5'b00100:
        casez_tmp_306 = rob_uop_3_4_ldst_val;
      5'b00101:
        casez_tmp_306 = rob_uop_3_5_ldst_val;
      5'b00110:
        casez_tmp_306 = rob_uop_3_6_ldst_val;
      5'b00111:
        casez_tmp_306 = rob_uop_3_7_ldst_val;
      5'b01000:
        casez_tmp_306 = rob_uop_3_8_ldst_val;
      5'b01001:
        casez_tmp_306 = rob_uop_3_9_ldst_val;
      5'b01010:
        casez_tmp_306 = rob_uop_3_10_ldst_val;
      5'b01011:
        casez_tmp_306 = rob_uop_3_11_ldst_val;
      5'b01100:
        casez_tmp_306 = rob_uop_3_12_ldst_val;
      5'b01101:
        casez_tmp_306 = rob_uop_3_13_ldst_val;
      5'b01110:
        casez_tmp_306 = rob_uop_3_14_ldst_val;
      5'b01111:
        casez_tmp_306 = rob_uop_3_15_ldst_val;
      5'b10000:
        casez_tmp_306 = rob_uop_3_16_ldst_val;
      5'b10001:
        casez_tmp_306 = rob_uop_3_17_ldst_val;
      5'b10010:
        casez_tmp_306 = rob_uop_3_18_ldst_val;
      5'b10011:
        casez_tmp_306 = rob_uop_3_19_ldst_val;
      5'b10100:
        casez_tmp_306 = rob_uop_3_20_ldst_val;
      5'b10101:
        casez_tmp_306 = rob_uop_3_21_ldst_val;
      5'b10110:
        casez_tmp_306 = rob_uop_3_22_ldst_val;
      5'b10111:
        casez_tmp_306 = rob_uop_3_23_ldst_val;
      5'b11000:
        casez_tmp_306 = rob_uop_3_24_ldst_val;
      5'b11001:
        casez_tmp_306 = rob_uop_3_25_ldst_val;
      5'b11010:
        casez_tmp_306 = rob_uop_3_26_ldst_val;
      5'b11011:
        casez_tmp_306 = rob_uop_3_27_ldst_val;
      5'b11100:
        casez_tmp_306 = rob_uop_3_28_ldst_val;
      5'b11101:
        casez_tmp_306 = rob_uop_3_29_ldst_val;
      5'b11110:
        casez_tmp_306 = rob_uop_3_30_ldst_val;
      default:
        casez_tmp_306 = rob_uop_3_31_ldst_val;
    endcase
  end // always @(*)
  reg         casez_tmp_307;
  always @(*) begin
    casez (io_wb_resps_9_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_307 = rob_val_3_0;
      5'b00001:
        casez_tmp_307 = rob_val_3_1;
      5'b00010:
        casez_tmp_307 = rob_val_3_2;
      5'b00011:
        casez_tmp_307 = rob_val_3_3;
      5'b00100:
        casez_tmp_307 = rob_val_3_4;
      5'b00101:
        casez_tmp_307 = rob_val_3_5;
      5'b00110:
        casez_tmp_307 = rob_val_3_6;
      5'b00111:
        casez_tmp_307 = rob_val_3_7;
      5'b01000:
        casez_tmp_307 = rob_val_3_8;
      5'b01001:
        casez_tmp_307 = rob_val_3_9;
      5'b01010:
        casez_tmp_307 = rob_val_3_10;
      5'b01011:
        casez_tmp_307 = rob_val_3_11;
      5'b01100:
        casez_tmp_307 = rob_val_3_12;
      5'b01101:
        casez_tmp_307 = rob_val_3_13;
      5'b01110:
        casez_tmp_307 = rob_val_3_14;
      5'b01111:
        casez_tmp_307 = rob_val_3_15;
      5'b10000:
        casez_tmp_307 = rob_val_3_16;
      5'b10001:
        casez_tmp_307 = rob_val_3_17;
      5'b10010:
        casez_tmp_307 = rob_val_3_18;
      5'b10011:
        casez_tmp_307 = rob_val_3_19;
      5'b10100:
        casez_tmp_307 = rob_val_3_20;
      5'b10101:
        casez_tmp_307 = rob_val_3_21;
      5'b10110:
        casez_tmp_307 = rob_val_3_22;
      5'b10111:
        casez_tmp_307 = rob_val_3_23;
      5'b11000:
        casez_tmp_307 = rob_val_3_24;
      5'b11001:
        casez_tmp_307 = rob_val_3_25;
      5'b11010:
        casez_tmp_307 = rob_val_3_26;
      5'b11011:
        casez_tmp_307 = rob_val_3_27;
      5'b11100:
        casez_tmp_307 = rob_val_3_28;
      5'b11101:
        casez_tmp_307 = rob_val_3_29;
      5'b11110:
        casez_tmp_307 = rob_val_3_30;
      default:
        casez_tmp_307 = rob_val_3_31;
    endcase
  end // always @(*)
  reg         casez_tmp_308;
  always @(*) begin
    casez (io_wb_resps_9_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_308 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_308 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_308 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_308 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_308 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_308 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_308 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_308 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_308 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_308 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_308 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_308 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_308 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_308 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_308 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_308 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_308 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_308 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_308 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_308 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_308 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_308 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_308 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_308 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_308 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_308 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_308 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_308 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_308 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_308 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_308 = rob_bsy_3_30;
      default:
        casez_tmp_308 = rob_bsy_3_31;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_309;
  always @(*) begin
    casez (io_wb_resps_9_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_309 = rob_uop_3_0_pdst;
      5'b00001:
        casez_tmp_309 = rob_uop_3_1_pdst;
      5'b00010:
        casez_tmp_309 = rob_uop_3_2_pdst;
      5'b00011:
        casez_tmp_309 = rob_uop_3_3_pdst;
      5'b00100:
        casez_tmp_309 = rob_uop_3_4_pdst;
      5'b00101:
        casez_tmp_309 = rob_uop_3_5_pdst;
      5'b00110:
        casez_tmp_309 = rob_uop_3_6_pdst;
      5'b00111:
        casez_tmp_309 = rob_uop_3_7_pdst;
      5'b01000:
        casez_tmp_309 = rob_uop_3_8_pdst;
      5'b01001:
        casez_tmp_309 = rob_uop_3_9_pdst;
      5'b01010:
        casez_tmp_309 = rob_uop_3_10_pdst;
      5'b01011:
        casez_tmp_309 = rob_uop_3_11_pdst;
      5'b01100:
        casez_tmp_309 = rob_uop_3_12_pdst;
      5'b01101:
        casez_tmp_309 = rob_uop_3_13_pdst;
      5'b01110:
        casez_tmp_309 = rob_uop_3_14_pdst;
      5'b01111:
        casez_tmp_309 = rob_uop_3_15_pdst;
      5'b10000:
        casez_tmp_309 = rob_uop_3_16_pdst;
      5'b10001:
        casez_tmp_309 = rob_uop_3_17_pdst;
      5'b10010:
        casez_tmp_309 = rob_uop_3_18_pdst;
      5'b10011:
        casez_tmp_309 = rob_uop_3_19_pdst;
      5'b10100:
        casez_tmp_309 = rob_uop_3_20_pdst;
      5'b10101:
        casez_tmp_309 = rob_uop_3_21_pdst;
      5'b10110:
        casez_tmp_309 = rob_uop_3_22_pdst;
      5'b10111:
        casez_tmp_309 = rob_uop_3_23_pdst;
      5'b11000:
        casez_tmp_309 = rob_uop_3_24_pdst;
      5'b11001:
        casez_tmp_309 = rob_uop_3_25_pdst;
      5'b11010:
        casez_tmp_309 = rob_uop_3_26_pdst;
      5'b11011:
        casez_tmp_309 = rob_uop_3_27_pdst;
      5'b11100:
        casez_tmp_309 = rob_uop_3_28_pdst;
      5'b11101:
        casez_tmp_309 = rob_uop_3_29_pdst;
      5'b11110:
        casez_tmp_309 = rob_uop_3_30_pdst;
      default:
        casez_tmp_309 = rob_uop_3_31_pdst;
    endcase
  end // always @(*)
  reg         casez_tmp_310;
  always @(*) begin
    casez (io_wb_resps_9_bits_uop_rob_idx[6:2])
      5'b00000:
        casez_tmp_310 = rob_uop_3_0_ldst_val;
      5'b00001:
        casez_tmp_310 = rob_uop_3_1_ldst_val;
      5'b00010:
        casez_tmp_310 = rob_uop_3_2_ldst_val;
      5'b00011:
        casez_tmp_310 = rob_uop_3_3_ldst_val;
      5'b00100:
        casez_tmp_310 = rob_uop_3_4_ldst_val;
      5'b00101:
        casez_tmp_310 = rob_uop_3_5_ldst_val;
      5'b00110:
        casez_tmp_310 = rob_uop_3_6_ldst_val;
      5'b00111:
        casez_tmp_310 = rob_uop_3_7_ldst_val;
      5'b01000:
        casez_tmp_310 = rob_uop_3_8_ldst_val;
      5'b01001:
        casez_tmp_310 = rob_uop_3_9_ldst_val;
      5'b01010:
        casez_tmp_310 = rob_uop_3_10_ldst_val;
      5'b01011:
        casez_tmp_310 = rob_uop_3_11_ldst_val;
      5'b01100:
        casez_tmp_310 = rob_uop_3_12_ldst_val;
      5'b01101:
        casez_tmp_310 = rob_uop_3_13_ldst_val;
      5'b01110:
        casez_tmp_310 = rob_uop_3_14_ldst_val;
      5'b01111:
        casez_tmp_310 = rob_uop_3_15_ldst_val;
      5'b10000:
        casez_tmp_310 = rob_uop_3_16_ldst_val;
      5'b10001:
        casez_tmp_310 = rob_uop_3_17_ldst_val;
      5'b10010:
        casez_tmp_310 = rob_uop_3_18_ldst_val;
      5'b10011:
        casez_tmp_310 = rob_uop_3_19_ldst_val;
      5'b10100:
        casez_tmp_310 = rob_uop_3_20_ldst_val;
      5'b10101:
        casez_tmp_310 = rob_uop_3_21_ldst_val;
      5'b10110:
        casez_tmp_310 = rob_uop_3_22_ldst_val;
      5'b10111:
        casez_tmp_310 = rob_uop_3_23_ldst_val;
      5'b11000:
        casez_tmp_310 = rob_uop_3_24_ldst_val;
      5'b11001:
        casez_tmp_310 = rob_uop_3_25_ldst_val;
      5'b11010:
        casez_tmp_310 = rob_uop_3_26_ldst_val;
      5'b11011:
        casez_tmp_310 = rob_uop_3_27_ldst_val;
      5'b11100:
        casez_tmp_310 = rob_uop_3_28_ldst_val;
      5'b11101:
        casez_tmp_310 = rob_uop_3_29_ldst_val;
      5'b11110:
        casez_tmp_310 = rob_uop_3_30_ldst_val;
      default:
        casez_tmp_310 = rob_uop_3_31_ldst_val;
    endcase
  end // always @(*)
  reg         block_commit_REG;
  reg         block_commit_REG_1;
  reg         block_commit_REG_2;
  wire        block_commit = rob_state != 2'h1 & rob_state != 2'h3 | block_commit_REG | block_commit_REG_2;
  assign will_commit_0 = can_commit_0 & ~can_throw_exception_0 & ~block_commit;
  wire        _GEN_65 = casez_tmp_7 & (~can_commit_0 | can_throw_exception_0) | block_commit;
  assign will_commit_1 = can_commit_1 & ~can_throw_exception_1 & ~_GEN_65;
  wire        _GEN_66 = casez_tmp_85 & (~can_commit_1 | can_throw_exception_1) | _GEN_65;
  assign will_commit_2 = can_commit_2 & ~can_throw_exception_2 & ~_GEN_66;
  wire        _GEN_67 = casez_tmp_163 & (~can_commit_2 | can_throw_exception_2) | _GEN_66;
  wire        exception_thrown = can_throw_exception_3 & ~_GEN_67 & ~will_commit_2 | can_throw_exception_2 & ~_GEN_66 & ~will_commit_1 | can_throw_exception_1 & ~_GEN_65 & ~will_commit_0 | can_throw_exception_0 & ~block_commit;
  assign will_commit_3 = casez_tmp_241 & ~casez_tmp_243 & ~io_csr_stall & ~can_throw_exception_3 & ~_GEN_67;
  wire        is_mini_exception = r_xcpt_uop_exc_cause == 64'h10 | r_xcpt_uop_exc_cause == 64'h11;
  wire [5:0]  com_xcpt_uop_ftq_idx = casez_tmp_7 ? casez_tmp_16 : casez_tmp_85 ? casez_tmp_94 : casez_tmp_163 ? casez_tmp_172 : casez_tmp_250;
  wire        com_xcpt_uop_edge_inst = casez_tmp_7 ? casez_tmp_17 : casez_tmp_85 ? casez_tmp_95 : casez_tmp_163 ? casez_tmp_173 : casez_tmp_251;
  wire [5:0]  com_xcpt_uop_pc_lob = casez_tmp_7 ? casez_tmp_18 : casez_tmp_85 ? casez_tmp_96 : casez_tmp_163 ? casez_tmp_174 : casez_tmp_252;
  wire        flush_commit_mask_0 = will_commit_0 & casez_tmp_25;
  wire        flush_commit_mask_1 = will_commit_1 & casez_tmp_103;
  wire        flush_commit_mask_2 = will_commit_2 & casez_tmp_181;
  wire        flush_commit_mask_3 = will_commit_3 & casez_tmp_259;
  wire        flush_commit = flush_commit_mask_0 | flush_commit_mask_1 | flush_commit_mask_2 | flush_commit_mask_3;
  wire        _io_flush_valid_output = exception_thrown | flush_commit;
  wire        _fflags_val_0_T = will_commit_0 & casez_tmp_29;
  wire        fflags_val_0 = _fflags_val_0_T & ~casez_tmp_23;
  wire        _fflags_val_1_T = will_commit_1 & casez_tmp_107;
  wire        fflags_val_1 = _fflags_val_1_T & ~casez_tmp_101;
  wire        _fflags_val_2_T = will_commit_2 & casez_tmp_185;
  wire        fflags_val_2 = _fflags_val_2_T & ~casez_tmp_179;
  wire        _fflags_val_3_T = will_commit_3 & casez_tmp_263;
  wire        fflags_val_3 = _fflags_val_3_T & ~casez_tmp_257;
  wire        enq_xcpts_0 = io_enq_valids_0 & io_enq_uops_0_exception;
  wire        enq_xcpts_1 = io_enq_valids_1 & io_enq_uops_1_exception;
  wire        enq_xcpts_2 = io_enq_valids_2 & io_enq_uops_2_exception;
  wire [1:0]  idx = enq_xcpts_0 ? 2'h0 : enq_xcpts_1 ? 2'h1 : {1'h1, ~enq_xcpts_2};
  reg  [19:0] casez_tmp_311;
  always @(*) begin
    casez (idx)
      2'b00:
        casez_tmp_311 = io_enq_uops_0_br_mask;
      2'b01:
        casez_tmp_311 = io_enq_uops_1_br_mask;
      2'b10:
        casez_tmp_311 = io_enq_uops_2_br_mask;
      default:
        casez_tmp_311 = io_enq_uops_3_br_mask;
    endcase
  end // always @(*)
  reg  [5:0]  casez_tmp_312;
  always @(*) begin
    casez (idx)
      2'b00:
        casez_tmp_312 = io_enq_uops_0_pc_lob;
      2'b01:
        casez_tmp_312 = io_enq_uops_1_pc_lob;
      2'b10:
        casez_tmp_312 = io_enq_uops_2_pc_lob;
      default:
        casez_tmp_312 = io_enq_uops_3_pc_lob;
    endcase
  end // always @(*)
  reg  [6:0]  casez_tmp_313;
  always @(*) begin
    casez (idx)
      2'b00:
        casez_tmp_313 = io_enq_uops_0_rob_idx;
      2'b01:
        casez_tmp_313 = io_enq_uops_1_rob_idx;
      2'b10:
        casez_tmp_313 = io_enq_uops_2_rob_idx;
      default:
        casez_tmp_313 = io_enq_uops_3_rob_idx;
    endcase
  end // always @(*)
  reg  [63:0] casez_tmp_314;
  always @(*) begin
    casez (idx)
      2'b00:
        casez_tmp_314 = io_enq_uops_0_exc_cause;
      2'b01:
        casez_tmp_314 = io_enq_uops_1_exc_cause;
      2'b10:
        casez_tmp_314 = io_enq_uops_2_exc_cause;
      default:
        casez_tmp_314 = io_enq_uops_3_exc_cause;
    endcase
  end // always @(*)
  reg         r_partial_row;
  wire        _empty_T = rob_head == rob_tail;
  wire        finished_committing_row = (|{will_commit_3, will_commit_2, will_commit_1, will_commit_0}) & ({will_commit_3, will_commit_2, will_commit_1, will_commit_0} ^ {casez_tmp_241, casez_tmp_163, casez_tmp_85, casez_tmp_7}) == 4'h0 & ~(r_partial_row & _empty_T & ~maybe_full);
  reg         pnr_maybe_at_tail;
  wire        _io_ready_T = rob_state == 2'h1;
  `ifndef SYNTHESIS
    wire [6:0] rob_pnr_idx = {rob_pnr, rob_pnr_lsb};
    wire       _GEN_68 = io_enq_valids_0 & ~reset;
    wire       _GEN_69 = _GEN_9 & ~reset;
    wire       _GEN_70 = _GEN_10 & ~reset;
    wire       _GEN_71 = _GEN_11 & ~reset;
    wire       _GEN_72 = ~reset & (will_commit_0 | will_commit_1 | will_commit_2 | will_commit_3) & (_io_commit_rbk_valids_0_output | _io_commit_rbk_valids_1_output | _io_commit_rbk_valids_2_output | _io_commit_rbk_valids_3_output);
    wire       _GEN_73 = io_enq_valids_1 & ~reset;
    wire       _GEN_74 = _GEN_27 & ~reset;
    wire       _GEN_75 = _GEN_28 & ~reset;
    wire       _GEN_76 = _GEN_29 & ~reset;
    wire       _GEN_77 = io_enq_valids_2 & ~reset;
    wire       _GEN_78 = _GEN_43 & ~reset;
    wire       _GEN_79 = _GEN_44 & ~reset;
    wire       _GEN_80 = _GEN_45 & ~reset;
    wire       _GEN_81 = io_enq_valids_3 & ~reset;
    wire       _GEN_82 = _GEN_59 & ~reset;
    wire       _GEN_83 = _GEN_60 & ~reset;
    wire       _GEN_84 = _GEN_61 & ~reset;
    wire       _GEN_85 = rob_pnr_idx < rob_head_idx;
    wire [2:0] _GEN_86 = {1'h0, {1'h0, flush_commit_mask_0} + {1'h0, flush_commit_mask_1}} + {1'h0, {1'h0, flush_commit_mask_2} + {1'h0, flush_commit_mask_3}};
    always @(posedge clock) begin
      if (_GEN_68 & casez_tmp) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] overwriting a valid entry.\n    at rob.scala:333 assert (rob_val(rob_tail) === false.B, \"[rob] overwriting a valid entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_68 & io_enq_uops_0_rob_idx[6:2] != rob_tail) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at rob.scala:334 assert ((io.enq_uops(w).rob_idx >> log2Ceil(coreWidth)) === rob_tail)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_69 & ~casez_tmp_0) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_69 & ~casez_tmp_1) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_70 & ~casez_tmp_2) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_70 & ~casez_tmp_3) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_71 & ~casez_tmp_4) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_71 & ~casez_tmp_5) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_14 & ~casez_tmp_6) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: An instruction marked as safe is causing an exception\n    at rob.scala:394 assert(rob_unsafe(GetRowIdx(io.lxcpt.bits.uop.rob_idx)),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_72) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: com_valids and rbk_valids are mutually exclusive\n    at rob.scala:434 assert (!(io.commit.valids.reduce(_||_) && io.commit.rbk_valids.reduce(_||_)),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN & ~casez_tmp_37) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (0) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN & ~casez_tmp_38) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (0) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN & casez_tmp_40 & casez_tmp_39 != io_wb_resps_0_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (0) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_0 & ~casez_tmp_41) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (1) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_0 & ~casez_tmp_42) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (1) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_0 & casez_tmp_44 & casez_tmp_43 != io_wb_resps_1_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (1) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_1 & ~casez_tmp_45) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (2) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_1 & ~casez_tmp_46) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (2) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_1 & casez_tmp_48 & casez_tmp_47 != io_wb_resps_2_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (2) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_2 & ~casez_tmp_49) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (3) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_2 & ~casez_tmp_50) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (3) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_2 & casez_tmp_52 & casez_tmp_51 != io_wb_resps_3_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (3) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_3 & ~casez_tmp_53) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (4) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_3 & ~casez_tmp_54) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (4) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_3 & casez_tmp_56 & casez_tmp_55 != io_wb_resps_4_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (4) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_4 & ~casez_tmp_57) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (5) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_4 & ~casez_tmp_58) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (5) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_4 & casez_tmp_60 & casez_tmp_59 != io_wb_resps_5_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (5) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_5 & ~casez_tmp_61) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (6) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_5 & ~casez_tmp_62) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (6) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_5 & casez_tmp_64 & casez_tmp_63 != io_wb_resps_6_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (6) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_6 & ~casez_tmp_65) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (7) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_6 & ~casez_tmp_66) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (7) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_6 & casez_tmp_68 & casez_tmp_67 != io_wb_resps_7_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (7) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_7 & ~casez_tmp_69) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (8) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_7 & ~casez_tmp_70) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (8) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_7 & casez_tmp_72 & casez_tmp_71 != io_wb_resps_8_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (8) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_8 & ~casez_tmp_73) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (9) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_8 & ~casez_tmp_74) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (9) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_8 & casez_tmp_76 & casez_tmp_75 != io_wb_resps_9_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (9) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_73 & casez_tmp_77) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] overwriting a valid entry.\n    at rob.scala:333 assert (rob_val(rob_tail) === false.B, \"[rob] overwriting a valid entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_73 & io_enq_uops_1_rob_idx[6:2] != rob_tail) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at rob.scala:334 assert ((io.enq_uops(w).rob_idx >> log2Ceil(coreWidth)) === rob_tail)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_74 & ~casez_tmp_78) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_74 & ~casez_tmp_79) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_75 & ~casez_tmp_80) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_75 & ~casez_tmp_81) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_76 & ~casez_tmp_82) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_76 & ~casez_tmp_83) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_31 & ~casez_tmp_84) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: An instruction marked as safe is causing an exception\n    at rob.scala:394 assert(rob_unsafe(GetRowIdx(io.lxcpt.bits.uop.rob_idx)),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_72) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: com_valids and rbk_valids are mutually exclusive\n    at rob.scala:434 assert (!(io.commit.valids.reduce(_||_) && io.commit.rbk_valids.reduce(_||_)),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_17 & ~casez_tmp_115) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (0) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_17 & ~casez_tmp_116) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (0) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_17 & casez_tmp_118 & casez_tmp_117 != io_wb_resps_0_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (0) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_18 & ~casez_tmp_119) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (1) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_18 & ~casez_tmp_120) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (1) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_18 & casez_tmp_122 & casez_tmp_121 != io_wb_resps_1_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (1) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_19 & ~casez_tmp_123) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (2) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_19 & ~casez_tmp_124) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (2) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_19 & casez_tmp_126 & casez_tmp_125 != io_wb_resps_2_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (2) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_20 & ~casez_tmp_127) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (3) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_20 & ~casez_tmp_128) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (3) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_20 & casez_tmp_130 & casez_tmp_129 != io_wb_resps_3_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (3) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_21 & ~casez_tmp_131) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (4) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_21 & ~casez_tmp_132) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (4) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_21 & casez_tmp_134 & casez_tmp_133 != io_wb_resps_4_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (4) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_22 & ~casez_tmp_135) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (5) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_22 & ~casez_tmp_136) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (5) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_22 & casez_tmp_138 & casez_tmp_137 != io_wb_resps_5_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (5) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_23 & ~casez_tmp_139) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (6) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_23 & ~casez_tmp_140) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (6) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_23 & casez_tmp_142 & casez_tmp_141 != io_wb_resps_6_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (6) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_24 & ~casez_tmp_143) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (7) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_24 & ~casez_tmp_144) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (7) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_24 & casez_tmp_146 & casez_tmp_145 != io_wb_resps_7_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (7) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_25 & ~casez_tmp_147) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (8) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_25 & ~casez_tmp_148) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (8) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_25 & casez_tmp_150 & casez_tmp_149 != io_wb_resps_8_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (8) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_26 & ~casez_tmp_151) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (9) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_26 & ~casez_tmp_152) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (9) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_26 & casez_tmp_154 & casez_tmp_153 != io_wb_resps_9_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (9) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_77 & casez_tmp_155) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] overwriting a valid entry.\n    at rob.scala:333 assert (rob_val(rob_tail) === false.B, \"[rob] overwriting a valid entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_77 & io_enq_uops_2_rob_idx[6:2] != rob_tail) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at rob.scala:334 assert ((io.enq_uops(w).rob_idx >> log2Ceil(coreWidth)) === rob_tail)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_78 & ~casez_tmp_156) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_78 & ~casez_tmp_157) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_79 & ~casez_tmp_158) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_79 & ~casez_tmp_159) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_80 & ~casez_tmp_160) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_80 & ~casez_tmp_161) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_47 & ~casez_tmp_162) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: An instruction marked as safe is causing an exception\n    at rob.scala:394 assert(rob_unsafe(GetRowIdx(io.lxcpt.bits.uop.rob_idx)),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_72) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: com_valids and rbk_valids are mutually exclusive\n    at rob.scala:434 assert (!(io.commit.valids.reduce(_||_) && io.commit.rbk_valids.reduce(_||_)),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_33 & ~casez_tmp_193) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (0) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_33 & ~casez_tmp_194) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (0) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_33 & casez_tmp_196 & casez_tmp_195 != io_wb_resps_0_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (0) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_34 & ~casez_tmp_197) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (1) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_34 & ~casez_tmp_198) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (1) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_34 & casez_tmp_200 & casez_tmp_199 != io_wb_resps_1_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (1) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_35 & ~casez_tmp_201) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (2) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_35 & ~casez_tmp_202) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (2) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_35 & casez_tmp_204 & casez_tmp_203 != io_wb_resps_2_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (2) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_36 & ~casez_tmp_205) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (3) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_36 & ~casez_tmp_206) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (3) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_36 & casez_tmp_208 & casez_tmp_207 != io_wb_resps_3_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (3) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_37 & ~casez_tmp_209) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (4) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_37 & ~casez_tmp_210) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (4) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_37 & casez_tmp_212 & casez_tmp_211 != io_wb_resps_4_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (4) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_38 & ~casez_tmp_213) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (5) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_38 & ~casez_tmp_214) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (5) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_38 & casez_tmp_216 & casez_tmp_215 != io_wb_resps_5_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (5) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_39 & ~casez_tmp_217) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (6) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_39 & ~casez_tmp_218) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (6) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_39 & casez_tmp_220 & casez_tmp_219 != io_wb_resps_6_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (6) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_40 & ~casez_tmp_221) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (7) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_40 & ~casez_tmp_222) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (7) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_40 & casez_tmp_224 & casez_tmp_223 != io_wb_resps_7_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (7) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_41 & ~casez_tmp_225) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (8) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_41 & ~casez_tmp_226) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (8) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_41 & casez_tmp_228 & casez_tmp_227 != io_wb_resps_8_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (8) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_42 & ~casez_tmp_229) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (9) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_42 & ~casez_tmp_230) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (9) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_42 & casez_tmp_232 & casez_tmp_231 != io_wb_resps_9_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (9) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_81 & casez_tmp_233) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] overwriting a valid entry.\n    at rob.scala:333 assert (rob_val(rob_tail) === false.B, \"[rob] overwriting a valid entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_81 & io_enq_uops_3_rob_idx[6:2] != rob_tail) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at rob.scala:334 assert ((io.enq_uops(w).rob_idx >> log2Ceil(coreWidth)) === rob_tail)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_82 & ~casez_tmp_234) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_82 & ~casez_tmp_235) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_83 & ~casez_tmp_236) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_83 & ~casez_tmp_237) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_84 & ~casez_tmp_238) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_84 & ~casez_tmp_239) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_63 & ~casez_tmp_240) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: An instruction marked as safe is causing an exception\n    at rob.scala:394 assert(rob_unsafe(GetRowIdx(io.lxcpt.bits.uop.rob_idx)),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (_GEN_72) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: com_valids and rbk_valids are mutually exclusive\n    at rob.scala:434 assert (!(io.commit.valids.reduce(_||_) && io.commit.rbk_valids.reduce(_||_)),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_49 & ~casez_tmp_271) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (0) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_49 & ~casez_tmp_272) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (0) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_49 & casez_tmp_274 & casez_tmp_273 != io_wb_resps_0_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (0) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_50 & ~casez_tmp_275) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (1) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_50 & ~casez_tmp_276) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (1) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_50 & casez_tmp_278 & casez_tmp_277 != io_wb_resps_1_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (1) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_51 & ~casez_tmp_279) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (2) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_51 & ~casez_tmp_280) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (2) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_51 & casez_tmp_282 & casez_tmp_281 != io_wb_resps_2_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (2) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_52 & ~casez_tmp_283) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (3) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_52 & ~casez_tmp_284) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (3) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_52 & casez_tmp_286 & casez_tmp_285 != io_wb_resps_3_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (3) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_53 & ~casez_tmp_287) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (4) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_53 & ~casez_tmp_288) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (4) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_53 & casez_tmp_290 & casez_tmp_289 != io_wb_resps_4_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (4) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_54 & ~casez_tmp_291) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (5) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_54 & ~casez_tmp_292) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (5) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_54 & casez_tmp_294 & casez_tmp_293 != io_wb_resps_5_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (5) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_55 & ~casez_tmp_295) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (6) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_55 & ~casez_tmp_296) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (6) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_55 & casez_tmp_298 & casez_tmp_297 != io_wb_resps_6_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (6) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_56 & ~casez_tmp_299) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (7) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_56 & ~casez_tmp_300) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (7) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_56 & casez_tmp_302 & casez_tmp_301 != io_wb_resps_7_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (7) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_57 & ~casez_tmp_303) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (8) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_57 & ~casez_tmp_304) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (8) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_57 & casez_tmp_306 & casez_tmp_305 != io_wb_resps_8_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (8) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_58 & ~casez_tmp_307) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (9) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_58 & ~casez_tmp_308) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (9) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _GEN_58 & casez_tmp_310 & casez_tmp_309 != io_wb_resps_9_bits_uop_pdst) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] writeback (9) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & (|(_GEN_86[2:1]))) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: [rob] Can't commit multiple flush_on_commit instructions on one cycle\n    at rob.scala:580 assert(!(PopCount(flush_commit_mask) > 1.U),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & will_commit_0 & ~casez_tmp_29 & (|casez_tmp_32)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Committed non-FP instruction has non-zero fflag bits.\n    at rob.scala:613 assert (!(io.commit.valids(w) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _fflags_val_0_T & (casez_tmp_22 | casez_tmp_23) & (|casez_tmp_32)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Committed FP load or store has non-zero fflag bits.\n    at rob.scala:617 assert (!(io.commit.valids(w) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & will_commit_1 & ~casez_tmp_107 & (|casez_tmp_110)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Committed non-FP instruction has non-zero fflag bits.\n    at rob.scala:613 assert (!(io.commit.valids(w) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _fflags_val_1_T & (casez_tmp_100 | casez_tmp_101) & (|casez_tmp_110)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Committed FP load or store has non-zero fflag bits.\n    at rob.scala:617 assert (!(io.commit.valids(w) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & will_commit_2 & ~casez_tmp_185 & (|casez_tmp_188)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Committed non-FP instruction has non-zero fflag bits.\n    at rob.scala:613 assert (!(io.commit.valids(w) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _fflags_val_2_T & (casez_tmp_178 | casez_tmp_179) & (|casez_tmp_188)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Committed FP load or store has non-zero fflag bits.\n    at rob.scala:617 assert (!(io.commit.valids(w) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & will_commit_3 & ~casez_tmp_263 & (|casez_tmp_266)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Committed non-FP instruction has non-zero fflag bits.\n    at rob.scala:613 assert (!(io.commit.valids(w) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & _fflags_val_3_T & (casez_tmp_256 | casez_tmp_257) & (|casez_tmp_266)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: Committed FP load or store has non-zero fflag bits.\n    at rob.scala:617 assert (!(io.commit.valids(w) &&\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & exception_thrown & ~r_xcpt_val) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: ROB trying to throw an exception, but it doesn't have a valid xcpt_cause\n    at rob.scala:667 assert (!(exception_thrown && !r_xcpt_val),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & empty & r_xcpt_val) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: ROB is empty, but believes it has an outstanding exception.\n    at rob.scala:670 assert (!(empty && r_xcpt_val),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & exception_thrown & r_xcpt_uop_rob_idx[6:2] != rob_head) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed: ROB is throwing an exception, but the stored exception information's rob_idx does not match the rob_head\n    at rob.scala:673 assert (!(will_throw_exception && (GetRowIdx(r_xcpt_uop.rob_idx) =/= rob_head)),\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & ~(_GEN_85 ^ rob_head_idx < rob_tail_idx ^ rob_pnr_idx >= rob_tail_idx | rob_pnr_idx == rob_tail_idx)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at rob.scala:749 assert(!IsOlder(rob_pnr_idx, rob_head_idx, rob_tail_idx) || rob_pnr_idx === rob_tail_idx)\n");
        if (`STOP_COND_)
          $fatal;
      end
      if (~reset & ~(rob_tail_idx < rob_head_idx ^ _GEN_85 ^ rob_tail_idx >= rob_pnr_idx | full)) begin
        if (`ASSERT_VERBOSE_COND_)
          $error("Assertion failed\n    at rob.scala:752 assert(!IsOlder(rob_tail_idx, rob_pnr_idx, rob_head_idx) || full)\n");
        if (`STOP_COND_)
          $fatal;
      end
    end // always @(posedge)
  `endif // not def SYNTHESIS
  wire        _GEN_87 = _io_commit_rollback_T_3 & (rob_tail != rob_head | maybe_full);
  wire        rob_deq = _GEN_87 | finished_committing_row;
  assign full = rob_tail == rob_head & maybe_full;
  assign empty = _empty_T & {casez_tmp_241, casez_tmp_163, casez_tmp_85, casez_tmp_7} == 4'h0;
  reg         REG;
  reg         REG_1;
  reg         REG_2;
  reg  [1:0]  casez_tmp_315;
  wire [1:0]  _GEN_88 = empty ? 2'h1 : rob_state;
  always @(*) begin
    casez (rob_state)
      2'b00:
        casez_tmp_315 = 2'h1;
      2'b01:
        casez_tmp_315 = REG_1 ? 2'h2 : io_enq_valids_3 & io_enq_uops_3_is_unique | io_enq_valids_2 & io_enq_uops_2_is_unique | io_enq_valids_1 & io_enq_uops_1_is_unique | io_enq_valids_0 & io_enq_uops_0_is_unique ? 2'h3 : rob_state;
      2'b10:
        casez_tmp_315 = _GEN_88;
      default:
        casez_tmp_315 = REG_2 ? 2'h2 : _GEN_88;
    endcase
  end // always @(*)
  reg         casez_tmp_316;
  always @(*) begin
    casez (casez_tmp_7 ? 2'h0 : casez_tmp_85 ? 2'h1 : {1'h1, ~casez_tmp_163})
      2'b00:
        casez_tmp_316 = casez_tmp_33;
      2'b01:
        casez_tmp_316 = casez_tmp_111;
      2'b10:
        casez_tmp_316 = casez_tmp_189;
      default:
        casez_tmp_316 = casez_tmp_267;
    endcase
  end // always @(*)
  reg         io_com_load_is_at_rob_head_REG;
  wire [2:0]  _GEN_89 = {io_enq_valids_2, io_enq_valids_1, io_enq_valids_0} | {io_enq_valids_3, io_enq_valids_2, io_enq_valids_1};
  wire [1:0]  _GEN_90 = _GEN_89[1:0] | {io_enq_valids_3, io_enq_valids_2};
  wire [2:0]  _rob_tail_lsb_T_8 = ~{_GEN_89[2], _GEN_90[1], _GEN_90[0] | io_enq_valids_3};
  wire [2:0]  _GEN_91 = {casez_tmp_155, casez_tmp_77, casez_tmp} | {casez_tmp_233, casez_tmp_155, casez_tmp_77};
  wire [1:0]  _GEN_92 = _GEN_91[1:0] | {casez_tmp_233, casez_tmp_155};
  wire        safe_to_inc = _io_ready_T | (&rob_state);
  wire        _GEN_93 = rob_head == 5'h0;
  wire        _GEN_94 = rob_head == 5'h1;
  wire        _GEN_95 = rob_head == 5'h2;
  wire        _GEN_96 = rob_head == 5'h3;
  wire        _GEN_97 = rob_head == 5'h4;
  wire        _GEN_98 = rob_head == 5'h5;
  wire        _GEN_99 = rob_head == 5'h6;
  wire        _GEN_100 = rob_head == 5'h7;
  wire        _GEN_101 = rob_head == 5'h8;
  wire        _GEN_102 = rob_head == 5'h9;
  wire        _GEN_103 = rob_head == 5'hA;
  wire        _GEN_104 = rob_head == 5'hB;
  wire        _GEN_105 = rob_head == 5'hC;
  wire        _GEN_106 = rob_head == 5'hD;
  wire        _GEN_107 = rob_head == 5'hE;
  wire        _GEN_108 = rob_head == 5'hF;
  wire        _GEN_109 = rob_head == 5'h10;
  wire        _GEN_110 = rob_head == 5'h11;
  wire        _GEN_111 = rob_head == 5'h12;
  wire        _GEN_112 = rob_head == 5'h13;
  wire        _GEN_113 = rob_head == 5'h14;
  wire        _GEN_114 = rob_head == 5'h15;
  wire        _GEN_115 = rob_head == 5'h16;
  wire        _GEN_116 = rob_head == 5'h17;
  wire        _GEN_117 = rob_head == 5'h18;
  wire        _GEN_118 = rob_head == 5'h19;
  wire        _GEN_119 = rob_head == 5'h1A;
  wire        _GEN_120 = rob_head == 5'h1B;
  wire        _GEN_121 = rob_head == 5'h1C;
  wire        _GEN_122 = rob_head == 5'h1D;
  wire        _GEN_123 = rob_head == 5'h1E;
  wire        rob_pnr_unsafe_0 = casez_tmp_36 & (casez_tmp_34 | casez_tmp_35);
  wire        rob_pnr_unsafe_1 = casez_tmp_114 & (casez_tmp_112 | casez_tmp_113);
  wire        rob_pnr_unsafe_2 = casez_tmp_192 & (casez_tmp_190 | casez_tmp_191);
  wire [2:0]  _rob_head_lsb_T_8 = casez_tmp_7 ? 3'h0 : casez_tmp_85 ? 3'h1 : casez_tmp_163 ? 3'h2 : {casez_tmp_241, 2'h0};
  wire        _do_inc_row_T_4 = rob_pnr != rob_tail;
  wire        do_inc_row = ~(rob_pnr_unsafe_0 | rob_pnr_unsafe_1 | rob_pnr_unsafe_2 | casez_tmp_270 & (casez_tmp_268 | casez_tmp_269)) & (_do_inc_row_T_4 | full & ~pnr_maybe_at_tail);
  wire [3:0]  _GEN_124 = {io_enq_valids_3, io_enq_valids_2, io_enq_valids_1, io_enq_valids_0};
  wire        _GEN_125 = _io_commit_rollback_T_3 & rob_tail == rob_head & ~maybe_full;
  wire        _GEN_126 = (|_GEN_124) & ~io_enq_partial_stall;
  wire [2:0]  _rob_pnr_lsb_T_16 = {rob_pnr_unsafe_2, rob_pnr_unsafe_1, rob_pnr_unsafe_0} | ~{_GEN_91[2], _GEN_92[1], _GEN_92[0] | casez_tmp_233};
  wire        _GEN_127 = rob_tail == 5'h0;
  wire        _GEN_128 = io_enq_valids_0 & _GEN_127;
  wire        _GEN_129 = rob_tail == 5'h1;
  wire        _GEN_130 = io_enq_valids_0 & _GEN_129;
  wire        _GEN_131 = rob_tail == 5'h2;
  wire        _GEN_132 = io_enq_valids_0 & _GEN_131;
  wire        _GEN_133 = rob_tail == 5'h3;
  wire        _GEN_134 = io_enq_valids_0 & _GEN_133;
  wire        _GEN_135 = rob_tail == 5'h4;
  wire        _GEN_136 = io_enq_valids_0 & _GEN_135;
  wire        _GEN_137 = rob_tail == 5'h5;
  wire        _GEN_138 = io_enq_valids_0 & _GEN_137;
  wire        _GEN_139 = rob_tail == 5'h6;
  wire        _GEN_140 = io_enq_valids_0 & _GEN_139;
  wire        _GEN_141 = rob_tail == 5'h7;
  wire        _GEN_142 = io_enq_valids_0 & _GEN_141;
  wire        _GEN_143 = rob_tail == 5'h8;
  wire        _GEN_144 = io_enq_valids_0 & _GEN_143;
  wire        _GEN_145 = rob_tail == 5'h9;
  wire        _GEN_146 = io_enq_valids_0 & _GEN_145;
  wire        _GEN_147 = rob_tail == 5'hA;
  wire        _GEN_148 = io_enq_valids_0 & _GEN_147;
  wire        _GEN_149 = rob_tail == 5'hB;
  wire        _GEN_150 = io_enq_valids_0 & _GEN_149;
  wire        _GEN_151 = rob_tail == 5'hC;
  wire        _GEN_152 = io_enq_valids_0 & _GEN_151;
  wire        _GEN_153 = rob_tail == 5'hD;
  wire        _GEN_154 = io_enq_valids_0 & _GEN_153;
  wire        _GEN_155 = rob_tail == 5'hE;
  wire        _GEN_156 = io_enq_valids_0 & _GEN_155;
  wire        _GEN_157 = rob_tail == 5'hF;
  wire        _GEN_158 = io_enq_valids_0 & _GEN_157;
  wire        _GEN_159 = rob_tail == 5'h10;
  wire        _GEN_160 = io_enq_valids_0 & _GEN_159;
  wire        _GEN_161 = rob_tail == 5'h11;
  wire        _GEN_162 = io_enq_valids_0 & _GEN_161;
  wire        _GEN_163 = rob_tail == 5'h12;
  wire        _GEN_164 = io_enq_valids_0 & _GEN_163;
  wire        _GEN_165 = rob_tail == 5'h13;
  wire        _GEN_166 = io_enq_valids_0 & _GEN_165;
  wire        _GEN_167 = rob_tail == 5'h14;
  wire        _GEN_168 = io_enq_valids_0 & _GEN_167;
  wire        _GEN_169 = rob_tail == 5'h15;
  wire        _GEN_170 = io_enq_valids_0 & _GEN_169;
  wire        _GEN_171 = rob_tail == 5'h16;
  wire        _GEN_172 = io_enq_valids_0 & _GEN_171;
  wire        _GEN_173 = rob_tail == 5'h17;
  wire        _GEN_174 = io_enq_valids_0 & _GEN_173;
  wire        _GEN_175 = rob_tail == 5'h18;
  wire        _GEN_176 = io_enq_valids_0 & _GEN_175;
  wire        _GEN_177 = rob_tail == 5'h19;
  wire        _GEN_178 = io_enq_valids_0 & _GEN_177;
  wire        _GEN_179 = rob_tail == 5'h1A;
  wire        _GEN_180 = io_enq_valids_0 & _GEN_179;
  wire        _GEN_181 = rob_tail == 5'h1B;
  wire        _GEN_182 = io_enq_valids_0 & _GEN_181;
  wire        _GEN_183 = rob_tail == 5'h1C;
  wire        _GEN_184 = io_enq_valids_0 & _GEN_183;
  wire        _GEN_185 = rob_tail == 5'h1D;
  wire        _GEN_186 = io_enq_valids_0 & _GEN_185;
  wire        _GEN_187 = rob_tail == 5'h1E;
  wire        _GEN_188 = io_enq_valids_0 & _GEN_187;
  wire        _GEN_189 = io_enq_valids_0 & (&rob_tail);
  wire        _rob_bsy_T = io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei;
  wire        _GEN_190 = _GEN_128 ? ~_rob_bsy_T : rob_bsy_0;
  wire        _GEN_191 = _GEN_130 ? ~_rob_bsy_T : rob_bsy_1;
  wire        _GEN_192 = _GEN_132 ? ~_rob_bsy_T : rob_bsy_2;
  wire        _GEN_193 = _GEN_134 ? ~_rob_bsy_T : rob_bsy_3;
  wire        _GEN_194 = _GEN_136 ? ~_rob_bsy_T : rob_bsy_4;
  wire        _GEN_195 = _GEN_138 ? ~_rob_bsy_T : rob_bsy_5;
  wire        _GEN_196 = _GEN_140 ? ~_rob_bsy_T : rob_bsy_6;
  wire        _GEN_197 = _GEN_142 ? ~_rob_bsy_T : rob_bsy_7;
  wire        _GEN_198 = _GEN_144 ? ~_rob_bsy_T : rob_bsy_8;
  wire        _GEN_199 = _GEN_146 ? ~_rob_bsy_T : rob_bsy_9;
  wire        _GEN_200 = _GEN_148 ? ~_rob_bsy_T : rob_bsy_10;
  wire        _GEN_201 = _GEN_150 ? ~_rob_bsy_T : rob_bsy_11;
  wire        _GEN_202 = _GEN_152 ? ~_rob_bsy_T : rob_bsy_12;
  wire        _GEN_203 = _GEN_154 ? ~_rob_bsy_T : rob_bsy_13;
  wire        _GEN_204 = _GEN_156 ? ~_rob_bsy_T : rob_bsy_14;
  wire        _GEN_205 = _GEN_158 ? ~_rob_bsy_T : rob_bsy_15;
  wire        _GEN_206 = _GEN_160 ? ~_rob_bsy_T : rob_bsy_16;
  wire        _GEN_207 = _GEN_162 ? ~_rob_bsy_T : rob_bsy_17;
  wire        _GEN_208 = _GEN_164 ? ~_rob_bsy_T : rob_bsy_18;
  wire        _GEN_209 = _GEN_166 ? ~_rob_bsy_T : rob_bsy_19;
  wire        _GEN_210 = _GEN_168 ? ~_rob_bsy_T : rob_bsy_20;
  wire        _GEN_211 = _GEN_170 ? ~_rob_bsy_T : rob_bsy_21;
  wire        _GEN_212 = _GEN_172 ? ~_rob_bsy_T : rob_bsy_22;
  wire        _GEN_213 = _GEN_174 ? ~_rob_bsy_T : rob_bsy_23;
  wire        _GEN_214 = _GEN_176 ? ~_rob_bsy_T : rob_bsy_24;
  wire        _GEN_215 = _GEN_178 ? ~_rob_bsy_T : rob_bsy_25;
  wire        _GEN_216 = _GEN_180 ? ~_rob_bsy_T : rob_bsy_26;
  wire        _GEN_217 = _GEN_182 ? ~_rob_bsy_T : rob_bsy_27;
  wire        _GEN_218 = _GEN_184 ? ~_rob_bsy_T : rob_bsy_28;
  wire        _GEN_219 = _GEN_186 ? ~_rob_bsy_T : rob_bsy_29;
  wire        _GEN_220 = _GEN_188 ? ~_rob_bsy_T : rob_bsy_30;
  wire        _GEN_221 = _GEN_189 ? ~_rob_bsy_T : rob_bsy_31;
  wire        _rob_unsafe_T_4 = io_enq_uops_0_uses_ldq | io_enq_uops_0_uses_stq & ~io_enq_uops_0_is_fence | io_enq_uops_0_is_br | io_enq_uops_0_is_jalr;
  wire        _GEN_222 = _GEN_128 ? _rob_unsafe_T_4 : rob_unsafe_0;
  wire        _GEN_223 = _GEN_130 ? _rob_unsafe_T_4 : rob_unsafe_1;
  wire        _GEN_224 = _GEN_132 ? _rob_unsafe_T_4 : rob_unsafe_2;
  wire        _GEN_225 = _GEN_134 ? _rob_unsafe_T_4 : rob_unsafe_3;
  wire        _GEN_226 = _GEN_136 ? _rob_unsafe_T_4 : rob_unsafe_4;
  wire        _GEN_227 = _GEN_138 ? _rob_unsafe_T_4 : rob_unsafe_5;
  wire        _GEN_228 = _GEN_140 ? _rob_unsafe_T_4 : rob_unsafe_6;
  wire        _GEN_229 = _GEN_142 ? _rob_unsafe_T_4 : rob_unsafe_7;
  wire        _GEN_230 = _GEN_144 ? _rob_unsafe_T_4 : rob_unsafe_8;
  wire        _GEN_231 = _GEN_146 ? _rob_unsafe_T_4 : rob_unsafe_9;
  wire        _GEN_232 = _GEN_148 ? _rob_unsafe_T_4 : rob_unsafe_10;
  wire        _GEN_233 = _GEN_150 ? _rob_unsafe_T_4 : rob_unsafe_11;
  wire        _GEN_234 = _GEN_152 ? _rob_unsafe_T_4 : rob_unsafe_12;
  wire        _GEN_235 = _GEN_154 ? _rob_unsafe_T_4 : rob_unsafe_13;
  wire        _GEN_236 = _GEN_156 ? _rob_unsafe_T_4 : rob_unsafe_14;
  wire        _GEN_237 = _GEN_158 ? _rob_unsafe_T_4 : rob_unsafe_15;
  wire        _GEN_238 = _GEN_160 ? _rob_unsafe_T_4 : rob_unsafe_16;
  wire        _GEN_239 = _GEN_162 ? _rob_unsafe_T_4 : rob_unsafe_17;
  wire        _GEN_240 = _GEN_164 ? _rob_unsafe_T_4 : rob_unsafe_18;
  wire        _GEN_241 = _GEN_166 ? _rob_unsafe_T_4 : rob_unsafe_19;
  wire        _GEN_242 = _GEN_168 ? _rob_unsafe_T_4 : rob_unsafe_20;
  wire        _GEN_243 = _GEN_170 ? _rob_unsafe_T_4 : rob_unsafe_21;
  wire        _GEN_244 = _GEN_172 ? _rob_unsafe_T_4 : rob_unsafe_22;
  wire        _GEN_245 = _GEN_174 ? _rob_unsafe_T_4 : rob_unsafe_23;
  wire        _GEN_246 = _GEN_176 ? _rob_unsafe_T_4 : rob_unsafe_24;
  wire        _GEN_247 = _GEN_178 ? _rob_unsafe_T_4 : rob_unsafe_25;
  wire        _GEN_248 = _GEN_180 ? _rob_unsafe_T_4 : rob_unsafe_26;
  wire        _GEN_249 = _GEN_182 ? _rob_unsafe_T_4 : rob_unsafe_27;
  wire        _GEN_250 = _GEN_184 ? _rob_unsafe_T_4 : rob_unsafe_28;
  wire        _GEN_251 = _GEN_186 ? _rob_unsafe_T_4 : rob_unsafe_29;
  wire        _GEN_252 = _GEN_188 ? _rob_unsafe_T_4 : rob_unsafe_30;
  wire        _GEN_253 = _GEN_189 ? _rob_unsafe_T_4 : rob_unsafe_31;
  wire        _GEN_254 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_255 = _GEN & _GEN_254;
  wire        _GEN_256 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_257 = _GEN & _GEN_256;
  wire        _GEN_258 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_259 = _GEN & _GEN_258;
  wire        _GEN_260 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_261 = _GEN & _GEN_260;
  wire        _GEN_262 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_263 = _GEN & _GEN_262;
  wire        _GEN_264 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_265 = _GEN & _GEN_264;
  wire        _GEN_266 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_267 = _GEN & _GEN_266;
  wire        _GEN_268 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_269 = _GEN & _GEN_268;
  wire        _GEN_270 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_271 = _GEN & _GEN_270;
  wire        _GEN_272 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_273 = _GEN & _GEN_272;
  wire        _GEN_274 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_275 = _GEN & _GEN_274;
  wire        _GEN_276 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_277 = _GEN & _GEN_276;
  wire        _GEN_278 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_279 = _GEN & _GEN_278;
  wire        _GEN_280 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_281 = _GEN & _GEN_280;
  wire        _GEN_282 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_283 = _GEN & _GEN_282;
  wire        _GEN_284 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_285 = _GEN & _GEN_284;
  wire        _GEN_286 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_287 = _GEN & _GEN_286;
  wire        _GEN_288 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_289 = _GEN & _GEN_288;
  wire        _GEN_290 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_291 = _GEN & _GEN_290;
  wire        _GEN_292 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_293 = _GEN & _GEN_292;
  wire        _GEN_294 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_295 = _GEN & _GEN_294;
  wire        _GEN_296 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_297 = _GEN & _GEN_296;
  wire        _GEN_298 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_299 = _GEN & _GEN_298;
  wire        _GEN_300 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_301 = _GEN & _GEN_300;
  wire        _GEN_302 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_303 = _GEN & _GEN_302;
  wire        _GEN_304 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_305 = _GEN & _GEN_304;
  wire        _GEN_306 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_307 = _GEN & _GEN_306;
  wire        _GEN_308 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_309 = _GEN & _GEN_308;
  wire        _GEN_310 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_311 = _GEN & _GEN_310;
  wire        _GEN_312 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_313 = _GEN & _GEN_312;
  wire        _GEN_314 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_315 = _GEN & _GEN_314;
  wire        _GEN_316 = _GEN & (&(io_wb_resps_0_bits_uop_rob_idx[6:2]));
  wire        _GEN_317 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_318 = _GEN_317 | _GEN_255;
  wire        _GEN_319 = _GEN_0 ? ~_GEN_318 & _GEN_190 : ~_GEN_255 & _GEN_190;
  wire        _GEN_320 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_321 = _GEN_320 | _GEN_257;
  wire        _GEN_322 = _GEN_0 ? ~_GEN_321 & _GEN_191 : ~_GEN_257 & _GEN_191;
  wire        _GEN_323 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_324 = _GEN_323 | _GEN_259;
  wire        _GEN_325 = _GEN_0 ? ~_GEN_324 & _GEN_192 : ~_GEN_259 & _GEN_192;
  wire        _GEN_326 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_327 = _GEN_326 | _GEN_261;
  wire        _GEN_328 = _GEN_0 ? ~_GEN_327 & _GEN_193 : ~_GEN_261 & _GEN_193;
  wire        _GEN_329 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_330 = _GEN_329 | _GEN_263;
  wire        _GEN_331 = _GEN_0 ? ~_GEN_330 & _GEN_194 : ~_GEN_263 & _GEN_194;
  wire        _GEN_332 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_333 = _GEN_332 | _GEN_265;
  wire        _GEN_334 = _GEN_0 ? ~_GEN_333 & _GEN_195 : ~_GEN_265 & _GEN_195;
  wire        _GEN_335 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_336 = _GEN_335 | _GEN_267;
  wire        _GEN_337 = _GEN_0 ? ~_GEN_336 & _GEN_196 : ~_GEN_267 & _GEN_196;
  wire        _GEN_338 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_339 = _GEN_338 | _GEN_269;
  wire        _GEN_340 = _GEN_0 ? ~_GEN_339 & _GEN_197 : ~_GEN_269 & _GEN_197;
  wire        _GEN_341 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_342 = _GEN_341 | _GEN_271;
  wire        _GEN_343 = _GEN_0 ? ~_GEN_342 & _GEN_198 : ~_GEN_271 & _GEN_198;
  wire        _GEN_344 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_345 = _GEN_344 | _GEN_273;
  wire        _GEN_346 = _GEN_0 ? ~_GEN_345 & _GEN_199 : ~_GEN_273 & _GEN_199;
  wire        _GEN_347 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_348 = _GEN_347 | _GEN_275;
  wire        _GEN_349 = _GEN_0 ? ~_GEN_348 & _GEN_200 : ~_GEN_275 & _GEN_200;
  wire        _GEN_350 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_351 = _GEN_350 | _GEN_277;
  wire        _GEN_352 = _GEN_0 ? ~_GEN_351 & _GEN_201 : ~_GEN_277 & _GEN_201;
  wire        _GEN_353 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_354 = _GEN_353 | _GEN_279;
  wire        _GEN_355 = _GEN_0 ? ~_GEN_354 & _GEN_202 : ~_GEN_279 & _GEN_202;
  wire        _GEN_356 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_357 = _GEN_356 | _GEN_281;
  wire        _GEN_358 = _GEN_0 ? ~_GEN_357 & _GEN_203 : ~_GEN_281 & _GEN_203;
  wire        _GEN_359 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_360 = _GEN_359 | _GEN_283;
  wire        _GEN_361 = _GEN_0 ? ~_GEN_360 & _GEN_204 : ~_GEN_283 & _GEN_204;
  wire        _GEN_362 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_363 = _GEN_362 | _GEN_285;
  wire        _GEN_364 = _GEN_0 ? ~_GEN_363 & _GEN_205 : ~_GEN_285 & _GEN_205;
  wire        _GEN_365 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_366 = _GEN_365 | _GEN_287;
  wire        _GEN_367 = _GEN_0 ? ~_GEN_366 & _GEN_206 : ~_GEN_287 & _GEN_206;
  wire        _GEN_368 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_369 = _GEN_368 | _GEN_289;
  wire        _GEN_370 = _GEN_0 ? ~_GEN_369 & _GEN_207 : ~_GEN_289 & _GEN_207;
  wire        _GEN_371 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_372 = _GEN_371 | _GEN_291;
  wire        _GEN_373 = _GEN_0 ? ~_GEN_372 & _GEN_208 : ~_GEN_291 & _GEN_208;
  wire        _GEN_374 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_375 = _GEN_374 | _GEN_293;
  wire        _GEN_376 = _GEN_0 ? ~_GEN_375 & _GEN_209 : ~_GEN_293 & _GEN_209;
  wire        _GEN_377 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_378 = _GEN_377 | _GEN_295;
  wire        _GEN_379 = _GEN_0 ? ~_GEN_378 & _GEN_210 : ~_GEN_295 & _GEN_210;
  wire        _GEN_380 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_381 = _GEN_380 | _GEN_297;
  wire        _GEN_382 = _GEN_0 ? ~_GEN_381 & _GEN_211 : ~_GEN_297 & _GEN_211;
  wire        _GEN_383 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_384 = _GEN_383 | _GEN_299;
  wire        _GEN_385 = _GEN_0 ? ~_GEN_384 & _GEN_212 : ~_GEN_299 & _GEN_212;
  wire        _GEN_386 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_387 = _GEN_386 | _GEN_301;
  wire        _GEN_388 = _GEN_0 ? ~_GEN_387 & _GEN_213 : ~_GEN_301 & _GEN_213;
  wire        _GEN_389 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_390 = _GEN_389 | _GEN_303;
  wire        _GEN_391 = _GEN_0 ? ~_GEN_390 & _GEN_214 : ~_GEN_303 & _GEN_214;
  wire        _GEN_392 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_393 = _GEN_392 | _GEN_305;
  wire        _GEN_394 = _GEN_0 ? ~_GEN_393 & _GEN_215 : ~_GEN_305 & _GEN_215;
  wire        _GEN_395 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_396 = _GEN_395 | _GEN_307;
  wire        _GEN_397 = _GEN_0 ? ~_GEN_396 & _GEN_216 : ~_GEN_307 & _GEN_216;
  wire        _GEN_398 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_399 = _GEN_398 | _GEN_309;
  wire        _GEN_400 = _GEN_0 ? ~_GEN_399 & _GEN_217 : ~_GEN_309 & _GEN_217;
  wire        _GEN_401 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_402 = _GEN_401 | _GEN_311;
  wire        _GEN_403 = _GEN_0 ? ~_GEN_402 & _GEN_218 : ~_GEN_311 & _GEN_218;
  wire        _GEN_404 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_405 = _GEN_404 | _GEN_313;
  wire        _GEN_406 = _GEN_0 ? ~_GEN_405 & _GEN_219 : ~_GEN_313 & _GEN_219;
  wire        _GEN_407 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_408 = _GEN_407 | _GEN_315;
  wire        _GEN_409 = _GEN_0 ? ~_GEN_408 & _GEN_220 : ~_GEN_315 & _GEN_220;
  wire        _GEN_410 = (&(io_wb_resps_1_bits_uop_rob_idx[6:2])) | _GEN_316;
  wire        _GEN_411 = _GEN_0 ? ~_GEN_410 & _GEN_221 : ~_GEN_316 & _GEN_221;
  wire        _GEN_412 = _GEN_0 ? ~_GEN_318 & _GEN_222 : ~_GEN_255 & _GEN_222;
  wire        _GEN_413 = _GEN_0 ? ~_GEN_321 & _GEN_223 : ~_GEN_257 & _GEN_223;
  wire        _GEN_414 = _GEN_0 ? ~_GEN_324 & _GEN_224 : ~_GEN_259 & _GEN_224;
  wire        _GEN_415 = _GEN_0 ? ~_GEN_327 & _GEN_225 : ~_GEN_261 & _GEN_225;
  wire        _GEN_416 = _GEN_0 ? ~_GEN_330 & _GEN_226 : ~_GEN_263 & _GEN_226;
  wire        _GEN_417 = _GEN_0 ? ~_GEN_333 & _GEN_227 : ~_GEN_265 & _GEN_227;
  wire        _GEN_418 = _GEN_0 ? ~_GEN_336 & _GEN_228 : ~_GEN_267 & _GEN_228;
  wire        _GEN_419 = _GEN_0 ? ~_GEN_339 & _GEN_229 : ~_GEN_269 & _GEN_229;
  wire        _GEN_420 = _GEN_0 ? ~_GEN_342 & _GEN_230 : ~_GEN_271 & _GEN_230;
  wire        _GEN_421 = _GEN_0 ? ~_GEN_345 & _GEN_231 : ~_GEN_273 & _GEN_231;
  wire        _GEN_422 = _GEN_0 ? ~_GEN_348 & _GEN_232 : ~_GEN_275 & _GEN_232;
  wire        _GEN_423 = _GEN_0 ? ~_GEN_351 & _GEN_233 : ~_GEN_277 & _GEN_233;
  wire        _GEN_424 = _GEN_0 ? ~_GEN_354 & _GEN_234 : ~_GEN_279 & _GEN_234;
  wire        _GEN_425 = _GEN_0 ? ~_GEN_357 & _GEN_235 : ~_GEN_281 & _GEN_235;
  wire        _GEN_426 = _GEN_0 ? ~_GEN_360 & _GEN_236 : ~_GEN_283 & _GEN_236;
  wire        _GEN_427 = _GEN_0 ? ~_GEN_363 & _GEN_237 : ~_GEN_285 & _GEN_237;
  wire        _GEN_428 = _GEN_0 ? ~_GEN_366 & _GEN_238 : ~_GEN_287 & _GEN_238;
  wire        _GEN_429 = _GEN_0 ? ~_GEN_369 & _GEN_239 : ~_GEN_289 & _GEN_239;
  wire        _GEN_430 = _GEN_0 ? ~_GEN_372 & _GEN_240 : ~_GEN_291 & _GEN_240;
  wire        _GEN_431 = _GEN_0 ? ~_GEN_375 & _GEN_241 : ~_GEN_293 & _GEN_241;
  wire        _GEN_432 = _GEN_0 ? ~_GEN_378 & _GEN_242 : ~_GEN_295 & _GEN_242;
  wire        _GEN_433 = _GEN_0 ? ~_GEN_381 & _GEN_243 : ~_GEN_297 & _GEN_243;
  wire        _GEN_434 = _GEN_0 ? ~_GEN_384 & _GEN_244 : ~_GEN_299 & _GEN_244;
  wire        _GEN_435 = _GEN_0 ? ~_GEN_387 & _GEN_245 : ~_GEN_301 & _GEN_245;
  wire        _GEN_436 = _GEN_0 ? ~_GEN_390 & _GEN_246 : ~_GEN_303 & _GEN_246;
  wire        _GEN_437 = _GEN_0 ? ~_GEN_393 & _GEN_247 : ~_GEN_305 & _GEN_247;
  wire        _GEN_438 = _GEN_0 ? ~_GEN_396 & _GEN_248 : ~_GEN_307 & _GEN_248;
  wire        _GEN_439 = _GEN_0 ? ~_GEN_399 & _GEN_249 : ~_GEN_309 & _GEN_249;
  wire        _GEN_440 = _GEN_0 ? ~_GEN_402 & _GEN_250 : ~_GEN_311 & _GEN_250;
  wire        _GEN_441 = _GEN_0 ? ~_GEN_405 & _GEN_251 : ~_GEN_313 & _GEN_251;
  wire        _GEN_442 = _GEN_0 ? ~_GEN_408 & _GEN_252 : ~_GEN_315 & _GEN_252;
  wire        _GEN_443 = _GEN_0 ? ~_GEN_410 & _GEN_253 : ~_GEN_316 & _GEN_253;
  wire        _GEN_444 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_445 = _GEN_1 & _GEN_444;
  wire        _GEN_446 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_447 = _GEN_1 & _GEN_446;
  wire        _GEN_448 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_449 = _GEN_1 & _GEN_448;
  wire        _GEN_450 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_451 = _GEN_1 & _GEN_450;
  wire        _GEN_452 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_453 = _GEN_1 & _GEN_452;
  wire        _GEN_454 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_455 = _GEN_1 & _GEN_454;
  wire        _GEN_456 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_457 = _GEN_1 & _GEN_456;
  wire        _GEN_458 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_459 = _GEN_1 & _GEN_458;
  wire        _GEN_460 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_461 = _GEN_1 & _GEN_460;
  wire        _GEN_462 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_463 = _GEN_1 & _GEN_462;
  wire        _GEN_464 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_465 = _GEN_1 & _GEN_464;
  wire        _GEN_466 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_467 = _GEN_1 & _GEN_466;
  wire        _GEN_468 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_469 = _GEN_1 & _GEN_468;
  wire        _GEN_470 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_471 = _GEN_1 & _GEN_470;
  wire        _GEN_472 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_473 = _GEN_1 & _GEN_472;
  wire        _GEN_474 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_475 = _GEN_1 & _GEN_474;
  wire        _GEN_476 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_477 = _GEN_1 & _GEN_476;
  wire        _GEN_478 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_479 = _GEN_1 & _GEN_478;
  wire        _GEN_480 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_481 = _GEN_1 & _GEN_480;
  wire        _GEN_482 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_483 = _GEN_1 & _GEN_482;
  wire        _GEN_484 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_485 = _GEN_1 & _GEN_484;
  wire        _GEN_486 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_487 = _GEN_1 & _GEN_486;
  wire        _GEN_488 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_489 = _GEN_1 & _GEN_488;
  wire        _GEN_490 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_491 = _GEN_1 & _GEN_490;
  wire        _GEN_492 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_493 = _GEN_1 & _GEN_492;
  wire        _GEN_494 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_495 = _GEN_1 & _GEN_494;
  wire        _GEN_496 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_497 = _GEN_1 & _GEN_496;
  wire        _GEN_498 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_499 = _GEN_1 & _GEN_498;
  wire        _GEN_500 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_501 = _GEN_1 & _GEN_500;
  wire        _GEN_502 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_503 = _GEN_1 & _GEN_502;
  wire        _GEN_504 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_505 = _GEN_1 & _GEN_504;
  wire        _GEN_506 = _GEN_1 & (&(io_wb_resps_2_bits_uop_rob_idx[6:2]));
  wire        _GEN_507 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_508 = _GEN_507 | _GEN_445;
  wire        _GEN_509 = _GEN_2 ? ~_GEN_508 & _GEN_319 : ~_GEN_445 & _GEN_319;
  wire        _GEN_510 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_511 = _GEN_510 | _GEN_447;
  wire        _GEN_512 = _GEN_2 ? ~_GEN_511 & _GEN_322 : ~_GEN_447 & _GEN_322;
  wire        _GEN_513 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_514 = _GEN_513 | _GEN_449;
  wire        _GEN_515 = _GEN_2 ? ~_GEN_514 & _GEN_325 : ~_GEN_449 & _GEN_325;
  wire        _GEN_516 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_517 = _GEN_516 | _GEN_451;
  wire        _GEN_518 = _GEN_2 ? ~_GEN_517 & _GEN_328 : ~_GEN_451 & _GEN_328;
  wire        _GEN_519 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_520 = _GEN_519 | _GEN_453;
  wire        _GEN_521 = _GEN_2 ? ~_GEN_520 & _GEN_331 : ~_GEN_453 & _GEN_331;
  wire        _GEN_522 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_523 = _GEN_522 | _GEN_455;
  wire        _GEN_524 = _GEN_2 ? ~_GEN_523 & _GEN_334 : ~_GEN_455 & _GEN_334;
  wire        _GEN_525 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_526 = _GEN_525 | _GEN_457;
  wire        _GEN_527 = _GEN_2 ? ~_GEN_526 & _GEN_337 : ~_GEN_457 & _GEN_337;
  wire        _GEN_528 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_529 = _GEN_528 | _GEN_459;
  wire        _GEN_530 = _GEN_2 ? ~_GEN_529 & _GEN_340 : ~_GEN_459 & _GEN_340;
  wire        _GEN_531 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_532 = _GEN_531 | _GEN_461;
  wire        _GEN_533 = _GEN_2 ? ~_GEN_532 & _GEN_343 : ~_GEN_461 & _GEN_343;
  wire        _GEN_534 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_535 = _GEN_534 | _GEN_463;
  wire        _GEN_536 = _GEN_2 ? ~_GEN_535 & _GEN_346 : ~_GEN_463 & _GEN_346;
  wire        _GEN_537 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_538 = _GEN_537 | _GEN_465;
  wire        _GEN_539 = _GEN_2 ? ~_GEN_538 & _GEN_349 : ~_GEN_465 & _GEN_349;
  wire        _GEN_540 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_541 = _GEN_540 | _GEN_467;
  wire        _GEN_542 = _GEN_2 ? ~_GEN_541 & _GEN_352 : ~_GEN_467 & _GEN_352;
  wire        _GEN_543 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_544 = _GEN_543 | _GEN_469;
  wire        _GEN_545 = _GEN_2 ? ~_GEN_544 & _GEN_355 : ~_GEN_469 & _GEN_355;
  wire        _GEN_546 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_547 = _GEN_546 | _GEN_471;
  wire        _GEN_548 = _GEN_2 ? ~_GEN_547 & _GEN_358 : ~_GEN_471 & _GEN_358;
  wire        _GEN_549 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_550 = _GEN_549 | _GEN_473;
  wire        _GEN_551 = _GEN_2 ? ~_GEN_550 & _GEN_361 : ~_GEN_473 & _GEN_361;
  wire        _GEN_552 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_553 = _GEN_552 | _GEN_475;
  wire        _GEN_554 = _GEN_2 ? ~_GEN_553 & _GEN_364 : ~_GEN_475 & _GEN_364;
  wire        _GEN_555 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_556 = _GEN_555 | _GEN_477;
  wire        _GEN_557 = _GEN_2 ? ~_GEN_556 & _GEN_367 : ~_GEN_477 & _GEN_367;
  wire        _GEN_558 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_559 = _GEN_558 | _GEN_479;
  wire        _GEN_560 = _GEN_2 ? ~_GEN_559 & _GEN_370 : ~_GEN_479 & _GEN_370;
  wire        _GEN_561 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_562 = _GEN_561 | _GEN_481;
  wire        _GEN_563 = _GEN_2 ? ~_GEN_562 & _GEN_373 : ~_GEN_481 & _GEN_373;
  wire        _GEN_564 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_565 = _GEN_564 | _GEN_483;
  wire        _GEN_566 = _GEN_2 ? ~_GEN_565 & _GEN_376 : ~_GEN_483 & _GEN_376;
  wire        _GEN_567 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_568 = _GEN_567 | _GEN_485;
  wire        _GEN_569 = _GEN_2 ? ~_GEN_568 & _GEN_379 : ~_GEN_485 & _GEN_379;
  wire        _GEN_570 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_571 = _GEN_570 | _GEN_487;
  wire        _GEN_572 = _GEN_2 ? ~_GEN_571 & _GEN_382 : ~_GEN_487 & _GEN_382;
  wire        _GEN_573 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_574 = _GEN_573 | _GEN_489;
  wire        _GEN_575 = _GEN_2 ? ~_GEN_574 & _GEN_385 : ~_GEN_489 & _GEN_385;
  wire        _GEN_576 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_577 = _GEN_576 | _GEN_491;
  wire        _GEN_578 = _GEN_2 ? ~_GEN_577 & _GEN_388 : ~_GEN_491 & _GEN_388;
  wire        _GEN_579 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_580 = _GEN_579 | _GEN_493;
  wire        _GEN_581 = _GEN_2 ? ~_GEN_580 & _GEN_391 : ~_GEN_493 & _GEN_391;
  wire        _GEN_582 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_583 = _GEN_582 | _GEN_495;
  wire        _GEN_584 = _GEN_2 ? ~_GEN_583 & _GEN_394 : ~_GEN_495 & _GEN_394;
  wire        _GEN_585 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_586 = _GEN_585 | _GEN_497;
  wire        _GEN_587 = _GEN_2 ? ~_GEN_586 & _GEN_397 : ~_GEN_497 & _GEN_397;
  wire        _GEN_588 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_589 = _GEN_588 | _GEN_499;
  wire        _GEN_590 = _GEN_2 ? ~_GEN_589 & _GEN_400 : ~_GEN_499 & _GEN_400;
  wire        _GEN_591 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_592 = _GEN_591 | _GEN_501;
  wire        _GEN_593 = _GEN_2 ? ~_GEN_592 & _GEN_403 : ~_GEN_501 & _GEN_403;
  wire        _GEN_594 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_595 = _GEN_594 | _GEN_503;
  wire        _GEN_596 = _GEN_2 ? ~_GEN_595 & _GEN_406 : ~_GEN_503 & _GEN_406;
  wire        _GEN_597 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_598 = _GEN_597 | _GEN_505;
  wire        _GEN_599 = _GEN_2 ? ~_GEN_598 & _GEN_409 : ~_GEN_505 & _GEN_409;
  wire        _GEN_600 = (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_506;
  wire        _GEN_601 = _GEN_2 ? ~_GEN_600 & _GEN_411 : ~_GEN_506 & _GEN_411;
  wire        _GEN_602 = _GEN_2 ? ~_GEN_508 & _GEN_412 : ~_GEN_445 & _GEN_412;
  wire        _GEN_603 = _GEN_2 ? ~_GEN_511 & _GEN_413 : ~_GEN_447 & _GEN_413;
  wire        _GEN_604 = _GEN_2 ? ~_GEN_514 & _GEN_414 : ~_GEN_449 & _GEN_414;
  wire        _GEN_605 = _GEN_2 ? ~_GEN_517 & _GEN_415 : ~_GEN_451 & _GEN_415;
  wire        _GEN_606 = _GEN_2 ? ~_GEN_520 & _GEN_416 : ~_GEN_453 & _GEN_416;
  wire        _GEN_607 = _GEN_2 ? ~_GEN_523 & _GEN_417 : ~_GEN_455 & _GEN_417;
  wire        _GEN_608 = _GEN_2 ? ~_GEN_526 & _GEN_418 : ~_GEN_457 & _GEN_418;
  wire        _GEN_609 = _GEN_2 ? ~_GEN_529 & _GEN_419 : ~_GEN_459 & _GEN_419;
  wire        _GEN_610 = _GEN_2 ? ~_GEN_532 & _GEN_420 : ~_GEN_461 & _GEN_420;
  wire        _GEN_611 = _GEN_2 ? ~_GEN_535 & _GEN_421 : ~_GEN_463 & _GEN_421;
  wire        _GEN_612 = _GEN_2 ? ~_GEN_538 & _GEN_422 : ~_GEN_465 & _GEN_422;
  wire        _GEN_613 = _GEN_2 ? ~_GEN_541 & _GEN_423 : ~_GEN_467 & _GEN_423;
  wire        _GEN_614 = _GEN_2 ? ~_GEN_544 & _GEN_424 : ~_GEN_469 & _GEN_424;
  wire        _GEN_615 = _GEN_2 ? ~_GEN_547 & _GEN_425 : ~_GEN_471 & _GEN_425;
  wire        _GEN_616 = _GEN_2 ? ~_GEN_550 & _GEN_426 : ~_GEN_473 & _GEN_426;
  wire        _GEN_617 = _GEN_2 ? ~_GEN_553 & _GEN_427 : ~_GEN_475 & _GEN_427;
  wire        _GEN_618 = _GEN_2 ? ~_GEN_556 & _GEN_428 : ~_GEN_477 & _GEN_428;
  wire        _GEN_619 = _GEN_2 ? ~_GEN_559 & _GEN_429 : ~_GEN_479 & _GEN_429;
  wire        _GEN_620 = _GEN_2 ? ~_GEN_562 & _GEN_430 : ~_GEN_481 & _GEN_430;
  wire        _GEN_621 = _GEN_2 ? ~_GEN_565 & _GEN_431 : ~_GEN_483 & _GEN_431;
  wire        _GEN_622 = _GEN_2 ? ~_GEN_568 & _GEN_432 : ~_GEN_485 & _GEN_432;
  wire        _GEN_623 = _GEN_2 ? ~_GEN_571 & _GEN_433 : ~_GEN_487 & _GEN_433;
  wire        _GEN_624 = _GEN_2 ? ~_GEN_574 & _GEN_434 : ~_GEN_489 & _GEN_434;
  wire        _GEN_625 = _GEN_2 ? ~_GEN_577 & _GEN_435 : ~_GEN_491 & _GEN_435;
  wire        _GEN_626 = _GEN_2 ? ~_GEN_580 & _GEN_436 : ~_GEN_493 & _GEN_436;
  wire        _GEN_627 = _GEN_2 ? ~_GEN_583 & _GEN_437 : ~_GEN_495 & _GEN_437;
  wire        _GEN_628 = _GEN_2 ? ~_GEN_586 & _GEN_438 : ~_GEN_497 & _GEN_438;
  wire        _GEN_629 = _GEN_2 ? ~_GEN_589 & _GEN_439 : ~_GEN_499 & _GEN_439;
  wire        _GEN_630 = _GEN_2 ? ~_GEN_592 & _GEN_440 : ~_GEN_501 & _GEN_440;
  wire        _GEN_631 = _GEN_2 ? ~_GEN_595 & _GEN_441 : ~_GEN_503 & _GEN_441;
  wire        _GEN_632 = _GEN_2 ? ~_GEN_598 & _GEN_442 : ~_GEN_505 & _GEN_442;
  wire        _GEN_633 = _GEN_2 ? ~_GEN_600 & _GEN_443 : ~_GEN_506 & _GEN_443;
  wire        _GEN_634 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_635 = _GEN_3 & _GEN_634;
  wire        _GEN_636 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_637 = _GEN_3 & _GEN_636;
  wire        _GEN_638 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_639 = _GEN_3 & _GEN_638;
  wire        _GEN_640 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_641 = _GEN_3 & _GEN_640;
  wire        _GEN_642 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_643 = _GEN_3 & _GEN_642;
  wire        _GEN_644 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_645 = _GEN_3 & _GEN_644;
  wire        _GEN_646 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_647 = _GEN_3 & _GEN_646;
  wire        _GEN_648 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_649 = _GEN_3 & _GEN_648;
  wire        _GEN_650 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_651 = _GEN_3 & _GEN_650;
  wire        _GEN_652 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_653 = _GEN_3 & _GEN_652;
  wire        _GEN_654 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_655 = _GEN_3 & _GEN_654;
  wire        _GEN_656 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_657 = _GEN_3 & _GEN_656;
  wire        _GEN_658 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_659 = _GEN_3 & _GEN_658;
  wire        _GEN_660 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_661 = _GEN_3 & _GEN_660;
  wire        _GEN_662 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_663 = _GEN_3 & _GEN_662;
  wire        _GEN_664 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_665 = _GEN_3 & _GEN_664;
  wire        _GEN_666 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_667 = _GEN_3 & _GEN_666;
  wire        _GEN_668 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_669 = _GEN_3 & _GEN_668;
  wire        _GEN_670 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_671 = _GEN_3 & _GEN_670;
  wire        _GEN_672 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_673 = _GEN_3 & _GEN_672;
  wire        _GEN_674 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_675 = _GEN_3 & _GEN_674;
  wire        _GEN_676 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_677 = _GEN_3 & _GEN_676;
  wire        _GEN_678 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_679 = _GEN_3 & _GEN_678;
  wire        _GEN_680 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_681 = _GEN_3 & _GEN_680;
  wire        _GEN_682 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_683 = _GEN_3 & _GEN_682;
  wire        _GEN_684 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_685 = _GEN_3 & _GEN_684;
  wire        _GEN_686 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_687 = _GEN_3 & _GEN_686;
  wire        _GEN_688 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_689 = _GEN_3 & _GEN_688;
  wire        _GEN_690 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_691 = _GEN_3 & _GEN_690;
  wire        _GEN_692 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_693 = _GEN_3 & _GEN_692;
  wire        _GEN_694 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_695 = _GEN_3 & _GEN_694;
  wire        _GEN_696 = _GEN_3 & (&(io_wb_resps_4_bits_uop_rob_idx[6:2]));
  wire        _GEN_697 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_698 = _GEN_697 | _GEN_635;
  wire        _GEN_699 = _GEN_4 ? ~_GEN_698 & _GEN_509 : ~_GEN_635 & _GEN_509;
  wire        _GEN_700 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_701 = _GEN_700 | _GEN_637;
  wire        _GEN_702 = _GEN_4 ? ~_GEN_701 & _GEN_512 : ~_GEN_637 & _GEN_512;
  wire        _GEN_703 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_704 = _GEN_703 | _GEN_639;
  wire        _GEN_705 = _GEN_4 ? ~_GEN_704 & _GEN_515 : ~_GEN_639 & _GEN_515;
  wire        _GEN_706 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_707 = _GEN_706 | _GEN_641;
  wire        _GEN_708 = _GEN_4 ? ~_GEN_707 & _GEN_518 : ~_GEN_641 & _GEN_518;
  wire        _GEN_709 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_710 = _GEN_709 | _GEN_643;
  wire        _GEN_711 = _GEN_4 ? ~_GEN_710 & _GEN_521 : ~_GEN_643 & _GEN_521;
  wire        _GEN_712 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_713 = _GEN_712 | _GEN_645;
  wire        _GEN_714 = _GEN_4 ? ~_GEN_713 & _GEN_524 : ~_GEN_645 & _GEN_524;
  wire        _GEN_715 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_716 = _GEN_715 | _GEN_647;
  wire        _GEN_717 = _GEN_4 ? ~_GEN_716 & _GEN_527 : ~_GEN_647 & _GEN_527;
  wire        _GEN_718 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_719 = _GEN_718 | _GEN_649;
  wire        _GEN_720 = _GEN_4 ? ~_GEN_719 & _GEN_530 : ~_GEN_649 & _GEN_530;
  wire        _GEN_721 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_722 = _GEN_721 | _GEN_651;
  wire        _GEN_723 = _GEN_4 ? ~_GEN_722 & _GEN_533 : ~_GEN_651 & _GEN_533;
  wire        _GEN_724 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_725 = _GEN_724 | _GEN_653;
  wire        _GEN_726 = _GEN_4 ? ~_GEN_725 & _GEN_536 : ~_GEN_653 & _GEN_536;
  wire        _GEN_727 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_728 = _GEN_727 | _GEN_655;
  wire        _GEN_729 = _GEN_4 ? ~_GEN_728 & _GEN_539 : ~_GEN_655 & _GEN_539;
  wire        _GEN_730 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_731 = _GEN_730 | _GEN_657;
  wire        _GEN_732 = _GEN_4 ? ~_GEN_731 & _GEN_542 : ~_GEN_657 & _GEN_542;
  wire        _GEN_733 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_734 = _GEN_733 | _GEN_659;
  wire        _GEN_735 = _GEN_4 ? ~_GEN_734 & _GEN_545 : ~_GEN_659 & _GEN_545;
  wire        _GEN_736 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_737 = _GEN_736 | _GEN_661;
  wire        _GEN_738 = _GEN_4 ? ~_GEN_737 & _GEN_548 : ~_GEN_661 & _GEN_548;
  wire        _GEN_739 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_740 = _GEN_739 | _GEN_663;
  wire        _GEN_741 = _GEN_4 ? ~_GEN_740 & _GEN_551 : ~_GEN_663 & _GEN_551;
  wire        _GEN_742 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_743 = _GEN_742 | _GEN_665;
  wire        _GEN_744 = _GEN_4 ? ~_GEN_743 & _GEN_554 : ~_GEN_665 & _GEN_554;
  wire        _GEN_745 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_746 = _GEN_745 | _GEN_667;
  wire        _GEN_747 = _GEN_4 ? ~_GEN_746 & _GEN_557 : ~_GEN_667 & _GEN_557;
  wire        _GEN_748 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_749 = _GEN_748 | _GEN_669;
  wire        _GEN_750 = _GEN_4 ? ~_GEN_749 & _GEN_560 : ~_GEN_669 & _GEN_560;
  wire        _GEN_751 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_752 = _GEN_751 | _GEN_671;
  wire        _GEN_753 = _GEN_4 ? ~_GEN_752 & _GEN_563 : ~_GEN_671 & _GEN_563;
  wire        _GEN_754 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_755 = _GEN_754 | _GEN_673;
  wire        _GEN_756 = _GEN_4 ? ~_GEN_755 & _GEN_566 : ~_GEN_673 & _GEN_566;
  wire        _GEN_757 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_758 = _GEN_757 | _GEN_675;
  wire        _GEN_759 = _GEN_4 ? ~_GEN_758 & _GEN_569 : ~_GEN_675 & _GEN_569;
  wire        _GEN_760 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_761 = _GEN_760 | _GEN_677;
  wire        _GEN_762 = _GEN_4 ? ~_GEN_761 & _GEN_572 : ~_GEN_677 & _GEN_572;
  wire        _GEN_763 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_764 = _GEN_763 | _GEN_679;
  wire        _GEN_765 = _GEN_4 ? ~_GEN_764 & _GEN_575 : ~_GEN_679 & _GEN_575;
  wire        _GEN_766 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_767 = _GEN_766 | _GEN_681;
  wire        _GEN_768 = _GEN_4 ? ~_GEN_767 & _GEN_578 : ~_GEN_681 & _GEN_578;
  wire        _GEN_769 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_770 = _GEN_769 | _GEN_683;
  wire        _GEN_771 = _GEN_4 ? ~_GEN_770 & _GEN_581 : ~_GEN_683 & _GEN_581;
  wire        _GEN_772 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_773 = _GEN_772 | _GEN_685;
  wire        _GEN_774 = _GEN_4 ? ~_GEN_773 & _GEN_584 : ~_GEN_685 & _GEN_584;
  wire        _GEN_775 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_776 = _GEN_775 | _GEN_687;
  wire        _GEN_777 = _GEN_4 ? ~_GEN_776 & _GEN_587 : ~_GEN_687 & _GEN_587;
  wire        _GEN_778 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_779 = _GEN_778 | _GEN_689;
  wire        _GEN_780 = _GEN_4 ? ~_GEN_779 & _GEN_590 : ~_GEN_689 & _GEN_590;
  wire        _GEN_781 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_782 = _GEN_781 | _GEN_691;
  wire        _GEN_783 = _GEN_4 ? ~_GEN_782 & _GEN_593 : ~_GEN_691 & _GEN_593;
  wire        _GEN_784 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_785 = _GEN_784 | _GEN_693;
  wire        _GEN_786 = _GEN_4 ? ~_GEN_785 & _GEN_596 : ~_GEN_693 & _GEN_596;
  wire        _GEN_787 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_788 = _GEN_787 | _GEN_695;
  wire        _GEN_789 = _GEN_4 ? ~_GEN_788 & _GEN_599 : ~_GEN_695 & _GEN_599;
  wire        _GEN_790 = (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_696;
  wire        _GEN_791 = _GEN_4 ? ~_GEN_790 & _GEN_601 : ~_GEN_696 & _GEN_601;
  wire        _GEN_792 = _GEN_4 ? ~_GEN_698 & _GEN_602 : ~_GEN_635 & _GEN_602;
  wire        _GEN_793 = _GEN_4 ? ~_GEN_701 & _GEN_603 : ~_GEN_637 & _GEN_603;
  wire        _GEN_794 = _GEN_4 ? ~_GEN_704 & _GEN_604 : ~_GEN_639 & _GEN_604;
  wire        _GEN_795 = _GEN_4 ? ~_GEN_707 & _GEN_605 : ~_GEN_641 & _GEN_605;
  wire        _GEN_796 = _GEN_4 ? ~_GEN_710 & _GEN_606 : ~_GEN_643 & _GEN_606;
  wire        _GEN_797 = _GEN_4 ? ~_GEN_713 & _GEN_607 : ~_GEN_645 & _GEN_607;
  wire        _GEN_798 = _GEN_4 ? ~_GEN_716 & _GEN_608 : ~_GEN_647 & _GEN_608;
  wire        _GEN_799 = _GEN_4 ? ~_GEN_719 & _GEN_609 : ~_GEN_649 & _GEN_609;
  wire        _GEN_800 = _GEN_4 ? ~_GEN_722 & _GEN_610 : ~_GEN_651 & _GEN_610;
  wire        _GEN_801 = _GEN_4 ? ~_GEN_725 & _GEN_611 : ~_GEN_653 & _GEN_611;
  wire        _GEN_802 = _GEN_4 ? ~_GEN_728 & _GEN_612 : ~_GEN_655 & _GEN_612;
  wire        _GEN_803 = _GEN_4 ? ~_GEN_731 & _GEN_613 : ~_GEN_657 & _GEN_613;
  wire        _GEN_804 = _GEN_4 ? ~_GEN_734 & _GEN_614 : ~_GEN_659 & _GEN_614;
  wire        _GEN_805 = _GEN_4 ? ~_GEN_737 & _GEN_615 : ~_GEN_661 & _GEN_615;
  wire        _GEN_806 = _GEN_4 ? ~_GEN_740 & _GEN_616 : ~_GEN_663 & _GEN_616;
  wire        _GEN_807 = _GEN_4 ? ~_GEN_743 & _GEN_617 : ~_GEN_665 & _GEN_617;
  wire        _GEN_808 = _GEN_4 ? ~_GEN_746 & _GEN_618 : ~_GEN_667 & _GEN_618;
  wire        _GEN_809 = _GEN_4 ? ~_GEN_749 & _GEN_619 : ~_GEN_669 & _GEN_619;
  wire        _GEN_810 = _GEN_4 ? ~_GEN_752 & _GEN_620 : ~_GEN_671 & _GEN_620;
  wire        _GEN_811 = _GEN_4 ? ~_GEN_755 & _GEN_621 : ~_GEN_673 & _GEN_621;
  wire        _GEN_812 = _GEN_4 ? ~_GEN_758 & _GEN_622 : ~_GEN_675 & _GEN_622;
  wire        _GEN_813 = _GEN_4 ? ~_GEN_761 & _GEN_623 : ~_GEN_677 & _GEN_623;
  wire        _GEN_814 = _GEN_4 ? ~_GEN_764 & _GEN_624 : ~_GEN_679 & _GEN_624;
  wire        _GEN_815 = _GEN_4 ? ~_GEN_767 & _GEN_625 : ~_GEN_681 & _GEN_625;
  wire        _GEN_816 = _GEN_4 ? ~_GEN_770 & _GEN_626 : ~_GEN_683 & _GEN_626;
  wire        _GEN_817 = _GEN_4 ? ~_GEN_773 & _GEN_627 : ~_GEN_685 & _GEN_627;
  wire        _GEN_818 = _GEN_4 ? ~_GEN_776 & _GEN_628 : ~_GEN_687 & _GEN_628;
  wire        _GEN_819 = _GEN_4 ? ~_GEN_779 & _GEN_629 : ~_GEN_689 & _GEN_629;
  wire        _GEN_820 = _GEN_4 ? ~_GEN_782 & _GEN_630 : ~_GEN_691 & _GEN_630;
  wire        _GEN_821 = _GEN_4 ? ~_GEN_785 & _GEN_631 : ~_GEN_693 & _GEN_631;
  wire        _GEN_822 = _GEN_4 ? ~_GEN_788 & _GEN_632 : ~_GEN_695 & _GEN_632;
  wire        _GEN_823 = _GEN_4 ? ~_GEN_790 & _GEN_633 : ~_GEN_696 & _GEN_633;
  wire        _GEN_824 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_825 = _GEN_5 & _GEN_824;
  wire        _GEN_826 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_827 = _GEN_5 & _GEN_826;
  wire        _GEN_828 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_829 = _GEN_5 & _GEN_828;
  wire        _GEN_830 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_831 = _GEN_5 & _GEN_830;
  wire        _GEN_832 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_833 = _GEN_5 & _GEN_832;
  wire        _GEN_834 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_835 = _GEN_5 & _GEN_834;
  wire        _GEN_836 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_837 = _GEN_5 & _GEN_836;
  wire        _GEN_838 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_839 = _GEN_5 & _GEN_838;
  wire        _GEN_840 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_841 = _GEN_5 & _GEN_840;
  wire        _GEN_842 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_843 = _GEN_5 & _GEN_842;
  wire        _GEN_844 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_845 = _GEN_5 & _GEN_844;
  wire        _GEN_846 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_847 = _GEN_5 & _GEN_846;
  wire        _GEN_848 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_849 = _GEN_5 & _GEN_848;
  wire        _GEN_850 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_851 = _GEN_5 & _GEN_850;
  wire        _GEN_852 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_853 = _GEN_5 & _GEN_852;
  wire        _GEN_854 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_855 = _GEN_5 & _GEN_854;
  wire        _GEN_856 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_857 = _GEN_5 & _GEN_856;
  wire        _GEN_858 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_859 = _GEN_5 & _GEN_858;
  wire        _GEN_860 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_861 = _GEN_5 & _GEN_860;
  wire        _GEN_862 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_863 = _GEN_5 & _GEN_862;
  wire        _GEN_864 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_865 = _GEN_5 & _GEN_864;
  wire        _GEN_866 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_867 = _GEN_5 & _GEN_866;
  wire        _GEN_868 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_869 = _GEN_5 & _GEN_868;
  wire        _GEN_870 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_871 = _GEN_5 & _GEN_870;
  wire        _GEN_872 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_873 = _GEN_5 & _GEN_872;
  wire        _GEN_874 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_875 = _GEN_5 & _GEN_874;
  wire        _GEN_876 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_877 = _GEN_5 & _GEN_876;
  wire        _GEN_878 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_879 = _GEN_5 & _GEN_878;
  wire        _GEN_880 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_881 = _GEN_5 & _GEN_880;
  wire        _GEN_882 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_883 = _GEN_5 & _GEN_882;
  wire        _GEN_884 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_885 = _GEN_5 & _GEN_884;
  wire        _GEN_886 = _GEN_5 & (&(io_wb_resps_6_bits_uop_rob_idx[6:2]));
  wire        _GEN_887 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_888 = _GEN_887 | _GEN_825;
  wire        _GEN_889 = _GEN_6 ? ~_GEN_888 & _GEN_699 : ~_GEN_825 & _GEN_699;
  wire        _GEN_890 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_891 = _GEN_890 | _GEN_827;
  wire        _GEN_892 = _GEN_6 ? ~_GEN_891 & _GEN_702 : ~_GEN_827 & _GEN_702;
  wire        _GEN_893 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_894 = _GEN_893 | _GEN_829;
  wire        _GEN_895 = _GEN_6 ? ~_GEN_894 & _GEN_705 : ~_GEN_829 & _GEN_705;
  wire        _GEN_896 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_897 = _GEN_896 | _GEN_831;
  wire        _GEN_898 = _GEN_6 ? ~_GEN_897 & _GEN_708 : ~_GEN_831 & _GEN_708;
  wire        _GEN_899 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_900 = _GEN_899 | _GEN_833;
  wire        _GEN_901 = _GEN_6 ? ~_GEN_900 & _GEN_711 : ~_GEN_833 & _GEN_711;
  wire        _GEN_902 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_903 = _GEN_902 | _GEN_835;
  wire        _GEN_904 = _GEN_6 ? ~_GEN_903 & _GEN_714 : ~_GEN_835 & _GEN_714;
  wire        _GEN_905 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_906 = _GEN_905 | _GEN_837;
  wire        _GEN_907 = _GEN_6 ? ~_GEN_906 & _GEN_717 : ~_GEN_837 & _GEN_717;
  wire        _GEN_908 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_909 = _GEN_908 | _GEN_839;
  wire        _GEN_910 = _GEN_6 ? ~_GEN_909 & _GEN_720 : ~_GEN_839 & _GEN_720;
  wire        _GEN_911 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_912 = _GEN_911 | _GEN_841;
  wire        _GEN_913 = _GEN_6 ? ~_GEN_912 & _GEN_723 : ~_GEN_841 & _GEN_723;
  wire        _GEN_914 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_915 = _GEN_914 | _GEN_843;
  wire        _GEN_916 = _GEN_6 ? ~_GEN_915 & _GEN_726 : ~_GEN_843 & _GEN_726;
  wire        _GEN_917 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_918 = _GEN_917 | _GEN_845;
  wire        _GEN_919 = _GEN_6 ? ~_GEN_918 & _GEN_729 : ~_GEN_845 & _GEN_729;
  wire        _GEN_920 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_921 = _GEN_920 | _GEN_847;
  wire        _GEN_922 = _GEN_6 ? ~_GEN_921 & _GEN_732 : ~_GEN_847 & _GEN_732;
  wire        _GEN_923 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_924 = _GEN_923 | _GEN_849;
  wire        _GEN_925 = _GEN_6 ? ~_GEN_924 & _GEN_735 : ~_GEN_849 & _GEN_735;
  wire        _GEN_926 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_927 = _GEN_926 | _GEN_851;
  wire        _GEN_928 = _GEN_6 ? ~_GEN_927 & _GEN_738 : ~_GEN_851 & _GEN_738;
  wire        _GEN_929 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_930 = _GEN_929 | _GEN_853;
  wire        _GEN_931 = _GEN_6 ? ~_GEN_930 & _GEN_741 : ~_GEN_853 & _GEN_741;
  wire        _GEN_932 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_933 = _GEN_932 | _GEN_855;
  wire        _GEN_934 = _GEN_6 ? ~_GEN_933 & _GEN_744 : ~_GEN_855 & _GEN_744;
  wire        _GEN_935 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_936 = _GEN_935 | _GEN_857;
  wire        _GEN_937 = _GEN_6 ? ~_GEN_936 & _GEN_747 : ~_GEN_857 & _GEN_747;
  wire        _GEN_938 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_939 = _GEN_938 | _GEN_859;
  wire        _GEN_940 = _GEN_6 ? ~_GEN_939 & _GEN_750 : ~_GEN_859 & _GEN_750;
  wire        _GEN_941 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_942 = _GEN_941 | _GEN_861;
  wire        _GEN_943 = _GEN_6 ? ~_GEN_942 & _GEN_753 : ~_GEN_861 & _GEN_753;
  wire        _GEN_944 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_945 = _GEN_944 | _GEN_863;
  wire        _GEN_946 = _GEN_6 ? ~_GEN_945 & _GEN_756 : ~_GEN_863 & _GEN_756;
  wire        _GEN_947 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_948 = _GEN_947 | _GEN_865;
  wire        _GEN_949 = _GEN_6 ? ~_GEN_948 & _GEN_759 : ~_GEN_865 & _GEN_759;
  wire        _GEN_950 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_951 = _GEN_950 | _GEN_867;
  wire        _GEN_952 = _GEN_6 ? ~_GEN_951 & _GEN_762 : ~_GEN_867 & _GEN_762;
  wire        _GEN_953 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_954 = _GEN_953 | _GEN_869;
  wire        _GEN_955 = _GEN_6 ? ~_GEN_954 & _GEN_765 : ~_GEN_869 & _GEN_765;
  wire        _GEN_956 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_957 = _GEN_956 | _GEN_871;
  wire        _GEN_958 = _GEN_6 ? ~_GEN_957 & _GEN_768 : ~_GEN_871 & _GEN_768;
  wire        _GEN_959 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_960 = _GEN_959 | _GEN_873;
  wire        _GEN_961 = _GEN_6 ? ~_GEN_960 & _GEN_771 : ~_GEN_873 & _GEN_771;
  wire        _GEN_962 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_963 = _GEN_962 | _GEN_875;
  wire        _GEN_964 = _GEN_6 ? ~_GEN_963 & _GEN_774 : ~_GEN_875 & _GEN_774;
  wire        _GEN_965 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_966 = _GEN_965 | _GEN_877;
  wire        _GEN_967 = _GEN_6 ? ~_GEN_966 & _GEN_777 : ~_GEN_877 & _GEN_777;
  wire        _GEN_968 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_969 = _GEN_968 | _GEN_879;
  wire        _GEN_970 = _GEN_6 ? ~_GEN_969 & _GEN_780 : ~_GEN_879 & _GEN_780;
  wire        _GEN_971 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_972 = _GEN_971 | _GEN_881;
  wire        _GEN_973 = _GEN_6 ? ~_GEN_972 & _GEN_783 : ~_GEN_881 & _GEN_783;
  wire        _GEN_974 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_975 = _GEN_974 | _GEN_883;
  wire        _GEN_976 = _GEN_6 ? ~_GEN_975 & _GEN_786 : ~_GEN_883 & _GEN_786;
  wire        _GEN_977 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_978 = _GEN_977 | _GEN_885;
  wire        _GEN_979 = _GEN_6 ? ~_GEN_978 & _GEN_789 : ~_GEN_885 & _GEN_789;
  wire        _GEN_980 = (&(io_wb_resps_7_bits_uop_rob_idx[6:2])) | _GEN_886;
  wire        _GEN_981 = _GEN_6 ? ~_GEN_980 & _GEN_791 : ~_GEN_886 & _GEN_791;
  wire        _GEN_982 = _GEN_6 ? ~_GEN_888 & _GEN_792 : ~_GEN_825 & _GEN_792;
  wire        _GEN_983 = _GEN_6 ? ~_GEN_891 & _GEN_793 : ~_GEN_827 & _GEN_793;
  wire        _GEN_984 = _GEN_6 ? ~_GEN_894 & _GEN_794 : ~_GEN_829 & _GEN_794;
  wire        _GEN_985 = _GEN_6 ? ~_GEN_897 & _GEN_795 : ~_GEN_831 & _GEN_795;
  wire        _GEN_986 = _GEN_6 ? ~_GEN_900 & _GEN_796 : ~_GEN_833 & _GEN_796;
  wire        _GEN_987 = _GEN_6 ? ~_GEN_903 & _GEN_797 : ~_GEN_835 & _GEN_797;
  wire        _GEN_988 = _GEN_6 ? ~_GEN_906 & _GEN_798 : ~_GEN_837 & _GEN_798;
  wire        _GEN_989 = _GEN_6 ? ~_GEN_909 & _GEN_799 : ~_GEN_839 & _GEN_799;
  wire        _GEN_990 = _GEN_6 ? ~_GEN_912 & _GEN_800 : ~_GEN_841 & _GEN_800;
  wire        _GEN_991 = _GEN_6 ? ~_GEN_915 & _GEN_801 : ~_GEN_843 & _GEN_801;
  wire        _GEN_992 = _GEN_6 ? ~_GEN_918 & _GEN_802 : ~_GEN_845 & _GEN_802;
  wire        _GEN_993 = _GEN_6 ? ~_GEN_921 & _GEN_803 : ~_GEN_847 & _GEN_803;
  wire        _GEN_994 = _GEN_6 ? ~_GEN_924 & _GEN_804 : ~_GEN_849 & _GEN_804;
  wire        _GEN_995 = _GEN_6 ? ~_GEN_927 & _GEN_805 : ~_GEN_851 & _GEN_805;
  wire        _GEN_996 = _GEN_6 ? ~_GEN_930 & _GEN_806 : ~_GEN_853 & _GEN_806;
  wire        _GEN_997 = _GEN_6 ? ~_GEN_933 & _GEN_807 : ~_GEN_855 & _GEN_807;
  wire        _GEN_998 = _GEN_6 ? ~_GEN_936 & _GEN_808 : ~_GEN_857 & _GEN_808;
  wire        _GEN_999 = _GEN_6 ? ~_GEN_939 & _GEN_809 : ~_GEN_859 & _GEN_809;
  wire        _GEN_1000 = _GEN_6 ? ~_GEN_942 & _GEN_810 : ~_GEN_861 & _GEN_810;
  wire        _GEN_1001 = _GEN_6 ? ~_GEN_945 & _GEN_811 : ~_GEN_863 & _GEN_811;
  wire        _GEN_1002 = _GEN_6 ? ~_GEN_948 & _GEN_812 : ~_GEN_865 & _GEN_812;
  wire        _GEN_1003 = _GEN_6 ? ~_GEN_951 & _GEN_813 : ~_GEN_867 & _GEN_813;
  wire        _GEN_1004 = _GEN_6 ? ~_GEN_954 & _GEN_814 : ~_GEN_869 & _GEN_814;
  wire        _GEN_1005 = _GEN_6 ? ~_GEN_957 & _GEN_815 : ~_GEN_871 & _GEN_815;
  wire        _GEN_1006 = _GEN_6 ? ~_GEN_960 & _GEN_816 : ~_GEN_873 & _GEN_816;
  wire        _GEN_1007 = _GEN_6 ? ~_GEN_963 & _GEN_817 : ~_GEN_875 & _GEN_817;
  wire        _GEN_1008 = _GEN_6 ? ~_GEN_966 & _GEN_818 : ~_GEN_877 & _GEN_818;
  wire        _GEN_1009 = _GEN_6 ? ~_GEN_969 & _GEN_819 : ~_GEN_879 & _GEN_819;
  wire        _GEN_1010 = _GEN_6 ? ~_GEN_972 & _GEN_820 : ~_GEN_881 & _GEN_820;
  wire        _GEN_1011 = _GEN_6 ? ~_GEN_975 & _GEN_821 : ~_GEN_883 & _GEN_821;
  wire        _GEN_1012 = _GEN_6 ? ~_GEN_978 & _GEN_822 : ~_GEN_885 & _GEN_822;
  wire        _GEN_1013 = _GEN_6 ? ~_GEN_980 & _GEN_823 : ~_GEN_886 & _GEN_823;
  wire        _GEN_1014 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_1015 = _GEN_7 & _GEN_1014;
  wire        _GEN_1016 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_1017 = _GEN_7 & _GEN_1016;
  wire        _GEN_1018 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_1019 = _GEN_7 & _GEN_1018;
  wire        _GEN_1020 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_1021 = _GEN_7 & _GEN_1020;
  wire        _GEN_1022 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_1023 = _GEN_7 & _GEN_1022;
  wire        _GEN_1024 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_1025 = _GEN_7 & _GEN_1024;
  wire        _GEN_1026 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_1027 = _GEN_7 & _GEN_1026;
  wire        _GEN_1028 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_1029 = _GEN_7 & _GEN_1028;
  wire        _GEN_1030 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_1031 = _GEN_7 & _GEN_1030;
  wire        _GEN_1032 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_1033 = _GEN_7 & _GEN_1032;
  wire        _GEN_1034 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_1035 = _GEN_7 & _GEN_1034;
  wire        _GEN_1036 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_1037 = _GEN_7 & _GEN_1036;
  wire        _GEN_1038 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_1039 = _GEN_7 & _GEN_1038;
  wire        _GEN_1040 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_1041 = _GEN_7 & _GEN_1040;
  wire        _GEN_1042 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_1043 = _GEN_7 & _GEN_1042;
  wire        _GEN_1044 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_1045 = _GEN_7 & _GEN_1044;
  wire        _GEN_1046 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_1047 = _GEN_7 & _GEN_1046;
  wire        _GEN_1048 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_1049 = _GEN_7 & _GEN_1048;
  wire        _GEN_1050 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_1051 = _GEN_7 & _GEN_1050;
  wire        _GEN_1052 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_1053 = _GEN_7 & _GEN_1052;
  wire        _GEN_1054 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_1055 = _GEN_7 & _GEN_1054;
  wire        _GEN_1056 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_1057 = _GEN_7 & _GEN_1056;
  wire        _GEN_1058 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_1059 = _GEN_7 & _GEN_1058;
  wire        _GEN_1060 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_1061 = _GEN_7 & _GEN_1060;
  wire        _GEN_1062 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_1063 = _GEN_7 & _GEN_1062;
  wire        _GEN_1064 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_1065 = _GEN_7 & _GEN_1064;
  wire        _GEN_1066 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_1067 = _GEN_7 & _GEN_1066;
  wire        _GEN_1068 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_1069 = _GEN_7 & _GEN_1068;
  wire        _GEN_1070 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_1071 = _GEN_7 & _GEN_1070;
  wire        _GEN_1072 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_1073 = _GEN_7 & _GEN_1072;
  wire        _GEN_1074 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_1075 = _GEN_7 & _GEN_1074;
  wire        _GEN_1076 = _GEN_7 & (&(io_wb_resps_8_bits_uop_rob_idx[6:2]));
  wire        _GEN_1077 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_1078 = _GEN_1077 | _GEN_1015;
  wire        _GEN_1079 = _GEN_8 ? ~_GEN_1078 & _GEN_889 : ~_GEN_1015 & _GEN_889;
  wire        _GEN_1080 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_1081 = _GEN_1080 | _GEN_1017;
  wire        _GEN_1082 = _GEN_8 ? ~_GEN_1081 & _GEN_892 : ~_GEN_1017 & _GEN_892;
  wire        _GEN_1083 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_1084 = _GEN_1083 | _GEN_1019;
  wire        _GEN_1085 = _GEN_8 ? ~_GEN_1084 & _GEN_895 : ~_GEN_1019 & _GEN_895;
  wire        _GEN_1086 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_1087 = _GEN_1086 | _GEN_1021;
  wire        _GEN_1088 = _GEN_8 ? ~_GEN_1087 & _GEN_898 : ~_GEN_1021 & _GEN_898;
  wire        _GEN_1089 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_1090 = _GEN_1089 | _GEN_1023;
  wire        _GEN_1091 = _GEN_8 ? ~_GEN_1090 & _GEN_901 : ~_GEN_1023 & _GEN_901;
  wire        _GEN_1092 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_1093 = _GEN_1092 | _GEN_1025;
  wire        _GEN_1094 = _GEN_8 ? ~_GEN_1093 & _GEN_904 : ~_GEN_1025 & _GEN_904;
  wire        _GEN_1095 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_1096 = _GEN_1095 | _GEN_1027;
  wire        _GEN_1097 = _GEN_8 ? ~_GEN_1096 & _GEN_907 : ~_GEN_1027 & _GEN_907;
  wire        _GEN_1098 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_1099 = _GEN_1098 | _GEN_1029;
  wire        _GEN_1100 = _GEN_8 ? ~_GEN_1099 & _GEN_910 : ~_GEN_1029 & _GEN_910;
  wire        _GEN_1101 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_1102 = _GEN_1101 | _GEN_1031;
  wire        _GEN_1103 = _GEN_8 ? ~_GEN_1102 & _GEN_913 : ~_GEN_1031 & _GEN_913;
  wire        _GEN_1104 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_1105 = _GEN_1104 | _GEN_1033;
  wire        _GEN_1106 = _GEN_8 ? ~_GEN_1105 & _GEN_916 : ~_GEN_1033 & _GEN_916;
  wire        _GEN_1107 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_1108 = _GEN_1107 | _GEN_1035;
  wire        _GEN_1109 = _GEN_8 ? ~_GEN_1108 & _GEN_919 : ~_GEN_1035 & _GEN_919;
  wire        _GEN_1110 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_1111 = _GEN_1110 | _GEN_1037;
  wire        _GEN_1112 = _GEN_8 ? ~_GEN_1111 & _GEN_922 : ~_GEN_1037 & _GEN_922;
  wire        _GEN_1113 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_1114 = _GEN_1113 | _GEN_1039;
  wire        _GEN_1115 = _GEN_8 ? ~_GEN_1114 & _GEN_925 : ~_GEN_1039 & _GEN_925;
  wire        _GEN_1116 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_1117 = _GEN_1116 | _GEN_1041;
  wire        _GEN_1118 = _GEN_8 ? ~_GEN_1117 & _GEN_928 : ~_GEN_1041 & _GEN_928;
  wire        _GEN_1119 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_1120 = _GEN_1119 | _GEN_1043;
  wire        _GEN_1121 = _GEN_8 ? ~_GEN_1120 & _GEN_931 : ~_GEN_1043 & _GEN_931;
  wire        _GEN_1122 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_1123 = _GEN_1122 | _GEN_1045;
  wire        _GEN_1124 = _GEN_8 ? ~_GEN_1123 & _GEN_934 : ~_GEN_1045 & _GEN_934;
  wire        _GEN_1125 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_1126 = _GEN_1125 | _GEN_1047;
  wire        _GEN_1127 = _GEN_8 ? ~_GEN_1126 & _GEN_937 : ~_GEN_1047 & _GEN_937;
  wire        _GEN_1128 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_1129 = _GEN_1128 | _GEN_1049;
  wire        _GEN_1130 = _GEN_8 ? ~_GEN_1129 & _GEN_940 : ~_GEN_1049 & _GEN_940;
  wire        _GEN_1131 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_1132 = _GEN_1131 | _GEN_1051;
  wire        _GEN_1133 = _GEN_8 ? ~_GEN_1132 & _GEN_943 : ~_GEN_1051 & _GEN_943;
  wire        _GEN_1134 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_1135 = _GEN_1134 | _GEN_1053;
  wire        _GEN_1136 = _GEN_8 ? ~_GEN_1135 & _GEN_946 : ~_GEN_1053 & _GEN_946;
  wire        _GEN_1137 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_1138 = _GEN_1137 | _GEN_1055;
  wire        _GEN_1139 = _GEN_8 ? ~_GEN_1138 & _GEN_949 : ~_GEN_1055 & _GEN_949;
  wire        _GEN_1140 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_1141 = _GEN_1140 | _GEN_1057;
  wire        _GEN_1142 = _GEN_8 ? ~_GEN_1141 & _GEN_952 : ~_GEN_1057 & _GEN_952;
  wire        _GEN_1143 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_1144 = _GEN_1143 | _GEN_1059;
  wire        _GEN_1145 = _GEN_8 ? ~_GEN_1144 & _GEN_955 : ~_GEN_1059 & _GEN_955;
  wire        _GEN_1146 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_1147 = _GEN_1146 | _GEN_1061;
  wire        _GEN_1148 = _GEN_8 ? ~_GEN_1147 & _GEN_958 : ~_GEN_1061 & _GEN_958;
  wire        _GEN_1149 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_1150 = _GEN_1149 | _GEN_1063;
  wire        _GEN_1151 = _GEN_8 ? ~_GEN_1150 & _GEN_961 : ~_GEN_1063 & _GEN_961;
  wire        _GEN_1152 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_1153 = _GEN_1152 | _GEN_1065;
  wire        _GEN_1154 = _GEN_8 ? ~_GEN_1153 & _GEN_964 : ~_GEN_1065 & _GEN_964;
  wire        _GEN_1155 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_1156 = _GEN_1155 | _GEN_1067;
  wire        _GEN_1157 = _GEN_8 ? ~_GEN_1156 & _GEN_967 : ~_GEN_1067 & _GEN_967;
  wire        _GEN_1158 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_1159 = _GEN_1158 | _GEN_1069;
  wire        _GEN_1160 = _GEN_8 ? ~_GEN_1159 & _GEN_970 : ~_GEN_1069 & _GEN_970;
  wire        _GEN_1161 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_1162 = _GEN_1161 | _GEN_1071;
  wire        _GEN_1163 = _GEN_8 ? ~_GEN_1162 & _GEN_973 : ~_GEN_1071 & _GEN_973;
  wire        _GEN_1164 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_1165 = _GEN_1164 | _GEN_1073;
  wire        _GEN_1166 = _GEN_8 ? ~_GEN_1165 & _GEN_976 : ~_GEN_1073 & _GEN_976;
  wire        _GEN_1167 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_1168 = _GEN_1167 | _GEN_1075;
  wire        _GEN_1169 = _GEN_8 ? ~_GEN_1168 & _GEN_979 : ~_GEN_1075 & _GEN_979;
  wire        _GEN_1170 = (&(io_wb_resps_9_bits_uop_rob_idx[6:2])) | _GEN_1076;
  wire        _GEN_1171 = _GEN_8 ? ~_GEN_1170 & _GEN_981 : ~_GEN_1076 & _GEN_981;
  wire        _GEN_1172 = _GEN_8 ? ~_GEN_1078 & _GEN_982 : ~_GEN_1015 & _GEN_982;
  wire        _GEN_1173 = _GEN_8 ? ~_GEN_1081 & _GEN_983 : ~_GEN_1017 & _GEN_983;
  wire        _GEN_1174 = _GEN_8 ? ~_GEN_1084 & _GEN_984 : ~_GEN_1019 & _GEN_984;
  wire        _GEN_1175 = _GEN_8 ? ~_GEN_1087 & _GEN_985 : ~_GEN_1021 & _GEN_985;
  wire        _GEN_1176 = _GEN_8 ? ~_GEN_1090 & _GEN_986 : ~_GEN_1023 & _GEN_986;
  wire        _GEN_1177 = _GEN_8 ? ~_GEN_1093 & _GEN_987 : ~_GEN_1025 & _GEN_987;
  wire        _GEN_1178 = _GEN_8 ? ~_GEN_1096 & _GEN_988 : ~_GEN_1027 & _GEN_988;
  wire        _GEN_1179 = _GEN_8 ? ~_GEN_1099 & _GEN_989 : ~_GEN_1029 & _GEN_989;
  wire        _GEN_1180 = _GEN_8 ? ~_GEN_1102 & _GEN_990 : ~_GEN_1031 & _GEN_990;
  wire        _GEN_1181 = _GEN_8 ? ~_GEN_1105 & _GEN_991 : ~_GEN_1033 & _GEN_991;
  wire        _GEN_1182 = _GEN_8 ? ~_GEN_1108 & _GEN_992 : ~_GEN_1035 & _GEN_992;
  wire        _GEN_1183 = _GEN_8 ? ~_GEN_1111 & _GEN_993 : ~_GEN_1037 & _GEN_993;
  wire        _GEN_1184 = _GEN_8 ? ~_GEN_1114 & _GEN_994 : ~_GEN_1039 & _GEN_994;
  wire        _GEN_1185 = _GEN_8 ? ~_GEN_1117 & _GEN_995 : ~_GEN_1041 & _GEN_995;
  wire        _GEN_1186 = _GEN_8 ? ~_GEN_1120 & _GEN_996 : ~_GEN_1043 & _GEN_996;
  wire        _GEN_1187 = _GEN_8 ? ~_GEN_1123 & _GEN_997 : ~_GEN_1045 & _GEN_997;
  wire        _GEN_1188 = _GEN_8 ? ~_GEN_1126 & _GEN_998 : ~_GEN_1047 & _GEN_998;
  wire        _GEN_1189 = _GEN_8 ? ~_GEN_1129 & _GEN_999 : ~_GEN_1049 & _GEN_999;
  wire        _GEN_1190 = _GEN_8 ? ~_GEN_1132 & _GEN_1000 : ~_GEN_1051 & _GEN_1000;
  wire        _GEN_1191 = _GEN_8 ? ~_GEN_1135 & _GEN_1001 : ~_GEN_1053 & _GEN_1001;
  wire        _GEN_1192 = _GEN_8 ? ~_GEN_1138 & _GEN_1002 : ~_GEN_1055 & _GEN_1002;
  wire        _GEN_1193 = _GEN_8 ? ~_GEN_1141 & _GEN_1003 : ~_GEN_1057 & _GEN_1003;
  wire        _GEN_1194 = _GEN_8 ? ~_GEN_1144 & _GEN_1004 : ~_GEN_1059 & _GEN_1004;
  wire        _GEN_1195 = _GEN_8 ? ~_GEN_1147 & _GEN_1005 : ~_GEN_1061 & _GEN_1005;
  wire        _GEN_1196 = _GEN_8 ? ~_GEN_1150 & _GEN_1006 : ~_GEN_1063 & _GEN_1006;
  wire        _GEN_1197 = _GEN_8 ? ~_GEN_1153 & _GEN_1007 : ~_GEN_1065 & _GEN_1007;
  wire        _GEN_1198 = _GEN_8 ? ~_GEN_1156 & _GEN_1008 : ~_GEN_1067 & _GEN_1008;
  wire        _GEN_1199 = _GEN_8 ? ~_GEN_1159 & _GEN_1009 : ~_GEN_1069 & _GEN_1009;
  wire        _GEN_1200 = _GEN_8 ? ~_GEN_1162 & _GEN_1010 : ~_GEN_1071 & _GEN_1010;
  wire        _GEN_1201 = _GEN_8 ? ~_GEN_1165 & _GEN_1011 : ~_GEN_1073 & _GEN_1011;
  wire        _GEN_1202 = _GEN_8 ? ~_GEN_1168 & _GEN_1012 : ~_GEN_1075 & _GEN_1012;
  wire        _GEN_1203 = _GEN_8 ? ~_GEN_1170 & _GEN_1013 : ~_GEN_1076 & _GEN_1013;
  wire        _GEN_1204 = io_lsu_clr_bsy_0_bits[6:2] == 5'h0;
  wire        _GEN_1205 = _GEN_9 & _GEN_1204;
  wire        _GEN_1206 = io_lsu_clr_bsy_0_bits[6:2] == 5'h1;
  wire        _GEN_1207 = _GEN_9 & _GEN_1206;
  wire        _GEN_1208 = io_lsu_clr_bsy_0_bits[6:2] == 5'h2;
  wire        _GEN_1209 = _GEN_9 & _GEN_1208;
  wire        _GEN_1210 = io_lsu_clr_bsy_0_bits[6:2] == 5'h3;
  wire        _GEN_1211 = _GEN_9 & _GEN_1210;
  wire        _GEN_1212 = io_lsu_clr_bsy_0_bits[6:2] == 5'h4;
  wire        _GEN_1213 = _GEN_9 & _GEN_1212;
  wire        _GEN_1214 = io_lsu_clr_bsy_0_bits[6:2] == 5'h5;
  wire        _GEN_1215 = _GEN_9 & _GEN_1214;
  wire        _GEN_1216 = io_lsu_clr_bsy_0_bits[6:2] == 5'h6;
  wire        _GEN_1217 = _GEN_9 & _GEN_1216;
  wire        _GEN_1218 = io_lsu_clr_bsy_0_bits[6:2] == 5'h7;
  wire        _GEN_1219 = _GEN_9 & _GEN_1218;
  wire        _GEN_1220 = io_lsu_clr_bsy_0_bits[6:2] == 5'h8;
  wire        _GEN_1221 = _GEN_9 & _GEN_1220;
  wire        _GEN_1222 = io_lsu_clr_bsy_0_bits[6:2] == 5'h9;
  wire        _GEN_1223 = _GEN_9 & _GEN_1222;
  wire        _GEN_1224 = io_lsu_clr_bsy_0_bits[6:2] == 5'hA;
  wire        _GEN_1225 = _GEN_9 & _GEN_1224;
  wire        _GEN_1226 = io_lsu_clr_bsy_0_bits[6:2] == 5'hB;
  wire        _GEN_1227 = _GEN_9 & _GEN_1226;
  wire        _GEN_1228 = io_lsu_clr_bsy_0_bits[6:2] == 5'hC;
  wire        _GEN_1229 = _GEN_9 & _GEN_1228;
  wire        _GEN_1230 = io_lsu_clr_bsy_0_bits[6:2] == 5'hD;
  wire        _GEN_1231 = _GEN_9 & _GEN_1230;
  wire        _GEN_1232 = io_lsu_clr_bsy_0_bits[6:2] == 5'hE;
  wire        _GEN_1233 = _GEN_9 & _GEN_1232;
  wire        _GEN_1234 = io_lsu_clr_bsy_0_bits[6:2] == 5'hF;
  wire        _GEN_1235 = _GEN_9 & _GEN_1234;
  wire        _GEN_1236 = io_lsu_clr_bsy_0_bits[6:2] == 5'h10;
  wire        _GEN_1237 = _GEN_9 & _GEN_1236;
  wire        _GEN_1238 = io_lsu_clr_bsy_0_bits[6:2] == 5'h11;
  wire        _GEN_1239 = _GEN_9 & _GEN_1238;
  wire        _GEN_1240 = io_lsu_clr_bsy_0_bits[6:2] == 5'h12;
  wire        _GEN_1241 = _GEN_9 & _GEN_1240;
  wire        _GEN_1242 = io_lsu_clr_bsy_0_bits[6:2] == 5'h13;
  wire        _GEN_1243 = _GEN_9 & _GEN_1242;
  wire        _GEN_1244 = io_lsu_clr_bsy_0_bits[6:2] == 5'h14;
  wire        _GEN_1245 = _GEN_9 & _GEN_1244;
  wire        _GEN_1246 = io_lsu_clr_bsy_0_bits[6:2] == 5'h15;
  wire        _GEN_1247 = _GEN_9 & _GEN_1246;
  wire        _GEN_1248 = io_lsu_clr_bsy_0_bits[6:2] == 5'h16;
  wire        _GEN_1249 = _GEN_9 & _GEN_1248;
  wire        _GEN_1250 = io_lsu_clr_bsy_0_bits[6:2] == 5'h17;
  wire        _GEN_1251 = _GEN_9 & _GEN_1250;
  wire        _GEN_1252 = io_lsu_clr_bsy_0_bits[6:2] == 5'h18;
  wire        _GEN_1253 = _GEN_9 & _GEN_1252;
  wire        _GEN_1254 = io_lsu_clr_bsy_0_bits[6:2] == 5'h19;
  wire        _GEN_1255 = _GEN_9 & _GEN_1254;
  wire        _GEN_1256 = io_lsu_clr_bsy_0_bits[6:2] == 5'h1A;
  wire        _GEN_1257 = _GEN_9 & _GEN_1256;
  wire        _GEN_1258 = io_lsu_clr_bsy_0_bits[6:2] == 5'h1B;
  wire        _GEN_1259 = _GEN_9 & _GEN_1258;
  wire        _GEN_1260 = io_lsu_clr_bsy_0_bits[6:2] == 5'h1C;
  wire        _GEN_1261 = _GEN_9 & _GEN_1260;
  wire        _GEN_1262 = io_lsu_clr_bsy_0_bits[6:2] == 5'h1D;
  wire        _GEN_1263 = _GEN_9 & _GEN_1262;
  wire        _GEN_1264 = io_lsu_clr_bsy_0_bits[6:2] == 5'h1E;
  wire        _GEN_1265 = _GEN_9 & _GEN_1264;
  wire        _GEN_1266 = _GEN_9 & (&(io_lsu_clr_bsy_0_bits[6:2]));
  wire        _GEN_1267 = io_lsu_clr_bsy_1_bits[6:2] == 5'h0;
  wire        _GEN_1268 = _GEN_1267 | _GEN_1205;
  wire        _GEN_1269 = io_lsu_clr_bsy_1_bits[6:2] == 5'h1;
  wire        _GEN_1270 = _GEN_1269 | _GEN_1207;
  wire        _GEN_1271 = io_lsu_clr_bsy_1_bits[6:2] == 5'h2;
  wire        _GEN_1272 = _GEN_1271 | _GEN_1209;
  wire        _GEN_1273 = io_lsu_clr_bsy_1_bits[6:2] == 5'h3;
  wire        _GEN_1274 = _GEN_1273 | _GEN_1211;
  wire        _GEN_1275 = io_lsu_clr_bsy_1_bits[6:2] == 5'h4;
  wire        _GEN_1276 = _GEN_1275 | _GEN_1213;
  wire        _GEN_1277 = io_lsu_clr_bsy_1_bits[6:2] == 5'h5;
  wire        _GEN_1278 = _GEN_1277 | _GEN_1215;
  wire        _GEN_1279 = io_lsu_clr_bsy_1_bits[6:2] == 5'h6;
  wire        _GEN_1280 = _GEN_1279 | _GEN_1217;
  wire        _GEN_1281 = io_lsu_clr_bsy_1_bits[6:2] == 5'h7;
  wire        _GEN_1282 = _GEN_1281 | _GEN_1219;
  wire        _GEN_1283 = io_lsu_clr_bsy_1_bits[6:2] == 5'h8;
  wire        _GEN_1284 = _GEN_1283 | _GEN_1221;
  wire        _GEN_1285 = io_lsu_clr_bsy_1_bits[6:2] == 5'h9;
  wire        _GEN_1286 = _GEN_1285 | _GEN_1223;
  wire        _GEN_1287 = io_lsu_clr_bsy_1_bits[6:2] == 5'hA;
  wire        _GEN_1288 = _GEN_1287 | _GEN_1225;
  wire        _GEN_1289 = io_lsu_clr_bsy_1_bits[6:2] == 5'hB;
  wire        _GEN_1290 = _GEN_1289 | _GEN_1227;
  wire        _GEN_1291 = io_lsu_clr_bsy_1_bits[6:2] == 5'hC;
  wire        _GEN_1292 = _GEN_1291 | _GEN_1229;
  wire        _GEN_1293 = io_lsu_clr_bsy_1_bits[6:2] == 5'hD;
  wire        _GEN_1294 = _GEN_1293 | _GEN_1231;
  wire        _GEN_1295 = io_lsu_clr_bsy_1_bits[6:2] == 5'hE;
  wire        _GEN_1296 = _GEN_1295 | _GEN_1233;
  wire        _GEN_1297 = io_lsu_clr_bsy_1_bits[6:2] == 5'hF;
  wire        _GEN_1298 = _GEN_1297 | _GEN_1235;
  wire        _GEN_1299 = io_lsu_clr_bsy_1_bits[6:2] == 5'h10;
  wire        _GEN_1300 = _GEN_1299 | _GEN_1237;
  wire        _GEN_1301 = io_lsu_clr_bsy_1_bits[6:2] == 5'h11;
  wire        _GEN_1302 = _GEN_1301 | _GEN_1239;
  wire        _GEN_1303 = io_lsu_clr_bsy_1_bits[6:2] == 5'h12;
  wire        _GEN_1304 = _GEN_1303 | _GEN_1241;
  wire        _GEN_1305 = io_lsu_clr_bsy_1_bits[6:2] == 5'h13;
  wire        _GEN_1306 = _GEN_1305 | _GEN_1243;
  wire        _GEN_1307 = io_lsu_clr_bsy_1_bits[6:2] == 5'h14;
  wire        _GEN_1308 = _GEN_1307 | _GEN_1245;
  wire        _GEN_1309 = io_lsu_clr_bsy_1_bits[6:2] == 5'h15;
  wire        _GEN_1310 = _GEN_1309 | _GEN_1247;
  wire        _GEN_1311 = io_lsu_clr_bsy_1_bits[6:2] == 5'h16;
  wire        _GEN_1312 = _GEN_1311 | _GEN_1249;
  wire        _GEN_1313 = io_lsu_clr_bsy_1_bits[6:2] == 5'h17;
  wire        _GEN_1314 = _GEN_1313 | _GEN_1251;
  wire        _GEN_1315 = io_lsu_clr_bsy_1_bits[6:2] == 5'h18;
  wire        _GEN_1316 = _GEN_1315 | _GEN_1253;
  wire        _GEN_1317 = io_lsu_clr_bsy_1_bits[6:2] == 5'h19;
  wire        _GEN_1318 = _GEN_1317 | _GEN_1255;
  wire        _GEN_1319 = io_lsu_clr_bsy_1_bits[6:2] == 5'h1A;
  wire        _GEN_1320 = _GEN_1319 | _GEN_1257;
  wire        _GEN_1321 = io_lsu_clr_bsy_1_bits[6:2] == 5'h1B;
  wire        _GEN_1322 = _GEN_1321 | _GEN_1259;
  wire        _GEN_1323 = io_lsu_clr_bsy_1_bits[6:2] == 5'h1C;
  wire        _GEN_1324 = _GEN_1323 | _GEN_1261;
  wire        _GEN_1325 = io_lsu_clr_bsy_1_bits[6:2] == 5'h1D;
  wire        _GEN_1326 = _GEN_1325 | _GEN_1263;
  wire        _GEN_1327 = io_lsu_clr_bsy_1_bits[6:2] == 5'h1E;
  wire        _GEN_1328 = _GEN_1327 | _GEN_1265;
  wire        _GEN_1329 = (&(io_lsu_clr_bsy_1_bits[6:2])) | _GEN_1266;
  wire        _GEN_1330 = io_lsu_clr_bsy_2_bits[6:2] == 5'h0;
  wire        _GEN_1331 = _GEN_11 & _GEN_1330;
  wire        _GEN_1332 = io_lsu_clr_bsy_2_bits[6:2] == 5'h1;
  wire        _GEN_1333 = _GEN_11 & _GEN_1332;
  wire        _GEN_1334 = io_lsu_clr_bsy_2_bits[6:2] == 5'h2;
  wire        _GEN_1335 = _GEN_11 & _GEN_1334;
  wire        _GEN_1336 = io_lsu_clr_bsy_2_bits[6:2] == 5'h3;
  wire        _GEN_1337 = _GEN_11 & _GEN_1336;
  wire        _GEN_1338 = io_lsu_clr_bsy_2_bits[6:2] == 5'h4;
  wire        _GEN_1339 = _GEN_11 & _GEN_1338;
  wire        _GEN_1340 = io_lsu_clr_bsy_2_bits[6:2] == 5'h5;
  wire        _GEN_1341 = _GEN_11 & _GEN_1340;
  wire        _GEN_1342 = io_lsu_clr_bsy_2_bits[6:2] == 5'h6;
  wire        _GEN_1343 = _GEN_11 & _GEN_1342;
  wire        _GEN_1344 = io_lsu_clr_bsy_2_bits[6:2] == 5'h7;
  wire        _GEN_1345 = _GEN_11 & _GEN_1344;
  wire        _GEN_1346 = io_lsu_clr_bsy_2_bits[6:2] == 5'h8;
  wire        _GEN_1347 = _GEN_11 & _GEN_1346;
  wire        _GEN_1348 = io_lsu_clr_bsy_2_bits[6:2] == 5'h9;
  wire        _GEN_1349 = _GEN_11 & _GEN_1348;
  wire        _GEN_1350 = io_lsu_clr_bsy_2_bits[6:2] == 5'hA;
  wire        _GEN_1351 = _GEN_11 & _GEN_1350;
  wire        _GEN_1352 = io_lsu_clr_bsy_2_bits[6:2] == 5'hB;
  wire        _GEN_1353 = _GEN_11 & _GEN_1352;
  wire        _GEN_1354 = io_lsu_clr_bsy_2_bits[6:2] == 5'hC;
  wire        _GEN_1355 = _GEN_11 & _GEN_1354;
  wire        _GEN_1356 = io_lsu_clr_bsy_2_bits[6:2] == 5'hD;
  wire        _GEN_1357 = _GEN_11 & _GEN_1356;
  wire        _GEN_1358 = io_lsu_clr_bsy_2_bits[6:2] == 5'hE;
  wire        _GEN_1359 = _GEN_11 & _GEN_1358;
  wire        _GEN_1360 = io_lsu_clr_bsy_2_bits[6:2] == 5'hF;
  wire        _GEN_1361 = _GEN_11 & _GEN_1360;
  wire        _GEN_1362 = io_lsu_clr_bsy_2_bits[6:2] == 5'h10;
  wire        _GEN_1363 = _GEN_11 & _GEN_1362;
  wire        _GEN_1364 = io_lsu_clr_bsy_2_bits[6:2] == 5'h11;
  wire        _GEN_1365 = _GEN_11 & _GEN_1364;
  wire        _GEN_1366 = io_lsu_clr_bsy_2_bits[6:2] == 5'h12;
  wire        _GEN_1367 = _GEN_11 & _GEN_1366;
  wire        _GEN_1368 = io_lsu_clr_bsy_2_bits[6:2] == 5'h13;
  wire        _GEN_1369 = _GEN_11 & _GEN_1368;
  wire        _GEN_1370 = io_lsu_clr_bsy_2_bits[6:2] == 5'h14;
  wire        _GEN_1371 = _GEN_11 & _GEN_1370;
  wire        _GEN_1372 = io_lsu_clr_bsy_2_bits[6:2] == 5'h15;
  wire        _GEN_1373 = _GEN_11 & _GEN_1372;
  wire        _GEN_1374 = io_lsu_clr_bsy_2_bits[6:2] == 5'h16;
  wire        _GEN_1375 = _GEN_11 & _GEN_1374;
  wire        _GEN_1376 = io_lsu_clr_bsy_2_bits[6:2] == 5'h17;
  wire        _GEN_1377 = _GEN_11 & _GEN_1376;
  wire        _GEN_1378 = io_lsu_clr_bsy_2_bits[6:2] == 5'h18;
  wire        _GEN_1379 = _GEN_11 & _GEN_1378;
  wire        _GEN_1380 = io_lsu_clr_bsy_2_bits[6:2] == 5'h19;
  wire        _GEN_1381 = _GEN_11 & _GEN_1380;
  wire        _GEN_1382 = io_lsu_clr_bsy_2_bits[6:2] == 5'h1A;
  wire        _GEN_1383 = _GEN_11 & _GEN_1382;
  wire        _GEN_1384 = io_lsu_clr_bsy_2_bits[6:2] == 5'h1B;
  wire        _GEN_1385 = _GEN_11 & _GEN_1384;
  wire        _GEN_1386 = io_lsu_clr_bsy_2_bits[6:2] == 5'h1C;
  wire        _GEN_1387 = _GEN_11 & _GEN_1386;
  wire        _GEN_1388 = io_lsu_clr_bsy_2_bits[6:2] == 5'h1D;
  wire        _GEN_1389 = _GEN_11 & _GEN_1388;
  wire        _GEN_1390 = io_lsu_clr_bsy_2_bits[6:2] == 5'h1E;
  wire        _GEN_1391 = _GEN_11 & _GEN_1390;
  wire        _GEN_1392 = _GEN_11 & (&(io_lsu_clr_bsy_2_bits[6:2]));
  wire        _GEN_1393 = io_fflags_0_valid & io_fflags_0_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_1394 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_1395 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_1396 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_1397 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_1398 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_1399 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_1400 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_1401 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_1402 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_1403 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_1404 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_1405 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_1406 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_1407 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_1408 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_1409 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_1410 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_1411 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_1412 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_1413 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_1414 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_1415 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_1416 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_1417 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_1418 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_1419 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_1420 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_1421 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_1422 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_1423 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_1424 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_1425 = io_fflags_2_valid & io_fflags_2_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_1426 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_1427 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_1428 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_1429 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_1430 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_1431 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_1432 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_1433 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_1434 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_1435 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_1436 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_1437 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_1438 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_1439 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_1440 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_1441 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_1442 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_1443 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_1444 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_1445 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_1446 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_1447 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_1448 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_1449 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_1450 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_1451 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_1452 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_1453 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_1454 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_1455 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_1456 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_1457 = io_fflags_3_valid & io_fflags_3_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_1458 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_1459 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_1460 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_1461 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_1462 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_1463 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_1464 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_1465 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_1466 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_1467 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_1468 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_1469 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_1470 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_1471 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_1472 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_1473 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_1474 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_1475 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_1476 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_1477 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_1478 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_1479 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_1480 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_1481 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_1482 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_1483 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_1484 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_1485 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_1486 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_1487 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_1488 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_1489 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_1490 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_1491 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_1492 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_1493 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_1494 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_1495 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_1496 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_1497 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_1498 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_1499 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_1500 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_1501 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_1502 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_1503 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_1504 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_1505 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_1506 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_1507 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_1508 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_1509 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_1510 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_1511 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_1512 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_1513 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_1514 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_1515 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_1516 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_1517 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_1518 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_1519 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_1520 = com_idx == 5'h0;
  wire        _GEN_1521 = rbk_row & _GEN_1520;
  wire        _GEN_1522 = com_idx == 5'h1;
  wire        _GEN_1523 = rbk_row & _GEN_1522;
  wire        _GEN_1524 = com_idx == 5'h2;
  wire        _GEN_1525 = rbk_row & _GEN_1524;
  wire        _GEN_1526 = com_idx == 5'h3;
  wire        _GEN_1527 = rbk_row & _GEN_1526;
  wire        _GEN_1528 = com_idx == 5'h4;
  wire        _GEN_1529 = rbk_row & _GEN_1528;
  wire        _GEN_1530 = com_idx == 5'h5;
  wire        _GEN_1531 = rbk_row & _GEN_1530;
  wire        _GEN_1532 = com_idx == 5'h6;
  wire        _GEN_1533 = rbk_row & _GEN_1532;
  wire        _GEN_1534 = com_idx == 5'h7;
  wire        _GEN_1535 = rbk_row & _GEN_1534;
  wire        _GEN_1536 = com_idx == 5'h8;
  wire        _GEN_1537 = rbk_row & _GEN_1536;
  wire        _GEN_1538 = com_idx == 5'h9;
  wire        _GEN_1539 = rbk_row & _GEN_1538;
  wire        _GEN_1540 = com_idx == 5'hA;
  wire        _GEN_1541 = rbk_row & _GEN_1540;
  wire        _GEN_1542 = com_idx == 5'hB;
  wire        _GEN_1543 = rbk_row & _GEN_1542;
  wire        _GEN_1544 = com_idx == 5'hC;
  wire        _GEN_1545 = rbk_row & _GEN_1544;
  wire        _GEN_1546 = com_idx == 5'hD;
  wire        _GEN_1547 = rbk_row & _GEN_1546;
  wire        _GEN_1548 = com_idx == 5'hE;
  wire        _GEN_1549 = rbk_row & _GEN_1548;
  wire        _GEN_1550 = com_idx == 5'hF;
  wire        _GEN_1551 = rbk_row & _GEN_1550;
  wire        _GEN_1552 = com_idx == 5'h10;
  wire        _GEN_1553 = rbk_row & _GEN_1552;
  wire        _GEN_1554 = com_idx == 5'h11;
  wire        _GEN_1555 = rbk_row & _GEN_1554;
  wire        _GEN_1556 = com_idx == 5'h12;
  wire        _GEN_1557 = rbk_row & _GEN_1556;
  wire        _GEN_1558 = com_idx == 5'h13;
  wire        _GEN_1559 = rbk_row & _GEN_1558;
  wire        _GEN_1560 = com_idx == 5'h14;
  wire        _GEN_1561 = rbk_row & _GEN_1560;
  wire        _GEN_1562 = com_idx == 5'h15;
  wire        _GEN_1563 = rbk_row & _GEN_1562;
  wire        _GEN_1564 = com_idx == 5'h16;
  wire        _GEN_1565 = rbk_row & _GEN_1564;
  wire        _GEN_1566 = com_idx == 5'h17;
  wire        _GEN_1567 = rbk_row & _GEN_1566;
  wire        _GEN_1568 = com_idx == 5'h18;
  wire        _GEN_1569 = rbk_row & _GEN_1568;
  wire        _GEN_1570 = com_idx == 5'h19;
  wire        _GEN_1571 = rbk_row & _GEN_1570;
  wire        _GEN_1572 = com_idx == 5'h1A;
  wire        _GEN_1573 = rbk_row & _GEN_1572;
  wire        _GEN_1574 = com_idx == 5'h1B;
  wire        _GEN_1575 = rbk_row & _GEN_1574;
  wire        _GEN_1576 = com_idx == 5'h1C;
  wire        _GEN_1577 = rbk_row & _GEN_1576;
  wire        _GEN_1578 = com_idx == 5'h1D;
  wire        _GEN_1579 = rbk_row & _GEN_1578;
  wire        _GEN_1580 = com_idx == 5'h1E;
  wire        _GEN_1581 = rbk_row & _GEN_1580;
  wire        _GEN_1582 = rbk_row & (&com_idx);
  wire [19:0] _GEN_1583 = io_brupdate_b1_mispredict_mask & rob_uop_0_br_mask;
  wire [19:0] _GEN_1584 = io_brupdate_b1_mispredict_mask & rob_uop_1_br_mask;
  wire [19:0] _GEN_1585 = io_brupdate_b1_mispredict_mask & rob_uop_2_br_mask;
  wire [19:0] _GEN_1586 = io_brupdate_b1_mispredict_mask & rob_uop_3_br_mask;
  wire [19:0] _GEN_1587 = io_brupdate_b1_mispredict_mask & rob_uop_4_br_mask;
  wire [19:0] _GEN_1588 = io_brupdate_b1_mispredict_mask & rob_uop_5_br_mask;
  wire [19:0] _GEN_1589 = io_brupdate_b1_mispredict_mask & rob_uop_6_br_mask;
  wire [19:0] _GEN_1590 = io_brupdate_b1_mispredict_mask & rob_uop_7_br_mask;
  wire [19:0] _GEN_1591 = io_brupdate_b1_mispredict_mask & rob_uop_8_br_mask;
  wire [19:0] _GEN_1592 = io_brupdate_b1_mispredict_mask & rob_uop_9_br_mask;
  wire [19:0] _GEN_1593 = io_brupdate_b1_mispredict_mask & rob_uop_10_br_mask;
  wire [19:0] _GEN_1594 = io_brupdate_b1_mispredict_mask & rob_uop_11_br_mask;
  wire [19:0] _GEN_1595 = io_brupdate_b1_mispredict_mask & rob_uop_12_br_mask;
  wire [19:0] _GEN_1596 = io_brupdate_b1_mispredict_mask & rob_uop_13_br_mask;
  wire [19:0] _GEN_1597 = io_brupdate_b1_mispredict_mask & rob_uop_14_br_mask;
  wire [19:0] _GEN_1598 = io_brupdate_b1_mispredict_mask & rob_uop_15_br_mask;
  wire [19:0] _GEN_1599 = io_brupdate_b1_mispredict_mask & rob_uop_16_br_mask;
  wire [19:0] _GEN_1600 = io_brupdate_b1_mispredict_mask & rob_uop_17_br_mask;
  wire [19:0] _GEN_1601 = io_brupdate_b1_mispredict_mask & rob_uop_18_br_mask;
  wire [19:0] _GEN_1602 = io_brupdate_b1_mispredict_mask & rob_uop_19_br_mask;
  wire [19:0] _GEN_1603 = io_brupdate_b1_mispredict_mask & rob_uop_20_br_mask;
  wire [19:0] _GEN_1604 = io_brupdate_b1_mispredict_mask & rob_uop_21_br_mask;
  wire [19:0] _GEN_1605 = io_brupdate_b1_mispredict_mask & rob_uop_22_br_mask;
  wire [19:0] _GEN_1606 = io_brupdate_b1_mispredict_mask & rob_uop_23_br_mask;
  wire [19:0] _GEN_1607 = io_brupdate_b1_mispredict_mask & rob_uop_24_br_mask;
  wire [19:0] _GEN_1608 = io_brupdate_b1_mispredict_mask & rob_uop_25_br_mask;
  wire [19:0] _GEN_1609 = io_brupdate_b1_mispredict_mask & rob_uop_26_br_mask;
  wire [19:0] _GEN_1610 = io_brupdate_b1_mispredict_mask & rob_uop_27_br_mask;
  wire [19:0] _GEN_1611 = io_brupdate_b1_mispredict_mask & rob_uop_28_br_mask;
  wire [19:0] _GEN_1612 = io_brupdate_b1_mispredict_mask & rob_uop_29_br_mask;
  wire [19:0] _GEN_1613 = io_brupdate_b1_mispredict_mask & rob_uop_30_br_mask;
  wire [19:0] _GEN_1614 = io_brupdate_b1_mispredict_mask & rob_uop_31_br_mask;
  wire        _GEN_1615 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_1616 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_1617 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_1618 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_1619 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_1620 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_1621 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_1622 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_1623 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_1624 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_1625 = io_brupdate_b2_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_1626 = io_brupdate_b2_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_1627 = io_brupdate_b2_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_1628 = io_brupdate_b2_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_1629 = io_brupdate_b2_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_1630 = io_brupdate_b2_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_1631 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_1632 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_1633 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_1634 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_1635 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_1636 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_1637 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_1638 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_1639 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_1640 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_1641 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_1642 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_1643 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_1644 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_1645 = io_brupdate_b2_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_1646 = io_enq_valids_1 & _GEN_127;
  wire        _GEN_1647 = io_enq_valids_1 & _GEN_129;
  wire        _GEN_1648 = io_enq_valids_1 & _GEN_131;
  wire        _GEN_1649 = io_enq_valids_1 & _GEN_133;
  wire        _GEN_1650 = io_enq_valids_1 & _GEN_135;
  wire        _GEN_1651 = io_enq_valids_1 & _GEN_137;
  wire        _GEN_1652 = io_enq_valids_1 & _GEN_139;
  wire        _GEN_1653 = io_enq_valids_1 & _GEN_141;
  wire        _GEN_1654 = io_enq_valids_1 & _GEN_143;
  wire        _GEN_1655 = io_enq_valids_1 & _GEN_145;
  wire        _GEN_1656 = io_enq_valids_1 & _GEN_147;
  wire        _GEN_1657 = io_enq_valids_1 & _GEN_149;
  wire        _GEN_1658 = io_enq_valids_1 & _GEN_151;
  wire        _GEN_1659 = io_enq_valids_1 & _GEN_153;
  wire        _GEN_1660 = io_enq_valids_1 & _GEN_155;
  wire        _GEN_1661 = io_enq_valids_1 & _GEN_157;
  wire        _GEN_1662 = io_enq_valids_1 & _GEN_159;
  wire        _GEN_1663 = io_enq_valids_1 & _GEN_161;
  wire        _GEN_1664 = io_enq_valids_1 & _GEN_163;
  wire        _GEN_1665 = io_enq_valids_1 & _GEN_165;
  wire        _GEN_1666 = io_enq_valids_1 & _GEN_167;
  wire        _GEN_1667 = io_enq_valids_1 & _GEN_169;
  wire        _GEN_1668 = io_enq_valids_1 & _GEN_171;
  wire        _GEN_1669 = io_enq_valids_1 & _GEN_173;
  wire        _GEN_1670 = io_enq_valids_1 & _GEN_175;
  wire        _GEN_1671 = io_enq_valids_1 & _GEN_177;
  wire        _GEN_1672 = io_enq_valids_1 & _GEN_179;
  wire        _GEN_1673 = io_enq_valids_1 & _GEN_181;
  wire        _GEN_1674 = io_enq_valids_1 & _GEN_183;
  wire        _GEN_1675 = io_enq_valids_1 & _GEN_185;
  wire        _GEN_1676 = io_enq_valids_1 & _GEN_187;
  wire        _GEN_1677 = io_enq_valids_1 & (&rob_tail);
  wire        _rob_bsy_T_2 = io_enq_uops_1_is_fence | io_enq_uops_1_is_fencei;
  wire        _GEN_1678 = _GEN_1646 ? ~_rob_bsy_T_2 : rob_bsy_1_0;
  wire        _GEN_1679 = _GEN_1647 ? ~_rob_bsy_T_2 : rob_bsy_1_1;
  wire        _GEN_1680 = _GEN_1648 ? ~_rob_bsy_T_2 : rob_bsy_1_2;
  wire        _GEN_1681 = _GEN_1649 ? ~_rob_bsy_T_2 : rob_bsy_1_3;
  wire        _GEN_1682 = _GEN_1650 ? ~_rob_bsy_T_2 : rob_bsy_1_4;
  wire        _GEN_1683 = _GEN_1651 ? ~_rob_bsy_T_2 : rob_bsy_1_5;
  wire        _GEN_1684 = _GEN_1652 ? ~_rob_bsy_T_2 : rob_bsy_1_6;
  wire        _GEN_1685 = _GEN_1653 ? ~_rob_bsy_T_2 : rob_bsy_1_7;
  wire        _GEN_1686 = _GEN_1654 ? ~_rob_bsy_T_2 : rob_bsy_1_8;
  wire        _GEN_1687 = _GEN_1655 ? ~_rob_bsy_T_2 : rob_bsy_1_9;
  wire        _GEN_1688 = _GEN_1656 ? ~_rob_bsy_T_2 : rob_bsy_1_10;
  wire        _GEN_1689 = _GEN_1657 ? ~_rob_bsy_T_2 : rob_bsy_1_11;
  wire        _GEN_1690 = _GEN_1658 ? ~_rob_bsy_T_2 : rob_bsy_1_12;
  wire        _GEN_1691 = _GEN_1659 ? ~_rob_bsy_T_2 : rob_bsy_1_13;
  wire        _GEN_1692 = _GEN_1660 ? ~_rob_bsy_T_2 : rob_bsy_1_14;
  wire        _GEN_1693 = _GEN_1661 ? ~_rob_bsy_T_2 : rob_bsy_1_15;
  wire        _GEN_1694 = _GEN_1662 ? ~_rob_bsy_T_2 : rob_bsy_1_16;
  wire        _GEN_1695 = _GEN_1663 ? ~_rob_bsy_T_2 : rob_bsy_1_17;
  wire        _GEN_1696 = _GEN_1664 ? ~_rob_bsy_T_2 : rob_bsy_1_18;
  wire        _GEN_1697 = _GEN_1665 ? ~_rob_bsy_T_2 : rob_bsy_1_19;
  wire        _GEN_1698 = _GEN_1666 ? ~_rob_bsy_T_2 : rob_bsy_1_20;
  wire        _GEN_1699 = _GEN_1667 ? ~_rob_bsy_T_2 : rob_bsy_1_21;
  wire        _GEN_1700 = _GEN_1668 ? ~_rob_bsy_T_2 : rob_bsy_1_22;
  wire        _GEN_1701 = _GEN_1669 ? ~_rob_bsy_T_2 : rob_bsy_1_23;
  wire        _GEN_1702 = _GEN_1670 ? ~_rob_bsy_T_2 : rob_bsy_1_24;
  wire        _GEN_1703 = _GEN_1671 ? ~_rob_bsy_T_2 : rob_bsy_1_25;
  wire        _GEN_1704 = _GEN_1672 ? ~_rob_bsy_T_2 : rob_bsy_1_26;
  wire        _GEN_1705 = _GEN_1673 ? ~_rob_bsy_T_2 : rob_bsy_1_27;
  wire        _GEN_1706 = _GEN_1674 ? ~_rob_bsy_T_2 : rob_bsy_1_28;
  wire        _GEN_1707 = _GEN_1675 ? ~_rob_bsy_T_2 : rob_bsy_1_29;
  wire        _GEN_1708 = _GEN_1676 ? ~_rob_bsy_T_2 : rob_bsy_1_30;
  wire        _GEN_1709 = _GEN_1677 ? ~_rob_bsy_T_2 : rob_bsy_1_31;
  wire        _rob_unsafe_T_9 = io_enq_uops_1_uses_ldq | io_enq_uops_1_uses_stq & ~io_enq_uops_1_is_fence | io_enq_uops_1_is_br | io_enq_uops_1_is_jalr;
  wire        _GEN_1710 = _GEN_1646 ? _rob_unsafe_T_9 : rob_unsafe_1_0;
  wire        _GEN_1711 = _GEN_1647 ? _rob_unsafe_T_9 : rob_unsafe_1_1;
  wire        _GEN_1712 = _GEN_1648 ? _rob_unsafe_T_9 : rob_unsafe_1_2;
  wire        _GEN_1713 = _GEN_1649 ? _rob_unsafe_T_9 : rob_unsafe_1_3;
  wire        _GEN_1714 = _GEN_1650 ? _rob_unsafe_T_9 : rob_unsafe_1_4;
  wire        _GEN_1715 = _GEN_1651 ? _rob_unsafe_T_9 : rob_unsafe_1_5;
  wire        _GEN_1716 = _GEN_1652 ? _rob_unsafe_T_9 : rob_unsafe_1_6;
  wire        _GEN_1717 = _GEN_1653 ? _rob_unsafe_T_9 : rob_unsafe_1_7;
  wire        _GEN_1718 = _GEN_1654 ? _rob_unsafe_T_9 : rob_unsafe_1_8;
  wire        _GEN_1719 = _GEN_1655 ? _rob_unsafe_T_9 : rob_unsafe_1_9;
  wire        _GEN_1720 = _GEN_1656 ? _rob_unsafe_T_9 : rob_unsafe_1_10;
  wire        _GEN_1721 = _GEN_1657 ? _rob_unsafe_T_9 : rob_unsafe_1_11;
  wire        _GEN_1722 = _GEN_1658 ? _rob_unsafe_T_9 : rob_unsafe_1_12;
  wire        _GEN_1723 = _GEN_1659 ? _rob_unsafe_T_9 : rob_unsafe_1_13;
  wire        _GEN_1724 = _GEN_1660 ? _rob_unsafe_T_9 : rob_unsafe_1_14;
  wire        _GEN_1725 = _GEN_1661 ? _rob_unsafe_T_9 : rob_unsafe_1_15;
  wire        _GEN_1726 = _GEN_1662 ? _rob_unsafe_T_9 : rob_unsafe_1_16;
  wire        _GEN_1727 = _GEN_1663 ? _rob_unsafe_T_9 : rob_unsafe_1_17;
  wire        _GEN_1728 = _GEN_1664 ? _rob_unsafe_T_9 : rob_unsafe_1_18;
  wire        _GEN_1729 = _GEN_1665 ? _rob_unsafe_T_9 : rob_unsafe_1_19;
  wire        _GEN_1730 = _GEN_1666 ? _rob_unsafe_T_9 : rob_unsafe_1_20;
  wire        _GEN_1731 = _GEN_1667 ? _rob_unsafe_T_9 : rob_unsafe_1_21;
  wire        _GEN_1732 = _GEN_1668 ? _rob_unsafe_T_9 : rob_unsafe_1_22;
  wire        _GEN_1733 = _GEN_1669 ? _rob_unsafe_T_9 : rob_unsafe_1_23;
  wire        _GEN_1734 = _GEN_1670 ? _rob_unsafe_T_9 : rob_unsafe_1_24;
  wire        _GEN_1735 = _GEN_1671 ? _rob_unsafe_T_9 : rob_unsafe_1_25;
  wire        _GEN_1736 = _GEN_1672 ? _rob_unsafe_T_9 : rob_unsafe_1_26;
  wire        _GEN_1737 = _GEN_1673 ? _rob_unsafe_T_9 : rob_unsafe_1_27;
  wire        _GEN_1738 = _GEN_1674 ? _rob_unsafe_T_9 : rob_unsafe_1_28;
  wire        _GEN_1739 = _GEN_1675 ? _rob_unsafe_T_9 : rob_unsafe_1_29;
  wire        _GEN_1740 = _GEN_1676 ? _rob_unsafe_T_9 : rob_unsafe_1_30;
  wire        _GEN_1741 = _GEN_1677 ? _rob_unsafe_T_9 : rob_unsafe_1_31;
  wire        _GEN_1742 = _GEN_17 & _GEN_254;
  wire        _GEN_1743 = _GEN_17 & _GEN_256;
  wire        _GEN_1744 = _GEN_17 & _GEN_258;
  wire        _GEN_1745 = _GEN_17 & _GEN_260;
  wire        _GEN_1746 = _GEN_17 & _GEN_262;
  wire        _GEN_1747 = _GEN_17 & _GEN_264;
  wire        _GEN_1748 = _GEN_17 & _GEN_266;
  wire        _GEN_1749 = _GEN_17 & _GEN_268;
  wire        _GEN_1750 = _GEN_17 & _GEN_270;
  wire        _GEN_1751 = _GEN_17 & _GEN_272;
  wire        _GEN_1752 = _GEN_17 & _GEN_274;
  wire        _GEN_1753 = _GEN_17 & _GEN_276;
  wire        _GEN_1754 = _GEN_17 & _GEN_278;
  wire        _GEN_1755 = _GEN_17 & _GEN_280;
  wire        _GEN_1756 = _GEN_17 & _GEN_282;
  wire        _GEN_1757 = _GEN_17 & _GEN_284;
  wire        _GEN_1758 = _GEN_17 & _GEN_286;
  wire        _GEN_1759 = _GEN_17 & _GEN_288;
  wire        _GEN_1760 = _GEN_17 & _GEN_290;
  wire        _GEN_1761 = _GEN_17 & _GEN_292;
  wire        _GEN_1762 = _GEN_17 & _GEN_294;
  wire        _GEN_1763 = _GEN_17 & _GEN_296;
  wire        _GEN_1764 = _GEN_17 & _GEN_298;
  wire        _GEN_1765 = _GEN_17 & _GEN_300;
  wire        _GEN_1766 = _GEN_17 & _GEN_302;
  wire        _GEN_1767 = _GEN_17 & _GEN_304;
  wire        _GEN_1768 = _GEN_17 & _GEN_306;
  wire        _GEN_1769 = _GEN_17 & _GEN_308;
  wire        _GEN_1770 = _GEN_17 & _GEN_310;
  wire        _GEN_1771 = _GEN_17 & _GEN_312;
  wire        _GEN_1772 = _GEN_17 & _GEN_314;
  wire        _GEN_1773 = _GEN_17 & (&(io_wb_resps_0_bits_uop_rob_idx[6:2]));
  wire        _GEN_1774 = _GEN_317 | _GEN_1742;
  wire        _GEN_1775 = _GEN_18 ? ~_GEN_1774 & _GEN_1678 : ~_GEN_1742 & _GEN_1678;
  wire        _GEN_1776 = _GEN_320 | _GEN_1743;
  wire        _GEN_1777 = _GEN_18 ? ~_GEN_1776 & _GEN_1679 : ~_GEN_1743 & _GEN_1679;
  wire        _GEN_1778 = _GEN_323 | _GEN_1744;
  wire        _GEN_1779 = _GEN_18 ? ~_GEN_1778 & _GEN_1680 : ~_GEN_1744 & _GEN_1680;
  wire        _GEN_1780 = _GEN_326 | _GEN_1745;
  wire        _GEN_1781 = _GEN_18 ? ~_GEN_1780 & _GEN_1681 : ~_GEN_1745 & _GEN_1681;
  wire        _GEN_1782 = _GEN_329 | _GEN_1746;
  wire        _GEN_1783 = _GEN_18 ? ~_GEN_1782 & _GEN_1682 : ~_GEN_1746 & _GEN_1682;
  wire        _GEN_1784 = _GEN_332 | _GEN_1747;
  wire        _GEN_1785 = _GEN_18 ? ~_GEN_1784 & _GEN_1683 : ~_GEN_1747 & _GEN_1683;
  wire        _GEN_1786 = _GEN_335 | _GEN_1748;
  wire        _GEN_1787 = _GEN_18 ? ~_GEN_1786 & _GEN_1684 : ~_GEN_1748 & _GEN_1684;
  wire        _GEN_1788 = _GEN_338 | _GEN_1749;
  wire        _GEN_1789 = _GEN_18 ? ~_GEN_1788 & _GEN_1685 : ~_GEN_1749 & _GEN_1685;
  wire        _GEN_1790 = _GEN_341 | _GEN_1750;
  wire        _GEN_1791 = _GEN_18 ? ~_GEN_1790 & _GEN_1686 : ~_GEN_1750 & _GEN_1686;
  wire        _GEN_1792 = _GEN_344 | _GEN_1751;
  wire        _GEN_1793 = _GEN_18 ? ~_GEN_1792 & _GEN_1687 : ~_GEN_1751 & _GEN_1687;
  wire        _GEN_1794 = _GEN_347 | _GEN_1752;
  wire        _GEN_1795 = _GEN_18 ? ~_GEN_1794 & _GEN_1688 : ~_GEN_1752 & _GEN_1688;
  wire        _GEN_1796 = _GEN_350 | _GEN_1753;
  wire        _GEN_1797 = _GEN_18 ? ~_GEN_1796 & _GEN_1689 : ~_GEN_1753 & _GEN_1689;
  wire        _GEN_1798 = _GEN_353 | _GEN_1754;
  wire        _GEN_1799 = _GEN_18 ? ~_GEN_1798 & _GEN_1690 : ~_GEN_1754 & _GEN_1690;
  wire        _GEN_1800 = _GEN_356 | _GEN_1755;
  wire        _GEN_1801 = _GEN_18 ? ~_GEN_1800 & _GEN_1691 : ~_GEN_1755 & _GEN_1691;
  wire        _GEN_1802 = _GEN_359 | _GEN_1756;
  wire        _GEN_1803 = _GEN_18 ? ~_GEN_1802 & _GEN_1692 : ~_GEN_1756 & _GEN_1692;
  wire        _GEN_1804 = _GEN_362 | _GEN_1757;
  wire        _GEN_1805 = _GEN_18 ? ~_GEN_1804 & _GEN_1693 : ~_GEN_1757 & _GEN_1693;
  wire        _GEN_1806 = _GEN_365 | _GEN_1758;
  wire        _GEN_1807 = _GEN_18 ? ~_GEN_1806 & _GEN_1694 : ~_GEN_1758 & _GEN_1694;
  wire        _GEN_1808 = _GEN_368 | _GEN_1759;
  wire        _GEN_1809 = _GEN_18 ? ~_GEN_1808 & _GEN_1695 : ~_GEN_1759 & _GEN_1695;
  wire        _GEN_1810 = _GEN_371 | _GEN_1760;
  wire        _GEN_1811 = _GEN_18 ? ~_GEN_1810 & _GEN_1696 : ~_GEN_1760 & _GEN_1696;
  wire        _GEN_1812 = _GEN_374 | _GEN_1761;
  wire        _GEN_1813 = _GEN_18 ? ~_GEN_1812 & _GEN_1697 : ~_GEN_1761 & _GEN_1697;
  wire        _GEN_1814 = _GEN_377 | _GEN_1762;
  wire        _GEN_1815 = _GEN_18 ? ~_GEN_1814 & _GEN_1698 : ~_GEN_1762 & _GEN_1698;
  wire        _GEN_1816 = _GEN_380 | _GEN_1763;
  wire        _GEN_1817 = _GEN_18 ? ~_GEN_1816 & _GEN_1699 : ~_GEN_1763 & _GEN_1699;
  wire        _GEN_1818 = _GEN_383 | _GEN_1764;
  wire        _GEN_1819 = _GEN_18 ? ~_GEN_1818 & _GEN_1700 : ~_GEN_1764 & _GEN_1700;
  wire        _GEN_1820 = _GEN_386 | _GEN_1765;
  wire        _GEN_1821 = _GEN_18 ? ~_GEN_1820 & _GEN_1701 : ~_GEN_1765 & _GEN_1701;
  wire        _GEN_1822 = _GEN_389 | _GEN_1766;
  wire        _GEN_1823 = _GEN_18 ? ~_GEN_1822 & _GEN_1702 : ~_GEN_1766 & _GEN_1702;
  wire        _GEN_1824 = _GEN_392 | _GEN_1767;
  wire        _GEN_1825 = _GEN_18 ? ~_GEN_1824 & _GEN_1703 : ~_GEN_1767 & _GEN_1703;
  wire        _GEN_1826 = _GEN_395 | _GEN_1768;
  wire        _GEN_1827 = _GEN_18 ? ~_GEN_1826 & _GEN_1704 : ~_GEN_1768 & _GEN_1704;
  wire        _GEN_1828 = _GEN_398 | _GEN_1769;
  wire        _GEN_1829 = _GEN_18 ? ~_GEN_1828 & _GEN_1705 : ~_GEN_1769 & _GEN_1705;
  wire        _GEN_1830 = _GEN_401 | _GEN_1770;
  wire        _GEN_1831 = _GEN_18 ? ~_GEN_1830 & _GEN_1706 : ~_GEN_1770 & _GEN_1706;
  wire        _GEN_1832 = _GEN_404 | _GEN_1771;
  wire        _GEN_1833 = _GEN_18 ? ~_GEN_1832 & _GEN_1707 : ~_GEN_1771 & _GEN_1707;
  wire        _GEN_1834 = _GEN_407 | _GEN_1772;
  wire        _GEN_1835 = _GEN_18 ? ~_GEN_1834 & _GEN_1708 : ~_GEN_1772 & _GEN_1708;
  wire        _GEN_1836 = (&(io_wb_resps_1_bits_uop_rob_idx[6:2])) | _GEN_1773;
  wire        _GEN_1837 = _GEN_18 ? ~_GEN_1836 & _GEN_1709 : ~_GEN_1773 & _GEN_1709;
  wire        _GEN_1838 = _GEN_18 ? ~_GEN_1774 & _GEN_1710 : ~_GEN_1742 & _GEN_1710;
  wire        _GEN_1839 = _GEN_18 ? ~_GEN_1776 & _GEN_1711 : ~_GEN_1743 & _GEN_1711;
  wire        _GEN_1840 = _GEN_18 ? ~_GEN_1778 & _GEN_1712 : ~_GEN_1744 & _GEN_1712;
  wire        _GEN_1841 = _GEN_18 ? ~_GEN_1780 & _GEN_1713 : ~_GEN_1745 & _GEN_1713;
  wire        _GEN_1842 = _GEN_18 ? ~_GEN_1782 & _GEN_1714 : ~_GEN_1746 & _GEN_1714;
  wire        _GEN_1843 = _GEN_18 ? ~_GEN_1784 & _GEN_1715 : ~_GEN_1747 & _GEN_1715;
  wire        _GEN_1844 = _GEN_18 ? ~_GEN_1786 & _GEN_1716 : ~_GEN_1748 & _GEN_1716;
  wire        _GEN_1845 = _GEN_18 ? ~_GEN_1788 & _GEN_1717 : ~_GEN_1749 & _GEN_1717;
  wire        _GEN_1846 = _GEN_18 ? ~_GEN_1790 & _GEN_1718 : ~_GEN_1750 & _GEN_1718;
  wire        _GEN_1847 = _GEN_18 ? ~_GEN_1792 & _GEN_1719 : ~_GEN_1751 & _GEN_1719;
  wire        _GEN_1848 = _GEN_18 ? ~_GEN_1794 & _GEN_1720 : ~_GEN_1752 & _GEN_1720;
  wire        _GEN_1849 = _GEN_18 ? ~_GEN_1796 & _GEN_1721 : ~_GEN_1753 & _GEN_1721;
  wire        _GEN_1850 = _GEN_18 ? ~_GEN_1798 & _GEN_1722 : ~_GEN_1754 & _GEN_1722;
  wire        _GEN_1851 = _GEN_18 ? ~_GEN_1800 & _GEN_1723 : ~_GEN_1755 & _GEN_1723;
  wire        _GEN_1852 = _GEN_18 ? ~_GEN_1802 & _GEN_1724 : ~_GEN_1756 & _GEN_1724;
  wire        _GEN_1853 = _GEN_18 ? ~_GEN_1804 & _GEN_1725 : ~_GEN_1757 & _GEN_1725;
  wire        _GEN_1854 = _GEN_18 ? ~_GEN_1806 & _GEN_1726 : ~_GEN_1758 & _GEN_1726;
  wire        _GEN_1855 = _GEN_18 ? ~_GEN_1808 & _GEN_1727 : ~_GEN_1759 & _GEN_1727;
  wire        _GEN_1856 = _GEN_18 ? ~_GEN_1810 & _GEN_1728 : ~_GEN_1760 & _GEN_1728;
  wire        _GEN_1857 = _GEN_18 ? ~_GEN_1812 & _GEN_1729 : ~_GEN_1761 & _GEN_1729;
  wire        _GEN_1858 = _GEN_18 ? ~_GEN_1814 & _GEN_1730 : ~_GEN_1762 & _GEN_1730;
  wire        _GEN_1859 = _GEN_18 ? ~_GEN_1816 & _GEN_1731 : ~_GEN_1763 & _GEN_1731;
  wire        _GEN_1860 = _GEN_18 ? ~_GEN_1818 & _GEN_1732 : ~_GEN_1764 & _GEN_1732;
  wire        _GEN_1861 = _GEN_18 ? ~_GEN_1820 & _GEN_1733 : ~_GEN_1765 & _GEN_1733;
  wire        _GEN_1862 = _GEN_18 ? ~_GEN_1822 & _GEN_1734 : ~_GEN_1766 & _GEN_1734;
  wire        _GEN_1863 = _GEN_18 ? ~_GEN_1824 & _GEN_1735 : ~_GEN_1767 & _GEN_1735;
  wire        _GEN_1864 = _GEN_18 ? ~_GEN_1826 & _GEN_1736 : ~_GEN_1768 & _GEN_1736;
  wire        _GEN_1865 = _GEN_18 ? ~_GEN_1828 & _GEN_1737 : ~_GEN_1769 & _GEN_1737;
  wire        _GEN_1866 = _GEN_18 ? ~_GEN_1830 & _GEN_1738 : ~_GEN_1770 & _GEN_1738;
  wire        _GEN_1867 = _GEN_18 ? ~_GEN_1832 & _GEN_1739 : ~_GEN_1771 & _GEN_1739;
  wire        _GEN_1868 = _GEN_18 ? ~_GEN_1834 & _GEN_1740 : ~_GEN_1772 & _GEN_1740;
  wire        _GEN_1869 = _GEN_18 ? ~_GEN_1836 & _GEN_1741 : ~_GEN_1773 & _GEN_1741;
  wire        _GEN_1870 = _GEN_19 & _GEN_444;
  wire        _GEN_1871 = _GEN_19 & _GEN_446;
  wire        _GEN_1872 = _GEN_19 & _GEN_448;
  wire        _GEN_1873 = _GEN_19 & _GEN_450;
  wire        _GEN_1874 = _GEN_19 & _GEN_452;
  wire        _GEN_1875 = _GEN_19 & _GEN_454;
  wire        _GEN_1876 = _GEN_19 & _GEN_456;
  wire        _GEN_1877 = _GEN_19 & _GEN_458;
  wire        _GEN_1878 = _GEN_19 & _GEN_460;
  wire        _GEN_1879 = _GEN_19 & _GEN_462;
  wire        _GEN_1880 = _GEN_19 & _GEN_464;
  wire        _GEN_1881 = _GEN_19 & _GEN_466;
  wire        _GEN_1882 = _GEN_19 & _GEN_468;
  wire        _GEN_1883 = _GEN_19 & _GEN_470;
  wire        _GEN_1884 = _GEN_19 & _GEN_472;
  wire        _GEN_1885 = _GEN_19 & _GEN_474;
  wire        _GEN_1886 = _GEN_19 & _GEN_476;
  wire        _GEN_1887 = _GEN_19 & _GEN_478;
  wire        _GEN_1888 = _GEN_19 & _GEN_480;
  wire        _GEN_1889 = _GEN_19 & _GEN_482;
  wire        _GEN_1890 = _GEN_19 & _GEN_484;
  wire        _GEN_1891 = _GEN_19 & _GEN_486;
  wire        _GEN_1892 = _GEN_19 & _GEN_488;
  wire        _GEN_1893 = _GEN_19 & _GEN_490;
  wire        _GEN_1894 = _GEN_19 & _GEN_492;
  wire        _GEN_1895 = _GEN_19 & _GEN_494;
  wire        _GEN_1896 = _GEN_19 & _GEN_496;
  wire        _GEN_1897 = _GEN_19 & _GEN_498;
  wire        _GEN_1898 = _GEN_19 & _GEN_500;
  wire        _GEN_1899 = _GEN_19 & _GEN_502;
  wire        _GEN_1900 = _GEN_19 & _GEN_504;
  wire        _GEN_1901 = _GEN_19 & (&(io_wb_resps_2_bits_uop_rob_idx[6:2]));
  wire        _GEN_1902 = _GEN_507 | _GEN_1870;
  wire        _GEN_1903 = _GEN_20 ? ~_GEN_1902 & _GEN_1775 : ~_GEN_1870 & _GEN_1775;
  wire        _GEN_1904 = _GEN_510 | _GEN_1871;
  wire        _GEN_1905 = _GEN_20 ? ~_GEN_1904 & _GEN_1777 : ~_GEN_1871 & _GEN_1777;
  wire        _GEN_1906 = _GEN_513 | _GEN_1872;
  wire        _GEN_1907 = _GEN_20 ? ~_GEN_1906 & _GEN_1779 : ~_GEN_1872 & _GEN_1779;
  wire        _GEN_1908 = _GEN_516 | _GEN_1873;
  wire        _GEN_1909 = _GEN_20 ? ~_GEN_1908 & _GEN_1781 : ~_GEN_1873 & _GEN_1781;
  wire        _GEN_1910 = _GEN_519 | _GEN_1874;
  wire        _GEN_1911 = _GEN_20 ? ~_GEN_1910 & _GEN_1783 : ~_GEN_1874 & _GEN_1783;
  wire        _GEN_1912 = _GEN_522 | _GEN_1875;
  wire        _GEN_1913 = _GEN_20 ? ~_GEN_1912 & _GEN_1785 : ~_GEN_1875 & _GEN_1785;
  wire        _GEN_1914 = _GEN_525 | _GEN_1876;
  wire        _GEN_1915 = _GEN_20 ? ~_GEN_1914 & _GEN_1787 : ~_GEN_1876 & _GEN_1787;
  wire        _GEN_1916 = _GEN_528 | _GEN_1877;
  wire        _GEN_1917 = _GEN_20 ? ~_GEN_1916 & _GEN_1789 : ~_GEN_1877 & _GEN_1789;
  wire        _GEN_1918 = _GEN_531 | _GEN_1878;
  wire        _GEN_1919 = _GEN_20 ? ~_GEN_1918 & _GEN_1791 : ~_GEN_1878 & _GEN_1791;
  wire        _GEN_1920 = _GEN_534 | _GEN_1879;
  wire        _GEN_1921 = _GEN_20 ? ~_GEN_1920 & _GEN_1793 : ~_GEN_1879 & _GEN_1793;
  wire        _GEN_1922 = _GEN_537 | _GEN_1880;
  wire        _GEN_1923 = _GEN_20 ? ~_GEN_1922 & _GEN_1795 : ~_GEN_1880 & _GEN_1795;
  wire        _GEN_1924 = _GEN_540 | _GEN_1881;
  wire        _GEN_1925 = _GEN_20 ? ~_GEN_1924 & _GEN_1797 : ~_GEN_1881 & _GEN_1797;
  wire        _GEN_1926 = _GEN_543 | _GEN_1882;
  wire        _GEN_1927 = _GEN_20 ? ~_GEN_1926 & _GEN_1799 : ~_GEN_1882 & _GEN_1799;
  wire        _GEN_1928 = _GEN_546 | _GEN_1883;
  wire        _GEN_1929 = _GEN_20 ? ~_GEN_1928 & _GEN_1801 : ~_GEN_1883 & _GEN_1801;
  wire        _GEN_1930 = _GEN_549 | _GEN_1884;
  wire        _GEN_1931 = _GEN_20 ? ~_GEN_1930 & _GEN_1803 : ~_GEN_1884 & _GEN_1803;
  wire        _GEN_1932 = _GEN_552 | _GEN_1885;
  wire        _GEN_1933 = _GEN_20 ? ~_GEN_1932 & _GEN_1805 : ~_GEN_1885 & _GEN_1805;
  wire        _GEN_1934 = _GEN_555 | _GEN_1886;
  wire        _GEN_1935 = _GEN_20 ? ~_GEN_1934 & _GEN_1807 : ~_GEN_1886 & _GEN_1807;
  wire        _GEN_1936 = _GEN_558 | _GEN_1887;
  wire        _GEN_1937 = _GEN_20 ? ~_GEN_1936 & _GEN_1809 : ~_GEN_1887 & _GEN_1809;
  wire        _GEN_1938 = _GEN_561 | _GEN_1888;
  wire        _GEN_1939 = _GEN_20 ? ~_GEN_1938 & _GEN_1811 : ~_GEN_1888 & _GEN_1811;
  wire        _GEN_1940 = _GEN_564 | _GEN_1889;
  wire        _GEN_1941 = _GEN_20 ? ~_GEN_1940 & _GEN_1813 : ~_GEN_1889 & _GEN_1813;
  wire        _GEN_1942 = _GEN_567 | _GEN_1890;
  wire        _GEN_1943 = _GEN_20 ? ~_GEN_1942 & _GEN_1815 : ~_GEN_1890 & _GEN_1815;
  wire        _GEN_1944 = _GEN_570 | _GEN_1891;
  wire        _GEN_1945 = _GEN_20 ? ~_GEN_1944 & _GEN_1817 : ~_GEN_1891 & _GEN_1817;
  wire        _GEN_1946 = _GEN_573 | _GEN_1892;
  wire        _GEN_1947 = _GEN_20 ? ~_GEN_1946 & _GEN_1819 : ~_GEN_1892 & _GEN_1819;
  wire        _GEN_1948 = _GEN_576 | _GEN_1893;
  wire        _GEN_1949 = _GEN_20 ? ~_GEN_1948 & _GEN_1821 : ~_GEN_1893 & _GEN_1821;
  wire        _GEN_1950 = _GEN_579 | _GEN_1894;
  wire        _GEN_1951 = _GEN_20 ? ~_GEN_1950 & _GEN_1823 : ~_GEN_1894 & _GEN_1823;
  wire        _GEN_1952 = _GEN_582 | _GEN_1895;
  wire        _GEN_1953 = _GEN_20 ? ~_GEN_1952 & _GEN_1825 : ~_GEN_1895 & _GEN_1825;
  wire        _GEN_1954 = _GEN_585 | _GEN_1896;
  wire        _GEN_1955 = _GEN_20 ? ~_GEN_1954 & _GEN_1827 : ~_GEN_1896 & _GEN_1827;
  wire        _GEN_1956 = _GEN_588 | _GEN_1897;
  wire        _GEN_1957 = _GEN_20 ? ~_GEN_1956 & _GEN_1829 : ~_GEN_1897 & _GEN_1829;
  wire        _GEN_1958 = _GEN_591 | _GEN_1898;
  wire        _GEN_1959 = _GEN_20 ? ~_GEN_1958 & _GEN_1831 : ~_GEN_1898 & _GEN_1831;
  wire        _GEN_1960 = _GEN_594 | _GEN_1899;
  wire        _GEN_1961 = _GEN_20 ? ~_GEN_1960 & _GEN_1833 : ~_GEN_1899 & _GEN_1833;
  wire        _GEN_1962 = _GEN_597 | _GEN_1900;
  wire        _GEN_1963 = _GEN_20 ? ~_GEN_1962 & _GEN_1835 : ~_GEN_1900 & _GEN_1835;
  wire        _GEN_1964 = (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_1901;
  wire        _GEN_1965 = _GEN_20 ? ~_GEN_1964 & _GEN_1837 : ~_GEN_1901 & _GEN_1837;
  wire        _GEN_1966 = _GEN_20 ? ~_GEN_1902 & _GEN_1838 : ~_GEN_1870 & _GEN_1838;
  wire        _GEN_1967 = _GEN_20 ? ~_GEN_1904 & _GEN_1839 : ~_GEN_1871 & _GEN_1839;
  wire        _GEN_1968 = _GEN_20 ? ~_GEN_1906 & _GEN_1840 : ~_GEN_1872 & _GEN_1840;
  wire        _GEN_1969 = _GEN_20 ? ~_GEN_1908 & _GEN_1841 : ~_GEN_1873 & _GEN_1841;
  wire        _GEN_1970 = _GEN_20 ? ~_GEN_1910 & _GEN_1842 : ~_GEN_1874 & _GEN_1842;
  wire        _GEN_1971 = _GEN_20 ? ~_GEN_1912 & _GEN_1843 : ~_GEN_1875 & _GEN_1843;
  wire        _GEN_1972 = _GEN_20 ? ~_GEN_1914 & _GEN_1844 : ~_GEN_1876 & _GEN_1844;
  wire        _GEN_1973 = _GEN_20 ? ~_GEN_1916 & _GEN_1845 : ~_GEN_1877 & _GEN_1845;
  wire        _GEN_1974 = _GEN_20 ? ~_GEN_1918 & _GEN_1846 : ~_GEN_1878 & _GEN_1846;
  wire        _GEN_1975 = _GEN_20 ? ~_GEN_1920 & _GEN_1847 : ~_GEN_1879 & _GEN_1847;
  wire        _GEN_1976 = _GEN_20 ? ~_GEN_1922 & _GEN_1848 : ~_GEN_1880 & _GEN_1848;
  wire        _GEN_1977 = _GEN_20 ? ~_GEN_1924 & _GEN_1849 : ~_GEN_1881 & _GEN_1849;
  wire        _GEN_1978 = _GEN_20 ? ~_GEN_1926 & _GEN_1850 : ~_GEN_1882 & _GEN_1850;
  wire        _GEN_1979 = _GEN_20 ? ~_GEN_1928 & _GEN_1851 : ~_GEN_1883 & _GEN_1851;
  wire        _GEN_1980 = _GEN_20 ? ~_GEN_1930 & _GEN_1852 : ~_GEN_1884 & _GEN_1852;
  wire        _GEN_1981 = _GEN_20 ? ~_GEN_1932 & _GEN_1853 : ~_GEN_1885 & _GEN_1853;
  wire        _GEN_1982 = _GEN_20 ? ~_GEN_1934 & _GEN_1854 : ~_GEN_1886 & _GEN_1854;
  wire        _GEN_1983 = _GEN_20 ? ~_GEN_1936 & _GEN_1855 : ~_GEN_1887 & _GEN_1855;
  wire        _GEN_1984 = _GEN_20 ? ~_GEN_1938 & _GEN_1856 : ~_GEN_1888 & _GEN_1856;
  wire        _GEN_1985 = _GEN_20 ? ~_GEN_1940 & _GEN_1857 : ~_GEN_1889 & _GEN_1857;
  wire        _GEN_1986 = _GEN_20 ? ~_GEN_1942 & _GEN_1858 : ~_GEN_1890 & _GEN_1858;
  wire        _GEN_1987 = _GEN_20 ? ~_GEN_1944 & _GEN_1859 : ~_GEN_1891 & _GEN_1859;
  wire        _GEN_1988 = _GEN_20 ? ~_GEN_1946 & _GEN_1860 : ~_GEN_1892 & _GEN_1860;
  wire        _GEN_1989 = _GEN_20 ? ~_GEN_1948 & _GEN_1861 : ~_GEN_1893 & _GEN_1861;
  wire        _GEN_1990 = _GEN_20 ? ~_GEN_1950 & _GEN_1862 : ~_GEN_1894 & _GEN_1862;
  wire        _GEN_1991 = _GEN_20 ? ~_GEN_1952 & _GEN_1863 : ~_GEN_1895 & _GEN_1863;
  wire        _GEN_1992 = _GEN_20 ? ~_GEN_1954 & _GEN_1864 : ~_GEN_1896 & _GEN_1864;
  wire        _GEN_1993 = _GEN_20 ? ~_GEN_1956 & _GEN_1865 : ~_GEN_1897 & _GEN_1865;
  wire        _GEN_1994 = _GEN_20 ? ~_GEN_1958 & _GEN_1866 : ~_GEN_1898 & _GEN_1866;
  wire        _GEN_1995 = _GEN_20 ? ~_GEN_1960 & _GEN_1867 : ~_GEN_1899 & _GEN_1867;
  wire        _GEN_1996 = _GEN_20 ? ~_GEN_1962 & _GEN_1868 : ~_GEN_1900 & _GEN_1868;
  wire        _GEN_1997 = _GEN_20 ? ~_GEN_1964 & _GEN_1869 : ~_GEN_1901 & _GEN_1869;
  wire        _GEN_1998 = _GEN_21 & _GEN_634;
  wire        _GEN_1999 = _GEN_21 & _GEN_636;
  wire        _GEN_2000 = _GEN_21 & _GEN_638;
  wire        _GEN_2001 = _GEN_21 & _GEN_640;
  wire        _GEN_2002 = _GEN_21 & _GEN_642;
  wire        _GEN_2003 = _GEN_21 & _GEN_644;
  wire        _GEN_2004 = _GEN_21 & _GEN_646;
  wire        _GEN_2005 = _GEN_21 & _GEN_648;
  wire        _GEN_2006 = _GEN_21 & _GEN_650;
  wire        _GEN_2007 = _GEN_21 & _GEN_652;
  wire        _GEN_2008 = _GEN_21 & _GEN_654;
  wire        _GEN_2009 = _GEN_21 & _GEN_656;
  wire        _GEN_2010 = _GEN_21 & _GEN_658;
  wire        _GEN_2011 = _GEN_21 & _GEN_660;
  wire        _GEN_2012 = _GEN_21 & _GEN_662;
  wire        _GEN_2013 = _GEN_21 & _GEN_664;
  wire        _GEN_2014 = _GEN_21 & _GEN_666;
  wire        _GEN_2015 = _GEN_21 & _GEN_668;
  wire        _GEN_2016 = _GEN_21 & _GEN_670;
  wire        _GEN_2017 = _GEN_21 & _GEN_672;
  wire        _GEN_2018 = _GEN_21 & _GEN_674;
  wire        _GEN_2019 = _GEN_21 & _GEN_676;
  wire        _GEN_2020 = _GEN_21 & _GEN_678;
  wire        _GEN_2021 = _GEN_21 & _GEN_680;
  wire        _GEN_2022 = _GEN_21 & _GEN_682;
  wire        _GEN_2023 = _GEN_21 & _GEN_684;
  wire        _GEN_2024 = _GEN_21 & _GEN_686;
  wire        _GEN_2025 = _GEN_21 & _GEN_688;
  wire        _GEN_2026 = _GEN_21 & _GEN_690;
  wire        _GEN_2027 = _GEN_21 & _GEN_692;
  wire        _GEN_2028 = _GEN_21 & _GEN_694;
  wire        _GEN_2029 = _GEN_21 & (&(io_wb_resps_4_bits_uop_rob_idx[6:2]));
  wire        _GEN_2030 = _GEN_697 | _GEN_1998;
  wire        _GEN_2031 = _GEN_22 ? ~_GEN_2030 & _GEN_1903 : ~_GEN_1998 & _GEN_1903;
  wire        _GEN_2032 = _GEN_700 | _GEN_1999;
  wire        _GEN_2033 = _GEN_22 ? ~_GEN_2032 & _GEN_1905 : ~_GEN_1999 & _GEN_1905;
  wire        _GEN_2034 = _GEN_703 | _GEN_2000;
  wire        _GEN_2035 = _GEN_22 ? ~_GEN_2034 & _GEN_1907 : ~_GEN_2000 & _GEN_1907;
  wire        _GEN_2036 = _GEN_706 | _GEN_2001;
  wire        _GEN_2037 = _GEN_22 ? ~_GEN_2036 & _GEN_1909 : ~_GEN_2001 & _GEN_1909;
  wire        _GEN_2038 = _GEN_709 | _GEN_2002;
  wire        _GEN_2039 = _GEN_22 ? ~_GEN_2038 & _GEN_1911 : ~_GEN_2002 & _GEN_1911;
  wire        _GEN_2040 = _GEN_712 | _GEN_2003;
  wire        _GEN_2041 = _GEN_22 ? ~_GEN_2040 & _GEN_1913 : ~_GEN_2003 & _GEN_1913;
  wire        _GEN_2042 = _GEN_715 | _GEN_2004;
  wire        _GEN_2043 = _GEN_22 ? ~_GEN_2042 & _GEN_1915 : ~_GEN_2004 & _GEN_1915;
  wire        _GEN_2044 = _GEN_718 | _GEN_2005;
  wire        _GEN_2045 = _GEN_22 ? ~_GEN_2044 & _GEN_1917 : ~_GEN_2005 & _GEN_1917;
  wire        _GEN_2046 = _GEN_721 | _GEN_2006;
  wire        _GEN_2047 = _GEN_22 ? ~_GEN_2046 & _GEN_1919 : ~_GEN_2006 & _GEN_1919;
  wire        _GEN_2048 = _GEN_724 | _GEN_2007;
  wire        _GEN_2049 = _GEN_22 ? ~_GEN_2048 & _GEN_1921 : ~_GEN_2007 & _GEN_1921;
  wire        _GEN_2050 = _GEN_727 | _GEN_2008;
  wire        _GEN_2051 = _GEN_22 ? ~_GEN_2050 & _GEN_1923 : ~_GEN_2008 & _GEN_1923;
  wire        _GEN_2052 = _GEN_730 | _GEN_2009;
  wire        _GEN_2053 = _GEN_22 ? ~_GEN_2052 & _GEN_1925 : ~_GEN_2009 & _GEN_1925;
  wire        _GEN_2054 = _GEN_733 | _GEN_2010;
  wire        _GEN_2055 = _GEN_22 ? ~_GEN_2054 & _GEN_1927 : ~_GEN_2010 & _GEN_1927;
  wire        _GEN_2056 = _GEN_736 | _GEN_2011;
  wire        _GEN_2057 = _GEN_22 ? ~_GEN_2056 & _GEN_1929 : ~_GEN_2011 & _GEN_1929;
  wire        _GEN_2058 = _GEN_739 | _GEN_2012;
  wire        _GEN_2059 = _GEN_22 ? ~_GEN_2058 & _GEN_1931 : ~_GEN_2012 & _GEN_1931;
  wire        _GEN_2060 = _GEN_742 | _GEN_2013;
  wire        _GEN_2061 = _GEN_22 ? ~_GEN_2060 & _GEN_1933 : ~_GEN_2013 & _GEN_1933;
  wire        _GEN_2062 = _GEN_745 | _GEN_2014;
  wire        _GEN_2063 = _GEN_22 ? ~_GEN_2062 & _GEN_1935 : ~_GEN_2014 & _GEN_1935;
  wire        _GEN_2064 = _GEN_748 | _GEN_2015;
  wire        _GEN_2065 = _GEN_22 ? ~_GEN_2064 & _GEN_1937 : ~_GEN_2015 & _GEN_1937;
  wire        _GEN_2066 = _GEN_751 | _GEN_2016;
  wire        _GEN_2067 = _GEN_22 ? ~_GEN_2066 & _GEN_1939 : ~_GEN_2016 & _GEN_1939;
  wire        _GEN_2068 = _GEN_754 | _GEN_2017;
  wire        _GEN_2069 = _GEN_22 ? ~_GEN_2068 & _GEN_1941 : ~_GEN_2017 & _GEN_1941;
  wire        _GEN_2070 = _GEN_757 | _GEN_2018;
  wire        _GEN_2071 = _GEN_22 ? ~_GEN_2070 & _GEN_1943 : ~_GEN_2018 & _GEN_1943;
  wire        _GEN_2072 = _GEN_760 | _GEN_2019;
  wire        _GEN_2073 = _GEN_22 ? ~_GEN_2072 & _GEN_1945 : ~_GEN_2019 & _GEN_1945;
  wire        _GEN_2074 = _GEN_763 | _GEN_2020;
  wire        _GEN_2075 = _GEN_22 ? ~_GEN_2074 & _GEN_1947 : ~_GEN_2020 & _GEN_1947;
  wire        _GEN_2076 = _GEN_766 | _GEN_2021;
  wire        _GEN_2077 = _GEN_22 ? ~_GEN_2076 & _GEN_1949 : ~_GEN_2021 & _GEN_1949;
  wire        _GEN_2078 = _GEN_769 | _GEN_2022;
  wire        _GEN_2079 = _GEN_22 ? ~_GEN_2078 & _GEN_1951 : ~_GEN_2022 & _GEN_1951;
  wire        _GEN_2080 = _GEN_772 | _GEN_2023;
  wire        _GEN_2081 = _GEN_22 ? ~_GEN_2080 & _GEN_1953 : ~_GEN_2023 & _GEN_1953;
  wire        _GEN_2082 = _GEN_775 | _GEN_2024;
  wire        _GEN_2083 = _GEN_22 ? ~_GEN_2082 & _GEN_1955 : ~_GEN_2024 & _GEN_1955;
  wire        _GEN_2084 = _GEN_778 | _GEN_2025;
  wire        _GEN_2085 = _GEN_22 ? ~_GEN_2084 & _GEN_1957 : ~_GEN_2025 & _GEN_1957;
  wire        _GEN_2086 = _GEN_781 | _GEN_2026;
  wire        _GEN_2087 = _GEN_22 ? ~_GEN_2086 & _GEN_1959 : ~_GEN_2026 & _GEN_1959;
  wire        _GEN_2088 = _GEN_784 | _GEN_2027;
  wire        _GEN_2089 = _GEN_22 ? ~_GEN_2088 & _GEN_1961 : ~_GEN_2027 & _GEN_1961;
  wire        _GEN_2090 = _GEN_787 | _GEN_2028;
  wire        _GEN_2091 = _GEN_22 ? ~_GEN_2090 & _GEN_1963 : ~_GEN_2028 & _GEN_1963;
  wire        _GEN_2092 = (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_2029;
  wire        _GEN_2093 = _GEN_22 ? ~_GEN_2092 & _GEN_1965 : ~_GEN_2029 & _GEN_1965;
  wire        _GEN_2094 = _GEN_22 ? ~_GEN_2030 & _GEN_1966 : ~_GEN_1998 & _GEN_1966;
  wire        _GEN_2095 = _GEN_22 ? ~_GEN_2032 & _GEN_1967 : ~_GEN_1999 & _GEN_1967;
  wire        _GEN_2096 = _GEN_22 ? ~_GEN_2034 & _GEN_1968 : ~_GEN_2000 & _GEN_1968;
  wire        _GEN_2097 = _GEN_22 ? ~_GEN_2036 & _GEN_1969 : ~_GEN_2001 & _GEN_1969;
  wire        _GEN_2098 = _GEN_22 ? ~_GEN_2038 & _GEN_1970 : ~_GEN_2002 & _GEN_1970;
  wire        _GEN_2099 = _GEN_22 ? ~_GEN_2040 & _GEN_1971 : ~_GEN_2003 & _GEN_1971;
  wire        _GEN_2100 = _GEN_22 ? ~_GEN_2042 & _GEN_1972 : ~_GEN_2004 & _GEN_1972;
  wire        _GEN_2101 = _GEN_22 ? ~_GEN_2044 & _GEN_1973 : ~_GEN_2005 & _GEN_1973;
  wire        _GEN_2102 = _GEN_22 ? ~_GEN_2046 & _GEN_1974 : ~_GEN_2006 & _GEN_1974;
  wire        _GEN_2103 = _GEN_22 ? ~_GEN_2048 & _GEN_1975 : ~_GEN_2007 & _GEN_1975;
  wire        _GEN_2104 = _GEN_22 ? ~_GEN_2050 & _GEN_1976 : ~_GEN_2008 & _GEN_1976;
  wire        _GEN_2105 = _GEN_22 ? ~_GEN_2052 & _GEN_1977 : ~_GEN_2009 & _GEN_1977;
  wire        _GEN_2106 = _GEN_22 ? ~_GEN_2054 & _GEN_1978 : ~_GEN_2010 & _GEN_1978;
  wire        _GEN_2107 = _GEN_22 ? ~_GEN_2056 & _GEN_1979 : ~_GEN_2011 & _GEN_1979;
  wire        _GEN_2108 = _GEN_22 ? ~_GEN_2058 & _GEN_1980 : ~_GEN_2012 & _GEN_1980;
  wire        _GEN_2109 = _GEN_22 ? ~_GEN_2060 & _GEN_1981 : ~_GEN_2013 & _GEN_1981;
  wire        _GEN_2110 = _GEN_22 ? ~_GEN_2062 & _GEN_1982 : ~_GEN_2014 & _GEN_1982;
  wire        _GEN_2111 = _GEN_22 ? ~_GEN_2064 & _GEN_1983 : ~_GEN_2015 & _GEN_1983;
  wire        _GEN_2112 = _GEN_22 ? ~_GEN_2066 & _GEN_1984 : ~_GEN_2016 & _GEN_1984;
  wire        _GEN_2113 = _GEN_22 ? ~_GEN_2068 & _GEN_1985 : ~_GEN_2017 & _GEN_1985;
  wire        _GEN_2114 = _GEN_22 ? ~_GEN_2070 & _GEN_1986 : ~_GEN_2018 & _GEN_1986;
  wire        _GEN_2115 = _GEN_22 ? ~_GEN_2072 & _GEN_1987 : ~_GEN_2019 & _GEN_1987;
  wire        _GEN_2116 = _GEN_22 ? ~_GEN_2074 & _GEN_1988 : ~_GEN_2020 & _GEN_1988;
  wire        _GEN_2117 = _GEN_22 ? ~_GEN_2076 & _GEN_1989 : ~_GEN_2021 & _GEN_1989;
  wire        _GEN_2118 = _GEN_22 ? ~_GEN_2078 & _GEN_1990 : ~_GEN_2022 & _GEN_1990;
  wire        _GEN_2119 = _GEN_22 ? ~_GEN_2080 & _GEN_1991 : ~_GEN_2023 & _GEN_1991;
  wire        _GEN_2120 = _GEN_22 ? ~_GEN_2082 & _GEN_1992 : ~_GEN_2024 & _GEN_1992;
  wire        _GEN_2121 = _GEN_22 ? ~_GEN_2084 & _GEN_1993 : ~_GEN_2025 & _GEN_1993;
  wire        _GEN_2122 = _GEN_22 ? ~_GEN_2086 & _GEN_1994 : ~_GEN_2026 & _GEN_1994;
  wire        _GEN_2123 = _GEN_22 ? ~_GEN_2088 & _GEN_1995 : ~_GEN_2027 & _GEN_1995;
  wire        _GEN_2124 = _GEN_22 ? ~_GEN_2090 & _GEN_1996 : ~_GEN_2028 & _GEN_1996;
  wire        _GEN_2125 = _GEN_22 ? ~_GEN_2092 & _GEN_1997 : ~_GEN_2029 & _GEN_1997;
  wire        _GEN_2126 = _GEN_23 & _GEN_824;
  wire        _GEN_2127 = _GEN_23 & _GEN_826;
  wire        _GEN_2128 = _GEN_23 & _GEN_828;
  wire        _GEN_2129 = _GEN_23 & _GEN_830;
  wire        _GEN_2130 = _GEN_23 & _GEN_832;
  wire        _GEN_2131 = _GEN_23 & _GEN_834;
  wire        _GEN_2132 = _GEN_23 & _GEN_836;
  wire        _GEN_2133 = _GEN_23 & _GEN_838;
  wire        _GEN_2134 = _GEN_23 & _GEN_840;
  wire        _GEN_2135 = _GEN_23 & _GEN_842;
  wire        _GEN_2136 = _GEN_23 & _GEN_844;
  wire        _GEN_2137 = _GEN_23 & _GEN_846;
  wire        _GEN_2138 = _GEN_23 & _GEN_848;
  wire        _GEN_2139 = _GEN_23 & _GEN_850;
  wire        _GEN_2140 = _GEN_23 & _GEN_852;
  wire        _GEN_2141 = _GEN_23 & _GEN_854;
  wire        _GEN_2142 = _GEN_23 & _GEN_856;
  wire        _GEN_2143 = _GEN_23 & _GEN_858;
  wire        _GEN_2144 = _GEN_23 & _GEN_860;
  wire        _GEN_2145 = _GEN_23 & _GEN_862;
  wire        _GEN_2146 = _GEN_23 & _GEN_864;
  wire        _GEN_2147 = _GEN_23 & _GEN_866;
  wire        _GEN_2148 = _GEN_23 & _GEN_868;
  wire        _GEN_2149 = _GEN_23 & _GEN_870;
  wire        _GEN_2150 = _GEN_23 & _GEN_872;
  wire        _GEN_2151 = _GEN_23 & _GEN_874;
  wire        _GEN_2152 = _GEN_23 & _GEN_876;
  wire        _GEN_2153 = _GEN_23 & _GEN_878;
  wire        _GEN_2154 = _GEN_23 & _GEN_880;
  wire        _GEN_2155 = _GEN_23 & _GEN_882;
  wire        _GEN_2156 = _GEN_23 & _GEN_884;
  wire        _GEN_2157 = _GEN_23 & (&(io_wb_resps_6_bits_uop_rob_idx[6:2]));
  wire        _GEN_2158 = _GEN_887 | _GEN_2126;
  wire        _GEN_2159 = _GEN_24 ? ~_GEN_2158 & _GEN_2031 : ~_GEN_2126 & _GEN_2031;
  wire        _GEN_2160 = _GEN_890 | _GEN_2127;
  wire        _GEN_2161 = _GEN_24 ? ~_GEN_2160 & _GEN_2033 : ~_GEN_2127 & _GEN_2033;
  wire        _GEN_2162 = _GEN_893 | _GEN_2128;
  wire        _GEN_2163 = _GEN_24 ? ~_GEN_2162 & _GEN_2035 : ~_GEN_2128 & _GEN_2035;
  wire        _GEN_2164 = _GEN_896 | _GEN_2129;
  wire        _GEN_2165 = _GEN_24 ? ~_GEN_2164 & _GEN_2037 : ~_GEN_2129 & _GEN_2037;
  wire        _GEN_2166 = _GEN_899 | _GEN_2130;
  wire        _GEN_2167 = _GEN_24 ? ~_GEN_2166 & _GEN_2039 : ~_GEN_2130 & _GEN_2039;
  wire        _GEN_2168 = _GEN_902 | _GEN_2131;
  wire        _GEN_2169 = _GEN_24 ? ~_GEN_2168 & _GEN_2041 : ~_GEN_2131 & _GEN_2041;
  wire        _GEN_2170 = _GEN_905 | _GEN_2132;
  wire        _GEN_2171 = _GEN_24 ? ~_GEN_2170 & _GEN_2043 : ~_GEN_2132 & _GEN_2043;
  wire        _GEN_2172 = _GEN_908 | _GEN_2133;
  wire        _GEN_2173 = _GEN_24 ? ~_GEN_2172 & _GEN_2045 : ~_GEN_2133 & _GEN_2045;
  wire        _GEN_2174 = _GEN_911 | _GEN_2134;
  wire        _GEN_2175 = _GEN_24 ? ~_GEN_2174 & _GEN_2047 : ~_GEN_2134 & _GEN_2047;
  wire        _GEN_2176 = _GEN_914 | _GEN_2135;
  wire        _GEN_2177 = _GEN_24 ? ~_GEN_2176 & _GEN_2049 : ~_GEN_2135 & _GEN_2049;
  wire        _GEN_2178 = _GEN_917 | _GEN_2136;
  wire        _GEN_2179 = _GEN_24 ? ~_GEN_2178 & _GEN_2051 : ~_GEN_2136 & _GEN_2051;
  wire        _GEN_2180 = _GEN_920 | _GEN_2137;
  wire        _GEN_2181 = _GEN_24 ? ~_GEN_2180 & _GEN_2053 : ~_GEN_2137 & _GEN_2053;
  wire        _GEN_2182 = _GEN_923 | _GEN_2138;
  wire        _GEN_2183 = _GEN_24 ? ~_GEN_2182 & _GEN_2055 : ~_GEN_2138 & _GEN_2055;
  wire        _GEN_2184 = _GEN_926 | _GEN_2139;
  wire        _GEN_2185 = _GEN_24 ? ~_GEN_2184 & _GEN_2057 : ~_GEN_2139 & _GEN_2057;
  wire        _GEN_2186 = _GEN_929 | _GEN_2140;
  wire        _GEN_2187 = _GEN_24 ? ~_GEN_2186 & _GEN_2059 : ~_GEN_2140 & _GEN_2059;
  wire        _GEN_2188 = _GEN_932 | _GEN_2141;
  wire        _GEN_2189 = _GEN_24 ? ~_GEN_2188 & _GEN_2061 : ~_GEN_2141 & _GEN_2061;
  wire        _GEN_2190 = _GEN_935 | _GEN_2142;
  wire        _GEN_2191 = _GEN_24 ? ~_GEN_2190 & _GEN_2063 : ~_GEN_2142 & _GEN_2063;
  wire        _GEN_2192 = _GEN_938 | _GEN_2143;
  wire        _GEN_2193 = _GEN_24 ? ~_GEN_2192 & _GEN_2065 : ~_GEN_2143 & _GEN_2065;
  wire        _GEN_2194 = _GEN_941 | _GEN_2144;
  wire        _GEN_2195 = _GEN_24 ? ~_GEN_2194 & _GEN_2067 : ~_GEN_2144 & _GEN_2067;
  wire        _GEN_2196 = _GEN_944 | _GEN_2145;
  wire        _GEN_2197 = _GEN_24 ? ~_GEN_2196 & _GEN_2069 : ~_GEN_2145 & _GEN_2069;
  wire        _GEN_2198 = _GEN_947 | _GEN_2146;
  wire        _GEN_2199 = _GEN_24 ? ~_GEN_2198 & _GEN_2071 : ~_GEN_2146 & _GEN_2071;
  wire        _GEN_2200 = _GEN_950 | _GEN_2147;
  wire        _GEN_2201 = _GEN_24 ? ~_GEN_2200 & _GEN_2073 : ~_GEN_2147 & _GEN_2073;
  wire        _GEN_2202 = _GEN_953 | _GEN_2148;
  wire        _GEN_2203 = _GEN_24 ? ~_GEN_2202 & _GEN_2075 : ~_GEN_2148 & _GEN_2075;
  wire        _GEN_2204 = _GEN_956 | _GEN_2149;
  wire        _GEN_2205 = _GEN_24 ? ~_GEN_2204 & _GEN_2077 : ~_GEN_2149 & _GEN_2077;
  wire        _GEN_2206 = _GEN_959 | _GEN_2150;
  wire        _GEN_2207 = _GEN_24 ? ~_GEN_2206 & _GEN_2079 : ~_GEN_2150 & _GEN_2079;
  wire        _GEN_2208 = _GEN_962 | _GEN_2151;
  wire        _GEN_2209 = _GEN_24 ? ~_GEN_2208 & _GEN_2081 : ~_GEN_2151 & _GEN_2081;
  wire        _GEN_2210 = _GEN_965 | _GEN_2152;
  wire        _GEN_2211 = _GEN_24 ? ~_GEN_2210 & _GEN_2083 : ~_GEN_2152 & _GEN_2083;
  wire        _GEN_2212 = _GEN_968 | _GEN_2153;
  wire        _GEN_2213 = _GEN_24 ? ~_GEN_2212 & _GEN_2085 : ~_GEN_2153 & _GEN_2085;
  wire        _GEN_2214 = _GEN_971 | _GEN_2154;
  wire        _GEN_2215 = _GEN_24 ? ~_GEN_2214 & _GEN_2087 : ~_GEN_2154 & _GEN_2087;
  wire        _GEN_2216 = _GEN_974 | _GEN_2155;
  wire        _GEN_2217 = _GEN_24 ? ~_GEN_2216 & _GEN_2089 : ~_GEN_2155 & _GEN_2089;
  wire        _GEN_2218 = _GEN_977 | _GEN_2156;
  wire        _GEN_2219 = _GEN_24 ? ~_GEN_2218 & _GEN_2091 : ~_GEN_2156 & _GEN_2091;
  wire        _GEN_2220 = (&(io_wb_resps_7_bits_uop_rob_idx[6:2])) | _GEN_2157;
  wire        _GEN_2221 = _GEN_24 ? ~_GEN_2220 & _GEN_2093 : ~_GEN_2157 & _GEN_2093;
  wire        _GEN_2222 = _GEN_24 ? ~_GEN_2158 & _GEN_2094 : ~_GEN_2126 & _GEN_2094;
  wire        _GEN_2223 = _GEN_24 ? ~_GEN_2160 & _GEN_2095 : ~_GEN_2127 & _GEN_2095;
  wire        _GEN_2224 = _GEN_24 ? ~_GEN_2162 & _GEN_2096 : ~_GEN_2128 & _GEN_2096;
  wire        _GEN_2225 = _GEN_24 ? ~_GEN_2164 & _GEN_2097 : ~_GEN_2129 & _GEN_2097;
  wire        _GEN_2226 = _GEN_24 ? ~_GEN_2166 & _GEN_2098 : ~_GEN_2130 & _GEN_2098;
  wire        _GEN_2227 = _GEN_24 ? ~_GEN_2168 & _GEN_2099 : ~_GEN_2131 & _GEN_2099;
  wire        _GEN_2228 = _GEN_24 ? ~_GEN_2170 & _GEN_2100 : ~_GEN_2132 & _GEN_2100;
  wire        _GEN_2229 = _GEN_24 ? ~_GEN_2172 & _GEN_2101 : ~_GEN_2133 & _GEN_2101;
  wire        _GEN_2230 = _GEN_24 ? ~_GEN_2174 & _GEN_2102 : ~_GEN_2134 & _GEN_2102;
  wire        _GEN_2231 = _GEN_24 ? ~_GEN_2176 & _GEN_2103 : ~_GEN_2135 & _GEN_2103;
  wire        _GEN_2232 = _GEN_24 ? ~_GEN_2178 & _GEN_2104 : ~_GEN_2136 & _GEN_2104;
  wire        _GEN_2233 = _GEN_24 ? ~_GEN_2180 & _GEN_2105 : ~_GEN_2137 & _GEN_2105;
  wire        _GEN_2234 = _GEN_24 ? ~_GEN_2182 & _GEN_2106 : ~_GEN_2138 & _GEN_2106;
  wire        _GEN_2235 = _GEN_24 ? ~_GEN_2184 & _GEN_2107 : ~_GEN_2139 & _GEN_2107;
  wire        _GEN_2236 = _GEN_24 ? ~_GEN_2186 & _GEN_2108 : ~_GEN_2140 & _GEN_2108;
  wire        _GEN_2237 = _GEN_24 ? ~_GEN_2188 & _GEN_2109 : ~_GEN_2141 & _GEN_2109;
  wire        _GEN_2238 = _GEN_24 ? ~_GEN_2190 & _GEN_2110 : ~_GEN_2142 & _GEN_2110;
  wire        _GEN_2239 = _GEN_24 ? ~_GEN_2192 & _GEN_2111 : ~_GEN_2143 & _GEN_2111;
  wire        _GEN_2240 = _GEN_24 ? ~_GEN_2194 & _GEN_2112 : ~_GEN_2144 & _GEN_2112;
  wire        _GEN_2241 = _GEN_24 ? ~_GEN_2196 & _GEN_2113 : ~_GEN_2145 & _GEN_2113;
  wire        _GEN_2242 = _GEN_24 ? ~_GEN_2198 & _GEN_2114 : ~_GEN_2146 & _GEN_2114;
  wire        _GEN_2243 = _GEN_24 ? ~_GEN_2200 & _GEN_2115 : ~_GEN_2147 & _GEN_2115;
  wire        _GEN_2244 = _GEN_24 ? ~_GEN_2202 & _GEN_2116 : ~_GEN_2148 & _GEN_2116;
  wire        _GEN_2245 = _GEN_24 ? ~_GEN_2204 & _GEN_2117 : ~_GEN_2149 & _GEN_2117;
  wire        _GEN_2246 = _GEN_24 ? ~_GEN_2206 & _GEN_2118 : ~_GEN_2150 & _GEN_2118;
  wire        _GEN_2247 = _GEN_24 ? ~_GEN_2208 & _GEN_2119 : ~_GEN_2151 & _GEN_2119;
  wire        _GEN_2248 = _GEN_24 ? ~_GEN_2210 & _GEN_2120 : ~_GEN_2152 & _GEN_2120;
  wire        _GEN_2249 = _GEN_24 ? ~_GEN_2212 & _GEN_2121 : ~_GEN_2153 & _GEN_2121;
  wire        _GEN_2250 = _GEN_24 ? ~_GEN_2214 & _GEN_2122 : ~_GEN_2154 & _GEN_2122;
  wire        _GEN_2251 = _GEN_24 ? ~_GEN_2216 & _GEN_2123 : ~_GEN_2155 & _GEN_2123;
  wire        _GEN_2252 = _GEN_24 ? ~_GEN_2218 & _GEN_2124 : ~_GEN_2156 & _GEN_2124;
  wire        _GEN_2253 = _GEN_24 ? ~_GEN_2220 & _GEN_2125 : ~_GEN_2157 & _GEN_2125;
  wire        _GEN_2254 = _GEN_25 & _GEN_1014;
  wire        _GEN_2255 = _GEN_25 & _GEN_1016;
  wire        _GEN_2256 = _GEN_25 & _GEN_1018;
  wire        _GEN_2257 = _GEN_25 & _GEN_1020;
  wire        _GEN_2258 = _GEN_25 & _GEN_1022;
  wire        _GEN_2259 = _GEN_25 & _GEN_1024;
  wire        _GEN_2260 = _GEN_25 & _GEN_1026;
  wire        _GEN_2261 = _GEN_25 & _GEN_1028;
  wire        _GEN_2262 = _GEN_25 & _GEN_1030;
  wire        _GEN_2263 = _GEN_25 & _GEN_1032;
  wire        _GEN_2264 = _GEN_25 & _GEN_1034;
  wire        _GEN_2265 = _GEN_25 & _GEN_1036;
  wire        _GEN_2266 = _GEN_25 & _GEN_1038;
  wire        _GEN_2267 = _GEN_25 & _GEN_1040;
  wire        _GEN_2268 = _GEN_25 & _GEN_1042;
  wire        _GEN_2269 = _GEN_25 & _GEN_1044;
  wire        _GEN_2270 = _GEN_25 & _GEN_1046;
  wire        _GEN_2271 = _GEN_25 & _GEN_1048;
  wire        _GEN_2272 = _GEN_25 & _GEN_1050;
  wire        _GEN_2273 = _GEN_25 & _GEN_1052;
  wire        _GEN_2274 = _GEN_25 & _GEN_1054;
  wire        _GEN_2275 = _GEN_25 & _GEN_1056;
  wire        _GEN_2276 = _GEN_25 & _GEN_1058;
  wire        _GEN_2277 = _GEN_25 & _GEN_1060;
  wire        _GEN_2278 = _GEN_25 & _GEN_1062;
  wire        _GEN_2279 = _GEN_25 & _GEN_1064;
  wire        _GEN_2280 = _GEN_25 & _GEN_1066;
  wire        _GEN_2281 = _GEN_25 & _GEN_1068;
  wire        _GEN_2282 = _GEN_25 & _GEN_1070;
  wire        _GEN_2283 = _GEN_25 & _GEN_1072;
  wire        _GEN_2284 = _GEN_25 & _GEN_1074;
  wire        _GEN_2285 = _GEN_25 & (&(io_wb_resps_8_bits_uop_rob_idx[6:2]));
  wire        _GEN_2286 = _GEN_1077 | _GEN_2254;
  wire        _GEN_2287 = _GEN_26 ? ~_GEN_2286 & _GEN_2159 : ~_GEN_2254 & _GEN_2159;
  wire        _GEN_2288 = _GEN_1080 | _GEN_2255;
  wire        _GEN_2289 = _GEN_26 ? ~_GEN_2288 & _GEN_2161 : ~_GEN_2255 & _GEN_2161;
  wire        _GEN_2290 = _GEN_1083 | _GEN_2256;
  wire        _GEN_2291 = _GEN_26 ? ~_GEN_2290 & _GEN_2163 : ~_GEN_2256 & _GEN_2163;
  wire        _GEN_2292 = _GEN_1086 | _GEN_2257;
  wire        _GEN_2293 = _GEN_26 ? ~_GEN_2292 & _GEN_2165 : ~_GEN_2257 & _GEN_2165;
  wire        _GEN_2294 = _GEN_1089 | _GEN_2258;
  wire        _GEN_2295 = _GEN_26 ? ~_GEN_2294 & _GEN_2167 : ~_GEN_2258 & _GEN_2167;
  wire        _GEN_2296 = _GEN_1092 | _GEN_2259;
  wire        _GEN_2297 = _GEN_26 ? ~_GEN_2296 & _GEN_2169 : ~_GEN_2259 & _GEN_2169;
  wire        _GEN_2298 = _GEN_1095 | _GEN_2260;
  wire        _GEN_2299 = _GEN_26 ? ~_GEN_2298 & _GEN_2171 : ~_GEN_2260 & _GEN_2171;
  wire        _GEN_2300 = _GEN_1098 | _GEN_2261;
  wire        _GEN_2301 = _GEN_26 ? ~_GEN_2300 & _GEN_2173 : ~_GEN_2261 & _GEN_2173;
  wire        _GEN_2302 = _GEN_1101 | _GEN_2262;
  wire        _GEN_2303 = _GEN_26 ? ~_GEN_2302 & _GEN_2175 : ~_GEN_2262 & _GEN_2175;
  wire        _GEN_2304 = _GEN_1104 | _GEN_2263;
  wire        _GEN_2305 = _GEN_26 ? ~_GEN_2304 & _GEN_2177 : ~_GEN_2263 & _GEN_2177;
  wire        _GEN_2306 = _GEN_1107 | _GEN_2264;
  wire        _GEN_2307 = _GEN_26 ? ~_GEN_2306 & _GEN_2179 : ~_GEN_2264 & _GEN_2179;
  wire        _GEN_2308 = _GEN_1110 | _GEN_2265;
  wire        _GEN_2309 = _GEN_26 ? ~_GEN_2308 & _GEN_2181 : ~_GEN_2265 & _GEN_2181;
  wire        _GEN_2310 = _GEN_1113 | _GEN_2266;
  wire        _GEN_2311 = _GEN_26 ? ~_GEN_2310 & _GEN_2183 : ~_GEN_2266 & _GEN_2183;
  wire        _GEN_2312 = _GEN_1116 | _GEN_2267;
  wire        _GEN_2313 = _GEN_26 ? ~_GEN_2312 & _GEN_2185 : ~_GEN_2267 & _GEN_2185;
  wire        _GEN_2314 = _GEN_1119 | _GEN_2268;
  wire        _GEN_2315 = _GEN_26 ? ~_GEN_2314 & _GEN_2187 : ~_GEN_2268 & _GEN_2187;
  wire        _GEN_2316 = _GEN_1122 | _GEN_2269;
  wire        _GEN_2317 = _GEN_26 ? ~_GEN_2316 & _GEN_2189 : ~_GEN_2269 & _GEN_2189;
  wire        _GEN_2318 = _GEN_1125 | _GEN_2270;
  wire        _GEN_2319 = _GEN_26 ? ~_GEN_2318 & _GEN_2191 : ~_GEN_2270 & _GEN_2191;
  wire        _GEN_2320 = _GEN_1128 | _GEN_2271;
  wire        _GEN_2321 = _GEN_26 ? ~_GEN_2320 & _GEN_2193 : ~_GEN_2271 & _GEN_2193;
  wire        _GEN_2322 = _GEN_1131 | _GEN_2272;
  wire        _GEN_2323 = _GEN_26 ? ~_GEN_2322 & _GEN_2195 : ~_GEN_2272 & _GEN_2195;
  wire        _GEN_2324 = _GEN_1134 | _GEN_2273;
  wire        _GEN_2325 = _GEN_26 ? ~_GEN_2324 & _GEN_2197 : ~_GEN_2273 & _GEN_2197;
  wire        _GEN_2326 = _GEN_1137 | _GEN_2274;
  wire        _GEN_2327 = _GEN_26 ? ~_GEN_2326 & _GEN_2199 : ~_GEN_2274 & _GEN_2199;
  wire        _GEN_2328 = _GEN_1140 | _GEN_2275;
  wire        _GEN_2329 = _GEN_26 ? ~_GEN_2328 & _GEN_2201 : ~_GEN_2275 & _GEN_2201;
  wire        _GEN_2330 = _GEN_1143 | _GEN_2276;
  wire        _GEN_2331 = _GEN_26 ? ~_GEN_2330 & _GEN_2203 : ~_GEN_2276 & _GEN_2203;
  wire        _GEN_2332 = _GEN_1146 | _GEN_2277;
  wire        _GEN_2333 = _GEN_26 ? ~_GEN_2332 & _GEN_2205 : ~_GEN_2277 & _GEN_2205;
  wire        _GEN_2334 = _GEN_1149 | _GEN_2278;
  wire        _GEN_2335 = _GEN_26 ? ~_GEN_2334 & _GEN_2207 : ~_GEN_2278 & _GEN_2207;
  wire        _GEN_2336 = _GEN_1152 | _GEN_2279;
  wire        _GEN_2337 = _GEN_26 ? ~_GEN_2336 & _GEN_2209 : ~_GEN_2279 & _GEN_2209;
  wire        _GEN_2338 = _GEN_1155 | _GEN_2280;
  wire        _GEN_2339 = _GEN_26 ? ~_GEN_2338 & _GEN_2211 : ~_GEN_2280 & _GEN_2211;
  wire        _GEN_2340 = _GEN_1158 | _GEN_2281;
  wire        _GEN_2341 = _GEN_26 ? ~_GEN_2340 & _GEN_2213 : ~_GEN_2281 & _GEN_2213;
  wire        _GEN_2342 = _GEN_1161 | _GEN_2282;
  wire        _GEN_2343 = _GEN_26 ? ~_GEN_2342 & _GEN_2215 : ~_GEN_2282 & _GEN_2215;
  wire        _GEN_2344 = _GEN_1164 | _GEN_2283;
  wire        _GEN_2345 = _GEN_26 ? ~_GEN_2344 & _GEN_2217 : ~_GEN_2283 & _GEN_2217;
  wire        _GEN_2346 = _GEN_1167 | _GEN_2284;
  wire        _GEN_2347 = _GEN_26 ? ~_GEN_2346 & _GEN_2219 : ~_GEN_2284 & _GEN_2219;
  wire        _GEN_2348 = (&(io_wb_resps_9_bits_uop_rob_idx[6:2])) | _GEN_2285;
  wire        _GEN_2349 = _GEN_26 ? ~_GEN_2348 & _GEN_2221 : ~_GEN_2285 & _GEN_2221;
  wire        _GEN_2350 = _GEN_26 ? ~_GEN_2286 & _GEN_2222 : ~_GEN_2254 & _GEN_2222;
  wire        _GEN_2351 = _GEN_26 ? ~_GEN_2288 & _GEN_2223 : ~_GEN_2255 & _GEN_2223;
  wire        _GEN_2352 = _GEN_26 ? ~_GEN_2290 & _GEN_2224 : ~_GEN_2256 & _GEN_2224;
  wire        _GEN_2353 = _GEN_26 ? ~_GEN_2292 & _GEN_2225 : ~_GEN_2257 & _GEN_2225;
  wire        _GEN_2354 = _GEN_26 ? ~_GEN_2294 & _GEN_2226 : ~_GEN_2258 & _GEN_2226;
  wire        _GEN_2355 = _GEN_26 ? ~_GEN_2296 & _GEN_2227 : ~_GEN_2259 & _GEN_2227;
  wire        _GEN_2356 = _GEN_26 ? ~_GEN_2298 & _GEN_2228 : ~_GEN_2260 & _GEN_2228;
  wire        _GEN_2357 = _GEN_26 ? ~_GEN_2300 & _GEN_2229 : ~_GEN_2261 & _GEN_2229;
  wire        _GEN_2358 = _GEN_26 ? ~_GEN_2302 & _GEN_2230 : ~_GEN_2262 & _GEN_2230;
  wire        _GEN_2359 = _GEN_26 ? ~_GEN_2304 & _GEN_2231 : ~_GEN_2263 & _GEN_2231;
  wire        _GEN_2360 = _GEN_26 ? ~_GEN_2306 & _GEN_2232 : ~_GEN_2264 & _GEN_2232;
  wire        _GEN_2361 = _GEN_26 ? ~_GEN_2308 & _GEN_2233 : ~_GEN_2265 & _GEN_2233;
  wire        _GEN_2362 = _GEN_26 ? ~_GEN_2310 & _GEN_2234 : ~_GEN_2266 & _GEN_2234;
  wire        _GEN_2363 = _GEN_26 ? ~_GEN_2312 & _GEN_2235 : ~_GEN_2267 & _GEN_2235;
  wire        _GEN_2364 = _GEN_26 ? ~_GEN_2314 & _GEN_2236 : ~_GEN_2268 & _GEN_2236;
  wire        _GEN_2365 = _GEN_26 ? ~_GEN_2316 & _GEN_2237 : ~_GEN_2269 & _GEN_2237;
  wire        _GEN_2366 = _GEN_26 ? ~_GEN_2318 & _GEN_2238 : ~_GEN_2270 & _GEN_2238;
  wire        _GEN_2367 = _GEN_26 ? ~_GEN_2320 & _GEN_2239 : ~_GEN_2271 & _GEN_2239;
  wire        _GEN_2368 = _GEN_26 ? ~_GEN_2322 & _GEN_2240 : ~_GEN_2272 & _GEN_2240;
  wire        _GEN_2369 = _GEN_26 ? ~_GEN_2324 & _GEN_2241 : ~_GEN_2273 & _GEN_2241;
  wire        _GEN_2370 = _GEN_26 ? ~_GEN_2326 & _GEN_2242 : ~_GEN_2274 & _GEN_2242;
  wire        _GEN_2371 = _GEN_26 ? ~_GEN_2328 & _GEN_2243 : ~_GEN_2275 & _GEN_2243;
  wire        _GEN_2372 = _GEN_26 ? ~_GEN_2330 & _GEN_2244 : ~_GEN_2276 & _GEN_2244;
  wire        _GEN_2373 = _GEN_26 ? ~_GEN_2332 & _GEN_2245 : ~_GEN_2277 & _GEN_2245;
  wire        _GEN_2374 = _GEN_26 ? ~_GEN_2334 & _GEN_2246 : ~_GEN_2278 & _GEN_2246;
  wire        _GEN_2375 = _GEN_26 ? ~_GEN_2336 & _GEN_2247 : ~_GEN_2279 & _GEN_2247;
  wire        _GEN_2376 = _GEN_26 ? ~_GEN_2338 & _GEN_2248 : ~_GEN_2280 & _GEN_2248;
  wire        _GEN_2377 = _GEN_26 ? ~_GEN_2340 & _GEN_2249 : ~_GEN_2281 & _GEN_2249;
  wire        _GEN_2378 = _GEN_26 ? ~_GEN_2342 & _GEN_2250 : ~_GEN_2282 & _GEN_2250;
  wire        _GEN_2379 = _GEN_26 ? ~_GEN_2344 & _GEN_2251 : ~_GEN_2283 & _GEN_2251;
  wire        _GEN_2380 = _GEN_26 ? ~_GEN_2346 & _GEN_2252 : ~_GEN_2284 & _GEN_2252;
  wire        _GEN_2381 = _GEN_26 ? ~_GEN_2348 & _GEN_2253 : ~_GEN_2285 & _GEN_2253;
  wire        _GEN_2382 = _GEN_27 & _GEN_1204;
  wire        _GEN_2383 = _GEN_27 & _GEN_1206;
  wire        _GEN_2384 = _GEN_27 & _GEN_1208;
  wire        _GEN_2385 = _GEN_27 & _GEN_1210;
  wire        _GEN_2386 = _GEN_27 & _GEN_1212;
  wire        _GEN_2387 = _GEN_27 & _GEN_1214;
  wire        _GEN_2388 = _GEN_27 & _GEN_1216;
  wire        _GEN_2389 = _GEN_27 & _GEN_1218;
  wire        _GEN_2390 = _GEN_27 & _GEN_1220;
  wire        _GEN_2391 = _GEN_27 & _GEN_1222;
  wire        _GEN_2392 = _GEN_27 & _GEN_1224;
  wire        _GEN_2393 = _GEN_27 & _GEN_1226;
  wire        _GEN_2394 = _GEN_27 & _GEN_1228;
  wire        _GEN_2395 = _GEN_27 & _GEN_1230;
  wire        _GEN_2396 = _GEN_27 & _GEN_1232;
  wire        _GEN_2397 = _GEN_27 & _GEN_1234;
  wire        _GEN_2398 = _GEN_27 & _GEN_1236;
  wire        _GEN_2399 = _GEN_27 & _GEN_1238;
  wire        _GEN_2400 = _GEN_27 & _GEN_1240;
  wire        _GEN_2401 = _GEN_27 & _GEN_1242;
  wire        _GEN_2402 = _GEN_27 & _GEN_1244;
  wire        _GEN_2403 = _GEN_27 & _GEN_1246;
  wire        _GEN_2404 = _GEN_27 & _GEN_1248;
  wire        _GEN_2405 = _GEN_27 & _GEN_1250;
  wire        _GEN_2406 = _GEN_27 & _GEN_1252;
  wire        _GEN_2407 = _GEN_27 & _GEN_1254;
  wire        _GEN_2408 = _GEN_27 & _GEN_1256;
  wire        _GEN_2409 = _GEN_27 & _GEN_1258;
  wire        _GEN_2410 = _GEN_27 & _GEN_1260;
  wire        _GEN_2411 = _GEN_27 & _GEN_1262;
  wire        _GEN_2412 = _GEN_27 & _GEN_1264;
  wire        _GEN_2413 = _GEN_27 & (&(io_lsu_clr_bsy_0_bits[6:2]));
  wire        _GEN_2414 = _GEN_1267 | _GEN_2382;
  wire        _GEN_2415 = _GEN_1269 | _GEN_2383;
  wire        _GEN_2416 = _GEN_1271 | _GEN_2384;
  wire        _GEN_2417 = _GEN_1273 | _GEN_2385;
  wire        _GEN_2418 = _GEN_1275 | _GEN_2386;
  wire        _GEN_2419 = _GEN_1277 | _GEN_2387;
  wire        _GEN_2420 = _GEN_1279 | _GEN_2388;
  wire        _GEN_2421 = _GEN_1281 | _GEN_2389;
  wire        _GEN_2422 = _GEN_1283 | _GEN_2390;
  wire        _GEN_2423 = _GEN_1285 | _GEN_2391;
  wire        _GEN_2424 = _GEN_1287 | _GEN_2392;
  wire        _GEN_2425 = _GEN_1289 | _GEN_2393;
  wire        _GEN_2426 = _GEN_1291 | _GEN_2394;
  wire        _GEN_2427 = _GEN_1293 | _GEN_2395;
  wire        _GEN_2428 = _GEN_1295 | _GEN_2396;
  wire        _GEN_2429 = _GEN_1297 | _GEN_2397;
  wire        _GEN_2430 = _GEN_1299 | _GEN_2398;
  wire        _GEN_2431 = _GEN_1301 | _GEN_2399;
  wire        _GEN_2432 = _GEN_1303 | _GEN_2400;
  wire        _GEN_2433 = _GEN_1305 | _GEN_2401;
  wire        _GEN_2434 = _GEN_1307 | _GEN_2402;
  wire        _GEN_2435 = _GEN_1309 | _GEN_2403;
  wire        _GEN_2436 = _GEN_1311 | _GEN_2404;
  wire        _GEN_2437 = _GEN_1313 | _GEN_2405;
  wire        _GEN_2438 = _GEN_1315 | _GEN_2406;
  wire        _GEN_2439 = _GEN_1317 | _GEN_2407;
  wire        _GEN_2440 = _GEN_1319 | _GEN_2408;
  wire        _GEN_2441 = _GEN_1321 | _GEN_2409;
  wire        _GEN_2442 = _GEN_1323 | _GEN_2410;
  wire        _GEN_2443 = _GEN_1325 | _GEN_2411;
  wire        _GEN_2444 = _GEN_1327 | _GEN_2412;
  wire        _GEN_2445 = (&(io_lsu_clr_bsy_1_bits[6:2])) | _GEN_2413;
  wire        _GEN_2446 = _GEN_29 & _GEN_1330;
  wire        _GEN_2447 = _GEN_29 & _GEN_1332;
  wire        _GEN_2448 = _GEN_29 & _GEN_1334;
  wire        _GEN_2449 = _GEN_29 & _GEN_1336;
  wire        _GEN_2450 = _GEN_29 & _GEN_1338;
  wire        _GEN_2451 = _GEN_29 & _GEN_1340;
  wire        _GEN_2452 = _GEN_29 & _GEN_1342;
  wire        _GEN_2453 = _GEN_29 & _GEN_1344;
  wire        _GEN_2454 = _GEN_29 & _GEN_1346;
  wire        _GEN_2455 = _GEN_29 & _GEN_1348;
  wire        _GEN_2456 = _GEN_29 & _GEN_1350;
  wire        _GEN_2457 = _GEN_29 & _GEN_1352;
  wire        _GEN_2458 = _GEN_29 & _GEN_1354;
  wire        _GEN_2459 = _GEN_29 & _GEN_1356;
  wire        _GEN_2460 = _GEN_29 & _GEN_1358;
  wire        _GEN_2461 = _GEN_29 & _GEN_1360;
  wire        _GEN_2462 = _GEN_29 & _GEN_1362;
  wire        _GEN_2463 = _GEN_29 & _GEN_1364;
  wire        _GEN_2464 = _GEN_29 & _GEN_1366;
  wire        _GEN_2465 = _GEN_29 & _GEN_1368;
  wire        _GEN_2466 = _GEN_29 & _GEN_1370;
  wire        _GEN_2467 = _GEN_29 & _GEN_1372;
  wire        _GEN_2468 = _GEN_29 & _GEN_1374;
  wire        _GEN_2469 = _GEN_29 & _GEN_1376;
  wire        _GEN_2470 = _GEN_29 & _GEN_1378;
  wire        _GEN_2471 = _GEN_29 & _GEN_1380;
  wire        _GEN_2472 = _GEN_29 & _GEN_1382;
  wire        _GEN_2473 = _GEN_29 & _GEN_1384;
  wire        _GEN_2474 = _GEN_29 & _GEN_1386;
  wire        _GEN_2475 = _GEN_29 & _GEN_1388;
  wire        _GEN_2476 = _GEN_29 & _GEN_1390;
  wire        _GEN_2477 = _GEN_29 & (&(io_lsu_clr_bsy_2_bits[6:2]));
  wire        _GEN_2478 = io_fflags_0_valid & io_fflags_0_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_2479 = io_fflags_2_valid & io_fflags_2_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_2480 = io_fflags_3_valid & io_fflags_3_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_2481 = rbk_row_1 & _GEN_1520;
  wire        _GEN_2482 = rbk_row_1 & _GEN_1522;
  wire        _GEN_2483 = rbk_row_1 & _GEN_1524;
  wire        _GEN_2484 = rbk_row_1 & _GEN_1526;
  wire        _GEN_2485 = rbk_row_1 & _GEN_1528;
  wire        _GEN_2486 = rbk_row_1 & _GEN_1530;
  wire        _GEN_2487 = rbk_row_1 & _GEN_1532;
  wire        _GEN_2488 = rbk_row_1 & _GEN_1534;
  wire        _GEN_2489 = rbk_row_1 & _GEN_1536;
  wire        _GEN_2490 = rbk_row_1 & _GEN_1538;
  wire        _GEN_2491 = rbk_row_1 & _GEN_1540;
  wire        _GEN_2492 = rbk_row_1 & _GEN_1542;
  wire        _GEN_2493 = rbk_row_1 & _GEN_1544;
  wire        _GEN_2494 = rbk_row_1 & _GEN_1546;
  wire        _GEN_2495 = rbk_row_1 & _GEN_1548;
  wire        _GEN_2496 = rbk_row_1 & _GEN_1550;
  wire        _GEN_2497 = rbk_row_1 & _GEN_1552;
  wire        _GEN_2498 = rbk_row_1 & _GEN_1554;
  wire        _GEN_2499 = rbk_row_1 & _GEN_1556;
  wire        _GEN_2500 = rbk_row_1 & _GEN_1558;
  wire        _GEN_2501 = rbk_row_1 & _GEN_1560;
  wire        _GEN_2502 = rbk_row_1 & _GEN_1562;
  wire        _GEN_2503 = rbk_row_1 & _GEN_1564;
  wire        _GEN_2504 = rbk_row_1 & _GEN_1566;
  wire        _GEN_2505 = rbk_row_1 & _GEN_1568;
  wire        _GEN_2506 = rbk_row_1 & _GEN_1570;
  wire        _GEN_2507 = rbk_row_1 & _GEN_1572;
  wire        _GEN_2508 = rbk_row_1 & _GEN_1574;
  wire        _GEN_2509 = rbk_row_1 & _GEN_1576;
  wire        _GEN_2510 = rbk_row_1 & _GEN_1578;
  wire        _GEN_2511 = rbk_row_1 & _GEN_1580;
  wire        _GEN_2512 = rbk_row_1 & (&com_idx);
  wire [19:0] _GEN_2513 = io_brupdate_b1_mispredict_mask & rob_uop_1_0_br_mask;
  wire [19:0] _GEN_2514 = io_brupdate_b1_mispredict_mask & rob_uop_1_1_br_mask;
  wire [19:0] _GEN_2515 = io_brupdate_b1_mispredict_mask & rob_uop_1_2_br_mask;
  wire [19:0] _GEN_2516 = io_brupdate_b1_mispredict_mask & rob_uop_1_3_br_mask;
  wire [19:0] _GEN_2517 = io_brupdate_b1_mispredict_mask & rob_uop_1_4_br_mask;
  wire [19:0] _GEN_2518 = io_brupdate_b1_mispredict_mask & rob_uop_1_5_br_mask;
  wire [19:0] _GEN_2519 = io_brupdate_b1_mispredict_mask & rob_uop_1_6_br_mask;
  wire [19:0] _GEN_2520 = io_brupdate_b1_mispredict_mask & rob_uop_1_7_br_mask;
  wire [19:0] _GEN_2521 = io_brupdate_b1_mispredict_mask & rob_uop_1_8_br_mask;
  wire [19:0] _GEN_2522 = io_brupdate_b1_mispredict_mask & rob_uop_1_9_br_mask;
  wire [19:0] _GEN_2523 = io_brupdate_b1_mispredict_mask & rob_uop_1_10_br_mask;
  wire [19:0] _GEN_2524 = io_brupdate_b1_mispredict_mask & rob_uop_1_11_br_mask;
  wire [19:0] _GEN_2525 = io_brupdate_b1_mispredict_mask & rob_uop_1_12_br_mask;
  wire [19:0] _GEN_2526 = io_brupdate_b1_mispredict_mask & rob_uop_1_13_br_mask;
  wire [19:0] _GEN_2527 = io_brupdate_b1_mispredict_mask & rob_uop_1_14_br_mask;
  wire [19:0] _GEN_2528 = io_brupdate_b1_mispredict_mask & rob_uop_1_15_br_mask;
  wire [19:0] _GEN_2529 = io_brupdate_b1_mispredict_mask & rob_uop_1_16_br_mask;
  wire [19:0] _GEN_2530 = io_brupdate_b1_mispredict_mask & rob_uop_1_17_br_mask;
  wire [19:0] _GEN_2531 = io_brupdate_b1_mispredict_mask & rob_uop_1_18_br_mask;
  wire [19:0] _GEN_2532 = io_brupdate_b1_mispredict_mask & rob_uop_1_19_br_mask;
  wire [19:0] _GEN_2533 = io_brupdate_b1_mispredict_mask & rob_uop_1_20_br_mask;
  wire [19:0] _GEN_2534 = io_brupdate_b1_mispredict_mask & rob_uop_1_21_br_mask;
  wire [19:0] _GEN_2535 = io_brupdate_b1_mispredict_mask & rob_uop_1_22_br_mask;
  wire [19:0] _GEN_2536 = io_brupdate_b1_mispredict_mask & rob_uop_1_23_br_mask;
  wire [19:0] _GEN_2537 = io_brupdate_b1_mispredict_mask & rob_uop_1_24_br_mask;
  wire [19:0] _GEN_2538 = io_brupdate_b1_mispredict_mask & rob_uop_1_25_br_mask;
  wire [19:0] _GEN_2539 = io_brupdate_b1_mispredict_mask & rob_uop_1_26_br_mask;
  wire [19:0] _GEN_2540 = io_brupdate_b1_mispredict_mask & rob_uop_1_27_br_mask;
  wire [19:0] _GEN_2541 = io_brupdate_b1_mispredict_mask & rob_uop_1_28_br_mask;
  wire [19:0] _GEN_2542 = io_brupdate_b1_mispredict_mask & rob_uop_1_29_br_mask;
  wire [19:0] _GEN_2543 = io_brupdate_b1_mispredict_mask & rob_uop_1_30_br_mask;
  wire [19:0] _GEN_2544 = io_brupdate_b1_mispredict_mask & rob_uop_1_31_br_mask;
  wire        _GEN_2545 = io_enq_valids_2 & _GEN_127;
  wire        _GEN_2546 = io_enq_valids_2 & _GEN_129;
  wire        _GEN_2547 = io_enq_valids_2 & _GEN_131;
  wire        _GEN_2548 = io_enq_valids_2 & _GEN_133;
  wire        _GEN_2549 = io_enq_valids_2 & _GEN_135;
  wire        _GEN_2550 = io_enq_valids_2 & _GEN_137;
  wire        _GEN_2551 = io_enq_valids_2 & _GEN_139;
  wire        _GEN_2552 = io_enq_valids_2 & _GEN_141;
  wire        _GEN_2553 = io_enq_valids_2 & _GEN_143;
  wire        _GEN_2554 = io_enq_valids_2 & _GEN_145;
  wire        _GEN_2555 = io_enq_valids_2 & _GEN_147;
  wire        _GEN_2556 = io_enq_valids_2 & _GEN_149;
  wire        _GEN_2557 = io_enq_valids_2 & _GEN_151;
  wire        _GEN_2558 = io_enq_valids_2 & _GEN_153;
  wire        _GEN_2559 = io_enq_valids_2 & _GEN_155;
  wire        _GEN_2560 = io_enq_valids_2 & _GEN_157;
  wire        _GEN_2561 = io_enq_valids_2 & _GEN_159;
  wire        _GEN_2562 = io_enq_valids_2 & _GEN_161;
  wire        _GEN_2563 = io_enq_valids_2 & _GEN_163;
  wire        _GEN_2564 = io_enq_valids_2 & _GEN_165;
  wire        _GEN_2565 = io_enq_valids_2 & _GEN_167;
  wire        _GEN_2566 = io_enq_valids_2 & _GEN_169;
  wire        _GEN_2567 = io_enq_valids_2 & _GEN_171;
  wire        _GEN_2568 = io_enq_valids_2 & _GEN_173;
  wire        _GEN_2569 = io_enq_valids_2 & _GEN_175;
  wire        _GEN_2570 = io_enq_valids_2 & _GEN_177;
  wire        _GEN_2571 = io_enq_valids_2 & _GEN_179;
  wire        _GEN_2572 = io_enq_valids_2 & _GEN_181;
  wire        _GEN_2573 = io_enq_valids_2 & _GEN_183;
  wire        _GEN_2574 = io_enq_valids_2 & _GEN_185;
  wire        _GEN_2575 = io_enq_valids_2 & _GEN_187;
  wire        _GEN_2576 = io_enq_valids_2 & (&rob_tail);
  wire        _rob_bsy_T_4 = io_enq_uops_2_is_fence | io_enq_uops_2_is_fencei;
  wire        _GEN_2577 = _GEN_2545 ? ~_rob_bsy_T_4 : rob_bsy_2_0;
  wire        _GEN_2578 = _GEN_2546 ? ~_rob_bsy_T_4 : rob_bsy_2_1;
  wire        _GEN_2579 = _GEN_2547 ? ~_rob_bsy_T_4 : rob_bsy_2_2;
  wire        _GEN_2580 = _GEN_2548 ? ~_rob_bsy_T_4 : rob_bsy_2_3;
  wire        _GEN_2581 = _GEN_2549 ? ~_rob_bsy_T_4 : rob_bsy_2_4;
  wire        _GEN_2582 = _GEN_2550 ? ~_rob_bsy_T_4 : rob_bsy_2_5;
  wire        _GEN_2583 = _GEN_2551 ? ~_rob_bsy_T_4 : rob_bsy_2_6;
  wire        _GEN_2584 = _GEN_2552 ? ~_rob_bsy_T_4 : rob_bsy_2_7;
  wire        _GEN_2585 = _GEN_2553 ? ~_rob_bsy_T_4 : rob_bsy_2_8;
  wire        _GEN_2586 = _GEN_2554 ? ~_rob_bsy_T_4 : rob_bsy_2_9;
  wire        _GEN_2587 = _GEN_2555 ? ~_rob_bsy_T_4 : rob_bsy_2_10;
  wire        _GEN_2588 = _GEN_2556 ? ~_rob_bsy_T_4 : rob_bsy_2_11;
  wire        _GEN_2589 = _GEN_2557 ? ~_rob_bsy_T_4 : rob_bsy_2_12;
  wire        _GEN_2590 = _GEN_2558 ? ~_rob_bsy_T_4 : rob_bsy_2_13;
  wire        _GEN_2591 = _GEN_2559 ? ~_rob_bsy_T_4 : rob_bsy_2_14;
  wire        _GEN_2592 = _GEN_2560 ? ~_rob_bsy_T_4 : rob_bsy_2_15;
  wire        _GEN_2593 = _GEN_2561 ? ~_rob_bsy_T_4 : rob_bsy_2_16;
  wire        _GEN_2594 = _GEN_2562 ? ~_rob_bsy_T_4 : rob_bsy_2_17;
  wire        _GEN_2595 = _GEN_2563 ? ~_rob_bsy_T_4 : rob_bsy_2_18;
  wire        _GEN_2596 = _GEN_2564 ? ~_rob_bsy_T_4 : rob_bsy_2_19;
  wire        _GEN_2597 = _GEN_2565 ? ~_rob_bsy_T_4 : rob_bsy_2_20;
  wire        _GEN_2598 = _GEN_2566 ? ~_rob_bsy_T_4 : rob_bsy_2_21;
  wire        _GEN_2599 = _GEN_2567 ? ~_rob_bsy_T_4 : rob_bsy_2_22;
  wire        _GEN_2600 = _GEN_2568 ? ~_rob_bsy_T_4 : rob_bsy_2_23;
  wire        _GEN_2601 = _GEN_2569 ? ~_rob_bsy_T_4 : rob_bsy_2_24;
  wire        _GEN_2602 = _GEN_2570 ? ~_rob_bsy_T_4 : rob_bsy_2_25;
  wire        _GEN_2603 = _GEN_2571 ? ~_rob_bsy_T_4 : rob_bsy_2_26;
  wire        _GEN_2604 = _GEN_2572 ? ~_rob_bsy_T_4 : rob_bsy_2_27;
  wire        _GEN_2605 = _GEN_2573 ? ~_rob_bsy_T_4 : rob_bsy_2_28;
  wire        _GEN_2606 = _GEN_2574 ? ~_rob_bsy_T_4 : rob_bsy_2_29;
  wire        _GEN_2607 = _GEN_2575 ? ~_rob_bsy_T_4 : rob_bsy_2_30;
  wire        _GEN_2608 = _GEN_2576 ? ~_rob_bsy_T_4 : rob_bsy_2_31;
  wire        _rob_unsafe_T_14 = io_enq_uops_2_uses_ldq | io_enq_uops_2_uses_stq & ~io_enq_uops_2_is_fence | io_enq_uops_2_is_br | io_enq_uops_2_is_jalr;
  wire        _GEN_2609 = _GEN_2545 ? _rob_unsafe_T_14 : rob_unsafe_2_0;
  wire        _GEN_2610 = _GEN_2546 ? _rob_unsafe_T_14 : rob_unsafe_2_1;
  wire        _GEN_2611 = _GEN_2547 ? _rob_unsafe_T_14 : rob_unsafe_2_2;
  wire        _GEN_2612 = _GEN_2548 ? _rob_unsafe_T_14 : rob_unsafe_2_3;
  wire        _GEN_2613 = _GEN_2549 ? _rob_unsafe_T_14 : rob_unsafe_2_4;
  wire        _GEN_2614 = _GEN_2550 ? _rob_unsafe_T_14 : rob_unsafe_2_5;
  wire        _GEN_2615 = _GEN_2551 ? _rob_unsafe_T_14 : rob_unsafe_2_6;
  wire        _GEN_2616 = _GEN_2552 ? _rob_unsafe_T_14 : rob_unsafe_2_7;
  wire        _GEN_2617 = _GEN_2553 ? _rob_unsafe_T_14 : rob_unsafe_2_8;
  wire        _GEN_2618 = _GEN_2554 ? _rob_unsafe_T_14 : rob_unsafe_2_9;
  wire        _GEN_2619 = _GEN_2555 ? _rob_unsafe_T_14 : rob_unsafe_2_10;
  wire        _GEN_2620 = _GEN_2556 ? _rob_unsafe_T_14 : rob_unsafe_2_11;
  wire        _GEN_2621 = _GEN_2557 ? _rob_unsafe_T_14 : rob_unsafe_2_12;
  wire        _GEN_2622 = _GEN_2558 ? _rob_unsafe_T_14 : rob_unsafe_2_13;
  wire        _GEN_2623 = _GEN_2559 ? _rob_unsafe_T_14 : rob_unsafe_2_14;
  wire        _GEN_2624 = _GEN_2560 ? _rob_unsafe_T_14 : rob_unsafe_2_15;
  wire        _GEN_2625 = _GEN_2561 ? _rob_unsafe_T_14 : rob_unsafe_2_16;
  wire        _GEN_2626 = _GEN_2562 ? _rob_unsafe_T_14 : rob_unsafe_2_17;
  wire        _GEN_2627 = _GEN_2563 ? _rob_unsafe_T_14 : rob_unsafe_2_18;
  wire        _GEN_2628 = _GEN_2564 ? _rob_unsafe_T_14 : rob_unsafe_2_19;
  wire        _GEN_2629 = _GEN_2565 ? _rob_unsafe_T_14 : rob_unsafe_2_20;
  wire        _GEN_2630 = _GEN_2566 ? _rob_unsafe_T_14 : rob_unsafe_2_21;
  wire        _GEN_2631 = _GEN_2567 ? _rob_unsafe_T_14 : rob_unsafe_2_22;
  wire        _GEN_2632 = _GEN_2568 ? _rob_unsafe_T_14 : rob_unsafe_2_23;
  wire        _GEN_2633 = _GEN_2569 ? _rob_unsafe_T_14 : rob_unsafe_2_24;
  wire        _GEN_2634 = _GEN_2570 ? _rob_unsafe_T_14 : rob_unsafe_2_25;
  wire        _GEN_2635 = _GEN_2571 ? _rob_unsafe_T_14 : rob_unsafe_2_26;
  wire        _GEN_2636 = _GEN_2572 ? _rob_unsafe_T_14 : rob_unsafe_2_27;
  wire        _GEN_2637 = _GEN_2573 ? _rob_unsafe_T_14 : rob_unsafe_2_28;
  wire        _GEN_2638 = _GEN_2574 ? _rob_unsafe_T_14 : rob_unsafe_2_29;
  wire        _GEN_2639 = _GEN_2575 ? _rob_unsafe_T_14 : rob_unsafe_2_30;
  wire        _GEN_2640 = _GEN_2576 ? _rob_unsafe_T_14 : rob_unsafe_2_31;
  wire        _GEN_2641 = _GEN_33 & _GEN_254;
  wire        _GEN_2642 = _GEN_33 & _GEN_256;
  wire        _GEN_2643 = _GEN_33 & _GEN_258;
  wire        _GEN_2644 = _GEN_33 & _GEN_260;
  wire        _GEN_2645 = _GEN_33 & _GEN_262;
  wire        _GEN_2646 = _GEN_33 & _GEN_264;
  wire        _GEN_2647 = _GEN_33 & _GEN_266;
  wire        _GEN_2648 = _GEN_33 & _GEN_268;
  wire        _GEN_2649 = _GEN_33 & _GEN_270;
  wire        _GEN_2650 = _GEN_33 & _GEN_272;
  wire        _GEN_2651 = _GEN_33 & _GEN_274;
  wire        _GEN_2652 = _GEN_33 & _GEN_276;
  wire        _GEN_2653 = _GEN_33 & _GEN_278;
  wire        _GEN_2654 = _GEN_33 & _GEN_280;
  wire        _GEN_2655 = _GEN_33 & _GEN_282;
  wire        _GEN_2656 = _GEN_33 & _GEN_284;
  wire        _GEN_2657 = _GEN_33 & _GEN_286;
  wire        _GEN_2658 = _GEN_33 & _GEN_288;
  wire        _GEN_2659 = _GEN_33 & _GEN_290;
  wire        _GEN_2660 = _GEN_33 & _GEN_292;
  wire        _GEN_2661 = _GEN_33 & _GEN_294;
  wire        _GEN_2662 = _GEN_33 & _GEN_296;
  wire        _GEN_2663 = _GEN_33 & _GEN_298;
  wire        _GEN_2664 = _GEN_33 & _GEN_300;
  wire        _GEN_2665 = _GEN_33 & _GEN_302;
  wire        _GEN_2666 = _GEN_33 & _GEN_304;
  wire        _GEN_2667 = _GEN_33 & _GEN_306;
  wire        _GEN_2668 = _GEN_33 & _GEN_308;
  wire        _GEN_2669 = _GEN_33 & _GEN_310;
  wire        _GEN_2670 = _GEN_33 & _GEN_312;
  wire        _GEN_2671 = _GEN_33 & _GEN_314;
  wire        _GEN_2672 = _GEN_33 & (&(io_wb_resps_0_bits_uop_rob_idx[6:2]));
  wire        _GEN_2673 = _GEN_317 | _GEN_2641;
  wire        _GEN_2674 = _GEN_34 ? ~_GEN_2673 & _GEN_2577 : ~_GEN_2641 & _GEN_2577;
  wire        _GEN_2675 = _GEN_320 | _GEN_2642;
  wire        _GEN_2676 = _GEN_34 ? ~_GEN_2675 & _GEN_2578 : ~_GEN_2642 & _GEN_2578;
  wire        _GEN_2677 = _GEN_323 | _GEN_2643;
  wire        _GEN_2678 = _GEN_34 ? ~_GEN_2677 & _GEN_2579 : ~_GEN_2643 & _GEN_2579;
  wire        _GEN_2679 = _GEN_326 | _GEN_2644;
  wire        _GEN_2680 = _GEN_34 ? ~_GEN_2679 & _GEN_2580 : ~_GEN_2644 & _GEN_2580;
  wire        _GEN_2681 = _GEN_329 | _GEN_2645;
  wire        _GEN_2682 = _GEN_34 ? ~_GEN_2681 & _GEN_2581 : ~_GEN_2645 & _GEN_2581;
  wire        _GEN_2683 = _GEN_332 | _GEN_2646;
  wire        _GEN_2684 = _GEN_34 ? ~_GEN_2683 & _GEN_2582 : ~_GEN_2646 & _GEN_2582;
  wire        _GEN_2685 = _GEN_335 | _GEN_2647;
  wire        _GEN_2686 = _GEN_34 ? ~_GEN_2685 & _GEN_2583 : ~_GEN_2647 & _GEN_2583;
  wire        _GEN_2687 = _GEN_338 | _GEN_2648;
  wire        _GEN_2688 = _GEN_34 ? ~_GEN_2687 & _GEN_2584 : ~_GEN_2648 & _GEN_2584;
  wire        _GEN_2689 = _GEN_341 | _GEN_2649;
  wire        _GEN_2690 = _GEN_34 ? ~_GEN_2689 & _GEN_2585 : ~_GEN_2649 & _GEN_2585;
  wire        _GEN_2691 = _GEN_344 | _GEN_2650;
  wire        _GEN_2692 = _GEN_34 ? ~_GEN_2691 & _GEN_2586 : ~_GEN_2650 & _GEN_2586;
  wire        _GEN_2693 = _GEN_347 | _GEN_2651;
  wire        _GEN_2694 = _GEN_34 ? ~_GEN_2693 & _GEN_2587 : ~_GEN_2651 & _GEN_2587;
  wire        _GEN_2695 = _GEN_350 | _GEN_2652;
  wire        _GEN_2696 = _GEN_34 ? ~_GEN_2695 & _GEN_2588 : ~_GEN_2652 & _GEN_2588;
  wire        _GEN_2697 = _GEN_353 | _GEN_2653;
  wire        _GEN_2698 = _GEN_34 ? ~_GEN_2697 & _GEN_2589 : ~_GEN_2653 & _GEN_2589;
  wire        _GEN_2699 = _GEN_356 | _GEN_2654;
  wire        _GEN_2700 = _GEN_34 ? ~_GEN_2699 & _GEN_2590 : ~_GEN_2654 & _GEN_2590;
  wire        _GEN_2701 = _GEN_359 | _GEN_2655;
  wire        _GEN_2702 = _GEN_34 ? ~_GEN_2701 & _GEN_2591 : ~_GEN_2655 & _GEN_2591;
  wire        _GEN_2703 = _GEN_362 | _GEN_2656;
  wire        _GEN_2704 = _GEN_34 ? ~_GEN_2703 & _GEN_2592 : ~_GEN_2656 & _GEN_2592;
  wire        _GEN_2705 = _GEN_365 | _GEN_2657;
  wire        _GEN_2706 = _GEN_34 ? ~_GEN_2705 & _GEN_2593 : ~_GEN_2657 & _GEN_2593;
  wire        _GEN_2707 = _GEN_368 | _GEN_2658;
  wire        _GEN_2708 = _GEN_34 ? ~_GEN_2707 & _GEN_2594 : ~_GEN_2658 & _GEN_2594;
  wire        _GEN_2709 = _GEN_371 | _GEN_2659;
  wire        _GEN_2710 = _GEN_34 ? ~_GEN_2709 & _GEN_2595 : ~_GEN_2659 & _GEN_2595;
  wire        _GEN_2711 = _GEN_374 | _GEN_2660;
  wire        _GEN_2712 = _GEN_34 ? ~_GEN_2711 & _GEN_2596 : ~_GEN_2660 & _GEN_2596;
  wire        _GEN_2713 = _GEN_377 | _GEN_2661;
  wire        _GEN_2714 = _GEN_34 ? ~_GEN_2713 & _GEN_2597 : ~_GEN_2661 & _GEN_2597;
  wire        _GEN_2715 = _GEN_380 | _GEN_2662;
  wire        _GEN_2716 = _GEN_34 ? ~_GEN_2715 & _GEN_2598 : ~_GEN_2662 & _GEN_2598;
  wire        _GEN_2717 = _GEN_383 | _GEN_2663;
  wire        _GEN_2718 = _GEN_34 ? ~_GEN_2717 & _GEN_2599 : ~_GEN_2663 & _GEN_2599;
  wire        _GEN_2719 = _GEN_386 | _GEN_2664;
  wire        _GEN_2720 = _GEN_34 ? ~_GEN_2719 & _GEN_2600 : ~_GEN_2664 & _GEN_2600;
  wire        _GEN_2721 = _GEN_389 | _GEN_2665;
  wire        _GEN_2722 = _GEN_34 ? ~_GEN_2721 & _GEN_2601 : ~_GEN_2665 & _GEN_2601;
  wire        _GEN_2723 = _GEN_392 | _GEN_2666;
  wire        _GEN_2724 = _GEN_34 ? ~_GEN_2723 & _GEN_2602 : ~_GEN_2666 & _GEN_2602;
  wire        _GEN_2725 = _GEN_395 | _GEN_2667;
  wire        _GEN_2726 = _GEN_34 ? ~_GEN_2725 & _GEN_2603 : ~_GEN_2667 & _GEN_2603;
  wire        _GEN_2727 = _GEN_398 | _GEN_2668;
  wire        _GEN_2728 = _GEN_34 ? ~_GEN_2727 & _GEN_2604 : ~_GEN_2668 & _GEN_2604;
  wire        _GEN_2729 = _GEN_401 | _GEN_2669;
  wire        _GEN_2730 = _GEN_34 ? ~_GEN_2729 & _GEN_2605 : ~_GEN_2669 & _GEN_2605;
  wire        _GEN_2731 = _GEN_404 | _GEN_2670;
  wire        _GEN_2732 = _GEN_34 ? ~_GEN_2731 & _GEN_2606 : ~_GEN_2670 & _GEN_2606;
  wire        _GEN_2733 = _GEN_407 | _GEN_2671;
  wire        _GEN_2734 = _GEN_34 ? ~_GEN_2733 & _GEN_2607 : ~_GEN_2671 & _GEN_2607;
  wire        _GEN_2735 = (&(io_wb_resps_1_bits_uop_rob_idx[6:2])) | _GEN_2672;
  wire        _GEN_2736 = _GEN_34 ? ~_GEN_2735 & _GEN_2608 : ~_GEN_2672 & _GEN_2608;
  wire        _GEN_2737 = _GEN_34 ? ~_GEN_2673 & _GEN_2609 : ~_GEN_2641 & _GEN_2609;
  wire        _GEN_2738 = _GEN_34 ? ~_GEN_2675 & _GEN_2610 : ~_GEN_2642 & _GEN_2610;
  wire        _GEN_2739 = _GEN_34 ? ~_GEN_2677 & _GEN_2611 : ~_GEN_2643 & _GEN_2611;
  wire        _GEN_2740 = _GEN_34 ? ~_GEN_2679 & _GEN_2612 : ~_GEN_2644 & _GEN_2612;
  wire        _GEN_2741 = _GEN_34 ? ~_GEN_2681 & _GEN_2613 : ~_GEN_2645 & _GEN_2613;
  wire        _GEN_2742 = _GEN_34 ? ~_GEN_2683 & _GEN_2614 : ~_GEN_2646 & _GEN_2614;
  wire        _GEN_2743 = _GEN_34 ? ~_GEN_2685 & _GEN_2615 : ~_GEN_2647 & _GEN_2615;
  wire        _GEN_2744 = _GEN_34 ? ~_GEN_2687 & _GEN_2616 : ~_GEN_2648 & _GEN_2616;
  wire        _GEN_2745 = _GEN_34 ? ~_GEN_2689 & _GEN_2617 : ~_GEN_2649 & _GEN_2617;
  wire        _GEN_2746 = _GEN_34 ? ~_GEN_2691 & _GEN_2618 : ~_GEN_2650 & _GEN_2618;
  wire        _GEN_2747 = _GEN_34 ? ~_GEN_2693 & _GEN_2619 : ~_GEN_2651 & _GEN_2619;
  wire        _GEN_2748 = _GEN_34 ? ~_GEN_2695 & _GEN_2620 : ~_GEN_2652 & _GEN_2620;
  wire        _GEN_2749 = _GEN_34 ? ~_GEN_2697 & _GEN_2621 : ~_GEN_2653 & _GEN_2621;
  wire        _GEN_2750 = _GEN_34 ? ~_GEN_2699 & _GEN_2622 : ~_GEN_2654 & _GEN_2622;
  wire        _GEN_2751 = _GEN_34 ? ~_GEN_2701 & _GEN_2623 : ~_GEN_2655 & _GEN_2623;
  wire        _GEN_2752 = _GEN_34 ? ~_GEN_2703 & _GEN_2624 : ~_GEN_2656 & _GEN_2624;
  wire        _GEN_2753 = _GEN_34 ? ~_GEN_2705 & _GEN_2625 : ~_GEN_2657 & _GEN_2625;
  wire        _GEN_2754 = _GEN_34 ? ~_GEN_2707 & _GEN_2626 : ~_GEN_2658 & _GEN_2626;
  wire        _GEN_2755 = _GEN_34 ? ~_GEN_2709 & _GEN_2627 : ~_GEN_2659 & _GEN_2627;
  wire        _GEN_2756 = _GEN_34 ? ~_GEN_2711 & _GEN_2628 : ~_GEN_2660 & _GEN_2628;
  wire        _GEN_2757 = _GEN_34 ? ~_GEN_2713 & _GEN_2629 : ~_GEN_2661 & _GEN_2629;
  wire        _GEN_2758 = _GEN_34 ? ~_GEN_2715 & _GEN_2630 : ~_GEN_2662 & _GEN_2630;
  wire        _GEN_2759 = _GEN_34 ? ~_GEN_2717 & _GEN_2631 : ~_GEN_2663 & _GEN_2631;
  wire        _GEN_2760 = _GEN_34 ? ~_GEN_2719 & _GEN_2632 : ~_GEN_2664 & _GEN_2632;
  wire        _GEN_2761 = _GEN_34 ? ~_GEN_2721 & _GEN_2633 : ~_GEN_2665 & _GEN_2633;
  wire        _GEN_2762 = _GEN_34 ? ~_GEN_2723 & _GEN_2634 : ~_GEN_2666 & _GEN_2634;
  wire        _GEN_2763 = _GEN_34 ? ~_GEN_2725 & _GEN_2635 : ~_GEN_2667 & _GEN_2635;
  wire        _GEN_2764 = _GEN_34 ? ~_GEN_2727 & _GEN_2636 : ~_GEN_2668 & _GEN_2636;
  wire        _GEN_2765 = _GEN_34 ? ~_GEN_2729 & _GEN_2637 : ~_GEN_2669 & _GEN_2637;
  wire        _GEN_2766 = _GEN_34 ? ~_GEN_2731 & _GEN_2638 : ~_GEN_2670 & _GEN_2638;
  wire        _GEN_2767 = _GEN_34 ? ~_GEN_2733 & _GEN_2639 : ~_GEN_2671 & _GEN_2639;
  wire        _GEN_2768 = _GEN_34 ? ~_GEN_2735 & _GEN_2640 : ~_GEN_2672 & _GEN_2640;
  wire        _GEN_2769 = _GEN_35 & _GEN_444;
  wire        _GEN_2770 = _GEN_35 & _GEN_446;
  wire        _GEN_2771 = _GEN_35 & _GEN_448;
  wire        _GEN_2772 = _GEN_35 & _GEN_450;
  wire        _GEN_2773 = _GEN_35 & _GEN_452;
  wire        _GEN_2774 = _GEN_35 & _GEN_454;
  wire        _GEN_2775 = _GEN_35 & _GEN_456;
  wire        _GEN_2776 = _GEN_35 & _GEN_458;
  wire        _GEN_2777 = _GEN_35 & _GEN_460;
  wire        _GEN_2778 = _GEN_35 & _GEN_462;
  wire        _GEN_2779 = _GEN_35 & _GEN_464;
  wire        _GEN_2780 = _GEN_35 & _GEN_466;
  wire        _GEN_2781 = _GEN_35 & _GEN_468;
  wire        _GEN_2782 = _GEN_35 & _GEN_470;
  wire        _GEN_2783 = _GEN_35 & _GEN_472;
  wire        _GEN_2784 = _GEN_35 & _GEN_474;
  wire        _GEN_2785 = _GEN_35 & _GEN_476;
  wire        _GEN_2786 = _GEN_35 & _GEN_478;
  wire        _GEN_2787 = _GEN_35 & _GEN_480;
  wire        _GEN_2788 = _GEN_35 & _GEN_482;
  wire        _GEN_2789 = _GEN_35 & _GEN_484;
  wire        _GEN_2790 = _GEN_35 & _GEN_486;
  wire        _GEN_2791 = _GEN_35 & _GEN_488;
  wire        _GEN_2792 = _GEN_35 & _GEN_490;
  wire        _GEN_2793 = _GEN_35 & _GEN_492;
  wire        _GEN_2794 = _GEN_35 & _GEN_494;
  wire        _GEN_2795 = _GEN_35 & _GEN_496;
  wire        _GEN_2796 = _GEN_35 & _GEN_498;
  wire        _GEN_2797 = _GEN_35 & _GEN_500;
  wire        _GEN_2798 = _GEN_35 & _GEN_502;
  wire        _GEN_2799 = _GEN_35 & _GEN_504;
  wire        _GEN_2800 = _GEN_35 & (&(io_wb_resps_2_bits_uop_rob_idx[6:2]));
  wire        _GEN_2801 = _GEN_507 | _GEN_2769;
  wire        _GEN_2802 = _GEN_36 ? ~_GEN_2801 & _GEN_2674 : ~_GEN_2769 & _GEN_2674;
  wire        _GEN_2803 = _GEN_510 | _GEN_2770;
  wire        _GEN_2804 = _GEN_36 ? ~_GEN_2803 & _GEN_2676 : ~_GEN_2770 & _GEN_2676;
  wire        _GEN_2805 = _GEN_513 | _GEN_2771;
  wire        _GEN_2806 = _GEN_36 ? ~_GEN_2805 & _GEN_2678 : ~_GEN_2771 & _GEN_2678;
  wire        _GEN_2807 = _GEN_516 | _GEN_2772;
  wire        _GEN_2808 = _GEN_36 ? ~_GEN_2807 & _GEN_2680 : ~_GEN_2772 & _GEN_2680;
  wire        _GEN_2809 = _GEN_519 | _GEN_2773;
  wire        _GEN_2810 = _GEN_36 ? ~_GEN_2809 & _GEN_2682 : ~_GEN_2773 & _GEN_2682;
  wire        _GEN_2811 = _GEN_522 | _GEN_2774;
  wire        _GEN_2812 = _GEN_36 ? ~_GEN_2811 & _GEN_2684 : ~_GEN_2774 & _GEN_2684;
  wire        _GEN_2813 = _GEN_525 | _GEN_2775;
  wire        _GEN_2814 = _GEN_36 ? ~_GEN_2813 & _GEN_2686 : ~_GEN_2775 & _GEN_2686;
  wire        _GEN_2815 = _GEN_528 | _GEN_2776;
  wire        _GEN_2816 = _GEN_36 ? ~_GEN_2815 & _GEN_2688 : ~_GEN_2776 & _GEN_2688;
  wire        _GEN_2817 = _GEN_531 | _GEN_2777;
  wire        _GEN_2818 = _GEN_36 ? ~_GEN_2817 & _GEN_2690 : ~_GEN_2777 & _GEN_2690;
  wire        _GEN_2819 = _GEN_534 | _GEN_2778;
  wire        _GEN_2820 = _GEN_36 ? ~_GEN_2819 & _GEN_2692 : ~_GEN_2778 & _GEN_2692;
  wire        _GEN_2821 = _GEN_537 | _GEN_2779;
  wire        _GEN_2822 = _GEN_36 ? ~_GEN_2821 & _GEN_2694 : ~_GEN_2779 & _GEN_2694;
  wire        _GEN_2823 = _GEN_540 | _GEN_2780;
  wire        _GEN_2824 = _GEN_36 ? ~_GEN_2823 & _GEN_2696 : ~_GEN_2780 & _GEN_2696;
  wire        _GEN_2825 = _GEN_543 | _GEN_2781;
  wire        _GEN_2826 = _GEN_36 ? ~_GEN_2825 & _GEN_2698 : ~_GEN_2781 & _GEN_2698;
  wire        _GEN_2827 = _GEN_546 | _GEN_2782;
  wire        _GEN_2828 = _GEN_36 ? ~_GEN_2827 & _GEN_2700 : ~_GEN_2782 & _GEN_2700;
  wire        _GEN_2829 = _GEN_549 | _GEN_2783;
  wire        _GEN_2830 = _GEN_36 ? ~_GEN_2829 & _GEN_2702 : ~_GEN_2783 & _GEN_2702;
  wire        _GEN_2831 = _GEN_552 | _GEN_2784;
  wire        _GEN_2832 = _GEN_36 ? ~_GEN_2831 & _GEN_2704 : ~_GEN_2784 & _GEN_2704;
  wire        _GEN_2833 = _GEN_555 | _GEN_2785;
  wire        _GEN_2834 = _GEN_36 ? ~_GEN_2833 & _GEN_2706 : ~_GEN_2785 & _GEN_2706;
  wire        _GEN_2835 = _GEN_558 | _GEN_2786;
  wire        _GEN_2836 = _GEN_36 ? ~_GEN_2835 & _GEN_2708 : ~_GEN_2786 & _GEN_2708;
  wire        _GEN_2837 = _GEN_561 | _GEN_2787;
  wire        _GEN_2838 = _GEN_36 ? ~_GEN_2837 & _GEN_2710 : ~_GEN_2787 & _GEN_2710;
  wire        _GEN_2839 = _GEN_564 | _GEN_2788;
  wire        _GEN_2840 = _GEN_36 ? ~_GEN_2839 & _GEN_2712 : ~_GEN_2788 & _GEN_2712;
  wire        _GEN_2841 = _GEN_567 | _GEN_2789;
  wire        _GEN_2842 = _GEN_36 ? ~_GEN_2841 & _GEN_2714 : ~_GEN_2789 & _GEN_2714;
  wire        _GEN_2843 = _GEN_570 | _GEN_2790;
  wire        _GEN_2844 = _GEN_36 ? ~_GEN_2843 & _GEN_2716 : ~_GEN_2790 & _GEN_2716;
  wire        _GEN_2845 = _GEN_573 | _GEN_2791;
  wire        _GEN_2846 = _GEN_36 ? ~_GEN_2845 & _GEN_2718 : ~_GEN_2791 & _GEN_2718;
  wire        _GEN_2847 = _GEN_576 | _GEN_2792;
  wire        _GEN_2848 = _GEN_36 ? ~_GEN_2847 & _GEN_2720 : ~_GEN_2792 & _GEN_2720;
  wire        _GEN_2849 = _GEN_579 | _GEN_2793;
  wire        _GEN_2850 = _GEN_36 ? ~_GEN_2849 & _GEN_2722 : ~_GEN_2793 & _GEN_2722;
  wire        _GEN_2851 = _GEN_582 | _GEN_2794;
  wire        _GEN_2852 = _GEN_36 ? ~_GEN_2851 & _GEN_2724 : ~_GEN_2794 & _GEN_2724;
  wire        _GEN_2853 = _GEN_585 | _GEN_2795;
  wire        _GEN_2854 = _GEN_36 ? ~_GEN_2853 & _GEN_2726 : ~_GEN_2795 & _GEN_2726;
  wire        _GEN_2855 = _GEN_588 | _GEN_2796;
  wire        _GEN_2856 = _GEN_36 ? ~_GEN_2855 & _GEN_2728 : ~_GEN_2796 & _GEN_2728;
  wire        _GEN_2857 = _GEN_591 | _GEN_2797;
  wire        _GEN_2858 = _GEN_36 ? ~_GEN_2857 & _GEN_2730 : ~_GEN_2797 & _GEN_2730;
  wire        _GEN_2859 = _GEN_594 | _GEN_2798;
  wire        _GEN_2860 = _GEN_36 ? ~_GEN_2859 & _GEN_2732 : ~_GEN_2798 & _GEN_2732;
  wire        _GEN_2861 = _GEN_597 | _GEN_2799;
  wire        _GEN_2862 = _GEN_36 ? ~_GEN_2861 & _GEN_2734 : ~_GEN_2799 & _GEN_2734;
  wire        _GEN_2863 = (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_2800;
  wire        _GEN_2864 = _GEN_36 ? ~_GEN_2863 & _GEN_2736 : ~_GEN_2800 & _GEN_2736;
  wire        _GEN_2865 = _GEN_36 ? ~_GEN_2801 & _GEN_2737 : ~_GEN_2769 & _GEN_2737;
  wire        _GEN_2866 = _GEN_36 ? ~_GEN_2803 & _GEN_2738 : ~_GEN_2770 & _GEN_2738;
  wire        _GEN_2867 = _GEN_36 ? ~_GEN_2805 & _GEN_2739 : ~_GEN_2771 & _GEN_2739;
  wire        _GEN_2868 = _GEN_36 ? ~_GEN_2807 & _GEN_2740 : ~_GEN_2772 & _GEN_2740;
  wire        _GEN_2869 = _GEN_36 ? ~_GEN_2809 & _GEN_2741 : ~_GEN_2773 & _GEN_2741;
  wire        _GEN_2870 = _GEN_36 ? ~_GEN_2811 & _GEN_2742 : ~_GEN_2774 & _GEN_2742;
  wire        _GEN_2871 = _GEN_36 ? ~_GEN_2813 & _GEN_2743 : ~_GEN_2775 & _GEN_2743;
  wire        _GEN_2872 = _GEN_36 ? ~_GEN_2815 & _GEN_2744 : ~_GEN_2776 & _GEN_2744;
  wire        _GEN_2873 = _GEN_36 ? ~_GEN_2817 & _GEN_2745 : ~_GEN_2777 & _GEN_2745;
  wire        _GEN_2874 = _GEN_36 ? ~_GEN_2819 & _GEN_2746 : ~_GEN_2778 & _GEN_2746;
  wire        _GEN_2875 = _GEN_36 ? ~_GEN_2821 & _GEN_2747 : ~_GEN_2779 & _GEN_2747;
  wire        _GEN_2876 = _GEN_36 ? ~_GEN_2823 & _GEN_2748 : ~_GEN_2780 & _GEN_2748;
  wire        _GEN_2877 = _GEN_36 ? ~_GEN_2825 & _GEN_2749 : ~_GEN_2781 & _GEN_2749;
  wire        _GEN_2878 = _GEN_36 ? ~_GEN_2827 & _GEN_2750 : ~_GEN_2782 & _GEN_2750;
  wire        _GEN_2879 = _GEN_36 ? ~_GEN_2829 & _GEN_2751 : ~_GEN_2783 & _GEN_2751;
  wire        _GEN_2880 = _GEN_36 ? ~_GEN_2831 & _GEN_2752 : ~_GEN_2784 & _GEN_2752;
  wire        _GEN_2881 = _GEN_36 ? ~_GEN_2833 & _GEN_2753 : ~_GEN_2785 & _GEN_2753;
  wire        _GEN_2882 = _GEN_36 ? ~_GEN_2835 & _GEN_2754 : ~_GEN_2786 & _GEN_2754;
  wire        _GEN_2883 = _GEN_36 ? ~_GEN_2837 & _GEN_2755 : ~_GEN_2787 & _GEN_2755;
  wire        _GEN_2884 = _GEN_36 ? ~_GEN_2839 & _GEN_2756 : ~_GEN_2788 & _GEN_2756;
  wire        _GEN_2885 = _GEN_36 ? ~_GEN_2841 & _GEN_2757 : ~_GEN_2789 & _GEN_2757;
  wire        _GEN_2886 = _GEN_36 ? ~_GEN_2843 & _GEN_2758 : ~_GEN_2790 & _GEN_2758;
  wire        _GEN_2887 = _GEN_36 ? ~_GEN_2845 & _GEN_2759 : ~_GEN_2791 & _GEN_2759;
  wire        _GEN_2888 = _GEN_36 ? ~_GEN_2847 & _GEN_2760 : ~_GEN_2792 & _GEN_2760;
  wire        _GEN_2889 = _GEN_36 ? ~_GEN_2849 & _GEN_2761 : ~_GEN_2793 & _GEN_2761;
  wire        _GEN_2890 = _GEN_36 ? ~_GEN_2851 & _GEN_2762 : ~_GEN_2794 & _GEN_2762;
  wire        _GEN_2891 = _GEN_36 ? ~_GEN_2853 & _GEN_2763 : ~_GEN_2795 & _GEN_2763;
  wire        _GEN_2892 = _GEN_36 ? ~_GEN_2855 & _GEN_2764 : ~_GEN_2796 & _GEN_2764;
  wire        _GEN_2893 = _GEN_36 ? ~_GEN_2857 & _GEN_2765 : ~_GEN_2797 & _GEN_2765;
  wire        _GEN_2894 = _GEN_36 ? ~_GEN_2859 & _GEN_2766 : ~_GEN_2798 & _GEN_2766;
  wire        _GEN_2895 = _GEN_36 ? ~_GEN_2861 & _GEN_2767 : ~_GEN_2799 & _GEN_2767;
  wire        _GEN_2896 = _GEN_36 ? ~_GEN_2863 & _GEN_2768 : ~_GEN_2800 & _GEN_2768;
  wire        _GEN_2897 = _GEN_37 & _GEN_634;
  wire        _GEN_2898 = _GEN_37 & _GEN_636;
  wire        _GEN_2899 = _GEN_37 & _GEN_638;
  wire        _GEN_2900 = _GEN_37 & _GEN_640;
  wire        _GEN_2901 = _GEN_37 & _GEN_642;
  wire        _GEN_2902 = _GEN_37 & _GEN_644;
  wire        _GEN_2903 = _GEN_37 & _GEN_646;
  wire        _GEN_2904 = _GEN_37 & _GEN_648;
  wire        _GEN_2905 = _GEN_37 & _GEN_650;
  wire        _GEN_2906 = _GEN_37 & _GEN_652;
  wire        _GEN_2907 = _GEN_37 & _GEN_654;
  wire        _GEN_2908 = _GEN_37 & _GEN_656;
  wire        _GEN_2909 = _GEN_37 & _GEN_658;
  wire        _GEN_2910 = _GEN_37 & _GEN_660;
  wire        _GEN_2911 = _GEN_37 & _GEN_662;
  wire        _GEN_2912 = _GEN_37 & _GEN_664;
  wire        _GEN_2913 = _GEN_37 & _GEN_666;
  wire        _GEN_2914 = _GEN_37 & _GEN_668;
  wire        _GEN_2915 = _GEN_37 & _GEN_670;
  wire        _GEN_2916 = _GEN_37 & _GEN_672;
  wire        _GEN_2917 = _GEN_37 & _GEN_674;
  wire        _GEN_2918 = _GEN_37 & _GEN_676;
  wire        _GEN_2919 = _GEN_37 & _GEN_678;
  wire        _GEN_2920 = _GEN_37 & _GEN_680;
  wire        _GEN_2921 = _GEN_37 & _GEN_682;
  wire        _GEN_2922 = _GEN_37 & _GEN_684;
  wire        _GEN_2923 = _GEN_37 & _GEN_686;
  wire        _GEN_2924 = _GEN_37 & _GEN_688;
  wire        _GEN_2925 = _GEN_37 & _GEN_690;
  wire        _GEN_2926 = _GEN_37 & _GEN_692;
  wire        _GEN_2927 = _GEN_37 & _GEN_694;
  wire        _GEN_2928 = _GEN_37 & (&(io_wb_resps_4_bits_uop_rob_idx[6:2]));
  wire        _GEN_2929 = _GEN_697 | _GEN_2897;
  wire        _GEN_2930 = _GEN_38 ? ~_GEN_2929 & _GEN_2802 : ~_GEN_2897 & _GEN_2802;
  wire        _GEN_2931 = _GEN_700 | _GEN_2898;
  wire        _GEN_2932 = _GEN_38 ? ~_GEN_2931 & _GEN_2804 : ~_GEN_2898 & _GEN_2804;
  wire        _GEN_2933 = _GEN_703 | _GEN_2899;
  wire        _GEN_2934 = _GEN_38 ? ~_GEN_2933 & _GEN_2806 : ~_GEN_2899 & _GEN_2806;
  wire        _GEN_2935 = _GEN_706 | _GEN_2900;
  wire        _GEN_2936 = _GEN_38 ? ~_GEN_2935 & _GEN_2808 : ~_GEN_2900 & _GEN_2808;
  wire        _GEN_2937 = _GEN_709 | _GEN_2901;
  wire        _GEN_2938 = _GEN_38 ? ~_GEN_2937 & _GEN_2810 : ~_GEN_2901 & _GEN_2810;
  wire        _GEN_2939 = _GEN_712 | _GEN_2902;
  wire        _GEN_2940 = _GEN_38 ? ~_GEN_2939 & _GEN_2812 : ~_GEN_2902 & _GEN_2812;
  wire        _GEN_2941 = _GEN_715 | _GEN_2903;
  wire        _GEN_2942 = _GEN_38 ? ~_GEN_2941 & _GEN_2814 : ~_GEN_2903 & _GEN_2814;
  wire        _GEN_2943 = _GEN_718 | _GEN_2904;
  wire        _GEN_2944 = _GEN_38 ? ~_GEN_2943 & _GEN_2816 : ~_GEN_2904 & _GEN_2816;
  wire        _GEN_2945 = _GEN_721 | _GEN_2905;
  wire        _GEN_2946 = _GEN_38 ? ~_GEN_2945 & _GEN_2818 : ~_GEN_2905 & _GEN_2818;
  wire        _GEN_2947 = _GEN_724 | _GEN_2906;
  wire        _GEN_2948 = _GEN_38 ? ~_GEN_2947 & _GEN_2820 : ~_GEN_2906 & _GEN_2820;
  wire        _GEN_2949 = _GEN_727 | _GEN_2907;
  wire        _GEN_2950 = _GEN_38 ? ~_GEN_2949 & _GEN_2822 : ~_GEN_2907 & _GEN_2822;
  wire        _GEN_2951 = _GEN_730 | _GEN_2908;
  wire        _GEN_2952 = _GEN_38 ? ~_GEN_2951 & _GEN_2824 : ~_GEN_2908 & _GEN_2824;
  wire        _GEN_2953 = _GEN_733 | _GEN_2909;
  wire        _GEN_2954 = _GEN_38 ? ~_GEN_2953 & _GEN_2826 : ~_GEN_2909 & _GEN_2826;
  wire        _GEN_2955 = _GEN_736 | _GEN_2910;
  wire        _GEN_2956 = _GEN_38 ? ~_GEN_2955 & _GEN_2828 : ~_GEN_2910 & _GEN_2828;
  wire        _GEN_2957 = _GEN_739 | _GEN_2911;
  wire        _GEN_2958 = _GEN_38 ? ~_GEN_2957 & _GEN_2830 : ~_GEN_2911 & _GEN_2830;
  wire        _GEN_2959 = _GEN_742 | _GEN_2912;
  wire        _GEN_2960 = _GEN_38 ? ~_GEN_2959 & _GEN_2832 : ~_GEN_2912 & _GEN_2832;
  wire        _GEN_2961 = _GEN_745 | _GEN_2913;
  wire        _GEN_2962 = _GEN_38 ? ~_GEN_2961 & _GEN_2834 : ~_GEN_2913 & _GEN_2834;
  wire        _GEN_2963 = _GEN_748 | _GEN_2914;
  wire        _GEN_2964 = _GEN_38 ? ~_GEN_2963 & _GEN_2836 : ~_GEN_2914 & _GEN_2836;
  wire        _GEN_2965 = _GEN_751 | _GEN_2915;
  wire        _GEN_2966 = _GEN_38 ? ~_GEN_2965 & _GEN_2838 : ~_GEN_2915 & _GEN_2838;
  wire        _GEN_2967 = _GEN_754 | _GEN_2916;
  wire        _GEN_2968 = _GEN_38 ? ~_GEN_2967 & _GEN_2840 : ~_GEN_2916 & _GEN_2840;
  wire        _GEN_2969 = _GEN_757 | _GEN_2917;
  wire        _GEN_2970 = _GEN_38 ? ~_GEN_2969 & _GEN_2842 : ~_GEN_2917 & _GEN_2842;
  wire        _GEN_2971 = _GEN_760 | _GEN_2918;
  wire        _GEN_2972 = _GEN_38 ? ~_GEN_2971 & _GEN_2844 : ~_GEN_2918 & _GEN_2844;
  wire        _GEN_2973 = _GEN_763 | _GEN_2919;
  wire        _GEN_2974 = _GEN_38 ? ~_GEN_2973 & _GEN_2846 : ~_GEN_2919 & _GEN_2846;
  wire        _GEN_2975 = _GEN_766 | _GEN_2920;
  wire        _GEN_2976 = _GEN_38 ? ~_GEN_2975 & _GEN_2848 : ~_GEN_2920 & _GEN_2848;
  wire        _GEN_2977 = _GEN_769 | _GEN_2921;
  wire        _GEN_2978 = _GEN_38 ? ~_GEN_2977 & _GEN_2850 : ~_GEN_2921 & _GEN_2850;
  wire        _GEN_2979 = _GEN_772 | _GEN_2922;
  wire        _GEN_2980 = _GEN_38 ? ~_GEN_2979 & _GEN_2852 : ~_GEN_2922 & _GEN_2852;
  wire        _GEN_2981 = _GEN_775 | _GEN_2923;
  wire        _GEN_2982 = _GEN_38 ? ~_GEN_2981 & _GEN_2854 : ~_GEN_2923 & _GEN_2854;
  wire        _GEN_2983 = _GEN_778 | _GEN_2924;
  wire        _GEN_2984 = _GEN_38 ? ~_GEN_2983 & _GEN_2856 : ~_GEN_2924 & _GEN_2856;
  wire        _GEN_2985 = _GEN_781 | _GEN_2925;
  wire        _GEN_2986 = _GEN_38 ? ~_GEN_2985 & _GEN_2858 : ~_GEN_2925 & _GEN_2858;
  wire        _GEN_2987 = _GEN_784 | _GEN_2926;
  wire        _GEN_2988 = _GEN_38 ? ~_GEN_2987 & _GEN_2860 : ~_GEN_2926 & _GEN_2860;
  wire        _GEN_2989 = _GEN_787 | _GEN_2927;
  wire        _GEN_2990 = _GEN_38 ? ~_GEN_2989 & _GEN_2862 : ~_GEN_2927 & _GEN_2862;
  wire        _GEN_2991 = (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_2928;
  wire        _GEN_2992 = _GEN_38 ? ~_GEN_2991 & _GEN_2864 : ~_GEN_2928 & _GEN_2864;
  wire        _GEN_2993 = _GEN_38 ? ~_GEN_2929 & _GEN_2865 : ~_GEN_2897 & _GEN_2865;
  wire        _GEN_2994 = _GEN_38 ? ~_GEN_2931 & _GEN_2866 : ~_GEN_2898 & _GEN_2866;
  wire        _GEN_2995 = _GEN_38 ? ~_GEN_2933 & _GEN_2867 : ~_GEN_2899 & _GEN_2867;
  wire        _GEN_2996 = _GEN_38 ? ~_GEN_2935 & _GEN_2868 : ~_GEN_2900 & _GEN_2868;
  wire        _GEN_2997 = _GEN_38 ? ~_GEN_2937 & _GEN_2869 : ~_GEN_2901 & _GEN_2869;
  wire        _GEN_2998 = _GEN_38 ? ~_GEN_2939 & _GEN_2870 : ~_GEN_2902 & _GEN_2870;
  wire        _GEN_2999 = _GEN_38 ? ~_GEN_2941 & _GEN_2871 : ~_GEN_2903 & _GEN_2871;
  wire        _GEN_3000 = _GEN_38 ? ~_GEN_2943 & _GEN_2872 : ~_GEN_2904 & _GEN_2872;
  wire        _GEN_3001 = _GEN_38 ? ~_GEN_2945 & _GEN_2873 : ~_GEN_2905 & _GEN_2873;
  wire        _GEN_3002 = _GEN_38 ? ~_GEN_2947 & _GEN_2874 : ~_GEN_2906 & _GEN_2874;
  wire        _GEN_3003 = _GEN_38 ? ~_GEN_2949 & _GEN_2875 : ~_GEN_2907 & _GEN_2875;
  wire        _GEN_3004 = _GEN_38 ? ~_GEN_2951 & _GEN_2876 : ~_GEN_2908 & _GEN_2876;
  wire        _GEN_3005 = _GEN_38 ? ~_GEN_2953 & _GEN_2877 : ~_GEN_2909 & _GEN_2877;
  wire        _GEN_3006 = _GEN_38 ? ~_GEN_2955 & _GEN_2878 : ~_GEN_2910 & _GEN_2878;
  wire        _GEN_3007 = _GEN_38 ? ~_GEN_2957 & _GEN_2879 : ~_GEN_2911 & _GEN_2879;
  wire        _GEN_3008 = _GEN_38 ? ~_GEN_2959 & _GEN_2880 : ~_GEN_2912 & _GEN_2880;
  wire        _GEN_3009 = _GEN_38 ? ~_GEN_2961 & _GEN_2881 : ~_GEN_2913 & _GEN_2881;
  wire        _GEN_3010 = _GEN_38 ? ~_GEN_2963 & _GEN_2882 : ~_GEN_2914 & _GEN_2882;
  wire        _GEN_3011 = _GEN_38 ? ~_GEN_2965 & _GEN_2883 : ~_GEN_2915 & _GEN_2883;
  wire        _GEN_3012 = _GEN_38 ? ~_GEN_2967 & _GEN_2884 : ~_GEN_2916 & _GEN_2884;
  wire        _GEN_3013 = _GEN_38 ? ~_GEN_2969 & _GEN_2885 : ~_GEN_2917 & _GEN_2885;
  wire        _GEN_3014 = _GEN_38 ? ~_GEN_2971 & _GEN_2886 : ~_GEN_2918 & _GEN_2886;
  wire        _GEN_3015 = _GEN_38 ? ~_GEN_2973 & _GEN_2887 : ~_GEN_2919 & _GEN_2887;
  wire        _GEN_3016 = _GEN_38 ? ~_GEN_2975 & _GEN_2888 : ~_GEN_2920 & _GEN_2888;
  wire        _GEN_3017 = _GEN_38 ? ~_GEN_2977 & _GEN_2889 : ~_GEN_2921 & _GEN_2889;
  wire        _GEN_3018 = _GEN_38 ? ~_GEN_2979 & _GEN_2890 : ~_GEN_2922 & _GEN_2890;
  wire        _GEN_3019 = _GEN_38 ? ~_GEN_2981 & _GEN_2891 : ~_GEN_2923 & _GEN_2891;
  wire        _GEN_3020 = _GEN_38 ? ~_GEN_2983 & _GEN_2892 : ~_GEN_2924 & _GEN_2892;
  wire        _GEN_3021 = _GEN_38 ? ~_GEN_2985 & _GEN_2893 : ~_GEN_2925 & _GEN_2893;
  wire        _GEN_3022 = _GEN_38 ? ~_GEN_2987 & _GEN_2894 : ~_GEN_2926 & _GEN_2894;
  wire        _GEN_3023 = _GEN_38 ? ~_GEN_2989 & _GEN_2895 : ~_GEN_2927 & _GEN_2895;
  wire        _GEN_3024 = _GEN_38 ? ~_GEN_2991 & _GEN_2896 : ~_GEN_2928 & _GEN_2896;
  wire        _GEN_3025 = _GEN_39 & _GEN_824;
  wire        _GEN_3026 = _GEN_39 & _GEN_826;
  wire        _GEN_3027 = _GEN_39 & _GEN_828;
  wire        _GEN_3028 = _GEN_39 & _GEN_830;
  wire        _GEN_3029 = _GEN_39 & _GEN_832;
  wire        _GEN_3030 = _GEN_39 & _GEN_834;
  wire        _GEN_3031 = _GEN_39 & _GEN_836;
  wire        _GEN_3032 = _GEN_39 & _GEN_838;
  wire        _GEN_3033 = _GEN_39 & _GEN_840;
  wire        _GEN_3034 = _GEN_39 & _GEN_842;
  wire        _GEN_3035 = _GEN_39 & _GEN_844;
  wire        _GEN_3036 = _GEN_39 & _GEN_846;
  wire        _GEN_3037 = _GEN_39 & _GEN_848;
  wire        _GEN_3038 = _GEN_39 & _GEN_850;
  wire        _GEN_3039 = _GEN_39 & _GEN_852;
  wire        _GEN_3040 = _GEN_39 & _GEN_854;
  wire        _GEN_3041 = _GEN_39 & _GEN_856;
  wire        _GEN_3042 = _GEN_39 & _GEN_858;
  wire        _GEN_3043 = _GEN_39 & _GEN_860;
  wire        _GEN_3044 = _GEN_39 & _GEN_862;
  wire        _GEN_3045 = _GEN_39 & _GEN_864;
  wire        _GEN_3046 = _GEN_39 & _GEN_866;
  wire        _GEN_3047 = _GEN_39 & _GEN_868;
  wire        _GEN_3048 = _GEN_39 & _GEN_870;
  wire        _GEN_3049 = _GEN_39 & _GEN_872;
  wire        _GEN_3050 = _GEN_39 & _GEN_874;
  wire        _GEN_3051 = _GEN_39 & _GEN_876;
  wire        _GEN_3052 = _GEN_39 & _GEN_878;
  wire        _GEN_3053 = _GEN_39 & _GEN_880;
  wire        _GEN_3054 = _GEN_39 & _GEN_882;
  wire        _GEN_3055 = _GEN_39 & _GEN_884;
  wire        _GEN_3056 = _GEN_39 & (&(io_wb_resps_6_bits_uop_rob_idx[6:2]));
  wire        _GEN_3057 = _GEN_887 | _GEN_3025;
  wire        _GEN_3058 = _GEN_40 ? ~_GEN_3057 & _GEN_2930 : ~_GEN_3025 & _GEN_2930;
  wire        _GEN_3059 = _GEN_890 | _GEN_3026;
  wire        _GEN_3060 = _GEN_40 ? ~_GEN_3059 & _GEN_2932 : ~_GEN_3026 & _GEN_2932;
  wire        _GEN_3061 = _GEN_893 | _GEN_3027;
  wire        _GEN_3062 = _GEN_40 ? ~_GEN_3061 & _GEN_2934 : ~_GEN_3027 & _GEN_2934;
  wire        _GEN_3063 = _GEN_896 | _GEN_3028;
  wire        _GEN_3064 = _GEN_40 ? ~_GEN_3063 & _GEN_2936 : ~_GEN_3028 & _GEN_2936;
  wire        _GEN_3065 = _GEN_899 | _GEN_3029;
  wire        _GEN_3066 = _GEN_40 ? ~_GEN_3065 & _GEN_2938 : ~_GEN_3029 & _GEN_2938;
  wire        _GEN_3067 = _GEN_902 | _GEN_3030;
  wire        _GEN_3068 = _GEN_40 ? ~_GEN_3067 & _GEN_2940 : ~_GEN_3030 & _GEN_2940;
  wire        _GEN_3069 = _GEN_905 | _GEN_3031;
  wire        _GEN_3070 = _GEN_40 ? ~_GEN_3069 & _GEN_2942 : ~_GEN_3031 & _GEN_2942;
  wire        _GEN_3071 = _GEN_908 | _GEN_3032;
  wire        _GEN_3072 = _GEN_40 ? ~_GEN_3071 & _GEN_2944 : ~_GEN_3032 & _GEN_2944;
  wire        _GEN_3073 = _GEN_911 | _GEN_3033;
  wire        _GEN_3074 = _GEN_40 ? ~_GEN_3073 & _GEN_2946 : ~_GEN_3033 & _GEN_2946;
  wire        _GEN_3075 = _GEN_914 | _GEN_3034;
  wire        _GEN_3076 = _GEN_40 ? ~_GEN_3075 & _GEN_2948 : ~_GEN_3034 & _GEN_2948;
  wire        _GEN_3077 = _GEN_917 | _GEN_3035;
  wire        _GEN_3078 = _GEN_40 ? ~_GEN_3077 & _GEN_2950 : ~_GEN_3035 & _GEN_2950;
  wire        _GEN_3079 = _GEN_920 | _GEN_3036;
  wire        _GEN_3080 = _GEN_40 ? ~_GEN_3079 & _GEN_2952 : ~_GEN_3036 & _GEN_2952;
  wire        _GEN_3081 = _GEN_923 | _GEN_3037;
  wire        _GEN_3082 = _GEN_40 ? ~_GEN_3081 & _GEN_2954 : ~_GEN_3037 & _GEN_2954;
  wire        _GEN_3083 = _GEN_926 | _GEN_3038;
  wire        _GEN_3084 = _GEN_40 ? ~_GEN_3083 & _GEN_2956 : ~_GEN_3038 & _GEN_2956;
  wire        _GEN_3085 = _GEN_929 | _GEN_3039;
  wire        _GEN_3086 = _GEN_40 ? ~_GEN_3085 & _GEN_2958 : ~_GEN_3039 & _GEN_2958;
  wire        _GEN_3087 = _GEN_932 | _GEN_3040;
  wire        _GEN_3088 = _GEN_40 ? ~_GEN_3087 & _GEN_2960 : ~_GEN_3040 & _GEN_2960;
  wire        _GEN_3089 = _GEN_935 | _GEN_3041;
  wire        _GEN_3090 = _GEN_40 ? ~_GEN_3089 & _GEN_2962 : ~_GEN_3041 & _GEN_2962;
  wire        _GEN_3091 = _GEN_938 | _GEN_3042;
  wire        _GEN_3092 = _GEN_40 ? ~_GEN_3091 & _GEN_2964 : ~_GEN_3042 & _GEN_2964;
  wire        _GEN_3093 = _GEN_941 | _GEN_3043;
  wire        _GEN_3094 = _GEN_40 ? ~_GEN_3093 & _GEN_2966 : ~_GEN_3043 & _GEN_2966;
  wire        _GEN_3095 = _GEN_944 | _GEN_3044;
  wire        _GEN_3096 = _GEN_40 ? ~_GEN_3095 & _GEN_2968 : ~_GEN_3044 & _GEN_2968;
  wire        _GEN_3097 = _GEN_947 | _GEN_3045;
  wire        _GEN_3098 = _GEN_40 ? ~_GEN_3097 & _GEN_2970 : ~_GEN_3045 & _GEN_2970;
  wire        _GEN_3099 = _GEN_950 | _GEN_3046;
  wire        _GEN_3100 = _GEN_40 ? ~_GEN_3099 & _GEN_2972 : ~_GEN_3046 & _GEN_2972;
  wire        _GEN_3101 = _GEN_953 | _GEN_3047;
  wire        _GEN_3102 = _GEN_40 ? ~_GEN_3101 & _GEN_2974 : ~_GEN_3047 & _GEN_2974;
  wire        _GEN_3103 = _GEN_956 | _GEN_3048;
  wire        _GEN_3104 = _GEN_40 ? ~_GEN_3103 & _GEN_2976 : ~_GEN_3048 & _GEN_2976;
  wire        _GEN_3105 = _GEN_959 | _GEN_3049;
  wire        _GEN_3106 = _GEN_40 ? ~_GEN_3105 & _GEN_2978 : ~_GEN_3049 & _GEN_2978;
  wire        _GEN_3107 = _GEN_962 | _GEN_3050;
  wire        _GEN_3108 = _GEN_40 ? ~_GEN_3107 & _GEN_2980 : ~_GEN_3050 & _GEN_2980;
  wire        _GEN_3109 = _GEN_965 | _GEN_3051;
  wire        _GEN_3110 = _GEN_40 ? ~_GEN_3109 & _GEN_2982 : ~_GEN_3051 & _GEN_2982;
  wire        _GEN_3111 = _GEN_968 | _GEN_3052;
  wire        _GEN_3112 = _GEN_40 ? ~_GEN_3111 & _GEN_2984 : ~_GEN_3052 & _GEN_2984;
  wire        _GEN_3113 = _GEN_971 | _GEN_3053;
  wire        _GEN_3114 = _GEN_40 ? ~_GEN_3113 & _GEN_2986 : ~_GEN_3053 & _GEN_2986;
  wire        _GEN_3115 = _GEN_974 | _GEN_3054;
  wire        _GEN_3116 = _GEN_40 ? ~_GEN_3115 & _GEN_2988 : ~_GEN_3054 & _GEN_2988;
  wire        _GEN_3117 = _GEN_977 | _GEN_3055;
  wire        _GEN_3118 = _GEN_40 ? ~_GEN_3117 & _GEN_2990 : ~_GEN_3055 & _GEN_2990;
  wire        _GEN_3119 = (&(io_wb_resps_7_bits_uop_rob_idx[6:2])) | _GEN_3056;
  wire        _GEN_3120 = _GEN_40 ? ~_GEN_3119 & _GEN_2992 : ~_GEN_3056 & _GEN_2992;
  wire        _GEN_3121 = _GEN_40 ? ~_GEN_3057 & _GEN_2993 : ~_GEN_3025 & _GEN_2993;
  wire        _GEN_3122 = _GEN_40 ? ~_GEN_3059 & _GEN_2994 : ~_GEN_3026 & _GEN_2994;
  wire        _GEN_3123 = _GEN_40 ? ~_GEN_3061 & _GEN_2995 : ~_GEN_3027 & _GEN_2995;
  wire        _GEN_3124 = _GEN_40 ? ~_GEN_3063 & _GEN_2996 : ~_GEN_3028 & _GEN_2996;
  wire        _GEN_3125 = _GEN_40 ? ~_GEN_3065 & _GEN_2997 : ~_GEN_3029 & _GEN_2997;
  wire        _GEN_3126 = _GEN_40 ? ~_GEN_3067 & _GEN_2998 : ~_GEN_3030 & _GEN_2998;
  wire        _GEN_3127 = _GEN_40 ? ~_GEN_3069 & _GEN_2999 : ~_GEN_3031 & _GEN_2999;
  wire        _GEN_3128 = _GEN_40 ? ~_GEN_3071 & _GEN_3000 : ~_GEN_3032 & _GEN_3000;
  wire        _GEN_3129 = _GEN_40 ? ~_GEN_3073 & _GEN_3001 : ~_GEN_3033 & _GEN_3001;
  wire        _GEN_3130 = _GEN_40 ? ~_GEN_3075 & _GEN_3002 : ~_GEN_3034 & _GEN_3002;
  wire        _GEN_3131 = _GEN_40 ? ~_GEN_3077 & _GEN_3003 : ~_GEN_3035 & _GEN_3003;
  wire        _GEN_3132 = _GEN_40 ? ~_GEN_3079 & _GEN_3004 : ~_GEN_3036 & _GEN_3004;
  wire        _GEN_3133 = _GEN_40 ? ~_GEN_3081 & _GEN_3005 : ~_GEN_3037 & _GEN_3005;
  wire        _GEN_3134 = _GEN_40 ? ~_GEN_3083 & _GEN_3006 : ~_GEN_3038 & _GEN_3006;
  wire        _GEN_3135 = _GEN_40 ? ~_GEN_3085 & _GEN_3007 : ~_GEN_3039 & _GEN_3007;
  wire        _GEN_3136 = _GEN_40 ? ~_GEN_3087 & _GEN_3008 : ~_GEN_3040 & _GEN_3008;
  wire        _GEN_3137 = _GEN_40 ? ~_GEN_3089 & _GEN_3009 : ~_GEN_3041 & _GEN_3009;
  wire        _GEN_3138 = _GEN_40 ? ~_GEN_3091 & _GEN_3010 : ~_GEN_3042 & _GEN_3010;
  wire        _GEN_3139 = _GEN_40 ? ~_GEN_3093 & _GEN_3011 : ~_GEN_3043 & _GEN_3011;
  wire        _GEN_3140 = _GEN_40 ? ~_GEN_3095 & _GEN_3012 : ~_GEN_3044 & _GEN_3012;
  wire        _GEN_3141 = _GEN_40 ? ~_GEN_3097 & _GEN_3013 : ~_GEN_3045 & _GEN_3013;
  wire        _GEN_3142 = _GEN_40 ? ~_GEN_3099 & _GEN_3014 : ~_GEN_3046 & _GEN_3014;
  wire        _GEN_3143 = _GEN_40 ? ~_GEN_3101 & _GEN_3015 : ~_GEN_3047 & _GEN_3015;
  wire        _GEN_3144 = _GEN_40 ? ~_GEN_3103 & _GEN_3016 : ~_GEN_3048 & _GEN_3016;
  wire        _GEN_3145 = _GEN_40 ? ~_GEN_3105 & _GEN_3017 : ~_GEN_3049 & _GEN_3017;
  wire        _GEN_3146 = _GEN_40 ? ~_GEN_3107 & _GEN_3018 : ~_GEN_3050 & _GEN_3018;
  wire        _GEN_3147 = _GEN_40 ? ~_GEN_3109 & _GEN_3019 : ~_GEN_3051 & _GEN_3019;
  wire        _GEN_3148 = _GEN_40 ? ~_GEN_3111 & _GEN_3020 : ~_GEN_3052 & _GEN_3020;
  wire        _GEN_3149 = _GEN_40 ? ~_GEN_3113 & _GEN_3021 : ~_GEN_3053 & _GEN_3021;
  wire        _GEN_3150 = _GEN_40 ? ~_GEN_3115 & _GEN_3022 : ~_GEN_3054 & _GEN_3022;
  wire        _GEN_3151 = _GEN_40 ? ~_GEN_3117 & _GEN_3023 : ~_GEN_3055 & _GEN_3023;
  wire        _GEN_3152 = _GEN_40 ? ~_GEN_3119 & _GEN_3024 : ~_GEN_3056 & _GEN_3024;
  wire        _GEN_3153 = _GEN_41 & _GEN_1014;
  wire        _GEN_3154 = _GEN_41 & _GEN_1016;
  wire        _GEN_3155 = _GEN_41 & _GEN_1018;
  wire        _GEN_3156 = _GEN_41 & _GEN_1020;
  wire        _GEN_3157 = _GEN_41 & _GEN_1022;
  wire        _GEN_3158 = _GEN_41 & _GEN_1024;
  wire        _GEN_3159 = _GEN_41 & _GEN_1026;
  wire        _GEN_3160 = _GEN_41 & _GEN_1028;
  wire        _GEN_3161 = _GEN_41 & _GEN_1030;
  wire        _GEN_3162 = _GEN_41 & _GEN_1032;
  wire        _GEN_3163 = _GEN_41 & _GEN_1034;
  wire        _GEN_3164 = _GEN_41 & _GEN_1036;
  wire        _GEN_3165 = _GEN_41 & _GEN_1038;
  wire        _GEN_3166 = _GEN_41 & _GEN_1040;
  wire        _GEN_3167 = _GEN_41 & _GEN_1042;
  wire        _GEN_3168 = _GEN_41 & _GEN_1044;
  wire        _GEN_3169 = _GEN_41 & _GEN_1046;
  wire        _GEN_3170 = _GEN_41 & _GEN_1048;
  wire        _GEN_3171 = _GEN_41 & _GEN_1050;
  wire        _GEN_3172 = _GEN_41 & _GEN_1052;
  wire        _GEN_3173 = _GEN_41 & _GEN_1054;
  wire        _GEN_3174 = _GEN_41 & _GEN_1056;
  wire        _GEN_3175 = _GEN_41 & _GEN_1058;
  wire        _GEN_3176 = _GEN_41 & _GEN_1060;
  wire        _GEN_3177 = _GEN_41 & _GEN_1062;
  wire        _GEN_3178 = _GEN_41 & _GEN_1064;
  wire        _GEN_3179 = _GEN_41 & _GEN_1066;
  wire        _GEN_3180 = _GEN_41 & _GEN_1068;
  wire        _GEN_3181 = _GEN_41 & _GEN_1070;
  wire        _GEN_3182 = _GEN_41 & _GEN_1072;
  wire        _GEN_3183 = _GEN_41 & _GEN_1074;
  wire        _GEN_3184 = _GEN_41 & (&(io_wb_resps_8_bits_uop_rob_idx[6:2]));
  wire        _GEN_3185 = _GEN_1077 | _GEN_3153;
  wire        _GEN_3186 = _GEN_42 ? ~_GEN_3185 & _GEN_3058 : ~_GEN_3153 & _GEN_3058;
  wire        _GEN_3187 = _GEN_1080 | _GEN_3154;
  wire        _GEN_3188 = _GEN_42 ? ~_GEN_3187 & _GEN_3060 : ~_GEN_3154 & _GEN_3060;
  wire        _GEN_3189 = _GEN_1083 | _GEN_3155;
  wire        _GEN_3190 = _GEN_42 ? ~_GEN_3189 & _GEN_3062 : ~_GEN_3155 & _GEN_3062;
  wire        _GEN_3191 = _GEN_1086 | _GEN_3156;
  wire        _GEN_3192 = _GEN_42 ? ~_GEN_3191 & _GEN_3064 : ~_GEN_3156 & _GEN_3064;
  wire        _GEN_3193 = _GEN_1089 | _GEN_3157;
  wire        _GEN_3194 = _GEN_42 ? ~_GEN_3193 & _GEN_3066 : ~_GEN_3157 & _GEN_3066;
  wire        _GEN_3195 = _GEN_1092 | _GEN_3158;
  wire        _GEN_3196 = _GEN_42 ? ~_GEN_3195 & _GEN_3068 : ~_GEN_3158 & _GEN_3068;
  wire        _GEN_3197 = _GEN_1095 | _GEN_3159;
  wire        _GEN_3198 = _GEN_42 ? ~_GEN_3197 & _GEN_3070 : ~_GEN_3159 & _GEN_3070;
  wire        _GEN_3199 = _GEN_1098 | _GEN_3160;
  wire        _GEN_3200 = _GEN_42 ? ~_GEN_3199 & _GEN_3072 : ~_GEN_3160 & _GEN_3072;
  wire        _GEN_3201 = _GEN_1101 | _GEN_3161;
  wire        _GEN_3202 = _GEN_42 ? ~_GEN_3201 & _GEN_3074 : ~_GEN_3161 & _GEN_3074;
  wire        _GEN_3203 = _GEN_1104 | _GEN_3162;
  wire        _GEN_3204 = _GEN_42 ? ~_GEN_3203 & _GEN_3076 : ~_GEN_3162 & _GEN_3076;
  wire        _GEN_3205 = _GEN_1107 | _GEN_3163;
  wire        _GEN_3206 = _GEN_42 ? ~_GEN_3205 & _GEN_3078 : ~_GEN_3163 & _GEN_3078;
  wire        _GEN_3207 = _GEN_1110 | _GEN_3164;
  wire        _GEN_3208 = _GEN_42 ? ~_GEN_3207 & _GEN_3080 : ~_GEN_3164 & _GEN_3080;
  wire        _GEN_3209 = _GEN_1113 | _GEN_3165;
  wire        _GEN_3210 = _GEN_42 ? ~_GEN_3209 & _GEN_3082 : ~_GEN_3165 & _GEN_3082;
  wire        _GEN_3211 = _GEN_1116 | _GEN_3166;
  wire        _GEN_3212 = _GEN_42 ? ~_GEN_3211 & _GEN_3084 : ~_GEN_3166 & _GEN_3084;
  wire        _GEN_3213 = _GEN_1119 | _GEN_3167;
  wire        _GEN_3214 = _GEN_42 ? ~_GEN_3213 & _GEN_3086 : ~_GEN_3167 & _GEN_3086;
  wire        _GEN_3215 = _GEN_1122 | _GEN_3168;
  wire        _GEN_3216 = _GEN_42 ? ~_GEN_3215 & _GEN_3088 : ~_GEN_3168 & _GEN_3088;
  wire        _GEN_3217 = _GEN_1125 | _GEN_3169;
  wire        _GEN_3218 = _GEN_42 ? ~_GEN_3217 & _GEN_3090 : ~_GEN_3169 & _GEN_3090;
  wire        _GEN_3219 = _GEN_1128 | _GEN_3170;
  wire        _GEN_3220 = _GEN_42 ? ~_GEN_3219 & _GEN_3092 : ~_GEN_3170 & _GEN_3092;
  wire        _GEN_3221 = _GEN_1131 | _GEN_3171;
  wire        _GEN_3222 = _GEN_42 ? ~_GEN_3221 & _GEN_3094 : ~_GEN_3171 & _GEN_3094;
  wire        _GEN_3223 = _GEN_1134 | _GEN_3172;
  wire        _GEN_3224 = _GEN_42 ? ~_GEN_3223 & _GEN_3096 : ~_GEN_3172 & _GEN_3096;
  wire        _GEN_3225 = _GEN_1137 | _GEN_3173;
  wire        _GEN_3226 = _GEN_42 ? ~_GEN_3225 & _GEN_3098 : ~_GEN_3173 & _GEN_3098;
  wire        _GEN_3227 = _GEN_1140 | _GEN_3174;
  wire        _GEN_3228 = _GEN_42 ? ~_GEN_3227 & _GEN_3100 : ~_GEN_3174 & _GEN_3100;
  wire        _GEN_3229 = _GEN_1143 | _GEN_3175;
  wire        _GEN_3230 = _GEN_42 ? ~_GEN_3229 & _GEN_3102 : ~_GEN_3175 & _GEN_3102;
  wire        _GEN_3231 = _GEN_1146 | _GEN_3176;
  wire        _GEN_3232 = _GEN_42 ? ~_GEN_3231 & _GEN_3104 : ~_GEN_3176 & _GEN_3104;
  wire        _GEN_3233 = _GEN_1149 | _GEN_3177;
  wire        _GEN_3234 = _GEN_42 ? ~_GEN_3233 & _GEN_3106 : ~_GEN_3177 & _GEN_3106;
  wire        _GEN_3235 = _GEN_1152 | _GEN_3178;
  wire        _GEN_3236 = _GEN_42 ? ~_GEN_3235 & _GEN_3108 : ~_GEN_3178 & _GEN_3108;
  wire        _GEN_3237 = _GEN_1155 | _GEN_3179;
  wire        _GEN_3238 = _GEN_42 ? ~_GEN_3237 & _GEN_3110 : ~_GEN_3179 & _GEN_3110;
  wire        _GEN_3239 = _GEN_1158 | _GEN_3180;
  wire        _GEN_3240 = _GEN_42 ? ~_GEN_3239 & _GEN_3112 : ~_GEN_3180 & _GEN_3112;
  wire        _GEN_3241 = _GEN_1161 | _GEN_3181;
  wire        _GEN_3242 = _GEN_42 ? ~_GEN_3241 & _GEN_3114 : ~_GEN_3181 & _GEN_3114;
  wire        _GEN_3243 = _GEN_1164 | _GEN_3182;
  wire        _GEN_3244 = _GEN_42 ? ~_GEN_3243 & _GEN_3116 : ~_GEN_3182 & _GEN_3116;
  wire        _GEN_3245 = _GEN_1167 | _GEN_3183;
  wire        _GEN_3246 = _GEN_42 ? ~_GEN_3245 & _GEN_3118 : ~_GEN_3183 & _GEN_3118;
  wire        _GEN_3247 = (&(io_wb_resps_9_bits_uop_rob_idx[6:2])) | _GEN_3184;
  wire        _GEN_3248 = _GEN_42 ? ~_GEN_3247 & _GEN_3120 : ~_GEN_3184 & _GEN_3120;
  wire        _GEN_3249 = _GEN_42 ? ~_GEN_3185 & _GEN_3121 : ~_GEN_3153 & _GEN_3121;
  wire        _GEN_3250 = _GEN_42 ? ~_GEN_3187 & _GEN_3122 : ~_GEN_3154 & _GEN_3122;
  wire        _GEN_3251 = _GEN_42 ? ~_GEN_3189 & _GEN_3123 : ~_GEN_3155 & _GEN_3123;
  wire        _GEN_3252 = _GEN_42 ? ~_GEN_3191 & _GEN_3124 : ~_GEN_3156 & _GEN_3124;
  wire        _GEN_3253 = _GEN_42 ? ~_GEN_3193 & _GEN_3125 : ~_GEN_3157 & _GEN_3125;
  wire        _GEN_3254 = _GEN_42 ? ~_GEN_3195 & _GEN_3126 : ~_GEN_3158 & _GEN_3126;
  wire        _GEN_3255 = _GEN_42 ? ~_GEN_3197 & _GEN_3127 : ~_GEN_3159 & _GEN_3127;
  wire        _GEN_3256 = _GEN_42 ? ~_GEN_3199 & _GEN_3128 : ~_GEN_3160 & _GEN_3128;
  wire        _GEN_3257 = _GEN_42 ? ~_GEN_3201 & _GEN_3129 : ~_GEN_3161 & _GEN_3129;
  wire        _GEN_3258 = _GEN_42 ? ~_GEN_3203 & _GEN_3130 : ~_GEN_3162 & _GEN_3130;
  wire        _GEN_3259 = _GEN_42 ? ~_GEN_3205 & _GEN_3131 : ~_GEN_3163 & _GEN_3131;
  wire        _GEN_3260 = _GEN_42 ? ~_GEN_3207 & _GEN_3132 : ~_GEN_3164 & _GEN_3132;
  wire        _GEN_3261 = _GEN_42 ? ~_GEN_3209 & _GEN_3133 : ~_GEN_3165 & _GEN_3133;
  wire        _GEN_3262 = _GEN_42 ? ~_GEN_3211 & _GEN_3134 : ~_GEN_3166 & _GEN_3134;
  wire        _GEN_3263 = _GEN_42 ? ~_GEN_3213 & _GEN_3135 : ~_GEN_3167 & _GEN_3135;
  wire        _GEN_3264 = _GEN_42 ? ~_GEN_3215 & _GEN_3136 : ~_GEN_3168 & _GEN_3136;
  wire        _GEN_3265 = _GEN_42 ? ~_GEN_3217 & _GEN_3137 : ~_GEN_3169 & _GEN_3137;
  wire        _GEN_3266 = _GEN_42 ? ~_GEN_3219 & _GEN_3138 : ~_GEN_3170 & _GEN_3138;
  wire        _GEN_3267 = _GEN_42 ? ~_GEN_3221 & _GEN_3139 : ~_GEN_3171 & _GEN_3139;
  wire        _GEN_3268 = _GEN_42 ? ~_GEN_3223 & _GEN_3140 : ~_GEN_3172 & _GEN_3140;
  wire        _GEN_3269 = _GEN_42 ? ~_GEN_3225 & _GEN_3141 : ~_GEN_3173 & _GEN_3141;
  wire        _GEN_3270 = _GEN_42 ? ~_GEN_3227 & _GEN_3142 : ~_GEN_3174 & _GEN_3142;
  wire        _GEN_3271 = _GEN_42 ? ~_GEN_3229 & _GEN_3143 : ~_GEN_3175 & _GEN_3143;
  wire        _GEN_3272 = _GEN_42 ? ~_GEN_3231 & _GEN_3144 : ~_GEN_3176 & _GEN_3144;
  wire        _GEN_3273 = _GEN_42 ? ~_GEN_3233 & _GEN_3145 : ~_GEN_3177 & _GEN_3145;
  wire        _GEN_3274 = _GEN_42 ? ~_GEN_3235 & _GEN_3146 : ~_GEN_3178 & _GEN_3146;
  wire        _GEN_3275 = _GEN_42 ? ~_GEN_3237 & _GEN_3147 : ~_GEN_3179 & _GEN_3147;
  wire        _GEN_3276 = _GEN_42 ? ~_GEN_3239 & _GEN_3148 : ~_GEN_3180 & _GEN_3148;
  wire        _GEN_3277 = _GEN_42 ? ~_GEN_3241 & _GEN_3149 : ~_GEN_3181 & _GEN_3149;
  wire        _GEN_3278 = _GEN_42 ? ~_GEN_3243 & _GEN_3150 : ~_GEN_3182 & _GEN_3150;
  wire        _GEN_3279 = _GEN_42 ? ~_GEN_3245 & _GEN_3151 : ~_GEN_3183 & _GEN_3151;
  wire        _GEN_3280 = _GEN_42 ? ~_GEN_3247 & _GEN_3152 : ~_GEN_3184 & _GEN_3152;
  wire        _GEN_3281 = _GEN_43 & _GEN_1204;
  wire        _GEN_3282 = _GEN_43 & _GEN_1206;
  wire        _GEN_3283 = _GEN_43 & _GEN_1208;
  wire        _GEN_3284 = _GEN_43 & _GEN_1210;
  wire        _GEN_3285 = _GEN_43 & _GEN_1212;
  wire        _GEN_3286 = _GEN_43 & _GEN_1214;
  wire        _GEN_3287 = _GEN_43 & _GEN_1216;
  wire        _GEN_3288 = _GEN_43 & _GEN_1218;
  wire        _GEN_3289 = _GEN_43 & _GEN_1220;
  wire        _GEN_3290 = _GEN_43 & _GEN_1222;
  wire        _GEN_3291 = _GEN_43 & _GEN_1224;
  wire        _GEN_3292 = _GEN_43 & _GEN_1226;
  wire        _GEN_3293 = _GEN_43 & _GEN_1228;
  wire        _GEN_3294 = _GEN_43 & _GEN_1230;
  wire        _GEN_3295 = _GEN_43 & _GEN_1232;
  wire        _GEN_3296 = _GEN_43 & _GEN_1234;
  wire        _GEN_3297 = _GEN_43 & _GEN_1236;
  wire        _GEN_3298 = _GEN_43 & _GEN_1238;
  wire        _GEN_3299 = _GEN_43 & _GEN_1240;
  wire        _GEN_3300 = _GEN_43 & _GEN_1242;
  wire        _GEN_3301 = _GEN_43 & _GEN_1244;
  wire        _GEN_3302 = _GEN_43 & _GEN_1246;
  wire        _GEN_3303 = _GEN_43 & _GEN_1248;
  wire        _GEN_3304 = _GEN_43 & _GEN_1250;
  wire        _GEN_3305 = _GEN_43 & _GEN_1252;
  wire        _GEN_3306 = _GEN_43 & _GEN_1254;
  wire        _GEN_3307 = _GEN_43 & _GEN_1256;
  wire        _GEN_3308 = _GEN_43 & _GEN_1258;
  wire        _GEN_3309 = _GEN_43 & _GEN_1260;
  wire        _GEN_3310 = _GEN_43 & _GEN_1262;
  wire        _GEN_3311 = _GEN_43 & _GEN_1264;
  wire        _GEN_3312 = _GEN_43 & (&(io_lsu_clr_bsy_0_bits[6:2]));
  wire        _GEN_3313 = _GEN_1267 | _GEN_3281;
  wire        _GEN_3314 = _GEN_1269 | _GEN_3282;
  wire        _GEN_3315 = _GEN_1271 | _GEN_3283;
  wire        _GEN_3316 = _GEN_1273 | _GEN_3284;
  wire        _GEN_3317 = _GEN_1275 | _GEN_3285;
  wire        _GEN_3318 = _GEN_1277 | _GEN_3286;
  wire        _GEN_3319 = _GEN_1279 | _GEN_3287;
  wire        _GEN_3320 = _GEN_1281 | _GEN_3288;
  wire        _GEN_3321 = _GEN_1283 | _GEN_3289;
  wire        _GEN_3322 = _GEN_1285 | _GEN_3290;
  wire        _GEN_3323 = _GEN_1287 | _GEN_3291;
  wire        _GEN_3324 = _GEN_1289 | _GEN_3292;
  wire        _GEN_3325 = _GEN_1291 | _GEN_3293;
  wire        _GEN_3326 = _GEN_1293 | _GEN_3294;
  wire        _GEN_3327 = _GEN_1295 | _GEN_3295;
  wire        _GEN_3328 = _GEN_1297 | _GEN_3296;
  wire        _GEN_3329 = _GEN_1299 | _GEN_3297;
  wire        _GEN_3330 = _GEN_1301 | _GEN_3298;
  wire        _GEN_3331 = _GEN_1303 | _GEN_3299;
  wire        _GEN_3332 = _GEN_1305 | _GEN_3300;
  wire        _GEN_3333 = _GEN_1307 | _GEN_3301;
  wire        _GEN_3334 = _GEN_1309 | _GEN_3302;
  wire        _GEN_3335 = _GEN_1311 | _GEN_3303;
  wire        _GEN_3336 = _GEN_1313 | _GEN_3304;
  wire        _GEN_3337 = _GEN_1315 | _GEN_3305;
  wire        _GEN_3338 = _GEN_1317 | _GEN_3306;
  wire        _GEN_3339 = _GEN_1319 | _GEN_3307;
  wire        _GEN_3340 = _GEN_1321 | _GEN_3308;
  wire        _GEN_3341 = _GEN_1323 | _GEN_3309;
  wire        _GEN_3342 = _GEN_1325 | _GEN_3310;
  wire        _GEN_3343 = _GEN_1327 | _GEN_3311;
  wire        _GEN_3344 = (&(io_lsu_clr_bsy_1_bits[6:2])) | _GEN_3312;
  wire        _GEN_3345 = _GEN_45 & _GEN_1330;
  wire        _GEN_3346 = _GEN_45 & _GEN_1332;
  wire        _GEN_3347 = _GEN_45 & _GEN_1334;
  wire        _GEN_3348 = _GEN_45 & _GEN_1336;
  wire        _GEN_3349 = _GEN_45 & _GEN_1338;
  wire        _GEN_3350 = _GEN_45 & _GEN_1340;
  wire        _GEN_3351 = _GEN_45 & _GEN_1342;
  wire        _GEN_3352 = _GEN_45 & _GEN_1344;
  wire        _GEN_3353 = _GEN_45 & _GEN_1346;
  wire        _GEN_3354 = _GEN_45 & _GEN_1348;
  wire        _GEN_3355 = _GEN_45 & _GEN_1350;
  wire        _GEN_3356 = _GEN_45 & _GEN_1352;
  wire        _GEN_3357 = _GEN_45 & _GEN_1354;
  wire        _GEN_3358 = _GEN_45 & _GEN_1356;
  wire        _GEN_3359 = _GEN_45 & _GEN_1358;
  wire        _GEN_3360 = _GEN_45 & _GEN_1360;
  wire        _GEN_3361 = _GEN_45 & _GEN_1362;
  wire        _GEN_3362 = _GEN_45 & _GEN_1364;
  wire        _GEN_3363 = _GEN_45 & _GEN_1366;
  wire        _GEN_3364 = _GEN_45 & _GEN_1368;
  wire        _GEN_3365 = _GEN_45 & _GEN_1370;
  wire        _GEN_3366 = _GEN_45 & _GEN_1372;
  wire        _GEN_3367 = _GEN_45 & _GEN_1374;
  wire        _GEN_3368 = _GEN_45 & _GEN_1376;
  wire        _GEN_3369 = _GEN_45 & _GEN_1378;
  wire        _GEN_3370 = _GEN_45 & _GEN_1380;
  wire        _GEN_3371 = _GEN_45 & _GEN_1382;
  wire        _GEN_3372 = _GEN_45 & _GEN_1384;
  wire        _GEN_3373 = _GEN_45 & _GEN_1386;
  wire        _GEN_3374 = _GEN_45 & _GEN_1388;
  wire        _GEN_3375 = _GEN_45 & _GEN_1390;
  wire        _GEN_3376 = _GEN_45 & (&(io_lsu_clr_bsy_2_bits[6:2]));
  wire        _GEN_3377 = io_fflags_0_valid & io_fflags_0_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_3378 = io_fflags_2_valid & io_fflags_2_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_3379 = io_fflags_3_valid & io_fflags_3_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_3380 = rbk_row_2 & _GEN_1520;
  wire        _GEN_3381 = rbk_row_2 & _GEN_1522;
  wire        _GEN_3382 = rbk_row_2 & _GEN_1524;
  wire        _GEN_3383 = rbk_row_2 & _GEN_1526;
  wire        _GEN_3384 = rbk_row_2 & _GEN_1528;
  wire        _GEN_3385 = rbk_row_2 & _GEN_1530;
  wire        _GEN_3386 = rbk_row_2 & _GEN_1532;
  wire        _GEN_3387 = rbk_row_2 & _GEN_1534;
  wire        _GEN_3388 = rbk_row_2 & _GEN_1536;
  wire        _GEN_3389 = rbk_row_2 & _GEN_1538;
  wire        _GEN_3390 = rbk_row_2 & _GEN_1540;
  wire        _GEN_3391 = rbk_row_2 & _GEN_1542;
  wire        _GEN_3392 = rbk_row_2 & _GEN_1544;
  wire        _GEN_3393 = rbk_row_2 & _GEN_1546;
  wire        _GEN_3394 = rbk_row_2 & _GEN_1548;
  wire        _GEN_3395 = rbk_row_2 & _GEN_1550;
  wire        _GEN_3396 = rbk_row_2 & _GEN_1552;
  wire        _GEN_3397 = rbk_row_2 & _GEN_1554;
  wire        _GEN_3398 = rbk_row_2 & _GEN_1556;
  wire        _GEN_3399 = rbk_row_2 & _GEN_1558;
  wire        _GEN_3400 = rbk_row_2 & _GEN_1560;
  wire        _GEN_3401 = rbk_row_2 & _GEN_1562;
  wire        _GEN_3402 = rbk_row_2 & _GEN_1564;
  wire        _GEN_3403 = rbk_row_2 & _GEN_1566;
  wire        _GEN_3404 = rbk_row_2 & _GEN_1568;
  wire        _GEN_3405 = rbk_row_2 & _GEN_1570;
  wire        _GEN_3406 = rbk_row_2 & _GEN_1572;
  wire        _GEN_3407 = rbk_row_2 & _GEN_1574;
  wire        _GEN_3408 = rbk_row_2 & _GEN_1576;
  wire        _GEN_3409 = rbk_row_2 & _GEN_1578;
  wire        _GEN_3410 = rbk_row_2 & _GEN_1580;
  wire        _GEN_3411 = rbk_row_2 & (&com_idx);
  wire [19:0] _GEN_3412 = io_brupdate_b1_mispredict_mask & rob_uop_2_0_br_mask;
  wire [19:0] _GEN_3413 = io_brupdate_b1_mispredict_mask & rob_uop_2_1_br_mask;
  wire [19:0] _GEN_3414 = io_brupdate_b1_mispredict_mask & rob_uop_2_2_br_mask;
  wire [19:0] _GEN_3415 = io_brupdate_b1_mispredict_mask & rob_uop_2_3_br_mask;
  wire [19:0] _GEN_3416 = io_brupdate_b1_mispredict_mask & rob_uop_2_4_br_mask;
  wire [19:0] _GEN_3417 = io_brupdate_b1_mispredict_mask & rob_uop_2_5_br_mask;
  wire [19:0] _GEN_3418 = io_brupdate_b1_mispredict_mask & rob_uop_2_6_br_mask;
  wire [19:0] _GEN_3419 = io_brupdate_b1_mispredict_mask & rob_uop_2_7_br_mask;
  wire [19:0] _GEN_3420 = io_brupdate_b1_mispredict_mask & rob_uop_2_8_br_mask;
  wire [19:0] _GEN_3421 = io_brupdate_b1_mispredict_mask & rob_uop_2_9_br_mask;
  wire [19:0] _GEN_3422 = io_brupdate_b1_mispredict_mask & rob_uop_2_10_br_mask;
  wire [19:0] _GEN_3423 = io_brupdate_b1_mispredict_mask & rob_uop_2_11_br_mask;
  wire [19:0] _GEN_3424 = io_brupdate_b1_mispredict_mask & rob_uop_2_12_br_mask;
  wire [19:0] _GEN_3425 = io_brupdate_b1_mispredict_mask & rob_uop_2_13_br_mask;
  wire [19:0] _GEN_3426 = io_brupdate_b1_mispredict_mask & rob_uop_2_14_br_mask;
  wire [19:0] _GEN_3427 = io_brupdate_b1_mispredict_mask & rob_uop_2_15_br_mask;
  wire [19:0] _GEN_3428 = io_brupdate_b1_mispredict_mask & rob_uop_2_16_br_mask;
  wire [19:0] _GEN_3429 = io_brupdate_b1_mispredict_mask & rob_uop_2_17_br_mask;
  wire [19:0] _GEN_3430 = io_brupdate_b1_mispredict_mask & rob_uop_2_18_br_mask;
  wire [19:0] _GEN_3431 = io_brupdate_b1_mispredict_mask & rob_uop_2_19_br_mask;
  wire [19:0] _GEN_3432 = io_brupdate_b1_mispredict_mask & rob_uop_2_20_br_mask;
  wire [19:0] _GEN_3433 = io_brupdate_b1_mispredict_mask & rob_uop_2_21_br_mask;
  wire [19:0] _GEN_3434 = io_brupdate_b1_mispredict_mask & rob_uop_2_22_br_mask;
  wire [19:0] _GEN_3435 = io_brupdate_b1_mispredict_mask & rob_uop_2_23_br_mask;
  wire [19:0] _GEN_3436 = io_brupdate_b1_mispredict_mask & rob_uop_2_24_br_mask;
  wire [19:0] _GEN_3437 = io_brupdate_b1_mispredict_mask & rob_uop_2_25_br_mask;
  wire [19:0] _GEN_3438 = io_brupdate_b1_mispredict_mask & rob_uop_2_26_br_mask;
  wire [19:0] _GEN_3439 = io_brupdate_b1_mispredict_mask & rob_uop_2_27_br_mask;
  wire [19:0] _GEN_3440 = io_brupdate_b1_mispredict_mask & rob_uop_2_28_br_mask;
  wire [19:0] _GEN_3441 = io_brupdate_b1_mispredict_mask & rob_uop_2_29_br_mask;
  wire [19:0] _GEN_3442 = io_brupdate_b1_mispredict_mask & rob_uop_2_30_br_mask;
  wire [19:0] _GEN_3443 = io_brupdate_b1_mispredict_mask & rob_uop_2_31_br_mask;
  wire        _GEN_3444 = io_enq_valids_3 & _GEN_127;
  wire        _GEN_3445 = io_enq_valids_3 & _GEN_129;
  wire        _GEN_3446 = io_enq_valids_3 & _GEN_131;
  wire        _GEN_3447 = io_enq_valids_3 & _GEN_133;
  wire        _GEN_3448 = io_enq_valids_3 & _GEN_135;
  wire        _GEN_3449 = io_enq_valids_3 & _GEN_137;
  wire        _GEN_3450 = io_enq_valids_3 & _GEN_139;
  wire        _GEN_3451 = io_enq_valids_3 & _GEN_141;
  wire        _GEN_3452 = io_enq_valids_3 & _GEN_143;
  wire        _GEN_3453 = io_enq_valids_3 & _GEN_145;
  wire        _GEN_3454 = io_enq_valids_3 & _GEN_147;
  wire        _GEN_3455 = io_enq_valids_3 & _GEN_149;
  wire        _GEN_3456 = io_enq_valids_3 & _GEN_151;
  wire        _GEN_3457 = io_enq_valids_3 & _GEN_153;
  wire        _GEN_3458 = io_enq_valids_3 & _GEN_155;
  wire        _GEN_3459 = io_enq_valids_3 & _GEN_157;
  wire        _GEN_3460 = io_enq_valids_3 & _GEN_159;
  wire        _GEN_3461 = io_enq_valids_3 & _GEN_161;
  wire        _GEN_3462 = io_enq_valids_3 & _GEN_163;
  wire        _GEN_3463 = io_enq_valids_3 & _GEN_165;
  wire        _GEN_3464 = io_enq_valids_3 & _GEN_167;
  wire        _GEN_3465 = io_enq_valids_3 & _GEN_169;
  wire        _GEN_3466 = io_enq_valids_3 & _GEN_171;
  wire        _GEN_3467 = io_enq_valids_3 & _GEN_173;
  wire        _GEN_3468 = io_enq_valids_3 & _GEN_175;
  wire        _GEN_3469 = io_enq_valids_3 & _GEN_177;
  wire        _GEN_3470 = io_enq_valids_3 & _GEN_179;
  wire        _GEN_3471 = io_enq_valids_3 & _GEN_181;
  wire        _GEN_3472 = io_enq_valids_3 & _GEN_183;
  wire        _GEN_3473 = io_enq_valids_3 & _GEN_185;
  wire        _GEN_3474 = io_enq_valids_3 & _GEN_187;
  wire        _GEN_3475 = io_enq_valids_3 & (&rob_tail);
  wire        _rob_bsy_T_6 = io_enq_uops_3_is_fence | io_enq_uops_3_is_fencei;
  wire        _GEN_3476 = _GEN_3444 ? ~_rob_bsy_T_6 : rob_bsy_3_0;
  wire        _GEN_3477 = _GEN_3445 ? ~_rob_bsy_T_6 : rob_bsy_3_1;
  wire        _GEN_3478 = _GEN_3446 ? ~_rob_bsy_T_6 : rob_bsy_3_2;
  wire        _GEN_3479 = _GEN_3447 ? ~_rob_bsy_T_6 : rob_bsy_3_3;
  wire        _GEN_3480 = _GEN_3448 ? ~_rob_bsy_T_6 : rob_bsy_3_4;
  wire        _GEN_3481 = _GEN_3449 ? ~_rob_bsy_T_6 : rob_bsy_3_5;
  wire        _GEN_3482 = _GEN_3450 ? ~_rob_bsy_T_6 : rob_bsy_3_6;
  wire        _GEN_3483 = _GEN_3451 ? ~_rob_bsy_T_6 : rob_bsy_3_7;
  wire        _GEN_3484 = _GEN_3452 ? ~_rob_bsy_T_6 : rob_bsy_3_8;
  wire        _GEN_3485 = _GEN_3453 ? ~_rob_bsy_T_6 : rob_bsy_3_9;
  wire        _GEN_3486 = _GEN_3454 ? ~_rob_bsy_T_6 : rob_bsy_3_10;
  wire        _GEN_3487 = _GEN_3455 ? ~_rob_bsy_T_6 : rob_bsy_3_11;
  wire        _GEN_3488 = _GEN_3456 ? ~_rob_bsy_T_6 : rob_bsy_3_12;
  wire        _GEN_3489 = _GEN_3457 ? ~_rob_bsy_T_6 : rob_bsy_3_13;
  wire        _GEN_3490 = _GEN_3458 ? ~_rob_bsy_T_6 : rob_bsy_3_14;
  wire        _GEN_3491 = _GEN_3459 ? ~_rob_bsy_T_6 : rob_bsy_3_15;
  wire        _GEN_3492 = _GEN_3460 ? ~_rob_bsy_T_6 : rob_bsy_3_16;
  wire        _GEN_3493 = _GEN_3461 ? ~_rob_bsy_T_6 : rob_bsy_3_17;
  wire        _GEN_3494 = _GEN_3462 ? ~_rob_bsy_T_6 : rob_bsy_3_18;
  wire        _GEN_3495 = _GEN_3463 ? ~_rob_bsy_T_6 : rob_bsy_3_19;
  wire        _GEN_3496 = _GEN_3464 ? ~_rob_bsy_T_6 : rob_bsy_3_20;
  wire        _GEN_3497 = _GEN_3465 ? ~_rob_bsy_T_6 : rob_bsy_3_21;
  wire        _GEN_3498 = _GEN_3466 ? ~_rob_bsy_T_6 : rob_bsy_3_22;
  wire        _GEN_3499 = _GEN_3467 ? ~_rob_bsy_T_6 : rob_bsy_3_23;
  wire        _GEN_3500 = _GEN_3468 ? ~_rob_bsy_T_6 : rob_bsy_3_24;
  wire        _GEN_3501 = _GEN_3469 ? ~_rob_bsy_T_6 : rob_bsy_3_25;
  wire        _GEN_3502 = _GEN_3470 ? ~_rob_bsy_T_6 : rob_bsy_3_26;
  wire        _GEN_3503 = _GEN_3471 ? ~_rob_bsy_T_6 : rob_bsy_3_27;
  wire        _GEN_3504 = _GEN_3472 ? ~_rob_bsy_T_6 : rob_bsy_3_28;
  wire        _GEN_3505 = _GEN_3473 ? ~_rob_bsy_T_6 : rob_bsy_3_29;
  wire        _GEN_3506 = _GEN_3474 ? ~_rob_bsy_T_6 : rob_bsy_3_30;
  wire        _GEN_3507 = _GEN_3475 ? ~_rob_bsy_T_6 : rob_bsy_3_31;
  wire        _rob_unsafe_T_19 = io_enq_uops_3_uses_ldq | io_enq_uops_3_uses_stq & ~io_enq_uops_3_is_fence | io_enq_uops_3_is_br | io_enq_uops_3_is_jalr;
  wire        _GEN_3508 = _GEN_3444 ? _rob_unsafe_T_19 : rob_unsafe_3_0;
  wire        _GEN_3509 = _GEN_3445 ? _rob_unsafe_T_19 : rob_unsafe_3_1;
  wire        _GEN_3510 = _GEN_3446 ? _rob_unsafe_T_19 : rob_unsafe_3_2;
  wire        _GEN_3511 = _GEN_3447 ? _rob_unsafe_T_19 : rob_unsafe_3_3;
  wire        _GEN_3512 = _GEN_3448 ? _rob_unsafe_T_19 : rob_unsafe_3_4;
  wire        _GEN_3513 = _GEN_3449 ? _rob_unsafe_T_19 : rob_unsafe_3_5;
  wire        _GEN_3514 = _GEN_3450 ? _rob_unsafe_T_19 : rob_unsafe_3_6;
  wire        _GEN_3515 = _GEN_3451 ? _rob_unsafe_T_19 : rob_unsafe_3_7;
  wire        _GEN_3516 = _GEN_3452 ? _rob_unsafe_T_19 : rob_unsafe_3_8;
  wire        _GEN_3517 = _GEN_3453 ? _rob_unsafe_T_19 : rob_unsafe_3_9;
  wire        _GEN_3518 = _GEN_3454 ? _rob_unsafe_T_19 : rob_unsafe_3_10;
  wire        _GEN_3519 = _GEN_3455 ? _rob_unsafe_T_19 : rob_unsafe_3_11;
  wire        _GEN_3520 = _GEN_3456 ? _rob_unsafe_T_19 : rob_unsafe_3_12;
  wire        _GEN_3521 = _GEN_3457 ? _rob_unsafe_T_19 : rob_unsafe_3_13;
  wire        _GEN_3522 = _GEN_3458 ? _rob_unsafe_T_19 : rob_unsafe_3_14;
  wire        _GEN_3523 = _GEN_3459 ? _rob_unsafe_T_19 : rob_unsafe_3_15;
  wire        _GEN_3524 = _GEN_3460 ? _rob_unsafe_T_19 : rob_unsafe_3_16;
  wire        _GEN_3525 = _GEN_3461 ? _rob_unsafe_T_19 : rob_unsafe_3_17;
  wire        _GEN_3526 = _GEN_3462 ? _rob_unsafe_T_19 : rob_unsafe_3_18;
  wire        _GEN_3527 = _GEN_3463 ? _rob_unsafe_T_19 : rob_unsafe_3_19;
  wire        _GEN_3528 = _GEN_3464 ? _rob_unsafe_T_19 : rob_unsafe_3_20;
  wire        _GEN_3529 = _GEN_3465 ? _rob_unsafe_T_19 : rob_unsafe_3_21;
  wire        _GEN_3530 = _GEN_3466 ? _rob_unsafe_T_19 : rob_unsafe_3_22;
  wire        _GEN_3531 = _GEN_3467 ? _rob_unsafe_T_19 : rob_unsafe_3_23;
  wire        _GEN_3532 = _GEN_3468 ? _rob_unsafe_T_19 : rob_unsafe_3_24;
  wire        _GEN_3533 = _GEN_3469 ? _rob_unsafe_T_19 : rob_unsafe_3_25;
  wire        _GEN_3534 = _GEN_3470 ? _rob_unsafe_T_19 : rob_unsafe_3_26;
  wire        _GEN_3535 = _GEN_3471 ? _rob_unsafe_T_19 : rob_unsafe_3_27;
  wire        _GEN_3536 = _GEN_3472 ? _rob_unsafe_T_19 : rob_unsafe_3_28;
  wire        _GEN_3537 = _GEN_3473 ? _rob_unsafe_T_19 : rob_unsafe_3_29;
  wire        _GEN_3538 = _GEN_3474 ? _rob_unsafe_T_19 : rob_unsafe_3_30;
  wire        _GEN_3539 = _GEN_3475 ? _rob_unsafe_T_19 : rob_unsafe_3_31;
  wire        _GEN_3540 = _GEN_49 & _GEN_254;
  wire        _GEN_3541 = _GEN_49 & _GEN_256;
  wire        _GEN_3542 = _GEN_49 & _GEN_258;
  wire        _GEN_3543 = _GEN_49 & _GEN_260;
  wire        _GEN_3544 = _GEN_49 & _GEN_262;
  wire        _GEN_3545 = _GEN_49 & _GEN_264;
  wire        _GEN_3546 = _GEN_49 & _GEN_266;
  wire        _GEN_3547 = _GEN_49 & _GEN_268;
  wire        _GEN_3548 = _GEN_49 & _GEN_270;
  wire        _GEN_3549 = _GEN_49 & _GEN_272;
  wire        _GEN_3550 = _GEN_49 & _GEN_274;
  wire        _GEN_3551 = _GEN_49 & _GEN_276;
  wire        _GEN_3552 = _GEN_49 & _GEN_278;
  wire        _GEN_3553 = _GEN_49 & _GEN_280;
  wire        _GEN_3554 = _GEN_49 & _GEN_282;
  wire        _GEN_3555 = _GEN_49 & _GEN_284;
  wire        _GEN_3556 = _GEN_49 & _GEN_286;
  wire        _GEN_3557 = _GEN_49 & _GEN_288;
  wire        _GEN_3558 = _GEN_49 & _GEN_290;
  wire        _GEN_3559 = _GEN_49 & _GEN_292;
  wire        _GEN_3560 = _GEN_49 & _GEN_294;
  wire        _GEN_3561 = _GEN_49 & _GEN_296;
  wire        _GEN_3562 = _GEN_49 & _GEN_298;
  wire        _GEN_3563 = _GEN_49 & _GEN_300;
  wire        _GEN_3564 = _GEN_49 & _GEN_302;
  wire        _GEN_3565 = _GEN_49 & _GEN_304;
  wire        _GEN_3566 = _GEN_49 & _GEN_306;
  wire        _GEN_3567 = _GEN_49 & _GEN_308;
  wire        _GEN_3568 = _GEN_49 & _GEN_310;
  wire        _GEN_3569 = _GEN_49 & _GEN_312;
  wire        _GEN_3570 = _GEN_49 & _GEN_314;
  wire        _GEN_3571 = _GEN_49 & (&(io_wb_resps_0_bits_uop_rob_idx[6:2]));
  wire        _GEN_3572 = _GEN_317 | _GEN_3540;
  wire        _GEN_3573 = _GEN_50 ? ~_GEN_3572 & _GEN_3476 : ~_GEN_3540 & _GEN_3476;
  wire        _GEN_3574 = _GEN_320 | _GEN_3541;
  wire        _GEN_3575 = _GEN_50 ? ~_GEN_3574 & _GEN_3477 : ~_GEN_3541 & _GEN_3477;
  wire        _GEN_3576 = _GEN_323 | _GEN_3542;
  wire        _GEN_3577 = _GEN_50 ? ~_GEN_3576 & _GEN_3478 : ~_GEN_3542 & _GEN_3478;
  wire        _GEN_3578 = _GEN_326 | _GEN_3543;
  wire        _GEN_3579 = _GEN_50 ? ~_GEN_3578 & _GEN_3479 : ~_GEN_3543 & _GEN_3479;
  wire        _GEN_3580 = _GEN_329 | _GEN_3544;
  wire        _GEN_3581 = _GEN_50 ? ~_GEN_3580 & _GEN_3480 : ~_GEN_3544 & _GEN_3480;
  wire        _GEN_3582 = _GEN_332 | _GEN_3545;
  wire        _GEN_3583 = _GEN_50 ? ~_GEN_3582 & _GEN_3481 : ~_GEN_3545 & _GEN_3481;
  wire        _GEN_3584 = _GEN_335 | _GEN_3546;
  wire        _GEN_3585 = _GEN_50 ? ~_GEN_3584 & _GEN_3482 : ~_GEN_3546 & _GEN_3482;
  wire        _GEN_3586 = _GEN_338 | _GEN_3547;
  wire        _GEN_3587 = _GEN_50 ? ~_GEN_3586 & _GEN_3483 : ~_GEN_3547 & _GEN_3483;
  wire        _GEN_3588 = _GEN_341 | _GEN_3548;
  wire        _GEN_3589 = _GEN_50 ? ~_GEN_3588 & _GEN_3484 : ~_GEN_3548 & _GEN_3484;
  wire        _GEN_3590 = _GEN_344 | _GEN_3549;
  wire        _GEN_3591 = _GEN_50 ? ~_GEN_3590 & _GEN_3485 : ~_GEN_3549 & _GEN_3485;
  wire        _GEN_3592 = _GEN_347 | _GEN_3550;
  wire        _GEN_3593 = _GEN_50 ? ~_GEN_3592 & _GEN_3486 : ~_GEN_3550 & _GEN_3486;
  wire        _GEN_3594 = _GEN_350 | _GEN_3551;
  wire        _GEN_3595 = _GEN_50 ? ~_GEN_3594 & _GEN_3487 : ~_GEN_3551 & _GEN_3487;
  wire        _GEN_3596 = _GEN_353 | _GEN_3552;
  wire        _GEN_3597 = _GEN_50 ? ~_GEN_3596 & _GEN_3488 : ~_GEN_3552 & _GEN_3488;
  wire        _GEN_3598 = _GEN_356 | _GEN_3553;
  wire        _GEN_3599 = _GEN_50 ? ~_GEN_3598 & _GEN_3489 : ~_GEN_3553 & _GEN_3489;
  wire        _GEN_3600 = _GEN_359 | _GEN_3554;
  wire        _GEN_3601 = _GEN_50 ? ~_GEN_3600 & _GEN_3490 : ~_GEN_3554 & _GEN_3490;
  wire        _GEN_3602 = _GEN_362 | _GEN_3555;
  wire        _GEN_3603 = _GEN_50 ? ~_GEN_3602 & _GEN_3491 : ~_GEN_3555 & _GEN_3491;
  wire        _GEN_3604 = _GEN_365 | _GEN_3556;
  wire        _GEN_3605 = _GEN_50 ? ~_GEN_3604 & _GEN_3492 : ~_GEN_3556 & _GEN_3492;
  wire        _GEN_3606 = _GEN_368 | _GEN_3557;
  wire        _GEN_3607 = _GEN_50 ? ~_GEN_3606 & _GEN_3493 : ~_GEN_3557 & _GEN_3493;
  wire        _GEN_3608 = _GEN_371 | _GEN_3558;
  wire        _GEN_3609 = _GEN_50 ? ~_GEN_3608 & _GEN_3494 : ~_GEN_3558 & _GEN_3494;
  wire        _GEN_3610 = _GEN_374 | _GEN_3559;
  wire        _GEN_3611 = _GEN_50 ? ~_GEN_3610 & _GEN_3495 : ~_GEN_3559 & _GEN_3495;
  wire        _GEN_3612 = _GEN_377 | _GEN_3560;
  wire        _GEN_3613 = _GEN_50 ? ~_GEN_3612 & _GEN_3496 : ~_GEN_3560 & _GEN_3496;
  wire        _GEN_3614 = _GEN_380 | _GEN_3561;
  wire        _GEN_3615 = _GEN_50 ? ~_GEN_3614 & _GEN_3497 : ~_GEN_3561 & _GEN_3497;
  wire        _GEN_3616 = _GEN_383 | _GEN_3562;
  wire        _GEN_3617 = _GEN_50 ? ~_GEN_3616 & _GEN_3498 : ~_GEN_3562 & _GEN_3498;
  wire        _GEN_3618 = _GEN_386 | _GEN_3563;
  wire        _GEN_3619 = _GEN_50 ? ~_GEN_3618 & _GEN_3499 : ~_GEN_3563 & _GEN_3499;
  wire        _GEN_3620 = _GEN_389 | _GEN_3564;
  wire        _GEN_3621 = _GEN_50 ? ~_GEN_3620 & _GEN_3500 : ~_GEN_3564 & _GEN_3500;
  wire        _GEN_3622 = _GEN_392 | _GEN_3565;
  wire        _GEN_3623 = _GEN_50 ? ~_GEN_3622 & _GEN_3501 : ~_GEN_3565 & _GEN_3501;
  wire        _GEN_3624 = _GEN_395 | _GEN_3566;
  wire        _GEN_3625 = _GEN_50 ? ~_GEN_3624 & _GEN_3502 : ~_GEN_3566 & _GEN_3502;
  wire        _GEN_3626 = _GEN_398 | _GEN_3567;
  wire        _GEN_3627 = _GEN_50 ? ~_GEN_3626 & _GEN_3503 : ~_GEN_3567 & _GEN_3503;
  wire        _GEN_3628 = _GEN_401 | _GEN_3568;
  wire        _GEN_3629 = _GEN_50 ? ~_GEN_3628 & _GEN_3504 : ~_GEN_3568 & _GEN_3504;
  wire        _GEN_3630 = _GEN_404 | _GEN_3569;
  wire        _GEN_3631 = _GEN_50 ? ~_GEN_3630 & _GEN_3505 : ~_GEN_3569 & _GEN_3505;
  wire        _GEN_3632 = _GEN_407 | _GEN_3570;
  wire        _GEN_3633 = _GEN_50 ? ~_GEN_3632 & _GEN_3506 : ~_GEN_3570 & _GEN_3506;
  wire        _GEN_3634 = (&(io_wb_resps_1_bits_uop_rob_idx[6:2])) | _GEN_3571;
  wire        _GEN_3635 = _GEN_50 ? ~_GEN_3634 & _GEN_3507 : ~_GEN_3571 & _GEN_3507;
  wire        _GEN_3636 = _GEN_50 ? ~_GEN_3572 & _GEN_3508 : ~_GEN_3540 & _GEN_3508;
  wire        _GEN_3637 = _GEN_50 ? ~_GEN_3574 & _GEN_3509 : ~_GEN_3541 & _GEN_3509;
  wire        _GEN_3638 = _GEN_50 ? ~_GEN_3576 & _GEN_3510 : ~_GEN_3542 & _GEN_3510;
  wire        _GEN_3639 = _GEN_50 ? ~_GEN_3578 & _GEN_3511 : ~_GEN_3543 & _GEN_3511;
  wire        _GEN_3640 = _GEN_50 ? ~_GEN_3580 & _GEN_3512 : ~_GEN_3544 & _GEN_3512;
  wire        _GEN_3641 = _GEN_50 ? ~_GEN_3582 & _GEN_3513 : ~_GEN_3545 & _GEN_3513;
  wire        _GEN_3642 = _GEN_50 ? ~_GEN_3584 & _GEN_3514 : ~_GEN_3546 & _GEN_3514;
  wire        _GEN_3643 = _GEN_50 ? ~_GEN_3586 & _GEN_3515 : ~_GEN_3547 & _GEN_3515;
  wire        _GEN_3644 = _GEN_50 ? ~_GEN_3588 & _GEN_3516 : ~_GEN_3548 & _GEN_3516;
  wire        _GEN_3645 = _GEN_50 ? ~_GEN_3590 & _GEN_3517 : ~_GEN_3549 & _GEN_3517;
  wire        _GEN_3646 = _GEN_50 ? ~_GEN_3592 & _GEN_3518 : ~_GEN_3550 & _GEN_3518;
  wire        _GEN_3647 = _GEN_50 ? ~_GEN_3594 & _GEN_3519 : ~_GEN_3551 & _GEN_3519;
  wire        _GEN_3648 = _GEN_50 ? ~_GEN_3596 & _GEN_3520 : ~_GEN_3552 & _GEN_3520;
  wire        _GEN_3649 = _GEN_50 ? ~_GEN_3598 & _GEN_3521 : ~_GEN_3553 & _GEN_3521;
  wire        _GEN_3650 = _GEN_50 ? ~_GEN_3600 & _GEN_3522 : ~_GEN_3554 & _GEN_3522;
  wire        _GEN_3651 = _GEN_50 ? ~_GEN_3602 & _GEN_3523 : ~_GEN_3555 & _GEN_3523;
  wire        _GEN_3652 = _GEN_50 ? ~_GEN_3604 & _GEN_3524 : ~_GEN_3556 & _GEN_3524;
  wire        _GEN_3653 = _GEN_50 ? ~_GEN_3606 & _GEN_3525 : ~_GEN_3557 & _GEN_3525;
  wire        _GEN_3654 = _GEN_50 ? ~_GEN_3608 & _GEN_3526 : ~_GEN_3558 & _GEN_3526;
  wire        _GEN_3655 = _GEN_50 ? ~_GEN_3610 & _GEN_3527 : ~_GEN_3559 & _GEN_3527;
  wire        _GEN_3656 = _GEN_50 ? ~_GEN_3612 & _GEN_3528 : ~_GEN_3560 & _GEN_3528;
  wire        _GEN_3657 = _GEN_50 ? ~_GEN_3614 & _GEN_3529 : ~_GEN_3561 & _GEN_3529;
  wire        _GEN_3658 = _GEN_50 ? ~_GEN_3616 & _GEN_3530 : ~_GEN_3562 & _GEN_3530;
  wire        _GEN_3659 = _GEN_50 ? ~_GEN_3618 & _GEN_3531 : ~_GEN_3563 & _GEN_3531;
  wire        _GEN_3660 = _GEN_50 ? ~_GEN_3620 & _GEN_3532 : ~_GEN_3564 & _GEN_3532;
  wire        _GEN_3661 = _GEN_50 ? ~_GEN_3622 & _GEN_3533 : ~_GEN_3565 & _GEN_3533;
  wire        _GEN_3662 = _GEN_50 ? ~_GEN_3624 & _GEN_3534 : ~_GEN_3566 & _GEN_3534;
  wire        _GEN_3663 = _GEN_50 ? ~_GEN_3626 & _GEN_3535 : ~_GEN_3567 & _GEN_3535;
  wire        _GEN_3664 = _GEN_50 ? ~_GEN_3628 & _GEN_3536 : ~_GEN_3568 & _GEN_3536;
  wire        _GEN_3665 = _GEN_50 ? ~_GEN_3630 & _GEN_3537 : ~_GEN_3569 & _GEN_3537;
  wire        _GEN_3666 = _GEN_50 ? ~_GEN_3632 & _GEN_3538 : ~_GEN_3570 & _GEN_3538;
  wire        _GEN_3667 = _GEN_50 ? ~_GEN_3634 & _GEN_3539 : ~_GEN_3571 & _GEN_3539;
  wire        _GEN_3668 = _GEN_51 & _GEN_444;
  wire        _GEN_3669 = _GEN_51 & _GEN_446;
  wire        _GEN_3670 = _GEN_51 & _GEN_448;
  wire        _GEN_3671 = _GEN_51 & _GEN_450;
  wire        _GEN_3672 = _GEN_51 & _GEN_452;
  wire        _GEN_3673 = _GEN_51 & _GEN_454;
  wire        _GEN_3674 = _GEN_51 & _GEN_456;
  wire        _GEN_3675 = _GEN_51 & _GEN_458;
  wire        _GEN_3676 = _GEN_51 & _GEN_460;
  wire        _GEN_3677 = _GEN_51 & _GEN_462;
  wire        _GEN_3678 = _GEN_51 & _GEN_464;
  wire        _GEN_3679 = _GEN_51 & _GEN_466;
  wire        _GEN_3680 = _GEN_51 & _GEN_468;
  wire        _GEN_3681 = _GEN_51 & _GEN_470;
  wire        _GEN_3682 = _GEN_51 & _GEN_472;
  wire        _GEN_3683 = _GEN_51 & _GEN_474;
  wire        _GEN_3684 = _GEN_51 & _GEN_476;
  wire        _GEN_3685 = _GEN_51 & _GEN_478;
  wire        _GEN_3686 = _GEN_51 & _GEN_480;
  wire        _GEN_3687 = _GEN_51 & _GEN_482;
  wire        _GEN_3688 = _GEN_51 & _GEN_484;
  wire        _GEN_3689 = _GEN_51 & _GEN_486;
  wire        _GEN_3690 = _GEN_51 & _GEN_488;
  wire        _GEN_3691 = _GEN_51 & _GEN_490;
  wire        _GEN_3692 = _GEN_51 & _GEN_492;
  wire        _GEN_3693 = _GEN_51 & _GEN_494;
  wire        _GEN_3694 = _GEN_51 & _GEN_496;
  wire        _GEN_3695 = _GEN_51 & _GEN_498;
  wire        _GEN_3696 = _GEN_51 & _GEN_500;
  wire        _GEN_3697 = _GEN_51 & _GEN_502;
  wire        _GEN_3698 = _GEN_51 & _GEN_504;
  wire        _GEN_3699 = _GEN_51 & (&(io_wb_resps_2_bits_uop_rob_idx[6:2]));
  wire        _GEN_3700 = _GEN_507 | _GEN_3668;
  wire        _GEN_3701 = _GEN_52 ? ~_GEN_3700 & _GEN_3573 : ~_GEN_3668 & _GEN_3573;
  wire        _GEN_3702 = _GEN_510 | _GEN_3669;
  wire        _GEN_3703 = _GEN_52 ? ~_GEN_3702 & _GEN_3575 : ~_GEN_3669 & _GEN_3575;
  wire        _GEN_3704 = _GEN_513 | _GEN_3670;
  wire        _GEN_3705 = _GEN_52 ? ~_GEN_3704 & _GEN_3577 : ~_GEN_3670 & _GEN_3577;
  wire        _GEN_3706 = _GEN_516 | _GEN_3671;
  wire        _GEN_3707 = _GEN_52 ? ~_GEN_3706 & _GEN_3579 : ~_GEN_3671 & _GEN_3579;
  wire        _GEN_3708 = _GEN_519 | _GEN_3672;
  wire        _GEN_3709 = _GEN_52 ? ~_GEN_3708 & _GEN_3581 : ~_GEN_3672 & _GEN_3581;
  wire        _GEN_3710 = _GEN_522 | _GEN_3673;
  wire        _GEN_3711 = _GEN_52 ? ~_GEN_3710 & _GEN_3583 : ~_GEN_3673 & _GEN_3583;
  wire        _GEN_3712 = _GEN_525 | _GEN_3674;
  wire        _GEN_3713 = _GEN_52 ? ~_GEN_3712 & _GEN_3585 : ~_GEN_3674 & _GEN_3585;
  wire        _GEN_3714 = _GEN_528 | _GEN_3675;
  wire        _GEN_3715 = _GEN_52 ? ~_GEN_3714 & _GEN_3587 : ~_GEN_3675 & _GEN_3587;
  wire        _GEN_3716 = _GEN_531 | _GEN_3676;
  wire        _GEN_3717 = _GEN_52 ? ~_GEN_3716 & _GEN_3589 : ~_GEN_3676 & _GEN_3589;
  wire        _GEN_3718 = _GEN_534 | _GEN_3677;
  wire        _GEN_3719 = _GEN_52 ? ~_GEN_3718 & _GEN_3591 : ~_GEN_3677 & _GEN_3591;
  wire        _GEN_3720 = _GEN_537 | _GEN_3678;
  wire        _GEN_3721 = _GEN_52 ? ~_GEN_3720 & _GEN_3593 : ~_GEN_3678 & _GEN_3593;
  wire        _GEN_3722 = _GEN_540 | _GEN_3679;
  wire        _GEN_3723 = _GEN_52 ? ~_GEN_3722 & _GEN_3595 : ~_GEN_3679 & _GEN_3595;
  wire        _GEN_3724 = _GEN_543 | _GEN_3680;
  wire        _GEN_3725 = _GEN_52 ? ~_GEN_3724 & _GEN_3597 : ~_GEN_3680 & _GEN_3597;
  wire        _GEN_3726 = _GEN_546 | _GEN_3681;
  wire        _GEN_3727 = _GEN_52 ? ~_GEN_3726 & _GEN_3599 : ~_GEN_3681 & _GEN_3599;
  wire        _GEN_3728 = _GEN_549 | _GEN_3682;
  wire        _GEN_3729 = _GEN_52 ? ~_GEN_3728 & _GEN_3601 : ~_GEN_3682 & _GEN_3601;
  wire        _GEN_3730 = _GEN_552 | _GEN_3683;
  wire        _GEN_3731 = _GEN_52 ? ~_GEN_3730 & _GEN_3603 : ~_GEN_3683 & _GEN_3603;
  wire        _GEN_3732 = _GEN_555 | _GEN_3684;
  wire        _GEN_3733 = _GEN_52 ? ~_GEN_3732 & _GEN_3605 : ~_GEN_3684 & _GEN_3605;
  wire        _GEN_3734 = _GEN_558 | _GEN_3685;
  wire        _GEN_3735 = _GEN_52 ? ~_GEN_3734 & _GEN_3607 : ~_GEN_3685 & _GEN_3607;
  wire        _GEN_3736 = _GEN_561 | _GEN_3686;
  wire        _GEN_3737 = _GEN_52 ? ~_GEN_3736 & _GEN_3609 : ~_GEN_3686 & _GEN_3609;
  wire        _GEN_3738 = _GEN_564 | _GEN_3687;
  wire        _GEN_3739 = _GEN_52 ? ~_GEN_3738 & _GEN_3611 : ~_GEN_3687 & _GEN_3611;
  wire        _GEN_3740 = _GEN_567 | _GEN_3688;
  wire        _GEN_3741 = _GEN_52 ? ~_GEN_3740 & _GEN_3613 : ~_GEN_3688 & _GEN_3613;
  wire        _GEN_3742 = _GEN_570 | _GEN_3689;
  wire        _GEN_3743 = _GEN_52 ? ~_GEN_3742 & _GEN_3615 : ~_GEN_3689 & _GEN_3615;
  wire        _GEN_3744 = _GEN_573 | _GEN_3690;
  wire        _GEN_3745 = _GEN_52 ? ~_GEN_3744 & _GEN_3617 : ~_GEN_3690 & _GEN_3617;
  wire        _GEN_3746 = _GEN_576 | _GEN_3691;
  wire        _GEN_3747 = _GEN_52 ? ~_GEN_3746 & _GEN_3619 : ~_GEN_3691 & _GEN_3619;
  wire        _GEN_3748 = _GEN_579 | _GEN_3692;
  wire        _GEN_3749 = _GEN_52 ? ~_GEN_3748 & _GEN_3621 : ~_GEN_3692 & _GEN_3621;
  wire        _GEN_3750 = _GEN_582 | _GEN_3693;
  wire        _GEN_3751 = _GEN_52 ? ~_GEN_3750 & _GEN_3623 : ~_GEN_3693 & _GEN_3623;
  wire        _GEN_3752 = _GEN_585 | _GEN_3694;
  wire        _GEN_3753 = _GEN_52 ? ~_GEN_3752 & _GEN_3625 : ~_GEN_3694 & _GEN_3625;
  wire        _GEN_3754 = _GEN_588 | _GEN_3695;
  wire        _GEN_3755 = _GEN_52 ? ~_GEN_3754 & _GEN_3627 : ~_GEN_3695 & _GEN_3627;
  wire        _GEN_3756 = _GEN_591 | _GEN_3696;
  wire        _GEN_3757 = _GEN_52 ? ~_GEN_3756 & _GEN_3629 : ~_GEN_3696 & _GEN_3629;
  wire        _GEN_3758 = _GEN_594 | _GEN_3697;
  wire        _GEN_3759 = _GEN_52 ? ~_GEN_3758 & _GEN_3631 : ~_GEN_3697 & _GEN_3631;
  wire        _GEN_3760 = _GEN_597 | _GEN_3698;
  wire        _GEN_3761 = _GEN_52 ? ~_GEN_3760 & _GEN_3633 : ~_GEN_3698 & _GEN_3633;
  wire        _GEN_3762 = (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_3699;
  wire        _GEN_3763 = _GEN_52 ? ~_GEN_3762 & _GEN_3635 : ~_GEN_3699 & _GEN_3635;
  wire        _GEN_3764 = _GEN_52 ? ~_GEN_3700 & _GEN_3636 : ~_GEN_3668 & _GEN_3636;
  wire        _GEN_3765 = _GEN_52 ? ~_GEN_3702 & _GEN_3637 : ~_GEN_3669 & _GEN_3637;
  wire        _GEN_3766 = _GEN_52 ? ~_GEN_3704 & _GEN_3638 : ~_GEN_3670 & _GEN_3638;
  wire        _GEN_3767 = _GEN_52 ? ~_GEN_3706 & _GEN_3639 : ~_GEN_3671 & _GEN_3639;
  wire        _GEN_3768 = _GEN_52 ? ~_GEN_3708 & _GEN_3640 : ~_GEN_3672 & _GEN_3640;
  wire        _GEN_3769 = _GEN_52 ? ~_GEN_3710 & _GEN_3641 : ~_GEN_3673 & _GEN_3641;
  wire        _GEN_3770 = _GEN_52 ? ~_GEN_3712 & _GEN_3642 : ~_GEN_3674 & _GEN_3642;
  wire        _GEN_3771 = _GEN_52 ? ~_GEN_3714 & _GEN_3643 : ~_GEN_3675 & _GEN_3643;
  wire        _GEN_3772 = _GEN_52 ? ~_GEN_3716 & _GEN_3644 : ~_GEN_3676 & _GEN_3644;
  wire        _GEN_3773 = _GEN_52 ? ~_GEN_3718 & _GEN_3645 : ~_GEN_3677 & _GEN_3645;
  wire        _GEN_3774 = _GEN_52 ? ~_GEN_3720 & _GEN_3646 : ~_GEN_3678 & _GEN_3646;
  wire        _GEN_3775 = _GEN_52 ? ~_GEN_3722 & _GEN_3647 : ~_GEN_3679 & _GEN_3647;
  wire        _GEN_3776 = _GEN_52 ? ~_GEN_3724 & _GEN_3648 : ~_GEN_3680 & _GEN_3648;
  wire        _GEN_3777 = _GEN_52 ? ~_GEN_3726 & _GEN_3649 : ~_GEN_3681 & _GEN_3649;
  wire        _GEN_3778 = _GEN_52 ? ~_GEN_3728 & _GEN_3650 : ~_GEN_3682 & _GEN_3650;
  wire        _GEN_3779 = _GEN_52 ? ~_GEN_3730 & _GEN_3651 : ~_GEN_3683 & _GEN_3651;
  wire        _GEN_3780 = _GEN_52 ? ~_GEN_3732 & _GEN_3652 : ~_GEN_3684 & _GEN_3652;
  wire        _GEN_3781 = _GEN_52 ? ~_GEN_3734 & _GEN_3653 : ~_GEN_3685 & _GEN_3653;
  wire        _GEN_3782 = _GEN_52 ? ~_GEN_3736 & _GEN_3654 : ~_GEN_3686 & _GEN_3654;
  wire        _GEN_3783 = _GEN_52 ? ~_GEN_3738 & _GEN_3655 : ~_GEN_3687 & _GEN_3655;
  wire        _GEN_3784 = _GEN_52 ? ~_GEN_3740 & _GEN_3656 : ~_GEN_3688 & _GEN_3656;
  wire        _GEN_3785 = _GEN_52 ? ~_GEN_3742 & _GEN_3657 : ~_GEN_3689 & _GEN_3657;
  wire        _GEN_3786 = _GEN_52 ? ~_GEN_3744 & _GEN_3658 : ~_GEN_3690 & _GEN_3658;
  wire        _GEN_3787 = _GEN_52 ? ~_GEN_3746 & _GEN_3659 : ~_GEN_3691 & _GEN_3659;
  wire        _GEN_3788 = _GEN_52 ? ~_GEN_3748 & _GEN_3660 : ~_GEN_3692 & _GEN_3660;
  wire        _GEN_3789 = _GEN_52 ? ~_GEN_3750 & _GEN_3661 : ~_GEN_3693 & _GEN_3661;
  wire        _GEN_3790 = _GEN_52 ? ~_GEN_3752 & _GEN_3662 : ~_GEN_3694 & _GEN_3662;
  wire        _GEN_3791 = _GEN_52 ? ~_GEN_3754 & _GEN_3663 : ~_GEN_3695 & _GEN_3663;
  wire        _GEN_3792 = _GEN_52 ? ~_GEN_3756 & _GEN_3664 : ~_GEN_3696 & _GEN_3664;
  wire        _GEN_3793 = _GEN_52 ? ~_GEN_3758 & _GEN_3665 : ~_GEN_3697 & _GEN_3665;
  wire        _GEN_3794 = _GEN_52 ? ~_GEN_3760 & _GEN_3666 : ~_GEN_3698 & _GEN_3666;
  wire        _GEN_3795 = _GEN_52 ? ~_GEN_3762 & _GEN_3667 : ~_GEN_3699 & _GEN_3667;
  wire        _GEN_3796 = _GEN_53 & _GEN_634;
  wire        _GEN_3797 = _GEN_53 & _GEN_636;
  wire        _GEN_3798 = _GEN_53 & _GEN_638;
  wire        _GEN_3799 = _GEN_53 & _GEN_640;
  wire        _GEN_3800 = _GEN_53 & _GEN_642;
  wire        _GEN_3801 = _GEN_53 & _GEN_644;
  wire        _GEN_3802 = _GEN_53 & _GEN_646;
  wire        _GEN_3803 = _GEN_53 & _GEN_648;
  wire        _GEN_3804 = _GEN_53 & _GEN_650;
  wire        _GEN_3805 = _GEN_53 & _GEN_652;
  wire        _GEN_3806 = _GEN_53 & _GEN_654;
  wire        _GEN_3807 = _GEN_53 & _GEN_656;
  wire        _GEN_3808 = _GEN_53 & _GEN_658;
  wire        _GEN_3809 = _GEN_53 & _GEN_660;
  wire        _GEN_3810 = _GEN_53 & _GEN_662;
  wire        _GEN_3811 = _GEN_53 & _GEN_664;
  wire        _GEN_3812 = _GEN_53 & _GEN_666;
  wire        _GEN_3813 = _GEN_53 & _GEN_668;
  wire        _GEN_3814 = _GEN_53 & _GEN_670;
  wire        _GEN_3815 = _GEN_53 & _GEN_672;
  wire        _GEN_3816 = _GEN_53 & _GEN_674;
  wire        _GEN_3817 = _GEN_53 & _GEN_676;
  wire        _GEN_3818 = _GEN_53 & _GEN_678;
  wire        _GEN_3819 = _GEN_53 & _GEN_680;
  wire        _GEN_3820 = _GEN_53 & _GEN_682;
  wire        _GEN_3821 = _GEN_53 & _GEN_684;
  wire        _GEN_3822 = _GEN_53 & _GEN_686;
  wire        _GEN_3823 = _GEN_53 & _GEN_688;
  wire        _GEN_3824 = _GEN_53 & _GEN_690;
  wire        _GEN_3825 = _GEN_53 & _GEN_692;
  wire        _GEN_3826 = _GEN_53 & _GEN_694;
  wire        _GEN_3827 = _GEN_53 & (&(io_wb_resps_4_bits_uop_rob_idx[6:2]));
  wire        _GEN_3828 = _GEN_697 | _GEN_3796;
  wire        _GEN_3829 = _GEN_54 ? ~_GEN_3828 & _GEN_3701 : ~_GEN_3796 & _GEN_3701;
  wire        _GEN_3830 = _GEN_700 | _GEN_3797;
  wire        _GEN_3831 = _GEN_54 ? ~_GEN_3830 & _GEN_3703 : ~_GEN_3797 & _GEN_3703;
  wire        _GEN_3832 = _GEN_703 | _GEN_3798;
  wire        _GEN_3833 = _GEN_54 ? ~_GEN_3832 & _GEN_3705 : ~_GEN_3798 & _GEN_3705;
  wire        _GEN_3834 = _GEN_706 | _GEN_3799;
  wire        _GEN_3835 = _GEN_54 ? ~_GEN_3834 & _GEN_3707 : ~_GEN_3799 & _GEN_3707;
  wire        _GEN_3836 = _GEN_709 | _GEN_3800;
  wire        _GEN_3837 = _GEN_54 ? ~_GEN_3836 & _GEN_3709 : ~_GEN_3800 & _GEN_3709;
  wire        _GEN_3838 = _GEN_712 | _GEN_3801;
  wire        _GEN_3839 = _GEN_54 ? ~_GEN_3838 & _GEN_3711 : ~_GEN_3801 & _GEN_3711;
  wire        _GEN_3840 = _GEN_715 | _GEN_3802;
  wire        _GEN_3841 = _GEN_54 ? ~_GEN_3840 & _GEN_3713 : ~_GEN_3802 & _GEN_3713;
  wire        _GEN_3842 = _GEN_718 | _GEN_3803;
  wire        _GEN_3843 = _GEN_54 ? ~_GEN_3842 & _GEN_3715 : ~_GEN_3803 & _GEN_3715;
  wire        _GEN_3844 = _GEN_721 | _GEN_3804;
  wire        _GEN_3845 = _GEN_54 ? ~_GEN_3844 & _GEN_3717 : ~_GEN_3804 & _GEN_3717;
  wire        _GEN_3846 = _GEN_724 | _GEN_3805;
  wire        _GEN_3847 = _GEN_54 ? ~_GEN_3846 & _GEN_3719 : ~_GEN_3805 & _GEN_3719;
  wire        _GEN_3848 = _GEN_727 | _GEN_3806;
  wire        _GEN_3849 = _GEN_54 ? ~_GEN_3848 & _GEN_3721 : ~_GEN_3806 & _GEN_3721;
  wire        _GEN_3850 = _GEN_730 | _GEN_3807;
  wire        _GEN_3851 = _GEN_54 ? ~_GEN_3850 & _GEN_3723 : ~_GEN_3807 & _GEN_3723;
  wire        _GEN_3852 = _GEN_733 | _GEN_3808;
  wire        _GEN_3853 = _GEN_54 ? ~_GEN_3852 & _GEN_3725 : ~_GEN_3808 & _GEN_3725;
  wire        _GEN_3854 = _GEN_736 | _GEN_3809;
  wire        _GEN_3855 = _GEN_54 ? ~_GEN_3854 & _GEN_3727 : ~_GEN_3809 & _GEN_3727;
  wire        _GEN_3856 = _GEN_739 | _GEN_3810;
  wire        _GEN_3857 = _GEN_54 ? ~_GEN_3856 & _GEN_3729 : ~_GEN_3810 & _GEN_3729;
  wire        _GEN_3858 = _GEN_742 | _GEN_3811;
  wire        _GEN_3859 = _GEN_54 ? ~_GEN_3858 & _GEN_3731 : ~_GEN_3811 & _GEN_3731;
  wire        _GEN_3860 = _GEN_745 | _GEN_3812;
  wire        _GEN_3861 = _GEN_54 ? ~_GEN_3860 & _GEN_3733 : ~_GEN_3812 & _GEN_3733;
  wire        _GEN_3862 = _GEN_748 | _GEN_3813;
  wire        _GEN_3863 = _GEN_54 ? ~_GEN_3862 & _GEN_3735 : ~_GEN_3813 & _GEN_3735;
  wire        _GEN_3864 = _GEN_751 | _GEN_3814;
  wire        _GEN_3865 = _GEN_54 ? ~_GEN_3864 & _GEN_3737 : ~_GEN_3814 & _GEN_3737;
  wire        _GEN_3866 = _GEN_754 | _GEN_3815;
  wire        _GEN_3867 = _GEN_54 ? ~_GEN_3866 & _GEN_3739 : ~_GEN_3815 & _GEN_3739;
  wire        _GEN_3868 = _GEN_757 | _GEN_3816;
  wire        _GEN_3869 = _GEN_54 ? ~_GEN_3868 & _GEN_3741 : ~_GEN_3816 & _GEN_3741;
  wire        _GEN_3870 = _GEN_760 | _GEN_3817;
  wire        _GEN_3871 = _GEN_54 ? ~_GEN_3870 & _GEN_3743 : ~_GEN_3817 & _GEN_3743;
  wire        _GEN_3872 = _GEN_763 | _GEN_3818;
  wire        _GEN_3873 = _GEN_54 ? ~_GEN_3872 & _GEN_3745 : ~_GEN_3818 & _GEN_3745;
  wire        _GEN_3874 = _GEN_766 | _GEN_3819;
  wire        _GEN_3875 = _GEN_54 ? ~_GEN_3874 & _GEN_3747 : ~_GEN_3819 & _GEN_3747;
  wire        _GEN_3876 = _GEN_769 | _GEN_3820;
  wire        _GEN_3877 = _GEN_54 ? ~_GEN_3876 & _GEN_3749 : ~_GEN_3820 & _GEN_3749;
  wire        _GEN_3878 = _GEN_772 | _GEN_3821;
  wire        _GEN_3879 = _GEN_54 ? ~_GEN_3878 & _GEN_3751 : ~_GEN_3821 & _GEN_3751;
  wire        _GEN_3880 = _GEN_775 | _GEN_3822;
  wire        _GEN_3881 = _GEN_54 ? ~_GEN_3880 & _GEN_3753 : ~_GEN_3822 & _GEN_3753;
  wire        _GEN_3882 = _GEN_778 | _GEN_3823;
  wire        _GEN_3883 = _GEN_54 ? ~_GEN_3882 & _GEN_3755 : ~_GEN_3823 & _GEN_3755;
  wire        _GEN_3884 = _GEN_781 | _GEN_3824;
  wire        _GEN_3885 = _GEN_54 ? ~_GEN_3884 & _GEN_3757 : ~_GEN_3824 & _GEN_3757;
  wire        _GEN_3886 = _GEN_784 | _GEN_3825;
  wire        _GEN_3887 = _GEN_54 ? ~_GEN_3886 & _GEN_3759 : ~_GEN_3825 & _GEN_3759;
  wire        _GEN_3888 = _GEN_787 | _GEN_3826;
  wire        _GEN_3889 = _GEN_54 ? ~_GEN_3888 & _GEN_3761 : ~_GEN_3826 & _GEN_3761;
  wire        _GEN_3890 = (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_3827;
  wire        _GEN_3891 = _GEN_54 ? ~_GEN_3890 & _GEN_3763 : ~_GEN_3827 & _GEN_3763;
  wire        _GEN_3892 = _GEN_54 ? ~_GEN_3828 & _GEN_3764 : ~_GEN_3796 & _GEN_3764;
  wire        _GEN_3893 = _GEN_54 ? ~_GEN_3830 & _GEN_3765 : ~_GEN_3797 & _GEN_3765;
  wire        _GEN_3894 = _GEN_54 ? ~_GEN_3832 & _GEN_3766 : ~_GEN_3798 & _GEN_3766;
  wire        _GEN_3895 = _GEN_54 ? ~_GEN_3834 & _GEN_3767 : ~_GEN_3799 & _GEN_3767;
  wire        _GEN_3896 = _GEN_54 ? ~_GEN_3836 & _GEN_3768 : ~_GEN_3800 & _GEN_3768;
  wire        _GEN_3897 = _GEN_54 ? ~_GEN_3838 & _GEN_3769 : ~_GEN_3801 & _GEN_3769;
  wire        _GEN_3898 = _GEN_54 ? ~_GEN_3840 & _GEN_3770 : ~_GEN_3802 & _GEN_3770;
  wire        _GEN_3899 = _GEN_54 ? ~_GEN_3842 & _GEN_3771 : ~_GEN_3803 & _GEN_3771;
  wire        _GEN_3900 = _GEN_54 ? ~_GEN_3844 & _GEN_3772 : ~_GEN_3804 & _GEN_3772;
  wire        _GEN_3901 = _GEN_54 ? ~_GEN_3846 & _GEN_3773 : ~_GEN_3805 & _GEN_3773;
  wire        _GEN_3902 = _GEN_54 ? ~_GEN_3848 & _GEN_3774 : ~_GEN_3806 & _GEN_3774;
  wire        _GEN_3903 = _GEN_54 ? ~_GEN_3850 & _GEN_3775 : ~_GEN_3807 & _GEN_3775;
  wire        _GEN_3904 = _GEN_54 ? ~_GEN_3852 & _GEN_3776 : ~_GEN_3808 & _GEN_3776;
  wire        _GEN_3905 = _GEN_54 ? ~_GEN_3854 & _GEN_3777 : ~_GEN_3809 & _GEN_3777;
  wire        _GEN_3906 = _GEN_54 ? ~_GEN_3856 & _GEN_3778 : ~_GEN_3810 & _GEN_3778;
  wire        _GEN_3907 = _GEN_54 ? ~_GEN_3858 & _GEN_3779 : ~_GEN_3811 & _GEN_3779;
  wire        _GEN_3908 = _GEN_54 ? ~_GEN_3860 & _GEN_3780 : ~_GEN_3812 & _GEN_3780;
  wire        _GEN_3909 = _GEN_54 ? ~_GEN_3862 & _GEN_3781 : ~_GEN_3813 & _GEN_3781;
  wire        _GEN_3910 = _GEN_54 ? ~_GEN_3864 & _GEN_3782 : ~_GEN_3814 & _GEN_3782;
  wire        _GEN_3911 = _GEN_54 ? ~_GEN_3866 & _GEN_3783 : ~_GEN_3815 & _GEN_3783;
  wire        _GEN_3912 = _GEN_54 ? ~_GEN_3868 & _GEN_3784 : ~_GEN_3816 & _GEN_3784;
  wire        _GEN_3913 = _GEN_54 ? ~_GEN_3870 & _GEN_3785 : ~_GEN_3817 & _GEN_3785;
  wire        _GEN_3914 = _GEN_54 ? ~_GEN_3872 & _GEN_3786 : ~_GEN_3818 & _GEN_3786;
  wire        _GEN_3915 = _GEN_54 ? ~_GEN_3874 & _GEN_3787 : ~_GEN_3819 & _GEN_3787;
  wire        _GEN_3916 = _GEN_54 ? ~_GEN_3876 & _GEN_3788 : ~_GEN_3820 & _GEN_3788;
  wire        _GEN_3917 = _GEN_54 ? ~_GEN_3878 & _GEN_3789 : ~_GEN_3821 & _GEN_3789;
  wire        _GEN_3918 = _GEN_54 ? ~_GEN_3880 & _GEN_3790 : ~_GEN_3822 & _GEN_3790;
  wire        _GEN_3919 = _GEN_54 ? ~_GEN_3882 & _GEN_3791 : ~_GEN_3823 & _GEN_3791;
  wire        _GEN_3920 = _GEN_54 ? ~_GEN_3884 & _GEN_3792 : ~_GEN_3824 & _GEN_3792;
  wire        _GEN_3921 = _GEN_54 ? ~_GEN_3886 & _GEN_3793 : ~_GEN_3825 & _GEN_3793;
  wire        _GEN_3922 = _GEN_54 ? ~_GEN_3888 & _GEN_3794 : ~_GEN_3826 & _GEN_3794;
  wire        _GEN_3923 = _GEN_54 ? ~_GEN_3890 & _GEN_3795 : ~_GEN_3827 & _GEN_3795;
  wire        _GEN_3924 = _GEN_55 & _GEN_824;
  wire        _GEN_3925 = _GEN_55 & _GEN_826;
  wire        _GEN_3926 = _GEN_55 & _GEN_828;
  wire        _GEN_3927 = _GEN_55 & _GEN_830;
  wire        _GEN_3928 = _GEN_55 & _GEN_832;
  wire        _GEN_3929 = _GEN_55 & _GEN_834;
  wire        _GEN_3930 = _GEN_55 & _GEN_836;
  wire        _GEN_3931 = _GEN_55 & _GEN_838;
  wire        _GEN_3932 = _GEN_55 & _GEN_840;
  wire        _GEN_3933 = _GEN_55 & _GEN_842;
  wire        _GEN_3934 = _GEN_55 & _GEN_844;
  wire        _GEN_3935 = _GEN_55 & _GEN_846;
  wire        _GEN_3936 = _GEN_55 & _GEN_848;
  wire        _GEN_3937 = _GEN_55 & _GEN_850;
  wire        _GEN_3938 = _GEN_55 & _GEN_852;
  wire        _GEN_3939 = _GEN_55 & _GEN_854;
  wire        _GEN_3940 = _GEN_55 & _GEN_856;
  wire        _GEN_3941 = _GEN_55 & _GEN_858;
  wire        _GEN_3942 = _GEN_55 & _GEN_860;
  wire        _GEN_3943 = _GEN_55 & _GEN_862;
  wire        _GEN_3944 = _GEN_55 & _GEN_864;
  wire        _GEN_3945 = _GEN_55 & _GEN_866;
  wire        _GEN_3946 = _GEN_55 & _GEN_868;
  wire        _GEN_3947 = _GEN_55 & _GEN_870;
  wire        _GEN_3948 = _GEN_55 & _GEN_872;
  wire        _GEN_3949 = _GEN_55 & _GEN_874;
  wire        _GEN_3950 = _GEN_55 & _GEN_876;
  wire        _GEN_3951 = _GEN_55 & _GEN_878;
  wire        _GEN_3952 = _GEN_55 & _GEN_880;
  wire        _GEN_3953 = _GEN_55 & _GEN_882;
  wire        _GEN_3954 = _GEN_55 & _GEN_884;
  wire        _GEN_3955 = _GEN_55 & (&(io_wb_resps_6_bits_uop_rob_idx[6:2]));
  wire        _GEN_3956 = _GEN_887 | _GEN_3924;
  wire        _GEN_3957 = _GEN_56 ? ~_GEN_3956 & _GEN_3829 : ~_GEN_3924 & _GEN_3829;
  wire        _GEN_3958 = _GEN_890 | _GEN_3925;
  wire        _GEN_3959 = _GEN_56 ? ~_GEN_3958 & _GEN_3831 : ~_GEN_3925 & _GEN_3831;
  wire        _GEN_3960 = _GEN_893 | _GEN_3926;
  wire        _GEN_3961 = _GEN_56 ? ~_GEN_3960 & _GEN_3833 : ~_GEN_3926 & _GEN_3833;
  wire        _GEN_3962 = _GEN_896 | _GEN_3927;
  wire        _GEN_3963 = _GEN_56 ? ~_GEN_3962 & _GEN_3835 : ~_GEN_3927 & _GEN_3835;
  wire        _GEN_3964 = _GEN_899 | _GEN_3928;
  wire        _GEN_3965 = _GEN_56 ? ~_GEN_3964 & _GEN_3837 : ~_GEN_3928 & _GEN_3837;
  wire        _GEN_3966 = _GEN_902 | _GEN_3929;
  wire        _GEN_3967 = _GEN_56 ? ~_GEN_3966 & _GEN_3839 : ~_GEN_3929 & _GEN_3839;
  wire        _GEN_3968 = _GEN_905 | _GEN_3930;
  wire        _GEN_3969 = _GEN_56 ? ~_GEN_3968 & _GEN_3841 : ~_GEN_3930 & _GEN_3841;
  wire        _GEN_3970 = _GEN_908 | _GEN_3931;
  wire        _GEN_3971 = _GEN_56 ? ~_GEN_3970 & _GEN_3843 : ~_GEN_3931 & _GEN_3843;
  wire        _GEN_3972 = _GEN_911 | _GEN_3932;
  wire        _GEN_3973 = _GEN_56 ? ~_GEN_3972 & _GEN_3845 : ~_GEN_3932 & _GEN_3845;
  wire        _GEN_3974 = _GEN_914 | _GEN_3933;
  wire        _GEN_3975 = _GEN_56 ? ~_GEN_3974 & _GEN_3847 : ~_GEN_3933 & _GEN_3847;
  wire        _GEN_3976 = _GEN_917 | _GEN_3934;
  wire        _GEN_3977 = _GEN_56 ? ~_GEN_3976 & _GEN_3849 : ~_GEN_3934 & _GEN_3849;
  wire        _GEN_3978 = _GEN_920 | _GEN_3935;
  wire        _GEN_3979 = _GEN_56 ? ~_GEN_3978 & _GEN_3851 : ~_GEN_3935 & _GEN_3851;
  wire        _GEN_3980 = _GEN_923 | _GEN_3936;
  wire        _GEN_3981 = _GEN_56 ? ~_GEN_3980 & _GEN_3853 : ~_GEN_3936 & _GEN_3853;
  wire        _GEN_3982 = _GEN_926 | _GEN_3937;
  wire        _GEN_3983 = _GEN_56 ? ~_GEN_3982 & _GEN_3855 : ~_GEN_3937 & _GEN_3855;
  wire        _GEN_3984 = _GEN_929 | _GEN_3938;
  wire        _GEN_3985 = _GEN_56 ? ~_GEN_3984 & _GEN_3857 : ~_GEN_3938 & _GEN_3857;
  wire        _GEN_3986 = _GEN_932 | _GEN_3939;
  wire        _GEN_3987 = _GEN_56 ? ~_GEN_3986 & _GEN_3859 : ~_GEN_3939 & _GEN_3859;
  wire        _GEN_3988 = _GEN_935 | _GEN_3940;
  wire        _GEN_3989 = _GEN_56 ? ~_GEN_3988 & _GEN_3861 : ~_GEN_3940 & _GEN_3861;
  wire        _GEN_3990 = _GEN_938 | _GEN_3941;
  wire        _GEN_3991 = _GEN_56 ? ~_GEN_3990 & _GEN_3863 : ~_GEN_3941 & _GEN_3863;
  wire        _GEN_3992 = _GEN_941 | _GEN_3942;
  wire        _GEN_3993 = _GEN_56 ? ~_GEN_3992 & _GEN_3865 : ~_GEN_3942 & _GEN_3865;
  wire        _GEN_3994 = _GEN_944 | _GEN_3943;
  wire        _GEN_3995 = _GEN_56 ? ~_GEN_3994 & _GEN_3867 : ~_GEN_3943 & _GEN_3867;
  wire        _GEN_3996 = _GEN_947 | _GEN_3944;
  wire        _GEN_3997 = _GEN_56 ? ~_GEN_3996 & _GEN_3869 : ~_GEN_3944 & _GEN_3869;
  wire        _GEN_3998 = _GEN_950 | _GEN_3945;
  wire        _GEN_3999 = _GEN_56 ? ~_GEN_3998 & _GEN_3871 : ~_GEN_3945 & _GEN_3871;
  wire        _GEN_4000 = _GEN_953 | _GEN_3946;
  wire        _GEN_4001 = _GEN_56 ? ~_GEN_4000 & _GEN_3873 : ~_GEN_3946 & _GEN_3873;
  wire        _GEN_4002 = _GEN_956 | _GEN_3947;
  wire        _GEN_4003 = _GEN_56 ? ~_GEN_4002 & _GEN_3875 : ~_GEN_3947 & _GEN_3875;
  wire        _GEN_4004 = _GEN_959 | _GEN_3948;
  wire        _GEN_4005 = _GEN_56 ? ~_GEN_4004 & _GEN_3877 : ~_GEN_3948 & _GEN_3877;
  wire        _GEN_4006 = _GEN_962 | _GEN_3949;
  wire        _GEN_4007 = _GEN_56 ? ~_GEN_4006 & _GEN_3879 : ~_GEN_3949 & _GEN_3879;
  wire        _GEN_4008 = _GEN_965 | _GEN_3950;
  wire        _GEN_4009 = _GEN_56 ? ~_GEN_4008 & _GEN_3881 : ~_GEN_3950 & _GEN_3881;
  wire        _GEN_4010 = _GEN_968 | _GEN_3951;
  wire        _GEN_4011 = _GEN_56 ? ~_GEN_4010 & _GEN_3883 : ~_GEN_3951 & _GEN_3883;
  wire        _GEN_4012 = _GEN_971 | _GEN_3952;
  wire        _GEN_4013 = _GEN_56 ? ~_GEN_4012 & _GEN_3885 : ~_GEN_3952 & _GEN_3885;
  wire        _GEN_4014 = _GEN_974 | _GEN_3953;
  wire        _GEN_4015 = _GEN_56 ? ~_GEN_4014 & _GEN_3887 : ~_GEN_3953 & _GEN_3887;
  wire        _GEN_4016 = _GEN_977 | _GEN_3954;
  wire        _GEN_4017 = _GEN_56 ? ~_GEN_4016 & _GEN_3889 : ~_GEN_3954 & _GEN_3889;
  wire        _GEN_4018 = (&(io_wb_resps_7_bits_uop_rob_idx[6:2])) | _GEN_3955;
  wire        _GEN_4019 = _GEN_56 ? ~_GEN_4018 & _GEN_3891 : ~_GEN_3955 & _GEN_3891;
  wire        _GEN_4020 = _GEN_56 ? ~_GEN_3956 & _GEN_3892 : ~_GEN_3924 & _GEN_3892;
  wire        _GEN_4021 = _GEN_56 ? ~_GEN_3958 & _GEN_3893 : ~_GEN_3925 & _GEN_3893;
  wire        _GEN_4022 = _GEN_56 ? ~_GEN_3960 & _GEN_3894 : ~_GEN_3926 & _GEN_3894;
  wire        _GEN_4023 = _GEN_56 ? ~_GEN_3962 & _GEN_3895 : ~_GEN_3927 & _GEN_3895;
  wire        _GEN_4024 = _GEN_56 ? ~_GEN_3964 & _GEN_3896 : ~_GEN_3928 & _GEN_3896;
  wire        _GEN_4025 = _GEN_56 ? ~_GEN_3966 & _GEN_3897 : ~_GEN_3929 & _GEN_3897;
  wire        _GEN_4026 = _GEN_56 ? ~_GEN_3968 & _GEN_3898 : ~_GEN_3930 & _GEN_3898;
  wire        _GEN_4027 = _GEN_56 ? ~_GEN_3970 & _GEN_3899 : ~_GEN_3931 & _GEN_3899;
  wire        _GEN_4028 = _GEN_56 ? ~_GEN_3972 & _GEN_3900 : ~_GEN_3932 & _GEN_3900;
  wire        _GEN_4029 = _GEN_56 ? ~_GEN_3974 & _GEN_3901 : ~_GEN_3933 & _GEN_3901;
  wire        _GEN_4030 = _GEN_56 ? ~_GEN_3976 & _GEN_3902 : ~_GEN_3934 & _GEN_3902;
  wire        _GEN_4031 = _GEN_56 ? ~_GEN_3978 & _GEN_3903 : ~_GEN_3935 & _GEN_3903;
  wire        _GEN_4032 = _GEN_56 ? ~_GEN_3980 & _GEN_3904 : ~_GEN_3936 & _GEN_3904;
  wire        _GEN_4033 = _GEN_56 ? ~_GEN_3982 & _GEN_3905 : ~_GEN_3937 & _GEN_3905;
  wire        _GEN_4034 = _GEN_56 ? ~_GEN_3984 & _GEN_3906 : ~_GEN_3938 & _GEN_3906;
  wire        _GEN_4035 = _GEN_56 ? ~_GEN_3986 & _GEN_3907 : ~_GEN_3939 & _GEN_3907;
  wire        _GEN_4036 = _GEN_56 ? ~_GEN_3988 & _GEN_3908 : ~_GEN_3940 & _GEN_3908;
  wire        _GEN_4037 = _GEN_56 ? ~_GEN_3990 & _GEN_3909 : ~_GEN_3941 & _GEN_3909;
  wire        _GEN_4038 = _GEN_56 ? ~_GEN_3992 & _GEN_3910 : ~_GEN_3942 & _GEN_3910;
  wire        _GEN_4039 = _GEN_56 ? ~_GEN_3994 & _GEN_3911 : ~_GEN_3943 & _GEN_3911;
  wire        _GEN_4040 = _GEN_56 ? ~_GEN_3996 & _GEN_3912 : ~_GEN_3944 & _GEN_3912;
  wire        _GEN_4041 = _GEN_56 ? ~_GEN_3998 & _GEN_3913 : ~_GEN_3945 & _GEN_3913;
  wire        _GEN_4042 = _GEN_56 ? ~_GEN_4000 & _GEN_3914 : ~_GEN_3946 & _GEN_3914;
  wire        _GEN_4043 = _GEN_56 ? ~_GEN_4002 & _GEN_3915 : ~_GEN_3947 & _GEN_3915;
  wire        _GEN_4044 = _GEN_56 ? ~_GEN_4004 & _GEN_3916 : ~_GEN_3948 & _GEN_3916;
  wire        _GEN_4045 = _GEN_56 ? ~_GEN_4006 & _GEN_3917 : ~_GEN_3949 & _GEN_3917;
  wire        _GEN_4046 = _GEN_56 ? ~_GEN_4008 & _GEN_3918 : ~_GEN_3950 & _GEN_3918;
  wire        _GEN_4047 = _GEN_56 ? ~_GEN_4010 & _GEN_3919 : ~_GEN_3951 & _GEN_3919;
  wire        _GEN_4048 = _GEN_56 ? ~_GEN_4012 & _GEN_3920 : ~_GEN_3952 & _GEN_3920;
  wire        _GEN_4049 = _GEN_56 ? ~_GEN_4014 & _GEN_3921 : ~_GEN_3953 & _GEN_3921;
  wire        _GEN_4050 = _GEN_56 ? ~_GEN_4016 & _GEN_3922 : ~_GEN_3954 & _GEN_3922;
  wire        _GEN_4051 = _GEN_56 ? ~_GEN_4018 & _GEN_3923 : ~_GEN_3955 & _GEN_3923;
  wire        _GEN_4052 = _GEN_57 & _GEN_1014;
  wire        _GEN_4053 = _GEN_57 & _GEN_1016;
  wire        _GEN_4054 = _GEN_57 & _GEN_1018;
  wire        _GEN_4055 = _GEN_57 & _GEN_1020;
  wire        _GEN_4056 = _GEN_57 & _GEN_1022;
  wire        _GEN_4057 = _GEN_57 & _GEN_1024;
  wire        _GEN_4058 = _GEN_57 & _GEN_1026;
  wire        _GEN_4059 = _GEN_57 & _GEN_1028;
  wire        _GEN_4060 = _GEN_57 & _GEN_1030;
  wire        _GEN_4061 = _GEN_57 & _GEN_1032;
  wire        _GEN_4062 = _GEN_57 & _GEN_1034;
  wire        _GEN_4063 = _GEN_57 & _GEN_1036;
  wire        _GEN_4064 = _GEN_57 & _GEN_1038;
  wire        _GEN_4065 = _GEN_57 & _GEN_1040;
  wire        _GEN_4066 = _GEN_57 & _GEN_1042;
  wire        _GEN_4067 = _GEN_57 & _GEN_1044;
  wire        _GEN_4068 = _GEN_57 & _GEN_1046;
  wire        _GEN_4069 = _GEN_57 & _GEN_1048;
  wire        _GEN_4070 = _GEN_57 & _GEN_1050;
  wire        _GEN_4071 = _GEN_57 & _GEN_1052;
  wire        _GEN_4072 = _GEN_57 & _GEN_1054;
  wire        _GEN_4073 = _GEN_57 & _GEN_1056;
  wire        _GEN_4074 = _GEN_57 & _GEN_1058;
  wire        _GEN_4075 = _GEN_57 & _GEN_1060;
  wire        _GEN_4076 = _GEN_57 & _GEN_1062;
  wire        _GEN_4077 = _GEN_57 & _GEN_1064;
  wire        _GEN_4078 = _GEN_57 & _GEN_1066;
  wire        _GEN_4079 = _GEN_57 & _GEN_1068;
  wire        _GEN_4080 = _GEN_57 & _GEN_1070;
  wire        _GEN_4081 = _GEN_57 & _GEN_1072;
  wire        _GEN_4082 = _GEN_57 & _GEN_1074;
  wire        _GEN_4083 = _GEN_57 & (&(io_wb_resps_8_bits_uop_rob_idx[6:2]));
  wire        _GEN_4084 = _GEN_1077 | _GEN_4052;
  wire        _GEN_4085 = _GEN_58 ? ~_GEN_4084 & _GEN_3957 : ~_GEN_4052 & _GEN_3957;
  wire        _GEN_4086 = _GEN_1080 | _GEN_4053;
  wire        _GEN_4087 = _GEN_58 ? ~_GEN_4086 & _GEN_3959 : ~_GEN_4053 & _GEN_3959;
  wire        _GEN_4088 = _GEN_1083 | _GEN_4054;
  wire        _GEN_4089 = _GEN_58 ? ~_GEN_4088 & _GEN_3961 : ~_GEN_4054 & _GEN_3961;
  wire        _GEN_4090 = _GEN_1086 | _GEN_4055;
  wire        _GEN_4091 = _GEN_58 ? ~_GEN_4090 & _GEN_3963 : ~_GEN_4055 & _GEN_3963;
  wire        _GEN_4092 = _GEN_1089 | _GEN_4056;
  wire        _GEN_4093 = _GEN_58 ? ~_GEN_4092 & _GEN_3965 : ~_GEN_4056 & _GEN_3965;
  wire        _GEN_4094 = _GEN_1092 | _GEN_4057;
  wire        _GEN_4095 = _GEN_58 ? ~_GEN_4094 & _GEN_3967 : ~_GEN_4057 & _GEN_3967;
  wire        _GEN_4096 = _GEN_1095 | _GEN_4058;
  wire        _GEN_4097 = _GEN_58 ? ~_GEN_4096 & _GEN_3969 : ~_GEN_4058 & _GEN_3969;
  wire        _GEN_4098 = _GEN_1098 | _GEN_4059;
  wire        _GEN_4099 = _GEN_58 ? ~_GEN_4098 & _GEN_3971 : ~_GEN_4059 & _GEN_3971;
  wire        _GEN_4100 = _GEN_1101 | _GEN_4060;
  wire        _GEN_4101 = _GEN_58 ? ~_GEN_4100 & _GEN_3973 : ~_GEN_4060 & _GEN_3973;
  wire        _GEN_4102 = _GEN_1104 | _GEN_4061;
  wire        _GEN_4103 = _GEN_58 ? ~_GEN_4102 & _GEN_3975 : ~_GEN_4061 & _GEN_3975;
  wire        _GEN_4104 = _GEN_1107 | _GEN_4062;
  wire        _GEN_4105 = _GEN_58 ? ~_GEN_4104 & _GEN_3977 : ~_GEN_4062 & _GEN_3977;
  wire        _GEN_4106 = _GEN_1110 | _GEN_4063;
  wire        _GEN_4107 = _GEN_58 ? ~_GEN_4106 & _GEN_3979 : ~_GEN_4063 & _GEN_3979;
  wire        _GEN_4108 = _GEN_1113 | _GEN_4064;
  wire        _GEN_4109 = _GEN_58 ? ~_GEN_4108 & _GEN_3981 : ~_GEN_4064 & _GEN_3981;
  wire        _GEN_4110 = _GEN_1116 | _GEN_4065;
  wire        _GEN_4111 = _GEN_58 ? ~_GEN_4110 & _GEN_3983 : ~_GEN_4065 & _GEN_3983;
  wire        _GEN_4112 = _GEN_1119 | _GEN_4066;
  wire        _GEN_4113 = _GEN_58 ? ~_GEN_4112 & _GEN_3985 : ~_GEN_4066 & _GEN_3985;
  wire        _GEN_4114 = _GEN_1122 | _GEN_4067;
  wire        _GEN_4115 = _GEN_58 ? ~_GEN_4114 & _GEN_3987 : ~_GEN_4067 & _GEN_3987;
  wire        _GEN_4116 = _GEN_1125 | _GEN_4068;
  wire        _GEN_4117 = _GEN_58 ? ~_GEN_4116 & _GEN_3989 : ~_GEN_4068 & _GEN_3989;
  wire        _GEN_4118 = _GEN_1128 | _GEN_4069;
  wire        _GEN_4119 = _GEN_58 ? ~_GEN_4118 & _GEN_3991 : ~_GEN_4069 & _GEN_3991;
  wire        _GEN_4120 = _GEN_1131 | _GEN_4070;
  wire        _GEN_4121 = _GEN_58 ? ~_GEN_4120 & _GEN_3993 : ~_GEN_4070 & _GEN_3993;
  wire        _GEN_4122 = _GEN_1134 | _GEN_4071;
  wire        _GEN_4123 = _GEN_58 ? ~_GEN_4122 & _GEN_3995 : ~_GEN_4071 & _GEN_3995;
  wire        _GEN_4124 = _GEN_1137 | _GEN_4072;
  wire        _GEN_4125 = _GEN_58 ? ~_GEN_4124 & _GEN_3997 : ~_GEN_4072 & _GEN_3997;
  wire        _GEN_4126 = _GEN_1140 | _GEN_4073;
  wire        _GEN_4127 = _GEN_58 ? ~_GEN_4126 & _GEN_3999 : ~_GEN_4073 & _GEN_3999;
  wire        _GEN_4128 = _GEN_1143 | _GEN_4074;
  wire        _GEN_4129 = _GEN_58 ? ~_GEN_4128 & _GEN_4001 : ~_GEN_4074 & _GEN_4001;
  wire        _GEN_4130 = _GEN_1146 | _GEN_4075;
  wire        _GEN_4131 = _GEN_58 ? ~_GEN_4130 & _GEN_4003 : ~_GEN_4075 & _GEN_4003;
  wire        _GEN_4132 = _GEN_1149 | _GEN_4076;
  wire        _GEN_4133 = _GEN_58 ? ~_GEN_4132 & _GEN_4005 : ~_GEN_4076 & _GEN_4005;
  wire        _GEN_4134 = _GEN_1152 | _GEN_4077;
  wire        _GEN_4135 = _GEN_58 ? ~_GEN_4134 & _GEN_4007 : ~_GEN_4077 & _GEN_4007;
  wire        _GEN_4136 = _GEN_1155 | _GEN_4078;
  wire        _GEN_4137 = _GEN_58 ? ~_GEN_4136 & _GEN_4009 : ~_GEN_4078 & _GEN_4009;
  wire        _GEN_4138 = _GEN_1158 | _GEN_4079;
  wire        _GEN_4139 = _GEN_58 ? ~_GEN_4138 & _GEN_4011 : ~_GEN_4079 & _GEN_4011;
  wire        _GEN_4140 = _GEN_1161 | _GEN_4080;
  wire        _GEN_4141 = _GEN_58 ? ~_GEN_4140 & _GEN_4013 : ~_GEN_4080 & _GEN_4013;
  wire        _GEN_4142 = _GEN_1164 | _GEN_4081;
  wire        _GEN_4143 = _GEN_58 ? ~_GEN_4142 & _GEN_4015 : ~_GEN_4081 & _GEN_4015;
  wire        _GEN_4144 = _GEN_1167 | _GEN_4082;
  wire        _GEN_4145 = _GEN_58 ? ~_GEN_4144 & _GEN_4017 : ~_GEN_4082 & _GEN_4017;
  wire        _GEN_4146 = (&(io_wb_resps_9_bits_uop_rob_idx[6:2])) | _GEN_4083;
  wire        _GEN_4147 = _GEN_58 ? ~_GEN_4146 & _GEN_4019 : ~_GEN_4083 & _GEN_4019;
  wire        _GEN_4148 = _GEN_58 ? ~_GEN_4084 & _GEN_4020 : ~_GEN_4052 & _GEN_4020;
  wire        _GEN_4149 = _GEN_58 ? ~_GEN_4086 & _GEN_4021 : ~_GEN_4053 & _GEN_4021;
  wire        _GEN_4150 = _GEN_58 ? ~_GEN_4088 & _GEN_4022 : ~_GEN_4054 & _GEN_4022;
  wire        _GEN_4151 = _GEN_58 ? ~_GEN_4090 & _GEN_4023 : ~_GEN_4055 & _GEN_4023;
  wire        _GEN_4152 = _GEN_58 ? ~_GEN_4092 & _GEN_4024 : ~_GEN_4056 & _GEN_4024;
  wire        _GEN_4153 = _GEN_58 ? ~_GEN_4094 & _GEN_4025 : ~_GEN_4057 & _GEN_4025;
  wire        _GEN_4154 = _GEN_58 ? ~_GEN_4096 & _GEN_4026 : ~_GEN_4058 & _GEN_4026;
  wire        _GEN_4155 = _GEN_58 ? ~_GEN_4098 & _GEN_4027 : ~_GEN_4059 & _GEN_4027;
  wire        _GEN_4156 = _GEN_58 ? ~_GEN_4100 & _GEN_4028 : ~_GEN_4060 & _GEN_4028;
  wire        _GEN_4157 = _GEN_58 ? ~_GEN_4102 & _GEN_4029 : ~_GEN_4061 & _GEN_4029;
  wire        _GEN_4158 = _GEN_58 ? ~_GEN_4104 & _GEN_4030 : ~_GEN_4062 & _GEN_4030;
  wire        _GEN_4159 = _GEN_58 ? ~_GEN_4106 & _GEN_4031 : ~_GEN_4063 & _GEN_4031;
  wire        _GEN_4160 = _GEN_58 ? ~_GEN_4108 & _GEN_4032 : ~_GEN_4064 & _GEN_4032;
  wire        _GEN_4161 = _GEN_58 ? ~_GEN_4110 & _GEN_4033 : ~_GEN_4065 & _GEN_4033;
  wire        _GEN_4162 = _GEN_58 ? ~_GEN_4112 & _GEN_4034 : ~_GEN_4066 & _GEN_4034;
  wire        _GEN_4163 = _GEN_58 ? ~_GEN_4114 & _GEN_4035 : ~_GEN_4067 & _GEN_4035;
  wire        _GEN_4164 = _GEN_58 ? ~_GEN_4116 & _GEN_4036 : ~_GEN_4068 & _GEN_4036;
  wire        _GEN_4165 = _GEN_58 ? ~_GEN_4118 & _GEN_4037 : ~_GEN_4069 & _GEN_4037;
  wire        _GEN_4166 = _GEN_58 ? ~_GEN_4120 & _GEN_4038 : ~_GEN_4070 & _GEN_4038;
  wire        _GEN_4167 = _GEN_58 ? ~_GEN_4122 & _GEN_4039 : ~_GEN_4071 & _GEN_4039;
  wire        _GEN_4168 = _GEN_58 ? ~_GEN_4124 & _GEN_4040 : ~_GEN_4072 & _GEN_4040;
  wire        _GEN_4169 = _GEN_58 ? ~_GEN_4126 & _GEN_4041 : ~_GEN_4073 & _GEN_4041;
  wire        _GEN_4170 = _GEN_58 ? ~_GEN_4128 & _GEN_4042 : ~_GEN_4074 & _GEN_4042;
  wire        _GEN_4171 = _GEN_58 ? ~_GEN_4130 & _GEN_4043 : ~_GEN_4075 & _GEN_4043;
  wire        _GEN_4172 = _GEN_58 ? ~_GEN_4132 & _GEN_4044 : ~_GEN_4076 & _GEN_4044;
  wire        _GEN_4173 = _GEN_58 ? ~_GEN_4134 & _GEN_4045 : ~_GEN_4077 & _GEN_4045;
  wire        _GEN_4174 = _GEN_58 ? ~_GEN_4136 & _GEN_4046 : ~_GEN_4078 & _GEN_4046;
  wire        _GEN_4175 = _GEN_58 ? ~_GEN_4138 & _GEN_4047 : ~_GEN_4079 & _GEN_4047;
  wire        _GEN_4176 = _GEN_58 ? ~_GEN_4140 & _GEN_4048 : ~_GEN_4080 & _GEN_4048;
  wire        _GEN_4177 = _GEN_58 ? ~_GEN_4142 & _GEN_4049 : ~_GEN_4081 & _GEN_4049;
  wire        _GEN_4178 = _GEN_58 ? ~_GEN_4144 & _GEN_4050 : ~_GEN_4082 & _GEN_4050;
  wire        _GEN_4179 = _GEN_58 ? ~_GEN_4146 & _GEN_4051 : ~_GEN_4083 & _GEN_4051;
  wire        _GEN_4180 = _GEN_59 & _GEN_1204;
  wire        _GEN_4181 = _GEN_59 & _GEN_1206;
  wire        _GEN_4182 = _GEN_59 & _GEN_1208;
  wire        _GEN_4183 = _GEN_59 & _GEN_1210;
  wire        _GEN_4184 = _GEN_59 & _GEN_1212;
  wire        _GEN_4185 = _GEN_59 & _GEN_1214;
  wire        _GEN_4186 = _GEN_59 & _GEN_1216;
  wire        _GEN_4187 = _GEN_59 & _GEN_1218;
  wire        _GEN_4188 = _GEN_59 & _GEN_1220;
  wire        _GEN_4189 = _GEN_59 & _GEN_1222;
  wire        _GEN_4190 = _GEN_59 & _GEN_1224;
  wire        _GEN_4191 = _GEN_59 & _GEN_1226;
  wire        _GEN_4192 = _GEN_59 & _GEN_1228;
  wire        _GEN_4193 = _GEN_59 & _GEN_1230;
  wire        _GEN_4194 = _GEN_59 & _GEN_1232;
  wire        _GEN_4195 = _GEN_59 & _GEN_1234;
  wire        _GEN_4196 = _GEN_59 & _GEN_1236;
  wire        _GEN_4197 = _GEN_59 & _GEN_1238;
  wire        _GEN_4198 = _GEN_59 & _GEN_1240;
  wire        _GEN_4199 = _GEN_59 & _GEN_1242;
  wire        _GEN_4200 = _GEN_59 & _GEN_1244;
  wire        _GEN_4201 = _GEN_59 & _GEN_1246;
  wire        _GEN_4202 = _GEN_59 & _GEN_1248;
  wire        _GEN_4203 = _GEN_59 & _GEN_1250;
  wire        _GEN_4204 = _GEN_59 & _GEN_1252;
  wire        _GEN_4205 = _GEN_59 & _GEN_1254;
  wire        _GEN_4206 = _GEN_59 & _GEN_1256;
  wire        _GEN_4207 = _GEN_59 & _GEN_1258;
  wire        _GEN_4208 = _GEN_59 & _GEN_1260;
  wire        _GEN_4209 = _GEN_59 & _GEN_1262;
  wire        _GEN_4210 = _GEN_59 & _GEN_1264;
  wire        _GEN_4211 = _GEN_59 & (&(io_lsu_clr_bsy_0_bits[6:2]));
  wire        _GEN_4212 = _GEN_1267 | _GEN_4180;
  wire        _GEN_4213 = _GEN_1269 | _GEN_4181;
  wire        _GEN_4214 = _GEN_1271 | _GEN_4182;
  wire        _GEN_4215 = _GEN_1273 | _GEN_4183;
  wire        _GEN_4216 = _GEN_1275 | _GEN_4184;
  wire        _GEN_4217 = _GEN_1277 | _GEN_4185;
  wire        _GEN_4218 = _GEN_1279 | _GEN_4186;
  wire        _GEN_4219 = _GEN_1281 | _GEN_4187;
  wire        _GEN_4220 = _GEN_1283 | _GEN_4188;
  wire        _GEN_4221 = _GEN_1285 | _GEN_4189;
  wire        _GEN_4222 = _GEN_1287 | _GEN_4190;
  wire        _GEN_4223 = _GEN_1289 | _GEN_4191;
  wire        _GEN_4224 = _GEN_1291 | _GEN_4192;
  wire        _GEN_4225 = _GEN_1293 | _GEN_4193;
  wire        _GEN_4226 = _GEN_1295 | _GEN_4194;
  wire        _GEN_4227 = _GEN_1297 | _GEN_4195;
  wire        _GEN_4228 = _GEN_1299 | _GEN_4196;
  wire        _GEN_4229 = _GEN_1301 | _GEN_4197;
  wire        _GEN_4230 = _GEN_1303 | _GEN_4198;
  wire        _GEN_4231 = _GEN_1305 | _GEN_4199;
  wire        _GEN_4232 = _GEN_1307 | _GEN_4200;
  wire        _GEN_4233 = _GEN_1309 | _GEN_4201;
  wire        _GEN_4234 = _GEN_1311 | _GEN_4202;
  wire        _GEN_4235 = _GEN_1313 | _GEN_4203;
  wire        _GEN_4236 = _GEN_1315 | _GEN_4204;
  wire        _GEN_4237 = _GEN_1317 | _GEN_4205;
  wire        _GEN_4238 = _GEN_1319 | _GEN_4206;
  wire        _GEN_4239 = _GEN_1321 | _GEN_4207;
  wire        _GEN_4240 = _GEN_1323 | _GEN_4208;
  wire        _GEN_4241 = _GEN_1325 | _GEN_4209;
  wire        _GEN_4242 = _GEN_1327 | _GEN_4210;
  wire        _GEN_4243 = (&(io_lsu_clr_bsy_1_bits[6:2])) | _GEN_4211;
  wire        _GEN_4244 = _GEN_61 & _GEN_1330;
  wire        _GEN_4245 = _GEN_61 & _GEN_1332;
  wire        _GEN_4246 = _GEN_61 & _GEN_1334;
  wire        _GEN_4247 = _GEN_61 & _GEN_1336;
  wire        _GEN_4248 = _GEN_61 & _GEN_1338;
  wire        _GEN_4249 = _GEN_61 & _GEN_1340;
  wire        _GEN_4250 = _GEN_61 & _GEN_1342;
  wire        _GEN_4251 = _GEN_61 & _GEN_1344;
  wire        _GEN_4252 = _GEN_61 & _GEN_1346;
  wire        _GEN_4253 = _GEN_61 & _GEN_1348;
  wire        _GEN_4254 = _GEN_61 & _GEN_1350;
  wire        _GEN_4255 = _GEN_61 & _GEN_1352;
  wire        _GEN_4256 = _GEN_61 & _GEN_1354;
  wire        _GEN_4257 = _GEN_61 & _GEN_1356;
  wire        _GEN_4258 = _GEN_61 & _GEN_1358;
  wire        _GEN_4259 = _GEN_61 & _GEN_1360;
  wire        _GEN_4260 = _GEN_61 & _GEN_1362;
  wire        _GEN_4261 = _GEN_61 & _GEN_1364;
  wire        _GEN_4262 = _GEN_61 & _GEN_1366;
  wire        _GEN_4263 = _GEN_61 & _GEN_1368;
  wire        _GEN_4264 = _GEN_61 & _GEN_1370;
  wire        _GEN_4265 = _GEN_61 & _GEN_1372;
  wire        _GEN_4266 = _GEN_61 & _GEN_1374;
  wire        _GEN_4267 = _GEN_61 & _GEN_1376;
  wire        _GEN_4268 = _GEN_61 & _GEN_1378;
  wire        _GEN_4269 = _GEN_61 & _GEN_1380;
  wire        _GEN_4270 = _GEN_61 & _GEN_1382;
  wire        _GEN_4271 = _GEN_61 & _GEN_1384;
  wire        _GEN_4272 = _GEN_61 & _GEN_1386;
  wire        _GEN_4273 = _GEN_61 & _GEN_1388;
  wire        _GEN_4274 = _GEN_61 & _GEN_1390;
  wire        _GEN_4275 = _GEN_61 & (&(io_lsu_clr_bsy_2_bits[6:2]));
  wire        _GEN_4276 = io_fflags_0_valid & (&(io_fflags_0_bits_uop_rob_idx[1:0]));
  wire        _GEN_4277 = io_fflags_2_valid & (&(io_fflags_2_bits_uop_rob_idx[1:0]));
  wire        _GEN_4278 = io_fflags_3_valid & (&(io_fflags_3_bits_uop_rob_idx[1:0]));
  wire        _GEN_4279 = rbk_row_3 & _GEN_1520;
  wire        _GEN_4280 = rbk_row_3 & _GEN_1522;
  wire        _GEN_4281 = rbk_row_3 & _GEN_1524;
  wire        _GEN_4282 = rbk_row_3 & _GEN_1526;
  wire        _GEN_4283 = rbk_row_3 & _GEN_1528;
  wire        _GEN_4284 = rbk_row_3 & _GEN_1530;
  wire        _GEN_4285 = rbk_row_3 & _GEN_1532;
  wire        _GEN_4286 = rbk_row_3 & _GEN_1534;
  wire        _GEN_4287 = rbk_row_3 & _GEN_1536;
  wire        _GEN_4288 = rbk_row_3 & _GEN_1538;
  wire        _GEN_4289 = rbk_row_3 & _GEN_1540;
  wire        _GEN_4290 = rbk_row_3 & _GEN_1542;
  wire        _GEN_4291 = rbk_row_3 & _GEN_1544;
  wire        _GEN_4292 = rbk_row_3 & _GEN_1546;
  wire        _GEN_4293 = rbk_row_3 & _GEN_1548;
  wire        _GEN_4294 = rbk_row_3 & _GEN_1550;
  wire        _GEN_4295 = rbk_row_3 & _GEN_1552;
  wire        _GEN_4296 = rbk_row_3 & _GEN_1554;
  wire        _GEN_4297 = rbk_row_3 & _GEN_1556;
  wire        _GEN_4298 = rbk_row_3 & _GEN_1558;
  wire        _GEN_4299 = rbk_row_3 & _GEN_1560;
  wire        _GEN_4300 = rbk_row_3 & _GEN_1562;
  wire        _GEN_4301 = rbk_row_3 & _GEN_1564;
  wire        _GEN_4302 = rbk_row_3 & _GEN_1566;
  wire        _GEN_4303 = rbk_row_3 & _GEN_1568;
  wire        _GEN_4304 = rbk_row_3 & _GEN_1570;
  wire        _GEN_4305 = rbk_row_3 & _GEN_1572;
  wire        _GEN_4306 = rbk_row_3 & _GEN_1574;
  wire        _GEN_4307 = rbk_row_3 & _GEN_1576;
  wire        _GEN_4308 = rbk_row_3 & _GEN_1578;
  wire        _GEN_4309 = rbk_row_3 & _GEN_1580;
  wire        _GEN_4310 = rbk_row_3 & (&com_idx);
  wire [19:0] _GEN_4311 = io_brupdate_b1_mispredict_mask & rob_uop_3_0_br_mask;
  wire [19:0] _GEN_4312 = io_brupdate_b1_mispredict_mask & rob_uop_3_1_br_mask;
  wire [19:0] _GEN_4313 = io_brupdate_b1_mispredict_mask & rob_uop_3_2_br_mask;
  wire [19:0] _GEN_4314 = io_brupdate_b1_mispredict_mask & rob_uop_3_3_br_mask;
  wire [19:0] _GEN_4315 = io_brupdate_b1_mispredict_mask & rob_uop_3_4_br_mask;
  wire [19:0] _GEN_4316 = io_brupdate_b1_mispredict_mask & rob_uop_3_5_br_mask;
  wire [19:0] _GEN_4317 = io_brupdate_b1_mispredict_mask & rob_uop_3_6_br_mask;
  wire [19:0] _GEN_4318 = io_brupdate_b1_mispredict_mask & rob_uop_3_7_br_mask;
  wire [19:0] _GEN_4319 = io_brupdate_b1_mispredict_mask & rob_uop_3_8_br_mask;
  wire [19:0] _GEN_4320 = io_brupdate_b1_mispredict_mask & rob_uop_3_9_br_mask;
  wire [19:0] _GEN_4321 = io_brupdate_b1_mispredict_mask & rob_uop_3_10_br_mask;
  wire [19:0] _GEN_4322 = io_brupdate_b1_mispredict_mask & rob_uop_3_11_br_mask;
  wire [19:0] _GEN_4323 = io_brupdate_b1_mispredict_mask & rob_uop_3_12_br_mask;
  wire [19:0] _GEN_4324 = io_brupdate_b1_mispredict_mask & rob_uop_3_13_br_mask;
  wire [19:0] _GEN_4325 = io_brupdate_b1_mispredict_mask & rob_uop_3_14_br_mask;
  wire [19:0] _GEN_4326 = io_brupdate_b1_mispredict_mask & rob_uop_3_15_br_mask;
  wire [19:0] _GEN_4327 = io_brupdate_b1_mispredict_mask & rob_uop_3_16_br_mask;
  wire [19:0] _GEN_4328 = io_brupdate_b1_mispredict_mask & rob_uop_3_17_br_mask;
  wire [19:0] _GEN_4329 = io_brupdate_b1_mispredict_mask & rob_uop_3_18_br_mask;
  wire [19:0] _GEN_4330 = io_brupdate_b1_mispredict_mask & rob_uop_3_19_br_mask;
  wire [19:0] _GEN_4331 = io_brupdate_b1_mispredict_mask & rob_uop_3_20_br_mask;
  wire [19:0] _GEN_4332 = io_brupdate_b1_mispredict_mask & rob_uop_3_21_br_mask;
  wire [19:0] _GEN_4333 = io_brupdate_b1_mispredict_mask & rob_uop_3_22_br_mask;
  wire [19:0] _GEN_4334 = io_brupdate_b1_mispredict_mask & rob_uop_3_23_br_mask;
  wire [19:0] _GEN_4335 = io_brupdate_b1_mispredict_mask & rob_uop_3_24_br_mask;
  wire [19:0] _GEN_4336 = io_brupdate_b1_mispredict_mask & rob_uop_3_25_br_mask;
  wire [19:0] _GEN_4337 = io_brupdate_b1_mispredict_mask & rob_uop_3_26_br_mask;
  wire [19:0] _GEN_4338 = io_brupdate_b1_mispredict_mask & rob_uop_3_27_br_mask;
  wire [19:0] _GEN_4339 = io_brupdate_b1_mispredict_mask & rob_uop_3_28_br_mask;
  wire [19:0] _GEN_4340 = io_brupdate_b1_mispredict_mask & rob_uop_3_29_br_mask;
  wire [19:0] _GEN_4341 = io_brupdate_b1_mispredict_mask & rob_uop_3_30_br_mask;
  wire [19:0] _GEN_4342 = io_brupdate_b1_mispredict_mask & rob_uop_3_31_br_mask;
  wire        _GEN_4343 = ~(_io_flush_valid_output | exception_thrown) & rob_state != 2'h2;
  wire        _GEN_4344 = ~r_xcpt_val | io_lxcpt_bits_uop_rob_idx < r_xcpt_uop_rob_idx ^ io_lxcpt_bits_uop_rob_idx < rob_head_idx ^ r_xcpt_uop_rob_idx < rob_head_idx;
  wire        _GEN_4345 = ~r_xcpt_val & (enq_xcpts_0 | enq_xcpts_1 | enq_xcpts_2 | io_enq_valids_3 & io_enq_uops_3_exception);
  wire [19:0] next_xcpt_uop_br_mask = _GEN_4343 ? (io_lxcpt_valid ? (_GEN_4344 ? io_lxcpt_bits_uop_br_mask : r_xcpt_uop_br_mask) : _GEN_4345 ? casez_tmp_311 : r_xcpt_uop_br_mask) : r_xcpt_uop_br_mask;
  wire        _GEN_4346 = _GEN_128 | rob_val_0;
  wire        _GEN_4347 = _GEN_130 | rob_val_1;
  wire        _GEN_4348 = _GEN_132 | rob_val_2;
  wire        _GEN_4349 = _GEN_134 | rob_val_3;
  wire        _GEN_4350 = _GEN_136 | rob_val_4;
  wire        _GEN_4351 = _GEN_138 | rob_val_5;
  wire        _GEN_4352 = _GEN_140 | rob_val_6;
  wire        _GEN_4353 = _GEN_142 | rob_val_7;
  wire        _GEN_4354 = _GEN_144 | rob_val_8;
  wire        _GEN_4355 = _GEN_146 | rob_val_9;
  wire        _GEN_4356 = _GEN_148 | rob_val_10;
  wire        _GEN_4357 = _GEN_150 | rob_val_11;
  wire        _GEN_4358 = _GEN_152 | rob_val_12;
  wire        _GEN_4359 = _GEN_154 | rob_val_13;
  wire        _GEN_4360 = _GEN_156 | rob_val_14;
  wire        _GEN_4361 = _GEN_158 | rob_val_15;
  wire        _GEN_4362 = _GEN_160 | rob_val_16;
  wire        _GEN_4363 = _GEN_162 | rob_val_17;
  wire        _GEN_4364 = _GEN_164 | rob_val_18;
  wire        _GEN_4365 = _GEN_166 | rob_val_19;
  wire        _GEN_4366 = _GEN_168 | rob_val_20;
  wire        _GEN_4367 = _GEN_170 | rob_val_21;
  wire        _GEN_4368 = _GEN_172 | rob_val_22;
  wire        _GEN_4369 = _GEN_174 | rob_val_23;
  wire        _GEN_4370 = _GEN_176 | rob_val_24;
  wire        _GEN_4371 = _GEN_178 | rob_val_25;
  wire        _GEN_4372 = _GEN_180 | rob_val_26;
  wire        _GEN_4373 = _GEN_182 | rob_val_27;
  wire        _GEN_4374 = _GEN_184 | rob_val_28;
  wire        _GEN_4375 = _GEN_186 | rob_val_29;
  wire        _GEN_4376 = _GEN_188 | rob_val_30;
  wire        _GEN_4377 = _GEN_189 | rob_val_31;
  wire        _GEN_4378 = _GEN_1646 | rob_val_1_0;
  wire        _GEN_4379 = _GEN_1647 | rob_val_1_1;
  wire        _GEN_4380 = _GEN_1648 | rob_val_1_2;
  wire        _GEN_4381 = _GEN_1649 | rob_val_1_3;
  wire        _GEN_4382 = _GEN_1650 | rob_val_1_4;
  wire        _GEN_4383 = _GEN_1651 | rob_val_1_5;
  wire        _GEN_4384 = _GEN_1652 | rob_val_1_6;
  wire        _GEN_4385 = _GEN_1653 | rob_val_1_7;
  wire        _GEN_4386 = _GEN_1654 | rob_val_1_8;
  wire        _GEN_4387 = _GEN_1655 | rob_val_1_9;
  wire        _GEN_4388 = _GEN_1656 | rob_val_1_10;
  wire        _GEN_4389 = _GEN_1657 | rob_val_1_11;
  wire        _GEN_4390 = _GEN_1658 | rob_val_1_12;
  wire        _GEN_4391 = _GEN_1659 | rob_val_1_13;
  wire        _GEN_4392 = _GEN_1660 | rob_val_1_14;
  wire        _GEN_4393 = _GEN_1661 | rob_val_1_15;
  wire        _GEN_4394 = _GEN_1662 | rob_val_1_16;
  wire        _GEN_4395 = _GEN_1663 | rob_val_1_17;
  wire        _GEN_4396 = _GEN_1664 | rob_val_1_18;
  wire        _GEN_4397 = _GEN_1665 | rob_val_1_19;
  wire        _GEN_4398 = _GEN_1666 | rob_val_1_20;
  wire        _GEN_4399 = _GEN_1667 | rob_val_1_21;
  wire        _GEN_4400 = _GEN_1668 | rob_val_1_22;
  wire        _GEN_4401 = _GEN_1669 | rob_val_1_23;
  wire        _GEN_4402 = _GEN_1670 | rob_val_1_24;
  wire        _GEN_4403 = _GEN_1671 | rob_val_1_25;
  wire        _GEN_4404 = _GEN_1672 | rob_val_1_26;
  wire        _GEN_4405 = _GEN_1673 | rob_val_1_27;
  wire        _GEN_4406 = _GEN_1674 | rob_val_1_28;
  wire        _GEN_4407 = _GEN_1675 | rob_val_1_29;
  wire        _GEN_4408 = _GEN_1676 | rob_val_1_30;
  wire        _GEN_4409 = _GEN_1677 | rob_val_1_31;
  wire        _GEN_4410 = _GEN_2545 | rob_val_2_0;
  wire        _GEN_4411 = _GEN_2546 | rob_val_2_1;
  wire        _GEN_4412 = _GEN_2547 | rob_val_2_2;
  wire        _GEN_4413 = _GEN_2548 | rob_val_2_3;
  wire        _GEN_4414 = _GEN_2549 | rob_val_2_4;
  wire        _GEN_4415 = _GEN_2550 | rob_val_2_5;
  wire        _GEN_4416 = _GEN_2551 | rob_val_2_6;
  wire        _GEN_4417 = _GEN_2552 | rob_val_2_7;
  wire        _GEN_4418 = _GEN_2553 | rob_val_2_8;
  wire        _GEN_4419 = _GEN_2554 | rob_val_2_9;
  wire        _GEN_4420 = _GEN_2555 | rob_val_2_10;
  wire        _GEN_4421 = _GEN_2556 | rob_val_2_11;
  wire        _GEN_4422 = _GEN_2557 | rob_val_2_12;
  wire        _GEN_4423 = _GEN_2558 | rob_val_2_13;
  wire        _GEN_4424 = _GEN_2559 | rob_val_2_14;
  wire        _GEN_4425 = _GEN_2560 | rob_val_2_15;
  wire        _GEN_4426 = _GEN_2561 | rob_val_2_16;
  wire        _GEN_4427 = _GEN_2562 | rob_val_2_17;
  wire        _GEN_4428 = _GEN_2563 | rob_val_2_18;
  wire        _GEN_4429 = _GEN_2564 | rob_val_2_19;
  wire        _GEN_4430 = _GEN_2565 | rob_val_2_20;
  wire        _GEN_4431 = _GEN_2566 | rob_val_2_21;
  wire        _GEN_4432 = _GEN_2567 | rob_val_2_22;
  wire        _GEN_4433 = _GEN_2568 | rob_val_2_23;
  wire        _GEN_4434 = _GEN_2569 | rob_val_2_24;
  wire        _GEN_4435 = _GEN_2570 | rob_val_2_25;
  wire        _GEN_4436 = _GEN_2571 | rob_val_2_26;
  wire        _GEN_4437 = _GEN_2572 | rob_val_2_27;
  wire        _GEN_4438 = _GEN_2573 | rob_val_2_28;
  wire        _GEN_4439 = _GEN_2574 | rob_val_2_29;
  wire        _GEN_4440 = _GEN_2575 | rob_val_2_30;
  wire        _GEN_4441 = _GEN_2576 | rob_val_2_31;
  wire        _GEN_4442 = _GEN_3444 | rob_val_3_0;
  wire        _GEN_4443 = _GEN_3445 | rob_val_3_1;
  wire        _GEN_4444 = _GEN_3446 | rob_val_3_2;
  wire        _GEN_4445 = _GEN_3447 | rob_val_3_3;
  wire        _GEN_4446 = _GEN_3448 | rob_val_3_4;
  wire        _GEN_4447 = _GEN_3449 | rob_val_3_5;
  wire        _GEN_4448 = _GEN_3450 | rob_val_3_6;
  wire        _GEN_4449 = _GEN_3451 | rob_val_3_7;
  wire        _GEN_4450 = _GEN_3452 | rob_val_3_8;
  wire        _GEN_4451 = _GEN_3453 | rob_val_3_9;
  wire        _GEN_4452 = _GEN_3454 | rob_val_3_10;
  wire        _GEN_4453 = _GEN_3455 | rob_val_3_11;
  wire        _GEN_4454 = _GEN_3456 | rob_val_3_12;
  wire        _GEN_4455 = _GEN_3457 | rob_val_3_13;
  wire        _GEN_4456 = _GEN_3458 | rob_val_3_14;
  wire        _GEN_4457 = _GEN_3459 | rob_val_3_15;
  wire        _GEN_4458 = _GEN_3460 | rob_val_3_16;
  wire        _GEN_4459 = _GEN_3461 | rob_val_3_17;
  wire        _GEN_4460 = _GEN_3462 | rob_val_3_18;
  wire        _GEN_4461 = _GEN_3463 | rob_val_3_19;
  wire        _GEN_4462 = _GEN_3464 | rob_val_3_20;
  wire        _GEN_4463 = _GEN_3465 | rob_val_3_21;
  wire        _GEN_4464 = _GEN_3466 | rob_val_3_22;
  wire        _GEN_4465 = _GEN_3467 | rob_val_3_23;
  wire        _GEN_4466 = _GEN_3468 | rob_val_3_24;
  wire        _GEN_4467 = _GEN_3469 | rob_val_3_25;
  wire        _GEN_4468 = _GEN_3470 | rob_val_3_26;
  wire        _GEN_4469 = _GEN_3471 | rob_val_3_27;
  wire        _GEN_4470 = _GEN_3472 | rob_val_3_28;
  wire        _GEN_4471 = _GEN_3473 | rob_val_3_29;
  wire        _GEN_4472 = _GEN_3474 | rob_val_3_30;
  wire        _GEN_4473 = _GEN_3475 | rob_val_3_31;
  always @(posedge clock) begin
    if (_GEN_14)
      assert__assert_8: assert(casez_tmp_6);
    if (_GEN_31)
      assert__assert_48: assert(casez_tmp_84);
    if (_GEN_47)
      assert__assert_88: assert(casez_tmp_162);
    if (_GEN_63)
      assert__assert_128: assert(casez_tmp_240);
    if (reset) begin
      rob_state <= 2'h0;
      rob_head <= 5'h0;
      rob_head_lsb <= 2'h0;
      rob_tail <= 5'h0;
      rob_tail_lsb <= 2'h0;
      rob_pnr <= 5'h0;
      rob_pnr_lsb <= 2'h0;
      maybe_full <= 1'h0;
      r_xcpt_val <= 1'h0;
      rob_val_0 <= 1'h0;
      rob_val_1 <= 1'h0;
      rob_val_2 <= 1'h0;
      rob_val_3 <= 1'h0;
      rob_val_4 <= 1'h0;
      rob_val_5 <= 1'h0;
      rob_val_6 <= 1'h0;
      rob_val_7 <= 1'h0;
      rob_val_8 <= 1'h0;
      rob_val_9 <= 1'h0;
      rob_val_10 <= 1'h0;
      rob_val_11 <= 1'h0;
      rob_val_12 <= 1'h0;
      rob_val_13 <= 1'h0;
      rob_val_14 <= 1'h0;
      rob_val_15 <= 1'h0;
      rob_val_16 <= 1'h0;
      rob_val_17 <= 1'h0;
      rob_val_18 <= 1'h0;
      rob_val_19 <= 1'h0;
      rob_val_20 <= 1'h0;
      rob_val_21 <= 1'h0;
      rob_val_22 <= 1'h0;
      rob_val_23 <= 1'h0;
      rob_val_24 <= 1'h0;
      rob_val_25 <= 1'h0;
      rob_val_26 <= 1'h0;
      rob_val_27 <= 1'h0;
      rob_val_28 <= 1'h0;
      rob_val_29 <= 1'h0;
      rob_val_30 <= 1'h0;
      rob_val_31 <= 1'h0;
      rob_val_1_0 <= 1'h0;
      rob_val_1_1 <= 1'h0;
      rob_val_1_2 <= 1'h0;
      rob_val_1_3 <= 1'h0;
      rob_val_1_4 <= 1'h0;
      rob_val_1_5 <= 1'h0;
      rob_val_1_6 <= 1'h0;
      rob_val_1_7 <= 1'h0;
      rob_val_1_8 <= 1'h0;
      rob_val_1_9 <= 1'h0;
      rob_val_1_10 <= 1'h0;
      rob_val_1_11 <= 1'h0;
      rob_val_1_12 <= 1'h0;
      rob_val_1_13 <= 1'h0;
      rob_val_1_14 <= 1'h0;
      rob_val_1_15 <= 1'h0;
      rob_val_1_16 <= 1'h0;
      rob_val_1_17 <= 1'h0;
      rob_val_1_18 <= 1'h0;
      rob_val_1_19 <= 1'h0;
      rob_val_1_20 <= 1'h0;
      rob_val_1_21 <= 1'h0;
      rob_val_1_22 <= 1'h0;
      rob_val_1_23 <= 1'h0;
      rob_val_1_24 <= 1'h0;
      rob_val_1_25 <= 1'h0;
      rob_val_1_26 <= 1'h0;
      rob_val_1_27 <= 1'h0;
      rob_val_1_28 <= 1'h0;
      rob_val_1_29 <= 1'h0;
      rob_val_1_30 <= 1'h0;
      rob_val_1_31 <= 1'h0;
      rob_val_2_0 <= 1'h0;
      rob_val_2_1 <= 1'h0;
      rob_val_2_2 <= 1'h0;
      rob_val_2_3 <= 1'h0;
      rob_val_2_4 <= 1'h0;
      rob_val_2_5 <= 1'h0;
      rob_val_2_6 <= 1'h0;
      rob_val_2_7 <= 1'h0;
      rob_val_2_8 <= 1'h0;
      rob_val_2_9 <= 1'h0;
      rob_val_2_10 <= 1'h0;
      rob_val_2_11 <= 1'h0;
      rob_val_2_12 <= 1'h0;
      rob_val_2_13 <= 1'h0;
      rob_val_2_14 <= 1'h0;
      rob_val_2_15 <= 1'h0;
      rob_val_2_16 <= 1'h0;
      rob_val_2_17 <= 1'h0;
      rob_val_2_18 <= 1'h0;
      rob_val_2_19 <= 1'h0;
      rob_val_2_20 <= 1'h0;
      rob_val_2_21 <= 1'h0;
      rob_val_2_22 <= 1'h0;
      rob_val_2_23 <= 1'h0;
      rob_val_2_24 <= 1'h0;
      rob_val_2_25 <= 1'h0;
      rob_val_2_26 <= 1'h0;
      rob_val_2_27 <= 1'h0;
      rob_val_2_28 <= 1'h0;
      rob_val_2_29 <= 1'h0;
      rob_val_2_30 <= 1'h0;
      rob_val_2_31 <= 1'h0;
      rob_val_3_0 <= 1'h0;
      rob_val_3_1 <= 1'h0;
      rob_val_3_2 <= 1'h0;
      rob_val_3_3 <= 1'h0;
      rob_val_3_4 <= 1'h0;
      rob_val_3_5 <= 1'h0;
      rob_val_3_6 <= 1'h0;
      rob_val_3_7 <= 1'h0;
      rob_val_3_8 <= 1'h0;
      rob_val_3_9 <= 1'h0;
      rob_val_3_10 <= 1'h0;
      rob_val_3_11 <= 1'h0;
      rob_val_3_12 <= 1'h0;
      rob_val_3_13 <= 1'h0;
      rob_val_3_14 <= 1'h0;
      rob_val_3_15 <= 1'h0;
      rob_val_3_16 <= 1'h0;
      rob_val_3_17 <= 1'h0;
      rob_val_3_18 <= 1'h0;
      rob_val_3_19 <= 1'h0;
      rob_val_3_20 <= 1'h0;
      rob_val_3_21 <= 1'h0;
      rob_val_3_22 <= 1'h0;
      rob_val_3_23 <= 1'h0;
      rob_val_3_24 <= 1'h0;
      rob_val_3_25 <= 1'h0;
      rob_val_3_26 <= 1'h0;
      rob_val_3_27 <= 1'h0;
      rob_val_3_28 <= 1'h0;
      rob_val_3_29 <= 1'h0;
      rob_val_3_30 <= 1'h0;
      rob_val_3_31 <= 1'h0;
      r_partial_row <= 1'h0;
      pnr_maybe_at_tail <= 1'h0;
    end
    else begin
      rob_state <= casez_tmp_315;
      if (finished_committing_row)
        rob_head <= rob_head + 5'h1;
      rob_head_lsb <= finished_committing_row ? 2'h0 : {|(_rob_head_lsb_T_8[2:1]), _rob_head_lsb_T_8[2] | _rob_head_lsb_T_8[0]};
      if (_GEN_87) begin
        rob_tail <= rob_tail - 5'h1;
        rob_tail_lsb <= 2'h3;
      end
      else if (_GEN_125)
        rob_tail_lsb <= rob_head_lsb;
      else begin
        if (io_brupdate_b2_mispredict)
          rob_tail <= io_brupdate_b2_uop_rob_idx[6:2] + 5'h1;
        else if (_GEN_126)
          rob_tail <= rob_tail + 5'h1;
        if (io_brupdate_b2_mispredict | _GEN_126)
          rob_tail_lsb <= 2'h0;
        else if ((|_GEN_124) & io_enq_partial_stall)
          rob_tail_lsb <= _rob_tail_lsb_T_8[0] ? 2'h0 : _rob_tail_lsb_T_8[1] ? 2'h1 : {1'h1, ~(_rob_tail_lsb_T_8[2])};
      end
      if (empty & (|_GEN_124)) begin
        rob_pnr <= rob_head;
        rob_pnr_lsb <= io_enq_valids_0 ? 2'h0 : io_enq_valids_1 ? 2'h1 : {1'h1, ~io_enq_valids_2};
      end
      else if (safe_to_inc & do_inc_row) begin
        rob_pnr <= rob_pnr + 5'h1;
        rob_pnr_lsb <= 2'h0;
      end
      else if (safe_to_inc & (_do_inc_row_T_4 | full & ~pnr_maybe_at_tail))
        rob_pnr_lsb <= rob_pnr_unsafe_0 ? 2'h0 : rob_pnr_unsafe_1 ? 2'h1 : {1'h1, ~rob_pnr_unsafe_2};
      else if (safe_to_inc & ~full & ~empty)
        rob_pnr_lsb <= _rob_pnr_lsb_T_16[0] ? 2'h0 : _rob_pnr_lsb_T_16[1] ? 2'h1 : {1'h1, ~(_rob_pnr_lsb_T_16[2])};
      else if (full & pnr_maybe_at_tail)
        rob_pnr_lsb <= 2'h0;
      maybe_full <= ~rob_deq & (~(_GEN_87 | _GEN_125 | io_brupdate_b2_mispredict) & _GEN_126 | maybe_full) | (|io_brupdate_b1_mispredict_mask);
      r_xcpt_val <= ~(_io_flush_valid_output | (|(io_brupdate_b1_mispredict_mask & next_xcpt_uop_br_mask))) & (_GEN_4343 ? (io_lxcpt_valid ? _GEN_4344 | r_xcpt_val : _GEN_4345 | r_xcpt_val) : r_xcpt_val);
      if (will_commit_0) begin
        rob_val_0 <= ~(_GEN_93 | (|_GEN_1583) | _GEN_1521) & _GEN_4346;
        rob_val_1 <= ~(_GEN_94 | (|_GEN_1584) | _GEN_1523) & _GEN_4347;
        rob_val_2 <= ~(_GEN_95 | (|_GEN_1585) | _GEN_1525) & _GEN_4348;
        rob_val_3 <= ~(_GEN_96 | (|_GEN_1586) | _GEN_1527) & _GEN_4349;
        rob_val_4 <= ~(_GEN_97 | (|_GEN_1587) | _GEN_1529) & _GEN_4350;
        rob_val_5 <= ~(_GEN_98 | (|_GEN_1588) | _GEN_1531) & _GEN_4351;
        rob_val_6 <= ~(_GEN_99 | (|_GEN_1589) | _GEN_1533) & _GEN_4352;
        rob_val_7 <= ~(_GEN_100 | (|_GEN_1590) | _GEN_1535) & _GEN_4353;
        rob_val_8 <= ~(_GEN_101 | (|_GEN_1591) | _GEN_1537) & _GEN_4354;
        rob_val_9 <= ~(_GEN_102 | (|_GEN_1592) | _GEN_1539) & _GEN_4355;
        rob_val_10 <= ~(_GEN_103 | (|_GEN_1593) | _GEN_1541) & _GEN_4356;
        rob_val_11 <= ~(_GEN_104 | (|_GEN_1594) | _GEN_1543) & _GEN_4357;
        rob_val_12 <= ~(_GEN_105 | (|_GEN_1595) | _GEN_1545) & _GEN_4358;
        rob_val_13 <= ~(_GEN_106 | (|_GEN_1596) | _GEN_1547) & _GEN_4359;
        rob_val_14 <= ~(_GEN_107 | (|_GEN_1597) | _GEN_1549) & _GEN_4360;
        rob_val_15 <= ~(_GEN_108 | (|_GEN_1598) | _GEN_1551) & _GEN_4361;
        rob_val_16 <= ~(_GEN_109 | (|_GEN_1599) | _GEN_1553) & _GEN_4362;
        rob_val_17 <= ~(_GEN_110 | (|_GEN_1600) | _GEN_1555) & _GEN_4363;
        rob_val_18 <= ~(_GEN_111 | (|_GEN_1601) | _GEN_1557) & _GEN_4364;
        rob_val_19 <= ~(_GEN_112 | (|_GEN_1602) | _GEN_1559) & _GEN_4365;
        rob_val_20 <= ~(_GEN_113 | (|_GEN_1603) | _GEN_1561) & _GEN_4366;
        rob_val_21 <= ~(_GEN_114 | (|_GEN_1604) | _GEN_1563) & _GEN_4367;
        rob_val_22 <= ~(_GEN_115 | (|_GEN_1605) | _GEN_1565) & _GEN_4368;
        rob_val_23 <= ~(_GEN_116 | (|_GEN_1606) | _GEN_1567) & _GEN_4369;
        rob_val_24 <= ~(_GEN_117 | (|_GEN_1607) | _GEN_1569) & _GEN_4370;
        rob_val_25 <= ~(_GEN_118 | (|_GEN_1608) | _GEN_1571) & _GEN_4371;
        rob_val_26 <= ~(_GEN_119 | (|_GEN_1609) | _GEN_1573) & _GEN_4372;
        rob_val_27 <= ~(_GEN_120 | (|_GEN_1610) | _GEN_1575) & _GEN_4373;
        rob_val_28 <= ~(_GEN_121 | (|_GEN_1611) | _GEN_1577) & _GEN_4374;
        rob_val_29 <= ~(_GEN_122 | (|_GEN_1612) | _GEN_1579) & _GEN_4375;
        rob_val_30 <= ~(_GEN_123 | (|_GEN_1613) | _GEN_1581) & _GEN_4376;
        rob_val_31 <= ~((&rob_head) | (|_GEN_1614) | _GEN_1582) & _GEN_4377;
      end
      else begin
        rob_val_0 <= ~((|_GEN_1583) | _GEN_1521) & _GEN_4346;
        rob_val_1 <= ~((|_GEN_1584) | _GEN_1523) & _GEN_4347;
        rob_val_2 <= ~((|_GEN_1585) | _GEN_1525) & _GEN_4348;
        rob_val_3 <= ~((|_GEN_1586) | _GEN_1527) & _GEN_4349;
        rob_val_4 <= ~((|_GEN_1587) | _GEN_1529) & _GEN_4350;
        rob_val_5 <= ~((|_GEN_1588) | _GEN_1531) & _GEN_4351;
        rob_val_6 <= ~((|_GEN_1589) | _GEN_1533) & _GEN_4352;
        rob_val_7 <= ~((|_GEN_1590) | _GEN_1535) & _GEN_4353;
        rob_val_8 <= ~((|_GEN_1591) | _GEN_1537) & _GEN_4354;
        rob_val_9 <= ~((|_GEN_1592) | _GEN_1539) & _GEN_4355;
        rob_val_10 <= ~((|_GEN_1593) | _GEN_1541) & _GEN_4356;
        rob_val_11 <= ~((|_GEN_1594) | _GEN_1543) & _GEN_4357;
        rob_val_12 <= ~((|_GEN_1595) | _GEN_1545) & _GEN_4358;
        rob_val_13 <= ~((|_GEN_1596) | _GEN_1547) & _GEN_4359;
        rob_val_14 <= ~((|_GEN_1597) | _GEN_1549) & _GEN_4360;
        rob_val_15 <= ~((|_GEN_1598) | _GEN_1551) & _GEN_4361;
        rob_val_16 <= ~((|_GEN_1599) | _GEN_1553) & _GEN_4362;
        rob_val_17 <= ~((|_GEN_1600) | _GEN_1555) & _GEN_4363;
        rob_val_18 <= ~((|_GEN_1601) | _GEN_1557) & _GEN_4364;
        rob_val_19 <= ~((|_GEN_1602) | _GEN_1559) & _GEN_4365;
        rob_val_20 <= ~((|_GEN_1603) | _GEN_1561) & _GEN_4366;
        rob_val_21 <= ~((|_GEN_1604) | _GEN_1563) & _GEN_4367;
        rob_val_22 <= ~((|_GEN_1605) | _GEN_1565) & _GEN_4368;
        rob_val_23 <= ~((|_GEN_1606) | _GEN_1567) & _GEN_4369;
        rob_val_24 <= ~((|_GEN_1607) | _GEN_1569) & _GEN_4370;
        rob_val_25 <= ~((|_GEN_1608) | _GEN_1571) & _GEN_4371;
        rob_val_26 <= ~((|_GEN_1609) | _GEN_1573) & _GEN_4372;
        rob_val_27 <= ~((|_GEN_1610) | _GEN_1575) & _GEN_4373;
        rob_val_28 <= ~((|_GEN_1611) | _GEN_1577) & _GEN_4374;
        rob_val_29 <= ~((|_GEN_1612) | _GEN_1579) & _GEN_4375;
        rob_val_30 <= ~((|_GEN_1613) | _GEN_1581) & _GEN_4376;
        rob_val_31 <= ~((|_GEN_1614) | _GEN_1582) & _GEN_4377;
      end
      if (will_commit_1) begin
        rob_val_1_0 <= ~(_GEN_93 | (|_GEN_2513) | _GEN_2481) & _GEN_4378;
        rob_val_1_1 <= ~(_GEN_94 | (|_GEN_2514) | _GEN_2482) & _GEN_4379;
        rob_val_1_2 <= ~(_GEN_95 | (|_GEN_2515) | _GEN_2483) & _GEN_4380;
        rob_val_1_3 <= ~(_GEN_96 | (|_GEN_2516) | _GEN_2484) & _GEN_4381;
        rob_val_1_4 <= ~(_GEN_97 | (|_GEN_2517) | _GEN_2485) & _GEN_4382;
        rob_val_1_5 <= ~(_GEN_98 | (|_GEN_2518) | _GEN_2486) & _GEN_4383;
        rob_val_1_6 <= ~(_GEN_99 | (|_GEN_2519) | _GEN_2487) & _GEN_4384;
        rob_val_1_7 <= ~(_GEN_100 | (|_GEN_2520) | _GEN_2488) & _GEN_4385;
        rob_val_1_8 <= ~(_GEN_101 | (|_GEN_2521) | _GEN_2489) & _GEN_4386;
        rob_val_1_9 <= ~(_GEN_102 | (|_GEN_2522) | _GEN_2490) & _GEN_4387;
        rob_val_1_10 <= ~(_GEN_103 | (|_GEN_2523) | _GEN_2491) & _GEN_4388;
        rob_val_1_11 <= ~(_GEN_104 | (|_GEN_2524) | _GEN_2492) & _GEN_4389;
        rob_val_1_12 <= ~(_GEN_105 | (|_GEN_2525) | _GEN_2493) & _GEN_4390;
        rob_val_1_13 <= ~(_GEN_106 | (|_GEN_2526) | _GEN_2494) & _GEN_4391;
        rob_val_1_14 <= ~(_GEN_107 | (|_GEN_2527) | _GEN_2495) & _GEN_4392;
        rob_val_1_15 <= ~(_GEN_108 | (|_GEN_2528) | _GEN_2496) & _GEN_4393;
        rob_val_1_16 <= ~(_GEN_109 | (|_GEN_2529) | _GEN_2497) & _GEN_4394;
        rob_val_1_17 <= ~(_GEN_110 | (|_GEN_2530) | _GEN_2498) & _GEN_4395;
        rob_val_1_18 <= ~(_GEN_111 | (|_GEN_2531) | _GEN_2499) & _GEN_4396;
        rob_val_1_19 <= ~(_GEN_112 | (|_GEN_2532) | _GEN_2500) & _GEN_4397;
        rob_val_1_20 <= ~(_GEN_113 | (|_GEN_2533) | _GEN_2501) & _GEN_4398;
        rob_val_1_21 <= ~(_GEN_114 | (|_GEN_2534) | _GEN_2502) & _GEN_4399;
        rob_val_1_22 <= ~(_GEN_115 | (|_GEN_2535) | _GEN_2503) & _GEN_4400;
        rob_val_1_23 <= ~(_GEN_116 | (|_GEN_2536) | _GEN_2504) & _GEN_4401;
        rob_val_1_24 <= ~(_GEN_117 | (|_GEN_2537) | _GEN_2505) & _GEN_4402;
        rob_val_1_25 <= ~(_GEN_118 | (|_GEN_2538) | _GEN_2506) & _GEN_4403;
        rob_val_1_26 <= ~(_GEN_119 | (|_GEN_2539) | _GEN_2507) & _GEN_4404;
        rob_val_1_27 <= ~(_GEN_120 | (|_GEN_2540) | _GEN_2508) & _GEN_4405;
        rob_val_1_28 <= ~(_GEN_121 | (|_GEN_2541) | _GEN_2509) & _GEN_4406;
        rob_val_1_29 <= ~(_GEN_122 | (|_GEN_2542) | _GEN_2510) & _GEN_4407;
        rob_val_1_30 <= ~(_GEN_123 | (|_GEN_2543) | _GEN_2511) & _GEN_4408;
        rob_val_1_31 <= ~((&rob_head) | (|_GEN_2544) | _GEN_2512) & _GEN_4409;
      end
      else begin
        rob_val_1_0 <= ~((|_GEN_2513) | _GEN_2481) & _GEN_4378;
        rob_val_1_1 <= ~((|_GEN_2514) | _GEN_2482) & _GEN_4379;
        rob_val_1_2 <= ~((|_GEN_2515) | _GEN_2483) & _GEN_4380;
        rob_val_1_3 <= ~((|_GEN_2516) | _GEN_2484) & _GEN_4381;
        rob_val_1_4 <= ~((|_GEN_2517) | _GEN_2485) & _GEN_4382;
        rob_val_1_5 <= ~((|_GEN_2518) | _GEN_2486) & _GEN_4383;
        rob_val_1_6 <= ~((|_GEN_2519) | _GEN_2487) & _GEN_4384;
        rob_val_1_7 <= ~((|_GEN_2520) | _GEN_2488) & _GEN_4385;
        rob_val_1_8 <= ~((|_GEN_2521) | _GEN_2489) & _GEN_4386;
        rob_val_1_9 <= ~((|_GEN_2522) | _GEN_2490) & _GEN_4387;
        rob_val_1_10 <= ~((|_GEN_2523) | _GEN_2491) & _GEN_4388;
        rob_val_1_11 <= ~((|_GEN_2524) | _GEN_2492) & _GEN_4389;
        rob_val_1_12 <= ~((|_GEN_2525) | _GEN_2493) & _GEN_4390;
        rob_val_1_13 <= ~((|_GEN_2526) | _GEN_2494) & _GEN_4391;
        rob_val_1_14 <= ~((|_GEN_2527) | _GEN_2495) & _GEN_4392;
        rob_val_1_15 <= ~((|_GEN_2528) | _GEN_2496) & _GEN_4393;
        rob_val_1_16 <= ~((|_GEN_2529) | _GEN_2497) & _GEN_4394;
        rob_val_1_17 <= ~((|_GEN_2530) | _GEN_2498) & _GEN_4395;
        rob_val_1_18 <= ~((|_GEN_2531) | _GEN_2499) & _GEN_4396;
        rob_val_1_19 <= ~((|_GEN_2532) | _GEN_2500) & _GEN_4397;
        rob_val_1_20 <= ~((|_GEN_2533) | _GEN_2501) & _GEN_4398;
        rob_val_1_21 <= ~((|_GEN_2534) | _GEN_2502) & _GEN_4399;
        rob_val_1_22 <= ~((|_GEN_2535) | _GEN_2503) & _GEN_4400;
        rob_val_1_23 <= ~((|_GEN_2536) | _GEN_2504) & _GEN_4401;
        rob_val_1_24 <= ~((|_GEN_2537) | _GEN_2505) & _GEN_4402;
        rob_val_1_25 <= ~((|_GEN_2538) | _GEN_2506) & _GEN_4403;
        rob_val_1_26 <= ~((|_GEN_2539) | _GEN_2507) & _GEN_4404;
        rob_val_1_27 <= ~((|_GEN_2540) | _GEN_2508) & _GEN_4405;
        rob_val_1_28 <= ~((|_GEN_2541) | _GEN_2509) & _GEN_4406;
        rob_val_1_29 <= ~((|_GEN_2542) | _GEN_2510) & _GEN_4407;
        rob_val_1_30 <= ~((|_GEN_2543) | _GEN_2511) & _GEN_4408;
        rob_val_1_31 <= ~((|_GEN_2544) | _GEN_2512) & _GEN_4409;
      end
      if (will_commit_2) begin
        rob_val_2_0 <= ~(_GEN_93 | (|_GEN_3412) | _GEN_3380) & _GEN_4410;
        rob_val_2_1 <= ~(_GEN_94 | (|_GEN_3413) | _GEN_3381) & _GEN_4411;
        rob_val_2_2 <= ~(_GEN_95 | (|_GEN_3414) | _GEN_3382) & _GEN_4412;
        rob_val_2_3 <= ~(_GEN_96 | (|_GEN_3415) | _GEN_3383) & _GEN_4413;
        rob_val_2_4 <= ~(_GEN_97 | (|_GEN_3416) | _GEN_3384) & _GEN_4414;
        rob_val_2_5 <= ~(_GEN_98 | (|_GEN_3417) | _GEN_3385) & _GEN_4415;
        rob_val_2_6 <= ~(_GEN_99 | (|_GEN_3418) | _GEN_3386) & _GEN_4416;
        rob_val_2_7 <= ~(_GEN_100 | (|_GEN_3419) | _GEN_3387) & _GEN_4417;
        rob_val_2_8 <= ~(_GEN_101 | (|_GEN_3420) | _GEN_3388) & _GEN_4418;
        rob_val_2_9 <= ~(_GEN_102 | (|_GEN_3421) | _GEN_3389) & _GEN_4419;
        rob_val_2_10 <= ~(_GEN_103 | (|_GEN_3422) | _GEN_3390) & _GEN_4420;
        rob_val_2_11 <= ~(_GEN_104 | (|_GEN_3423) | _GEN_3391) & _GEN_4421;
        rob_val_2_12 <= ~(_GEN_105 | (|_GEN_3424) | _GEN_3392) & _GEN_4422;
        rob_val_2_13 <= ~(_GEN_106 | (|_GEN_3425) | _GEN_3393) & _GEN_4423;
        rob_val_2_14 <= ~(_GEN_107 | (|_GEN_3426) | _GEN_3394) & _GEN_4424;
        rob_val_2_15 <= ~(_GEN_108 | (|_GEN_3427) | _GEN_3395) & _GEN_4425;
        rob_val_2_16 <= ~(_GEN_109 | (|_GEN_3428) | _GEN_3396) & _GEN_4426;
        rob_val_2_17 <= ~(_GEN_110 | (|_GEN_3429) | _GEN_3397) & _GEN_4427;
        rob_val_2_18 <= ~(_GEN_111 | (|_GEN_3430) | _GEN_3398) & _GEN_4428;
        rob_val_2_19 <= ~(_GEN_112 | (|_GEN_3431) | _GEN_3399) & _GEN_4429;
        rob_val_2_20 <= ~(_GEN_113 | (|_GEN_3432) | _GEN_3400) & _GEN_4430;
        rob_val_2_21 <= ~(_GEN_114 | (|_GEN_3433) | _GEN_3401) & _GEN_4431;
        rob_val_2_22 <= ~(_GEN_115 | (|_GEN_3434) | _GEN_3402) & _GEN_4432;
        rob_val_2_23 <= ~(_GEN_116 | (|_GEN_3435) | _GEN_3403) & _GEN_4433;
        rob_val_2_24 <= ~(_GEN_117 | (|_GEN_3436) | _GEN_3404) & _GEN_4434;
        rob_val_2_25 <= ~(_GEN_118 | (|_GEN_3437) | _GEN_3405) & _GEN_4435;
        rob_val_2_26 <= ~(_GEN_119 | (|_GEN_3438) | _GEN_3406) & _GEN_4436;
        rob_val_2_27 <= ~(_GEN_120 | (|_GEN_3439) | _GEN_3407) & _GEN_4437;
        rob_val_2_28 <= ~(_GEN_121 | (|_GEN_3440) | _GEN_3408) & _GEN_4438;
        rob_val_2_29 <= ~(_GEN_122 | (|_GEN_3441) | _GEN_3409) & _GEN_4439;
        rob_val_2_30 <= ~(_GEN_123 | (|_GEN_3442) | _GEN_3410) & _GEN_4440;
        rob_val_2_31 <= ~((&rob_head) | (|_GEN_3443) | _GEN_3411) & _GEN_4441;
      end
      else begin
        rob_val_2_0 <= ~((|_GEN_3412) | _GEN_3380) & _GEN_4410;
        rob_val_2_1 <= ~((|_GEN_3413) | _GEN_3381) & _GEN_4411;
        rob_val_2_2 <= ~((|_GEN_3414) | _GEN_3382) & _GEN_4412;
        rob_val_2_3 <= ~((|_GEN_3415) | _GEN_3383) & _GEN_4413;
        rob_val_2_4 <= ~((|_GEN_3416) | _GEN_3384) & _GEN_4414;
        rob_val_2_5 <= ~((|_GEN_3417) | _GEN_3385) & _GEN_4415;
        rob_val_2_6 <= ~((|_GEN_3418) | _GEN_3386) & _GEN_4416;
        rob_val_2_7 <= ~((|_GEN_3419) | _GEN_3387) & _GEN_4417;
        rob_val_2_8 <= ~((|_GEN_3420) | _GEN_3388) & _GEN_4418;
        rob_val_2_9 <= ~((|_GEN_3421) | _GEN_3389) & _GEN_4419;
        rob_val_2_10 <= ~((|_GEN_3422) | _GEN_3390) & _GEN_4420;
        rob_val_2_11 <= ~((|_GEN_3423) | _GEN_3391) & _GEN_4421;
        rob_val_2_12 <= ~((|_GEN_3424) | _GEN_3392) & _GEN_4422;
        rob_val_2_13 <= ~((|_GEN_3425) | _GEN_3393) & _GEN_4423;
        rob_val_2_14 <= ~((|_GEN_3426) | _GEN_3394) & _GEN_4424;
        rob_val_2_15 <= ~((|_GEN_3427) | _GEN_3395) & _GEN_4425;
        rob_val_2_16 <= ~((|_GEN_3428) | _GEN_3396) & _GEN_4426;
        rob_val_2_17 <= ~((|_GEN_3429) | _GEN_3397) & _GEN_4427;
        rob_val_2_18 <= ~((|_GEN_3430) | _GEN_3398) & _GEN_4428;
        rob_val_2_19 <= ~((|_GEN_3431) | _GEN_3399) & _GEN_4429;
        rob_val_2_20 <= ~((|_GEN_3432) | _GEN_3400) & _GEN_4430;
        rob_val_2_21 <= ~((|_GEN_3433) | _GEN_3401) & _GEN_4431;
        rob_val_2_22 <= ~((|_GEN_3434) | _GEN_3402) & _GEN_4432;
        rob_val_2_23 <= ~((|_GEN_3435) | _GEN_3403) & _GEN_4433;
        rob_val_2_24 <= ~((|_GEN_3436) | _GEN_3404) & _GEN_4434;
        rob_val_2_25 <= ~((|_GEN_3437) | _GEN_3405) & _GEN_4435;
        rob_val_2_26 <= ~((|_GEN_3438) | _GEN_3406) & _GEN_4436;
        rob_val_2_27 <= ~((|_GEN_3439) | _GEN_3407) & _GEN_4437;
        rob_val_2_28 <= ~((|_GEN_3440) | _GEN_3408) & _GEN_4438;
        rob_val_2_29 <= ~((|_GEN_3441) | _GEN_3409) & _GEN_4439;
        rob_val_2_30 <= ~((|_GEN_3442) | _GEN_3410) & _GEN_4440;
        rob_val_2_31 <= ~((|_GEN_3443) | _GEN_3411) & _GEN_4441;
      end
      if (will_commit_3) begin
        rob_val_3_0 <= ~(_GEN_93 | (|_GEN_4311) | _GEN_4279) & _GEN_4442;
        rob_val_3_1 <= ~(_GEN_94 | (|_GEN_4312) | _GEN_4280) & _GEN_4443;
        rob_val_3_2 <= ~(_GEN_95 | (|_GEN_4313) | _GEN_4281) & _GEN_4444;
        rob_val_3_3 <= ~(_GEN_96 | (|_GEN_4314) | _GEN_4282) & _GEN_4445;
        rob_val_3_4 <= ~(_GEN_97 | (|_GEN_4315) | _GEN_4283) & _GEN_4446;
        rob_val_3_5 <= ~(_GEN_98 | (|_GEN_4316) | _GEN_4284) & _GEN_4447;
        rob_val_3_6 <= ~(_GEN_99 | (|_GEN_4317) | _GEN_4285) & _GEN_4448;
        rob_val_3_7 <= ~(_GEN_100 | (|_GEN_4318) | _GEN_4286) & _GEN_4449;
        rob_val_3_8 <= ~(_GEN_101 | (|_GEN_4319) | _GEN_4287) & _GEN_4450;
        rob_val_3_9 <= ~(_GEN_102 | (|_GEN_4320) | _GEN_4288) & _GEN_4451;
        rob_val_3_10 <= ~(_GEN_103 | (|_GEN_4321) | _GEN_4289) & _GEN_4452;
        rob_val_3_11 <= ~(_GEN_104 | (|_GEN_4322) | _GEN_4290) & _GEN_4453;
        rob_val_3_12 <= ~(_GEN_105 | (|_GEN_4323) | _GEN_4291) & _GEN_4454;
        rob_val_3_13 <= ~(_GEN_106 | (|_GEN_4324) | _GEN_4292) & _GEN_4455;
        rob_val_3_14 <= ~(_GEN_107 | (|_GEN_4325) | _GEN_4293) & _GEN_4456;
        rob_val_3_15 <= ~(_GEN_108 | (|_GEN_4326) | _GEN_4294) & _GEN_4457;
        rob_val_3_16 <= ~(_GEN_109 | (|_GEN_4327) | _GEN_4295) & _GEN_4458;
        rob_val_3_17 <= ~(_GEN_110 | (|_GEN_4328) | _GEN_4296) & _GEN_4459;
        rob_val_3_18 <= ~(_GEN_111 | (|_GEN_4329) | _GEN_4297) & _GEN_4460;
        rob_val_3_19 <= ~(_GEN_112 | (|_GEN_4330) | _GEN_4298) & _GEN_4461;
        rob_val_3_20 <= ~(_GEN_113 | (|_GEN_4331) | _GEN_4299) & _GEN_4462;
        rob_val_3_21 <= ~(_GEN_114 | (|_GEN_4332) | _GEN_4300) & _GEN_4463;
        rob_val_3_22 <= ~(_GEN_115 | (|_GEN_4333) | _GEN_4301) & _GEN_4464;
        rob_val_3_23 <= ~(_GEN_116 | (|_GEN_4334) | _GEN_4302) & _GEN_4465;
        rob_val_3_24 <= ~(_GEN_117 | (|_GEN_4335) | _GEN_4303) & _GEN_4466;
        rob_val_3_25 <= ~(_GEN_118 | (|_GEN_4336) | _GEN_4304) & _GEN_4467;
        rob_val_3_26 <= ~(_GEN_119 | (|_GEN_4337) | _GEN_4305) & _GEN_4468;
        rob_val_3_27 <= ~(_GEN_120 | (|_GEN_4338) | _GEN_4306) & _GEN_4469;
        rob_val_3_28 <= ~(_GEN_121 | (|_GEN_4339) | _GEN_4307) & _GEN_4470;
        rob_val_3_29 <= ~(_GEN_122 | (|_GEN_4340) | _GEN_4308) & _GEN_4471;
        rob_val_3_30 <= ~(_GEN_123 | (|_GEN_4341) | _GEN_4309) & _GEN_4472;
        rob_val_3_31 <= ~((&rob_head) | (|_GEN_4342) | _GEN_4310) & _GEN_4473;
      end
      else begin
        rob_val_3_0 <= ~((|_GEN_4311) | _GEN_4279) & _GEN_4442;
        rob_val_3_1 <= ~((|_GEN_4312) | _GEN_4280) & _GEN_4443;
        rob_val_3_2 <= ~((|_GEN_4313) | _GEN_4281) & _GEN_4444;
        rob_val_3_3 <= ~((|_GEN_4314) | _GEN_4282) & _GEN_4445;
        rob_val_3_4 <= ~((|_GEN_4315) | _GEN_4283) & _GEN_4446;
        rob_val_3_5 <= ~((|_GEN_4316) | _GEN_4284) & _GEN_4447;
        rob_val_3_6 <= ~((|_GEN_4317) | _GEN_4285) & _GEN_4448;
        rob_val_3_7 <= ~((|_GEN_4318) | _GEN_4286) & _GEN_4449;
        rob_val_3_8 <= ~((|_GEN_4319) | _GEN_4287) & _GEN_4450;
        rob_val_3_9 <= ~((|_GEN_4320) | _GEN_4288) & _GEN_4451;
        rob_val_3_10 <= ~((|_GEN_4321) | _GEN_4289) & _GEN_4452;
        rob_val_3_11 <= ~((|_GEN_4322) | _GEN_4290) & _GEN_4453;
        rob_val_3_12 <= ~((|_GEN_4323) | _GEN_4291) & _GEN_4454;
        rob_val_3_13 <= ~((|_GEN_4324) | _GEN_4292) & _GEN_4455;
        rob_val_3_14 <= ~((|_GEN_4325) | _GEN_4293) & _GEN_4456;
        rob_val_3_15 <= ~((|_GEN_4326) | _GEN_4294) & _GEN_4457;
        rob_val_3_16 <= ~((|_GEN_4327) | _GEN_4295) & _GEN_4458;
        rob_val_3_17 <= ~((|_GEN_4328) | _GEN_4296) & _GEN_4459;
        rob_val_3_18 <= ~((|_GEN_4329) | _GEN_4297) & _GEN_4460;
        rob_val_3_19 <= ~((|_GEN_4330) | _GEN_4298) & _GEN_4461;
        rob_val_3_20 <= ~((|_GEN_4331) | _GEN_4299) & _GEN_4462;
        rob_val_3_21 <= ~((|_GEN_4332) | _GEN_4300) & _GEN_4463;
        rob_val_3_22 <= ~((|_GEN_4333) | _GEN_4301) & _GEN_4464;
        rob_val_3_23 <= ~((|_GEN_4334) | _GEN_4302) & _GEN_4465;
        rob_val_3_24 <= ~((|_GEN_4335) | _GEN_4303) & _GEN_4466;
        rob_val_3_25 <= ~((|_GEN_4336) | _GEN_4304) & _GEN_4467;
        rob_val_3_26 <= ~((|_GEN_4337) | _GEN_4305) & _GEN_4468;
        rob_val_3_27 <= ~((|_GEN_4338) | _GEN_4306) & _GEN_4469;
        rob_val_3_28 <= ~((|_GEN_4339) | _GEN_4307) & _GEN_4470;
        rob_val_3_29 <= ~((|_GEN_4340) | _GEN_4308) & _GEN_4471;
        rob_val_3_30 <= ~((|_GEN_4341) | _GEN_4309) & _GEN_4472;
        rob_val_3_31 <= ~((|_GEN_4342) | _GEN_4310) & _GEN_4473;
      end
      if (io_enq_valids_0 | io_enq_valids_1 | io_enq_valids_2 | io_enq_valids_3)
        r_partial_row <= io_enq_partial_stall;
      pnr_maybe_at_tail <= ~rob_deq & (do_inc_row | pnr_maybe_at_tail);
    end
    r_xcpt_uop_br_mask <= next_xcpt_uop_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_4343) begin
      if (io_lxcpt_valid) begin
        if (_GEN_4344) begin
          r_xcpt_uop_rob_idx <= io_lxcpt_bits_uop_rob_idx;
          r_xcpt_uop_exc_cause <= {59'h0, io_lxcpt_bits_cause};
          r_xcpt_badvaddr <= io_lxcpt_bits_badvaddr;
        end
      end
      else if (_GEN_4345) begin
        r_xcpt_uop_rob_idx <= casez_tmp_313;
        r_xcpt_uop_exc_cause <= casez_tmp_314;
        r_xcpt_badvaddr <= {io_xcpt_fetch_pc[39:6], casez_tmp_312};
      end
    end
    if (_GEN_1457 & _GEN_1458)
      rob_fflags_0_0 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1426)
      rob_fflags_0_0 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1394)
      rob_fflags_0_0 <= io_fflags_0_bits_flags;
    else if (_GEN_128)
      rob_fflags_0_0 <= 5'h0;
    if (_GEN_1457 & _GEN_1459)
      rob_fflags_0_1 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1427)
      rob_fflags_0_1 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1395)
      rob_fflags_0_1 <= io_fflags_0_bits_flags;
    else if (_GEN_130)
      rob_fflags_0_1 <= 5'h0;
    if (_GEN_1457 & _GEN_1460)
      rob_fflags_0_2 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1428)
      rob_fflags_0_2 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1396)
      rob_fflags_0_2 <= io_fflags_0_bits_flags;
    else if (_GEN_132)
      rob_fflags_0_2 <= 5'h0;
    if (_GEN_1457 & _GEN_1461)
      rob_fflags_0_3 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1429)
      rob_fflags_0_3 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1397)
      rob_fflags_0_3 <= io_fflags_0_bits_flags;
    else if (_GEN_134)
      rob_fflags_0_3 <= 5'h0;
    if (_GEN_1457 & _GEN_1462)
      rob_fflags_0_4 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1430)
      rob_fflags_0_4 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1398)
      rob_fflags_0_4 <= io_fflags_0_bits_flags;
    else if (_GEN_136)
      rob_fflags_0_4 <= 5'h0;
    if (_GEN_1457 & _GEN_1463)
      rob_fflags_0_5 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1431)
      rob_fflags_0_5 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1399)
      rob_fflags_0_5 <= io_fflags_0_bits_flags;
    else if (_GEN_138)
      rob_fflags_0_5 <= 5'h0;
    if (_GEN_1457 & _GEN_1464)
      rob_fflags_0_6 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1432)
      rob_fflags_0_6 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1400)
      rob_fflags_0_6 <= io_fflags_0_bits_flags;
    else if (_GEN_140)
      rob_fflags_0_6 <= 5'h0;
    if (_GEN_1457 & _GEN_1465)
      rob_fflags_0_7 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1433)
      rob_fflags_0_7 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1401)
      rob_fflags_0_7 <= io_fflags_0_bits_flags;
    else if (_GEN_142)
      rob_fflags_0_7 <= 5'h0;
    if (_GEN_1457 & _GEN_1466)
      rob_fflags_0_8 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1434)
      rob_fflags_0_8 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1402)
      rob_fflags_0_8 <= io_fflags_0_bits_flags;
    else if (_GEN_144)
      rob_fflags_0_8 <= 5'h0;
    if (_GEN_1457 & _GEN_1467)
      rob_fflags_0_9 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1435)
      rob_fflags_0_9 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1403)
      rob_fflags_0_9 <= io_fflags_0_bits_flags;
    else if (_GEN_146)
      rob_fflags_0_9 <= 5'h0;
    if (_GEN_1457 & _GEN_1468)
      rob_fflags_0_10 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1436)
      rob_fflags_0_10 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1404)
      rob_fflags_0_10 <= io_fflags_0_bits_flags;
    else if (_GEN_148)
      rob_fflags_0_10 <= 5'h0;
    if (_GEN_1457 & _GEN_1469)
      rob_fflags_0_11 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1437)
      rob_fflags_0_11 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1405)
      rob_fflags_0_11 <= io_fflags_0_bits_flags;
    else if (_GEN_150)
      rob_fflags_0_11 <= 5'h0;
    if (_GEN_1457 & _GEN_1470)
      rob_fflags_0_12 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1438)
      rob_fflags_0_12 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1406)
      rob_fflags_0_12 <= io_fflags_0_bits_flags;
    else if (_GEN_152)
      rob_fflags_0_12 <= 5'h0;
    if (_GEN_1457 & _GEN_1471)
      rob_fflags_0_13 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1439)
      rob_fflags_0_13 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1407)
      rob_fflags_0_13 <= io_fflags_0_bits_flags;
    else if (_GEN_154)
      rob_fflags_0_13 <= 5'h0;
    if (_GEN_1457 & _GEN_1472)
      rob_fflags_0_14 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1440)
      rob_fflags_0_14 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1408)
      rob_fflags_0_14 <= io_fflags_0_bits_flags;
    else if (_GEN_156)
      rob_fflags_0_14 <= 5'h0;
    if (_GEN_1457 & _GEN_1473)
      rob_fflags_0_15 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1441)
      rob_fflags_0_15 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1409)
      rob_fflags_0_15 <= io_fflags_0_bits_flags;
    else if (_GEN_158)
      rob_fflags_0_15 <= 5'h0;
    if (_GEN_1457 & _GEN_1474)
      rob_fflags_0_16 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1442)
      rob_fflags_0_16 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1410)
      rob_fflags_0_16 <= io_fflags_0_bits_flags;
    else if (_GEN_160)
      rob_fflags_0_16 <= 5'h0;
    if (_GEN_1457 & _GEN_1475)
      rob_fflags_0_17 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1443)
      rob_fflags_0_17 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1411)
      rob_fflags_0_17 <= io_fflags_0_bits_flags;
    else if (_GEN_162)
      rob_fflags_0_17 <= 5'h0;
    if (_GEN_1457 & _GEN_1476)
      rob_fflags_0_18 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1444)
      rob_fflags_0_18 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1412)
      rob_fflags_0_18 <= io_fflags_0_bits_flags;
    else if (_GEN_164)
      rob_fflags_0_18 <= 5'h0;
    if (_GEN_1457 & _GEN_1477)
      rob_fflags_0_19 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1445)
      rob_fflags_0_19 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1413)
      rob_fflags_0_19 <= io_fflags_0_bits_flags;
    else if (_GEN_166)
      rob_fflags_0_19 <= 5'h0;
    if (_GEN_1457 & _GEN_1478)
      rob_fflags_0_20 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1446)
      rob_fflags_0_20 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1414)
      rob_fflags_0_20 <= io_fflags_0_bits_flags;
    else if (_GEN_168)
      rob_fflags_0_20 <= 5'h0;
    if (_GEN_1457 & _GEN_1479)
      rob_fflags_0_21 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1447)
      rob_fflags_0_21 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1415)
      rob_fflags_0_21 <= io_fflags_0_bits_flags;
    else if (_GEN_170)
      rob_fflags_0_21 <= 5'h0;
    if (_GEN_1457 & _GEN_1480)
      rob_fflags_0_22 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1448)
      rob_fflags_0_22 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1416)
      rob_fflags_0_22 <= io_fflags_0_bits_flags;
    else if (_GEN_172)
      rob_fflags_0_22 <= 5'h0;
    if (_GEN_1457 & _GEN_1481)
      rob_fflags_0_23 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1449)
      rob_fflags_0_23 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1417)
      rob_fflags_0_23 <= io_fflags_0_bits_flags;
    else if (_GEN_174)
      rob_fflags_0_23 <= 5'h0;
    if (_GEN_1457 & _GEN_1482)
      rob_fflags_0_24 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1450)
      rob_fflags_0_24 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1418)
      rob_fflags_0_24 <= io_fflags_0_bits_flags;
    else if (_GEN_176)
      rob_fflags_0_24 <= 5'h0;
    if (_GEN_1457 & _GEN_1483)
      rob_fflags_0_25 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1451)
      rob_fflags_0_25 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1419)
      rob_fflags_0_25 <= io_fflags_0_bits_flags;
    else if (_GEN_178)
      rob_fflags_0_25 <= 5'h0;
    if (_GEN_1457 & _GEN_1484)
      rob_fflags_0_26 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1452)
      rob_fflags_0_26 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1420)
      rob_fflags_0_26 <= io_fflags_0_bits_flags;
    else if (_GEN_180)
      rob_fflags_0_26 <= 5'h0;
    if (_GEN_1457 & _GEN_1485)
      rob_fflags_0_27 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1453)
      rob_fflags_0_27 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1421)
      rob_fflags_0_27 <= io_fflags_0_bits_flags;
    else if (_GEN_182)
      rob_fflags_0_27 <= 5'h0;
    if (_GEN_1457 & _GEN_1486)
      rob_fflags_0_28 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1454)
      rob_fflags_0_28 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1422)
      rob_fflags_0_28 <= io_fflags_0_bits_flags;
    else if (_GEN_184)
      rob_fflags_0_28 <= 5'h0;
    if (_GEN_1457 & _GEN_1487)
      rob_fflags_0_29 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1455)
      rob_fflags_0_29 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1423)
      rob_fflags_0_29 <= io_fflags_0_bits_flags;
    else if (_GEN_186)
      rob_fflags_0_29 <= 5'h0;
    if (_GEN_1457 & _GEN_1488)
      rob_fflags_0_30 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & _GEN_1456)
      rob_fflags_0_30 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & _GEN_1424)
      rob_fflags_0_30 <= io_fflags_0_bits_flags;
    else if (_GEN_188)
      rob_fflags_0_30 <= 5'h0;
    if (_GEN_1457 & (&(io_fflags_3_bits_uop_rob_idx[6:2])))
      rob_fflags_0_31 <= io_fflags_3_bits_flags;
    else if (_GEN_1425 & (&(io_fflags_2_bits_uop_rob_idx[6:2])))
      rob_fflags_0_31 <= io_fflags_2_bits_flags;
    else if (_GEN_1393 & (&(io_fflags_0_bits_uop_rob_idx[6:2])))
      rob_fflags_0_31 <= io_fflags_0_bits_flags;
    else if (_GEN_189)
      rob_fflags_0_31 <= 5'h0;
    if (_GEN_2480 & _GEN_1458)
      rob_fflags_1_0 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1426)
      rob_fflags_1_0 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1394)
      rob_fflags_1_0 <= io_fflags_0_bits_flags;
    else if (_GEN_1646)
      rob_fflags_1_0 <= 5'h0;
    if (_GEN_2480 & _GEN_1459)
      rob_fflags_1_1 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1427)
      rob_fflags_1_1 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1395)
      rob_fflags_1_1 <= io_fflags_0_bits_flags;
    else if (_GEN_1647)
      rob_fflags_1_1 <= 5'h0;
    if (_GEN_2480 & _GEN_1460)
      rob_fflags_1_2 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1428)
      rob_fflags_1_2 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1396)
      rob_fflags_1_2 <= io_fflags_0_bits_flags;
    else if (_GEN_1648)
      rob_fflags_1_2 <= 5'h0;
    if (_GEN_2480 & _GEN_1461)
      rob_fflags_1_3 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1429)
      rob_fflags_1_3 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1397)
      rob_fflags_1_3 <= io_fflags_0_bits_flags;
    else if (_GEN_1649)
      rob_fflags_1_3 <= 5'h0;
    if (_GEN_2480 & _GEN_1462)
      rob_fflags_1_4 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1430)
      rob_fflags_1_4 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1398)
      rob_fflags_1_4 <= io_fflags_0_bits_flags;
    else if (_GEN_1650)
      rob_fflags_1_4 <= 5'h0;
    if (_GEN_2480 & _GEN_1463)
      rob_fflags_1_5 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1431)
      rob_fflags_1_5 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1399)
      rob_fflags_1_5 <= io_fflags_0_bits_flags;
    else if (_GEN_1651)
      rob_fflags_1_5 <= 5'h0;
    if (_GEN_2480 & _GEN_1464)
      rob_fflags_1_6 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1432)
      rob_fflags_1_6 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1400)
      rob_fflags_1_6 <= io_fflags_0_bits_flags;
    else if (_GEN_1652)
      rob_fflags_1_6 <= 5'h0;
    if (_GEN_2480 & _GEN_1465)
      rob_fflags_1_7 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1433)
      rob_fflags_1_7 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1401)
      rob_fflags_1_7 <= io_fflags_0_bits_flags;
    else if (_GEN_1653)
      rob_fflags_1_7 <= 5'h0;
    if (_GEN_2480 & _GEN_1466)
      rob_fflags_1_8 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1434)
      rob_fflags_1_8 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1402)
      rob_fflags_1_8 <= io_fflags_0_bits_flags;
    else if (_GEN_1654)
      rob_fflags_1_8 <= 5'h0;
    if (_GEN_2480 & _GEN_1467)
      rob_fflags_1_9 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1435)
      rob_fflags_1_9 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1403)
      rob_fflags_1_9 <= io_fflags_0_bits_flags;
    else if (_GEN_1655)
      rob_fflags_1_9 <= 5'h0;
    if (_GEN_2480 & _GEN_1468)
      rob_fflags_1_10 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1436)
      rob_fflags_1_10 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1404)
      rob_fflags_1_10 <= io_fflags_0_bits_flags;
    else if (_GEN_1656)
      rob_fflags_1_10 <= 5'h0;
    if (_GEN_2480 & _GEN_1469)
      rob_fflags_1_11 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1437)
      rob_fflags_1_11 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1405)
      rob_fflags_1_11 <= io_fflags_0_bits_flags;
    else if (_GEN_1657)
      rob_fflags_1_11 <= 5'h0;
    if (_GEN_2480 & _GEN_1470)
      rob_fflags_1_12 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1438)
      rob_fflags_1_12 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1406)
      rob_fflags_1_12 <= io_fflags_0_bits_flags;
    else if (_GEN_1658)
      rob_fflags_1_12 <= 5'h0;
    if (_GEN_2480 & _GEN_1471)
      rob_fflags_1_13 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1439)
      rob_fflags_1_13 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1407)
      rob_fflags_1_13 <= io_fflags_0_bits_flags;
    else if (_GEN_1659)
      rob_fflags_1_13 <= 5'h0;
    if (_GEN_2480 & _GEN_1472)
      rob_fflags_1_14 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1440)
      rob_fflags_1_14 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1408)
      rob_fflags_1_14 <= io_fflags_0_bits_flags;
    else if (_GEN_1660)
      rob_fflags_1_14 <= 5'h0;
    if (_GEN_2480 & _GEN_1473)
      rob_fflags_1_15 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1441)
      rob_fflags_1_15 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1409)
      rob_fflags_1_15 <= io_fflags_0_bits_flags;
    else if (_GEN_1661)
      rob_fflags_1_15 <= 5'h0;
    if (_GEN_2480 & _GEN_1474)
      rob_fflags_1_16 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1442)
      rob_fflags_1_16 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1410)
      rob_fflags_1_16 <= io_fflags_0_bits_flags;
    else if (_GEN_1662)
      rob_fflags_1_16 <= 5'h0;
    if (_GEN_2480 & _GEN_1475)
      rob_fflags_1_17 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1443)
      rob_fflags_1_17 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1411)
      rob_fflags_1_17 <= io_fflags_0_bits_flags;
    else if (_GEN_1663)
      rob_fflags_1_17 <= 5'h0;
    if (_GEN_2480 & _GEN_1476)
      rob_fflags_1_18 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1444)
      rob_fflags_1_18 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1412)
      rob_fflags_1_18 <= io_fflags_0_bits_flags;
    else if (_GEN_1664)
      rob_fflags_1_18 <= 5'h0;
    if (_GEN_2480 & _GEN_1477)
      rob_fflags_1_19 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1445)
      rob_fflags_1_19 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1413)
      rob_fflags_1_19 <= io_fflags_0_bits_flags;
    else if (_GEN_1665)
      rob_fflags_1_19 <= 5'h0;
    if (_GEN_2480 & _GEN_1478)
      rob_fflags_1_20 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1446)
      rob_fflags_1_20 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1414)
      rob_fflags_1_20 <= io_fflags_0_bits_flags;
    else if (_GEN_1666)
      rob_fflags_1_20 <= 5'h0;
    if (_GEN_2480 & _GEN_1479)
      rob_fflags_1_21 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1447)
      rob_fflags_1_21 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1415)
      rob_fflags_1_21 <= io_fflags_0_bits_flags;
    else if (_GEN_1667)
      rob_fflags_1_21 <= 5'h0;
    if (_GEN_2480 & _GEN_1480)
      rob_fflags_1_22 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1448)
      rob_fflags_1_22 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1416)
      rob_fflags_1_22 <= io_fflags_0_bits_flags;
    else if (_GEN_1668)
      rob_fflags_1_22 <= 5'h0;
    if (_GEN_2480 & _GEN_1481)
      rob_fflags_1_23 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1449)
      rob_fflags_1_23 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1417)
      rob_fflags_1_23 <= io_fflags_0_bits_flags;
    else if (_GEN_1669)
      rob_fflags_1_23 <= 5'h0;
    if (_GEN_2480 & _GEN_1482)
      rob_fflags_1_24 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1450)
      rob_fflags_1_24 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1418)
      rob_fflags_1_24 <= io_fflags_0_bits_flags;
    else if (_GEN_1670)
      rob_fflags_1_24 <= 5'h0;
    if (_GEN_2480 & _GEN_1483)
      rob_fflags_1_25 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1451)
      rob_fflags_1_25 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1419)
      rob_fflags_1_25 <= io_fflags_0_bits_flags;
    else if (_GEN_1671)
      rob_fflags_1_25 <= 5'h0;
    if (_GEN_2480 & _GEN_1484)
      rob_fflags_1_26 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1452)
      rob_fflags_1_26 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1420)
      rob_fflags_1_26 <= io_fflags_0_bits_flags;
    else if (_GEN_1672)
      rob_fflags_1_26 <= 5'h0;
    if (_GEN_2480 & _GEN_1485)
      rob_fflags_1_27 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1453)
      rob_fflags_1_27 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1421)
      rob_fflags_1_27 <= io_fflags_0_bits_flags;
    else if (_GEN_1673)
      rob_fflags_1_27 <= 5'h0;
    if (_GEN_2480 & _GEN_1486)
      rob_fflags_1_28 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1454)
      rob_fflags_1_28 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1422)
      rob_fflags_1_28 <= io_fflags_0_bits_flags;
    else if (_GEN_1674)
      rob_fflags_1_28 <= 5'h0;
    if (_GEN_2480 & _GEN_1487)
      rob_fflags_1_29 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1455)
      rob_fflags_1_29 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1423)
      rob_fflags_1_29 <= io_fflags_0_bits_flags;
    else if (_GEN_1675)
      rob_fflags_1_29 <= 5'h0;
    if (_GEN_2480 & _GEN_1488)
      rob_fflags_1_30 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & _GEN_1456)
      rob_fflags_1_30 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & _GEN_1424)
      rob_fflags_1_30 <= io_fflags_0_bits_flags;
    else if (_GEN_1676)
      rob_fflags_1_30 <= 5'h0;
    if (_GEN_2480 & (&(io_fflags_3_bits_uop_rob_idx[6:2])))
      rob_fflags_1_31 <= io_fflags_3_bits_flags;
    else if (_GEN_2479 & (&(io_fflags_2_bits_uop_rob_idx[6:2])))
      rob_fflags_1_31 <= io_fflags_2_bits_flags;
    else if (_GEN_2478 & (&(io_fflags_0_bits_uop_rob_idx[6:2])))
      rob_fflags_1_31 <= io_fflags_0_bits_flags;
    else if (_GEN_1677)
      rob_fflags_1_31 <= 5'h0;
    if (_GEN_3379 & _GEN_1458)
      rob_fflags_2_0 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1426)
      rob_fflags_2_0 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1394)
      rob_fflags_2_0 <= io_fflags_0_bits_flags;
    else if (_GEN_2545)
      rob_fflags_2_0 <= 5'h0;
    if (_GEN_3379 & _GEN_1459)
      rob_fflags_2_1 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1427)
      rob_fflags_2_1 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1395)
      rob_fflags_2_1 <= io_fflags_0_bits_flags;
    else if (_GEN_2546)
      rob_fflags_2_1 <= 5'h0;
    if (_GEN_3379 & _GEN_1460)
      rob_fflags_2_2 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1428)
      rob_fflags_2_2 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1396)
      rob_fflags_2_2 <= io_fflags_0_bits_flags;
    else if (_GEN_2547)
      rob_fflags_2_2 <= 5'h0;
    if (_GEN_3379 & _GEN_1461)
      rob_fflags_2_3 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1429)
      rob_fflags_2_3 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1397)
      rob_fflags_2_3 <= io_fflags_0_bits_flags;
    else if (_GEN_2548)
      rob_fflags_2_3 <= 5'h0;
    if (_GEN_3379 & _GEN_1462)
      rob_fflags_2_4 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1430)
      rob_fflags_2_4 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1398)
      rob_fflags_2_4 <= io_fflags_0_bits_flags;
    else if (_GEN_2549)
      rob_fflags_2_4 <= 5'h0;
    if (_GEN_3379 & _GEN_1463)
      rob_fflags_2_5 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1431)
      rob_fflags_2_5 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1399)
      rob_fflags_2_5 <= io_fflags_0_bits_flags;
    else if (_GEN_2550)
      rob_fflags_2_5 <= 5'h0;
    if (_GEN_3379 & _GEN_1464)
      rob_fflags_2_6 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1432)
      rob_fflags_2_6 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1400)
      rob_fflags_2_6 <= io_fflags_0_bits_flags;
    else if (_GEN_2551)
      rob_fflags_2_6 <= 5'h0;
    if (_GEN_3379 & _GEN_1465)
      rob_fflags_2_7 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1433)
      rob_fflags_2_7 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1401)
      rob_fflags_2_7 <= io_fflags_0_bits_flags;
    else if (_GEN_2552)
      rob_fflags_2_7 <= 5'h0;
    if (_GEN_3379 & _GEN_1466)
      rob_fflags_2_8 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1434)
      rob_fflags_2_8 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1402)
      rob_fflags_2_8 <= io_fflags_0_bits_flags;
    else if (_GEN_2553)
      rob_fflags_2_8 <= 5'h0;
    if (_GEN_3379 & _GEN_1467)
      rob_fflags_2_9 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1435)
      rob_fflags_2_9 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1403)
      rob_fflags_2_9 <= io_fflags_0_bits_flags;
    else if (_GEN_2554)
      rob_fflags_2_9 <= 5'h0;
    if (_GEN_3379 & _GEN_1468)
      rob_fflags_2_10 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1436)
      rob_fflags_2_10 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1404)
      rob_fflags_2_10 <= io_fflags_0_bits_flags;
    else if (_GEN_2555)
      rob_fflags_2_10 <= 5'h0;
    if (_GEN_3379 & _GEN_1469)
      rob_fflags_2_11 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1437)
      rob_fflags_2_11 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1405)
      rob_fflags_2_11 <= io_fflags_0_bits_flags;
    else if (_GEN_2556)
      rob_fflags_2_11 <= 5'h0;
    if (_GEN_3379 & _GEN_1470)
      rob_fflags_2_12 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1438)
      rob_fflags_2_12 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1406)
      rob_fflags_2_12 <= io_fflags_0_bits_flags;
    else if (_GEN_2557)
      rob_fflags_2_12 <= 5'h0;
    if (_GEN_3379 & _GEN_1471)
      rob_fflags_2_13 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1439)
      rob_fflags_2_13 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1407)
      rob_fflags_2_13 <= io_fflags_0_bits_flags;
    else if (_GEN_2558)
      rob_fflags_2_13 <= 5'h0;
    if (_GEN_3379 & _GEN_1472)
      rob_fflags_2_14 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1440)
      rob_fflags_2_14 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1408)
      rob_fflags_2_14 <= io_fflags_0_bits_flags;
    else if (_GEN_2559)
      rob_fflags_2_14 <= 5'h0;
    if (_GEN_3379 & _GEN_1473)
      rob_fflags_2_15 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1441)
      rob_fflags_2_15 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1409)
      rob_fflags_2_15 <= io_fflags_0_bits_flags;
    else if (_GEN_2560)
      rob_fflags_2_15 <= 5'h0;
    if (_GEN_3379 & _GEN_1474)
      rob_fflags_2_16 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1442)
      rob_fflags_2_16 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1410)
      rob_fflags_2_16 <= io_fflags_0_bits_flags;
    else if (_GEN_2561)
      rob_fflags_2_16 <= 5'h0;
    if (_GEN_3379 & _GEN_1475)
      rob_fflags_2_17 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1443)
      rob_fflags_2_17 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1411)
      rob_fflags_2_17 <= io_fflags_0_bits_flags;
    else if (_GEN_2562)
      rob_fflags_2_17 <= 5'h0;
    if (_GEN_3379 & _GEN_1476)
      rob_fflags_2_18 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1444)
      rob_fflags_2_18 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1412)
      rob_fflags_2_18 <= io_fflags_0_bits_flags;
    else if (_GEN_2563)
      rob_fflags_2_18 <= 5'h0;
    if (_GEN_3379 & _GEN_1477)
      rob_fflags_2_19 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1445)
      rob_fflags_2_19 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1413)
      rob_fflags_2_19 <= io_fflags_0_bits_flags;
    else if (_GEN_2564)
      rob_fflags_2_19 <= 5'h0;
    if (_GEN_3379 & _GEN_1478)
      rob_fflags_2_20 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1446)
      rob_fflags_2_20 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1414)
      rob_fflags_2_20 <= io_fflags_0_bits_flags;
    else if (_GEN_2565)
      rob_fflags_2_20 <= 5'h0;
    if (_GEN_3379 & _GEN_1479)
      rob_fflags_2_21 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1447)
      rob_fflags_2_21 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1415)
      rob_fflags_2_21 <= io_fflags_0_bits_flags;
    else if (_GEN_2566)
      rob_fflags_2_21 <= 5'h0;
    if (_GEN_3379 & _GEN_1480)
      rob_fflags_2_22 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1448)
      rob_fflags_2_22 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1416)
      rob_fflags_2_22 <= io_fflags_0_bits_flags;
    else if (_GEN_2567)
      rob_fflags_2_22 <= 5'h0;
    if (_GEN_3379 & _GEN_1481)
      rob_fflags_2_23 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1449)
      rob_fflags_2_23 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1417)
      rob_fflags_2_23 <= io_fflags_0_bits_flags;
    else if (_GEN_2568)
      rob_fflags_2_23 <= 5'h0;
    if (_GEN_3379 & _GEN_1482)
      rob_fflags_2_24 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1450)
      rob_fflags_2_24 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1418)
      rob_fflags_2_24 <= io_fflags_0_bits_flags;
    else if (_GEN_2569)
      rob_fflags_2_24 <= 5'h0;
    if (_GEN_3379 & _GEN_1483)
      rob_fflags_2_25 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1451)
      rob_fflags_2_25 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1419)
      rob_fflags_2_25 <= io_fflags_0_bits_flags;
    else if (_GEN_2570)
      rob_fflags_2_25 <= 5'h0;
    if (_GEN_3379 & _GEN_1484)
      rob_fflags_2_26 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1452)
      rob_fflags_2_26 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1420)
      rob_fflags_2_26 <= io_fflags_0_bits_flags;
    else if (_GEN_2571)
      rob_fflags_2_26 <= 5'h0;
    if (_GEN_3379 & _GEN_1485)
      rob_fflags_2_27 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1453)
      rob_fflags_2_27 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1421)
      rob_fflags_2_27 <= io_fflags_0_bits_flags;
    else if (_GEN_2572)
      rob_fflags_2_27 <= 5'h0;
    if (_GEN_3379 & _GEN_1486)
      rob_fflags_2_28 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1454)
      rob_fflags_2_28 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1422)
      rob_fflags_2_28 <= io_fflags_0_bits_flags;
    else if (_GEN_2573)
      rob_fflags_2_28 <= 5'h0;
    if (_GEN_3379 & _GEN_1487)
      rob_fflags_2_29 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1455)
      rob_fflags_2_29 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1423)
      rob_fflags_2_29 <= io_fflags_0_bits_flags;
    else if (_GEN_2574)
      rob_fflags_2_29 <= 5'h0;
    if (_GEN_3379 & _GEN_1488)
      rob_fflags_2_30 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & _GEN_1456)
      rob_fflags_2_30 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & _GEN_1424)
      rob_fflags_2_30 <= io_fflags_0_bits_flags;
    else if (_GEN_2575)
      rob_fflags_2_30 <= 5'h0;
    if (_GEN_3379 & (&(io_fflags_3_bits_uop_rob_idx[6:2])))
      rob_fflags_2_31 <= io_fflags_3_bits_flags;
    else if (_GEN_3378 & (&(io_fflags_2_bits_uop_rob_idx[6:2])))
      rob_fflags_2_31 <= io_fflags_2_bits_flags;
    else if (_GEN_3377 & (&(io_fflags_0_bits_uop_rob_idx[6:2])))
      rob_fflags_2_31 <= io_fflags_0_bits_flags;
    else if (_GEN_2576)
      rob_fflags_2_31 <= 5'h0;
    if (_GEN_4278 & _GEN_1458)
      rob_fflags_3_0 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1426)
      rob_fflags_3_0 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1394)
      rob_fflags_3_0 <= io_fflags_0_bits_flags;
    else if (_GEN_3444)
      rob_fflags_3_0 <= 5'h0;
    if (_GEN_4278 & _GEN_1459)
      rob_fflags_3_1 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1427)
      rob_fflags_3_1 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1395)
      rob_fflags_3_1 <= io_fflags_0_bits_flags;
    else if (_GEN_3445)
      rob_fflags_3_1 <= 5'h0;
    if (_GEN_4278 & _GEN_1460)
      rob_fflags_3_2 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1428)
      rob_fflags_3_2 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1396)
      rob_fflags_3_2 <= io_fflags_0_bits_flags;
    else if (_GEN_3446)
      rob_fflags_3_2 <= 5'h0;
    if (_GEN_4278 & _GEN_1461)
      rob_fflags_3_3 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1429)
      rob_fflags_3_3 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1397)
      rob_fflags_3_3 <= io_fflags_0_bits_flags;
    else if (_GEN_3447)
      rob_fflags_3_3 <= 5'h0;
    if (_GEN_4278 & _GEN_1462)
      rob_fflags_3_4 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1430)
      rob_fflags_3_4 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1398)
      rob_fflags_3_4 <= io_fflags_0_bits_flags;
    else if (_GEN_3448)
      rob_fflags_3_4 <= 5'h0;
    if (_GEN_4278 & _GEN_1463)
      rob_fflags_3_5 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1431)
      rob_fflags_3_5 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1399)
      rob_fflags_3_5 <= io_fflags_0_bits_flags;
    else if (_GEN_3449)
      rob_fflags_3_5 <= 5'h0;
    if (_GEN_4278 & _GEN_1464)
      rob_fflags_3_6 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1432)
      rob_fflags_3_6 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1400)
      rob_fflags_3_6 <= io_fflags_0_bits_flags;
    else if (_GEN_3450)
      rob_fflags_3_6 <= 5'h0;
    if (_GEN_4278 & _GEN_1465)
      rob_fflags_3_7 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1433)
      rob_fflags_3_7 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1401)
      rob_fflags_3_7 <= io_fflags_0_bits_flags;
    else if (_GEN_3451)
      rob_fflags_3_7 <= 5'h0;
    if (_GEN_4278 & _GEN_1466)
      rob_fflags_3_8 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1434)
      rob_fflags_3_8 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1402)
      rob_fflags_3_8 <= io_fflags_0_bits_flags;
    else if (_GEN_3452)
      rob_fflags_3_8 <= 5'h0;
    if (_GEN_4278 & _GEN_1467)
      rob_fflags_3_9 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1435)
      rob_fflags_3_9 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1403)
      rob_fflags_3_9 <= io_fflags_0_bits_flags;
    else if (_GEN_3453)
      rob_fflags_3_9 <= 5'h0;
    if (_GEN_4278 & _GEN_1468)
      rob_fflags_3_10 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1436)
      rob_fflags_3_10 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1404)
      rob_fflags_3_10 <= io_fflags_0_bits_flags;
    else if (_GEN_3454)
      rob_fflags_3_10 <= 5'h0;
    if (_GEN_4278 & _GEN_1469)
      rob_fflags_3_11 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1437)
      rob_fflags_3_11 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1405)
      rob_fflags_3_11 <= io_fflags_0_bits_flags;
    else if (_GEN_3455)
      rob_fflags_3_11 <= 5'h0;
    if (_GEN_4278 & _GEN_1470)
      rob_fflags_3_12 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1438)
      rob_fflags_3_12 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1406)
      rob_fflags_3_12 <= io_fflags_0_bits_flags;
    else if (_GEN_3456)
      rob_fflags_3_12 <= 5'h0;
    if (_GEN_4278 & _GEN_1471)
      rob_fflags_3_13 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1439)
      rob_fflags_3_13 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1407)
      rob_fflags_3_13 <= io_fflags_0_bits_flags;
    else if (_GEN_3457)
      rob_fflags_3_13 <= 5'h0;
    if (_GEN_4278 & _GEN_1472)
      rob_fflags_3_14 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1440)
      rob_fflags_3_14 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1408)
      rob_fflags_3_14 <= io_fflags_0_bits_flags;
    else if (_GEN_3458)
      rob_fflags_3_14 <= 5'h0;
    if (_GEN_4278 & _GEN_1473)
      rob_fflags_3_15 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1441)
      rob_fflags_3_15 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1409)
      rob_fflags_3_15 <= io_fflags_0_bits_flags;
    else if (_GEN_3459)
      rob_fflags_3_15 <= 5'h0;
    if (_GEN_4278 & _GEN_1474)
      rob_fflags_3_16 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1442)
      rob_fflags_3_16 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1410)
      rob_fflags_3_16 <= io_fflags_0_bits_flags;
    else if (_GEN_3460)
      rob_fflags_3_16 <= 5'h0;
    if (_GEN_4278 & _GEN_1475)
      rob_fflags_3_17 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1443)
      rob_fflags_3_17 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1411)
      rob_fflags_3_17 <= io_fflags_0_bits_flags;
    else if (_GEN_3461)
      rob_fflags_3_17 <= 5'h0;
    if (_GEN_4278 & _GEN_1476)
      rob_fflags_3_18 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1444)
      rob_fflags_3_18 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1412)
      rob_fflags_3_18 <= io_fflags_0_bits_flags;
    else if (_GEN_3462)
      rob_fflags_3_18 <= 5'h0;
    if (_GEN_4278 & _GEN_1477)
      rob_fflags_3_19 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1445)
      rob_fflags_3_19 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1413)
      rob_fflags_3_19 <= io_fflags_0_bits_flags;
    else if (_GEN_3463)
      rob_fflags_3_19 <= 5'h0;
    if (_GEN_4278 & _GEN_1478)
      rob_fflags_3_20 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1446)
      rob_fflags_3_20 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1414)
      rob_fflags_3_20 <= io_fflags_0_bits_flags;
    else if (_GEN_3464)
      rob_fflags_3_20 <= 5'h0;
    if (_GEN_4278 & _GEN_1479)
      rob_fflags_3_21 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1447)
      rob_fflags_3_21 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1415)
      rob_fflags_3_21 <= io_fflags_0_bits_flags;
    else if (_GEN_3465)
      rob_fflags_3_21 <= 5'h0;
    if (_GEN_4278 & _GEN_1480)
      rob_fflags_3_22 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1448)
      rob_fflags_3_22 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1416)
      rob_fflags_3_22 <= io_fflags_0_bits_flags;
    else if (_GEN_3466)
      rob_fflags_3_22 <= 5'h0;
    if (_GEN_4278 & _GEN_1481)
      rob_fflags_3_23 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1449)
      rob_fflags_3_23 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1417)
      rob_fflags_3_23 <= io_fflags_0_bits_flags;
    else if (_GEN_3467)
      rob_fflags_3_23 <= 5'h0;
    if (_GEN_4278 & _GEN_1482)
      rob_fflags_3_24 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1450)
      rob_fflags_3_24 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1418)
      rob_fflags_3_24 <= io_fflags_0_bits_flags;
    else if (_GEN_3468)
      rob_fflags_3_24 <= 5'h0;
    if (_GEN_4278 & _GEN_1483)
      rob_fflags_3_25 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1451)
      rob_fflags_3_25 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1419)
      rob_fflags_3_25 <= io_fflags_0_bits_flags;
    else if (_GEN_3469)
      rob_fflags_3_25 <= 5'h0;
    if (_GEN_4278 & _GEN_1484)
      rob_fflags_3_26 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1452)
      rob_fflags_3_26 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1420)
      rob_fflags_3_26 <= io_fflags_0_bits_flags;
    else if (_GEN_3470)
      rob_fflags_3_26 <= 5'h0;
    if (_GEN_4278 & _GEN_1485)
      rob_fflags_3_27 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1453)
      rob_fflags_3_27 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1421)
      rob_fflags_3_27 <= io_fflags_0_bits_flags;
    else if (_GEN_3471)
      rob_fflags_3_27 <= 5'h0;
    if (_GEN_4278 & _GEN_1486)
      rob_fflags_3_28 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1454)
      rob_fflags_3_28 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1422)
      rob_fflags_3_28 <= io_fflags_0_bits_flags;
    else if (_GEN_3472)
      rob_fflags_3_28 <= 5'h0;
    if (_GEN_4278 & _GEN_1487)
      rob_fflags_3_29 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1455)
      rob_fflags_3_29 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1423)
      rob_fflags_3_29 <= io_fflags_0_bits_flags;
    else if (_GEN_3473)
      rob_fflags_3_29 <= 5'h0;
    if (_GEN_4278 & _GEN_1488)
      rob_fflags_3_30 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & _GEN_1456)
      rob_fflags_3_30 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & _GEN_1424)
      rob_fflags_3_30 <= io_fflags_0_bits_flags;
    else if (_GEN_3474)
      rob_fflags_3_30 <= 5'h0;
    if (_GEN_4278 & (&(io_fflags_3_bits_uop_rob_idx[6:2])))
      rob_fflags_3_31 <= io_fflags_3_bits_flags;
    else if (_GEN_4277 & (&(io_fflags_2_bits_uop_rob_idx[6:2])))
      rob_fflags_3_31 <= io_fflags_2_bits_flags;
    else if (_GEN_4276 & (&(io_fflags_0_bits_uop_rob_idx[6:2])))
      rob_fflags_3_31 <= io_fflags_0_bits_flags;
    else if (_GEN_3475)
      rob_fflags_3_31 <= 5'h0;
    rob_bsy_0 <= ~_GEN_1331 & (_GEN_10 ? ~_GEN_1268 & _GEN_1079 : ~_GEN_1205 & _GEN_1079);
    rob_bsy_1 <= ~_GEN_1333 & (_GEN_10 ? ~_GEN_1270 & _GEN_1082 : ~_GEN_1207 & _GEN_1082);
    rob_bsy_2 <= ~_GEN_1335 & (_GEN_10 ? ~_GEN_1272 & _GEN_1085 : ~_GEN_1209 & _GEN_1085);
    rob_bsy_3 <= ~_GEN_1337 & (_GEN_10 ? ~_GEN_1274 & _GEN_1088 : ~_GEN_1211 & _GEN_1088);
    rob_bsy_4 <= ~_GEN_1339 & (_GEN_10 ? ~_GEN_1276 & _GEN_1091 : ~_GEN_1213 & _GEN_1091);
    rob_bsy_5 <= ~_GEN_1341 & (_GEN_10 ? ~_GEN_1278 & _GEN_1094 : ~_GEN_1215 & _GEN_1094);
    rob_bsy_6 <= ~_GEN_1343 & (_GEN_10 ? ~_GEN_1280 & _GEN_1097 : ~_GEN_1217 & _GEN_1097);
    rob_bsy_7 <= ~_GEN_1345 & (_GEN_10 ? ~_GEN_1282 & _GEN_1100 : ~_GEN_1219 & _GEN_1100);
    rob_bsy_8 <= ~_GEN_1347 & (_GEN_10 ? ~_GEN_1284 & _GEN_1103 : ~_GEN_1221 & _GEN_1103);
    rob_bsy_9 <= ~_GEN_1349 & (_GEN_10 ? ~_GEN_1286 & _GEN_1106 : ~_GEN_1223 & _GEN_1106);
    rob_bsy_10 <= ~_GEN_1351 & (_GEN_10 ? ~_GEN_1288 & _GEN_1109 : ~_GEN_1225 & _GEN_1109);
    rob_bsy_11 <= ~_GEN_1353 & (_GEN_10 ? ~_GEN_1290 & _GEN_1112 : ~_GEN_1227 & _GEN_1112);
    rob_bsy_12 <= ~_GEN_1355 & (_GEN_10 ? ~_GEN_1292 & _GEN_1115 : ~_GEN_1229 & _GEN_1115);
    rob_bsy_13 <= ~_GEN_1357 & (_GEN_10 ? ~_GEN_1294 & _GEN_1118 : ~_GEN_1231 & _GEN_1118);
    rob_bsy_14 <= ~_GEN_1359 & (_GEN_10 ? ~_GEN_1296 & _GEN_1121 : ~_GEN_1233 & _GEN_1121);
    rob_bsy_15 <= ~_GEN_1361 & (_GEN_10 ? ~_GEN_1298 & _GEN_1124 : ~_GEN_1235 & _GEN_1124);
    rob_bsy_16 <= ~_GEN_1363 & (_GEN_10 ? ~_GEN_1300 & _GEN_1127 : ~_GEN_1237 & _GEN_1127);
    rob_bsy_17 <= ~_GEN_1365 & (_GEN_10 ? ~_GEN_1302 & _GEN_1130 : ~_GEN_1239 & _GEN_1130);
    rob_bsy_18 <= ~_GEN_1367 & (_GEN_10 ? ~_GEN_1304 & _GEN_1133 : ~_GEN_1241 & _GEN_1133);
    rob_bsy_19 <= ~_GEN_1369 & (_GEN_10 ? ~_GEN_1306 & _GEN_1136 : ~_GEN_1243 & _GEN_1136);
    rob_bsy_20 <= ~_GEN_1371 & (_GEN_10 ? ~_GEN_1308 & _GEN_1139 : ~_GEN_1245 & _GEN_1139);
    rob_bsy_21 <= ~_GEN_1373 & (_GEN_10 ? ~_GEN_1310 & _GEN_1142 : ~_GEN_1247 & _GEN_1142);
    rob_bsy_22 <= ~_GEN_1375 & (_GEN_10 ? ~_GEN_1312 & _GEN_1145 : ~_GEN_1249 & _GEN_1145);
    rob_bsy_23 <= ~_GEN_1377 & (_GEN_10 ? ~_GEN_1314 & _GEN_1148 : ~_GEN_1251 & _GEN_1148);
    rob_bsy_24 <= ~_GEN_1379 & (_GEN_10 ? ~_GEN_1316 & _GEN_1151 : ~_GEN_1253 & _GEN_1151);
    rob_bsy_25 <= ~_GEN_1381 & (_GEN_10 ? ~_GEN_1318 & _GEN_1154 : ~_GEN_1255 & _GEN_1154);
    rob_bsy_26 <= ~_GEN_1383 & (_GEN_10 ? ~_GEN_1320 & _GEN_1157 : ~_GEN_1257 & _GEN_1157);
    rob_bsy_27 <= ~_GEN_1385 & (_GEN_10 ? ~_GEN_1322 & _GEN_1160 : ~_GEN_1259 & _GEN_1160);
    rob_bsy_28 <= ~_GEN_1387 & (_GEN_10 ? ~_GEN_1324 & _GEN_1163 : ~_GEN_1261 & _GEN_1163);
    rob_bsy_29 <= ~_GEN_1389 & (_GEN_10 ? ~_GEN_1326 & _GEN_1166 : ~_GEN_1263 & _GEN_1166);
    rob_bsy_30 <= ~_GEN_1391 & (_GEN_10 ? ~_GEN_1328 & _GEN_1169 : ~_GEN_1265 & _GEN_1169);
    rob_bsy_31 <= ~_GEN_1392 & (_GEN_10 ? ~_GEN_1329 & _GEN_1171 : ~_GEN_1266 & _GEN_1171);
    rob_unsafe_0 <= ~_GEN_1331 & (_GEN_10 ? ~_GEN_1268 & _GEN_1172 : ~_GEN_1205 & _GEN_1172);
    rob_unsafe_1 <= ~_GEN_1333 & (_GEN_10 ? ~_GEN_1270 & _GEN_1173 : ~_GEN_1207 & _GEN_1173);
    rob_unsafe_2 <= ~_GEN_1335 & (_GEN_10 ? ~_GEN_1272 & _GEN_1174 : ~_GEN_1209 & _GEN_1174);
    rob_unsafe_3 <= ~_GEN_1337 & (_GEN_10 ? ~_GEN_1274 & _GEN_1175 : ~_GEN_1211 & _GEN_1175);
    rob_unsafe_4 <= ~_GEN_1339 & (_GEN_10 ? ~_GEN_1276 & _GEN_1176 : ~_GEN_1213 & _GEN_1176);
    rob_unsafe_5 <= ~_GEN_1341 & (_GEN_10 ? ~_GEN_1278 & _GEN_1177 : ~_GEN_1215 & _GEN_1177);
    rob_unsafe_6 <= ~_GEN_1343 & (_GEN_10 ? ~_GEN_1280 & _GEN_1178 : ~_GEN_1217 & _GEN_1178);
    rob_unsafe_7 <= ~_GEN_1345 & (_GEN_10 ? ~_GEN_1282 & _GEN_1179 : ~_GEN_1219 & _GEN_1179);
    rob_unsafe_8 <= ~_GEN_1347 & (_GEN_10 ? ~_GEN_1284 & _GEN_1180 : ~_GEN_1221 & _GEN_1180);
    rob_unsafe_9 <= ~_GEN_1349 & (_GEN_10 ? ~_GEN_1286 & _GEN_1181 : ~_GEN_1223 & _GEN_1181);
    rob_unsafe_10 <= ~_GEN_1351 & (_GEN_10 ? ~_GEN_1288 & _GEN_1182 : ~_GEN_1225 & _GEN_1182);
    rob_unsafe_11 <= ~_GEN_1353 & (_GEN_10 ? ~_GEN_1290 & _GEN_1183 : ~_GEN_1227 & _GEN_1183);
    rob_unsafe_12 <= ~_GEN_1355 & (_GEN_10 ? ~_GEN_1292 & _GEN_1184 : ~_GEN_1229 & _GEN_1184);
    rob_unsafe_13 <= ~_GEN_1357 & (_GEN_10 ? ~_GEN_1294 & _GEN_1185 : ~_GEN_1231 & _GEN_1185);
    rob_unsafe_14 <= ~_GEN_1359 & (_GEN_10 ? ~_GEN_1296 & _GEN_1186 : ~_GEN_1233 & _GEN_1186);
    rob_unsafe_15 <= ~_GEN_1361 & (_GEN_10 ? ~_GEN_1298 & _GEN_1187 : ~_GEN_1235 & _GEN_1187);
    rob_unsafe_16 <= ~_GEN_1363 & (_GEN_10 ? ~_GEN_1300 & _GEN_1188 : ~_GEN_1237 & _GEN_1188);
    rob_unsafe_17 <= ~_GEN_1365 & (_GEN_10 ? ~_GEN_1302 & _GEN_1189 : ~_GEN_1239 & _GEN_1189);
    rob_unsafe_18 <= ~_GEN_1367 & (_GEN_10 ? ~_GEN_1304 & _GEN_1190 : ~_GEN_1241 & _GEN_1190);
    rob_unsafe_19 <= ~_GEN_1369 & (_GEN_10 ? ~_GEN_1306 & _GEN_1191 : ~_GEN_1243 & _GEN_1191);
    rob_unsafe_20 <= ~_GEN_1371 & (_GEN_10 ? ~_GEN_1308 & _GEN_1192 : ~_GEN_1245 & _GEN_1192);
    rob_unsafe_21 <= ~_GEN_1373 & (_GEN_10 ? ~_GEN_1310 & _GEN_1193 : ~_GEN_1247 & _GEN_1193);
    rob_unsafe_22 <= ~_GEN_1375 & (_GEN_10 ? ~_GEN_1312 & _GEN_1194 : ~_GEN_1249 & _GEN_1194);
    rob_unsafe_23 <= ~_GEN_1377 & (_GEN_10 ? ~_GEN_1314 & _GEN_1195 : ~_GEN_1251 & _GEN_1195);
    rob_unsafe_24 <= ~_GEN_1379 & (_GEN_10 ? ~_GEN_1316 & _GEN_1196 : ~_GEN_1253 & _GEN_1196);
    rob_unsafe_25 <= ~_GEN_1381 & (_GEN_10 ? ~_GEN_1318 & _GEN_1197 : ~_GEN_1255 & _GEN_1197);
    rob_unsafe_26 <= ~_GEN_1383 & (_GEN_10 ? ~_GEN_1320 & _GEN_1198 : ~_GEN_1257 & _GEN_1198);
    rob_unsafe_27 <= ~_GEN_1385 & (_GEN_10 ? ~_GEN_1322 & _GEN_1199 : ~_GEN_1259 & _GEN_1199);
    rob_unsafe_28 <= ~_GEN_1387 & (_GEN_10 ? ~_GEN_1324 & _GEN_1200 : ~_GEN_1261 & _GEN_1200);
    rob_unsafe_29 <= ~_GEN_1389 & (_GEN_10 ? ~_GEN_1326 & _GEN_1201 : ~_GEN_1263 & _GEN_1201);
    rob_unsafe_30 <= ~_GEN_1391 & (_GEN_10 ? ~_GEN_1328 & _GEN_1202 : ~_GEN_1265 & _GEN_1202);
    rob_unsafe_31 <= ~_GEN_1392 & (_GEN_10 ? ~_GEN_1329 & _GEN_1203 : ~_GEN_1266 & _GEN_1203);
    if (_GEN_128) begin
      rob_uop_0_uopc <= io_enq_uops_0_uopc;
      rob_uop_0_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_0_is_br <= io_enq_uops_0_is_br;
      rob_uop_0_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_0_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_0_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_0_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_0_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_0_pdst <= io_enq_uops_0_pdst;
      rob_uop_0_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_0_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_0_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_0_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_0_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_0_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_0_ldst <= io_enq_uops_0_ldst;
      rob_uop_0_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_0_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_0_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1583) | ~rob_val_0) begin
      if (_GEN_128)
        rob_uop_0_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_0_br_mask <= rob_uop_0_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1615)
      rob_uop_0_debug_fsrc <= 2'h3;
    else if (_GEN_128)
      rob_uop_0_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_130) begin
      rob_uop_1_uopc <= io_enq_uops_0_uopc;
      rob_uop_1_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_1_is_br <= io_enq_uops_0_is_br;
      rob_uop_1_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_1_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_1_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_1_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_1_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_1_pdst <= io_enq_uops_0_pdst;
      rob_uop_1_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_1_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_1_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_1_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_1_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_1_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_1_ldst <= io_enq_uops_0_ldst;
      rob_uop_1_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_1_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_1_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1584) | ~rob_val_1) begin
      if (_GEN_130)
        rob_uop_1_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_1_br_mask <= rob_uop_1_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1616)
      rob_uop_1_debug_fsrc <= 2'h3;
    else if (_GEN_130)
      rob_uop_1_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_132) begin
      rob_uop_2_uopc <= io_enq_uops_0_uopc;
      rob_uop_2_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_2_is_br <= io_enq_uops_0_is_br;
      rob_uop_2_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_2_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_2_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_2_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_2_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_2_pdst <= io_enq_uops_0_pdst;
      rob_uop_2_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_2_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_2_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_2_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_2_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_2_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_2_ldst <= io_enq_uops_0_ldst;
      rob_uop_2_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_2_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_2_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1585) | ~rob_val_2) begin
      if (_GEN_132)
        rob_uop_2_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_2_br_mask <= rob_uop_2_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1617)
      rob_uop_2_debug_fsrc <= 2'h3;
    else if (_GEN_132)
      rob_uop_2_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_134) begin
      rob_uop_3_uopc <= io_enq_uops_0_uopc;
      rob_uop_3_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_3_is_br <= io_enq_uops_0_is_br;
      rob_uop_3_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_3_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_3_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_3_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_3_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_3_pdst <= io_enq_uops_0_pdst;
      rob_uop_3_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_3_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_3_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_3_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_3_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_3_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_3_ldst <= io_enq_uops_0_ldst;
      rob_uop_3_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_3_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_3_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1586) | ~rob_val_3) begin
      if (_GEN_134)
        rob_uop_3_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_3_br_mask <= rob_uop_3_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1618)
      rob_uop_3_debug_fsrc <= 2'h3;
    else if (_GEN_134)
      rob_uop_3_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_136) begin
      rob_uop_4_uopc <= io_enq_uops_0_uopc;
      rob_uop_4_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_4_is_br <= io_enq_uops_0_is_br;
      rob_uop_4_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_4_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_4_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_4_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_4_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_4_pdst <= io_enq_uops_0_pdst;
      rob_uop_4_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_4_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_4_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_4_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_4_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_4_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_4_ldst <= io_enq_uops_0_ldst;
      rob_uop_4_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_4_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_4_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1587) | ~rob_val_4) begin
      if (_GEN_136)
        rob_uop_4_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_4_br_mask <= rob_uop_4_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1619)
      rob_uop_4_debug_fsrc <= 2'h3;
    else if (_GEN_136)
      rob_uop_4_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_138) begin
      rob_uop_5_uopc <= io_enq_uops_0_uopc;
      rob_uop_5_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_5_is_br <= io_enq_uops_0_is_br;
      rob_uop_5_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_5_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_5_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_5_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_5_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_5_pdst <= io_enq_uops_0_pdst;
      rob_uop_5_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_5_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_5_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_5_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_5_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_5_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_5_ldst <= io_enq_uops_0_ldst;
      rob_uop_5_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_5_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_5_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1588) | ~rob_val_5) begin
      if (_GEN_138)
        rob_uop_5_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_5_br_mask <= rob_uop_5_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1620)
      rob_uop_5_debug_fsrc <= 2'h3;
    else if (_GEN_138)
      rob_uop_5_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_140) begin
      rob_uop_6_uopc <= io_enq_uops_0_uopc;
      rob_uop_6_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_6_is_br <= io_enq_uops_0_is_br;
      rob_uop_6_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_6_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_6_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_6_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_6_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_6_pdst <= io_enq_uops_0_pdst;
      rob_uop_6_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_6_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_6_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_6_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_6_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_6_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_6_ldst <= io_enq_uops_0_ldst;
      rob_uop_6_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_6_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_6_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1589) | ~rob_val_6) begin
      if (_GEN_140)
        rob_uop_6_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_6_br_mask <= rob_uop_6_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1621)
      rob_uop_6_debug_fsrc <= 2'h3;
    else if (_GEN_140)
      rob_uop_6_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_142) begin
      rob_uop_7_uopc <= io_enq_uops_0_uopc;
      rob_uop_7_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_7_is_br <= io_enq_uops_0_is_br;
      rob_uop_7_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_7_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_7_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_7_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_7_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_7_pdst <= io_enq_uops_0_pdst;
      rob_uop_7_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_7_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_7_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_7_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_7_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_7_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_7_ldst <= io_enq_uops_0_ldst;
      rob_uop_7_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_7_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_7_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1590) | ~rob_val_7) begin
      if (_GEN_142)
        rob_uop_7_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_7_br_mask <= rob_uop_7_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1622)
      rob_uop_7_debug_fsrc <= 2'h3;
    else if (_GEN_142)
      rob_uop_7_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_144) begin
      rob_uop_8_uopc <= io_enq_uops_0_uopc;
      rob_uop_8_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_8_is_br <= io_enq_uops_0_is_br;
      rob_uop_8_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_8_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_8_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_8_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_8_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_8_pdst <= io_enq_uops_0_pdst;
      rob_uop_8_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_8_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_8_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_8_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_8_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_8_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_8_ldst <= io_enq_uops_0_ldst;
      rob_uop_8_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_8_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_8_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1591) | ~rob_val_8) begin
      if (_GEN_144)
        rob_uop_8_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_8_br_mask <= rob_uop_8_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1623)
      rob_uop_8_debug_fsrc <= 2'h3;
    else if (_GEN_144)
      rob_uop_8_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_146) begin
      rob_uop_9_uopc <= io_enq_uops_0_uopc;
      rob_uop_9_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_9_is_br <= io_enq_uops_0_is_br;
      rob_uop_9_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_9_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_9_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_9_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_9_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_9_pdst <= io_enq_uops_0_pdst;
      rob_uop_9_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_9_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_9_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_9_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_9_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_9_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_9_ldst <= io_enq_uops_0_ldst;
      rob_uop_9_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_9_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_9_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1592) | ~rob_val_9) begin
      if (_GEN_146)
        rob_uop_9_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_9_br_mask <= rob_uop_9_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1624)
      rob_uop_9_debug_fsrc <= 2'h3;
    else if (_GEN_146)
      rob_uop_9_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_148) begin
      rob_uop_10_uopc <= io_enq_uops_0_uopc;
      rob_uop_10_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_10_is_br <= io_enq_uops_0_is_br;
      rob_uop_10_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_10_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_10_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_10_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_10_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_10_pdst <= io_enq_uops_0_pdst;
      rob_uop_10_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_10_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_10_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_10_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_10_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_10_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_10_ldst <= io_enq_uops_0_ldst;
      rob_uop_10_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_10_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_10_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1593) | ~rob_val_10) begin
      if (_GEN_148)
        rob_uop_10_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_10_br_mask <= rob_uop_10_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1625)
      rob_uop_10_debug_fsrc <= 2'h3;
    else if (_GEN_148)
      rob_uop_10_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_150) begin
      rob_uop_11_uopc <= io_enq_uops_0_uopc;
      rob_uop_11_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_11_is_br <= io_enq_uops_0_is_br;
      rob_uop_11_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_11_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_11_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_11_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_11_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_11_pdst <= io_enq_uops_0_pdst;
      rob_uop_11_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_11_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_11_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_11_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_11_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_11_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_11_ldst <= io_enq_uops_0_ldst;
      rob_uop_11_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_11_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_11_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1594) | ~rob_val_11) begin
      if (_GEN_150)
        rob_uop_11_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_11_br_mask <= rob_uop_11_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1626)
      rob_uop_11_debug_fsrc <= 2'h3;
    else if (_GEN_150)
      rob_uop_11_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_152) begin
      rob_uop_12_uopc <= io_enq_uops_0_uopc;
      rob_uop_12_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_12_is_br <= io_enq_uops_0_is_br;
      rob_uop_12_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_12_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_12_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_12_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_12_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_12_pdst <= io_enq_uops_0_pdst;
      rob_uop_12_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_12_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_12_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_12_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_12_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_12_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_12_ldst <= io_enq_uops_0_ldst;
      rob_uop_12_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_12_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_12_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1595) | ~rob_val_12) begin
      if (_GEN_152)
        rob_uop_12_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_12_br_mask <= rob_uop_12_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1627)
      rob_uop_12_debug_fsrc <= 2'h3;
    else if (_GEN_152)
      rob_uop_12_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_154) begin
      rob_uop_13_uopc <= io_enq_uops_0_uopc;
      rob_uop_13_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_13_is_br <= io_enq_uops_0_is_br;
      rob_uop_13_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_13_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_13_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_13_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_13_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_13_pdst <= io_enq_uops_0_pdst;
      rob_uop_13_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_13_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_13_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_13_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_13_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_13_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_13_ldst <= io_enq_uops_0_ldst;
      rob_uop_13_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_13_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_13_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1596) | ~rob_val_13) begin
      if (_GEN_154)
        rob_uop_13_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_13_br_mask <= rob_uop_13_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1628)
      rob_uop_13_debug_fsrc <= 2'h3;
    else if (_GEN_154)
      rob_uop_13_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_156) begin
      rob_uop_14_uopc <= io_enq_uops_0_uopc;
      rob_uop_14_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_14_is_br <= io_enq_uops_0_is_br;
      rob_uop_14_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_14_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_14_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_14_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_14_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_14_pdst <= io_enq_uops_0_pdst;
      rob_uop_14_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_14_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_14_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_14_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_14_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_14_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_14_ldst <= io_enq_uops_0_ldst;
      rob_uop_14_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_14_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_14_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1597) | ~rob_val_14) begin
      if (_GEN_156)
        rob_uop_14_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_14_br_mask <= rob_uop_14_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1629)
      rob_uop_14_debug_fsrc <= 2'h3;
    else if (_GEN_156)
      rob_uop_14_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_158) begin
      rob_uop_15_uopc <= io_enq_uops_0_uopc;
      rob_uop_15_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_15_is_br <= io_enq_uops_0_is_br;
      rob_uop_15_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_15_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_15_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_15_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_15_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_15_pdst <= io_enq_uops_0_pdst;
      rob_uop_15_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_15_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_15_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_15_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_15_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_15_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_15_ldst <= io_enq_uops_0_ldst;
      rob_uop_15_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_15_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_15_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1598) | ~rob_val_15) begin
      if (_GEN_158)
        rob_uop_15_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_15_br_mask <= rob_uop_15_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1630)
      rob_uop_15_debug_fsrc <= 2'h3;
    else if (_GEN_158)
      rob_uop_15_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_160) begin
      rob_uop_16_uopc <= io_enq_uops_0_uopc;
      rob_uop_16_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_16_is_br <= io_enq_uops_0_is_br;
      rob_uop_16_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_16_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_16_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_16_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_16_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_16_pdst <= io_enq_uops_0_pdst;
      rob_uop_16_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_16_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_16_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_16_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_16_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_16_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_16_ldst <= io_enq_uops_0_ldst;
      rob_uop_16_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_16_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_16_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1599) | ~rob_val_16) begin
      if (_GEN_160)
        rob_uop_16_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_16_br_mask <= rob_uop_16_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1631)
      rob_uop_16_debug_fsrc <= 2'h3;
    else if (_GEN_160)
      rob_uop_16_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_162) begin
      rob_uop_17_uopc <= io_enq_uops_0_uopc;
      rob_uop_17_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_17_is_br <= io_enq_uops_0_is_br;
      rob_uop_17_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_17_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_17_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_17_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_17_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_17_pdst <= io_enq_uops_0_pdst;
      rob_uop_17_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_17_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_17_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_17_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_17_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_17_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_17_ldst <= io_enq_uops_0_ldst;
      rob_uop_17_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_17_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_17_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1600) | ~rob_val_17) begin
      if (_GEN_162)
        rob_uop_17_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_17_br_mask <= rob_uop_17_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1632)
      rob_uop_17_debug_fsrc <= 2'h3;
    else if (_GEN_162)
      rob_uop_17_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_164) begin
      rob_uop_18_uopc <= io_enq_uops_0_uopc;
      rob_uop_18_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_18_is_br <= io_enq_uops_0_is_br;
      rob_uop_18_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_18_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_18_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_18_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_18_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_18_pdst <= io_enq_uops_0_pdst;
      rob_uop_18_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_18_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_18_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_18_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_18_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_18_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_18_ldst <= io_enq_uops_0_ldst;
      rob_uop_18_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_18_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_18_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1601) | ~rob_val_18) begin
      if (_GEN_164)
        rob_uop_18_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_18_br_mask <= rob_uop_18_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1633)
      rob_uop_18_debug_fsrc <= 2'h3;
    else if (_GEN_164)
      rob_uop_18_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_166) begin
      rob_uop_19_uopc <= io_enq_uops_0_uopc;
      rob_uop_19_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_19_is_br <= io_enq_uops_0_is_br;
      rob_uop_19_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_19_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_19_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_19_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_19_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_19_pdst <= io_enq_uops_0_pdst;
      rob_uop_19_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_19_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_19_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_19_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_19_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_19_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_19_ldst <= io_enq_uops_0_ldst;
      rob_uop_19_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_19_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_19_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1602) | ~rob_val_19) begin
      if (_GEN_166)
        rob_uop_19_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_19_br_mask <= rob_uop_19_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1634)
      rob_uop_19_debug_fsrc <= 2'h3;
    else if (_GEN_166)
      rob_uop_19_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_168) begin
      rob_uop_20_uopc <= io_enq_uops_0_uopc;
      rob_uop_20_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_20_is_br <= io_enq_uops_0_is_br;
      rob_uop_20_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_20_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_20_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_20_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_20_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_20_pdst <= io_enq_uops_0_pdst;
      rob_uop_20_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_20_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_20_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_20_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_20_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_20_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_20_ldst <= io_enq_uops_0_ldst;
      rob_uop_20_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_20_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_20_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1603) | ~rob_val_20) begin
      if (_GEN_168)
        rob_uop_20_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_20_br_mask <= rob_uop_20_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1635)
      rob_uop_20_debug_fsrc <= 2'h3;
    else if (_GEN_168)
      rob_uop_20_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_170) begin
      rob_uop_21_uopc <= io_enq_uops_0_uopc;
      rob_uop_21_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_21_is_br <= io_enq_uops_0_is_br;
      rob_uop_21_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_21_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_21_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_21_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_21_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_21_pdst <= io_enq_uops_0_pdst;
      rob_uop_21_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_21_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_21_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_21_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_21_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_21_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_21_ldst <= io_enq_uops_0_ldst;
      rob_uop_21_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_21_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_21_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1604) | ~rob_val_21) begin
      if (_GEN_170)
        rob_uop_21_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_21_br_mask <= rob_uop_21_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1636)
      rob_uop_21_debug_fsrc <= 2'h3;
    else if (_GEN_170)
      rob_uop_21_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_172) begin
      rob_uop_22_uopc <= io_enq_uops_0_uopc;
      rob_uop_22_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_22_is_br <= io_enq_uops_0_is_br;
      rob_uop_22_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_22_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_22_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_22_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_22_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_22_pdst <= io_enq_uops_0_pdst;
      rob_uop_22_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_22_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_22_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_22_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_22_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_22_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_22_ldst <= io_enq_uops_0_ldst;
      rob_uop_22_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_22_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_22_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1605) | ~rob_val_22) begin
      if (_GEN_172)
        rob_uop_22_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_22_br_mask <= rob_uop_22_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1637)
      rob_uop_22_debug_fsrc <= 2'h3;
    else if (_GEN_172)
      rob_uop_22_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_174) begin
      rob_uop_23_uopc <= io_enq_uops_0_uopc;
      rob_uop_23_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_23_is_br <= io_enq_uops_0_is_br;
      rob_uop_23_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_23_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_23_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_23_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_23_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_23_pdst <= io_enq_uops_0_pdst;
      rob_uop_23_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_23_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_23_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_23_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_23_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_23_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_23_ldst <= io_enq_uops_0_ldst;
      rob_uop_23_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_23_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_23_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1606) | ~rob_val_23) begin
      if (_GEN_174)
        rob_uop_23_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_23_br_mask <= rob_uop_23_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1638)
      rob_uop_23_debug_fsrc <= 2'h3;
    else if (_GEN_174)
      rob_uop_23_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_176) begin
      rob_uop_24_uopc <= io_enq_uops_0_uopc;
      rob_uop_24_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_24_is_br <= io_enq_uops_0_is_br;
      rob_uop_24_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_24_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_24_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_24_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_24_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_24_pdst <= io_enq_uops_0_pdst;
      rob_uop_24_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_24_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_24_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_24_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_24_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_24_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_24_ldst <= io_enq_uops_0_ldst;
      rob_uop_24_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_24_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_24_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1607) | ~rob_val_24) begin
      if (_GEN_176)
        rob_uop_24_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_24_br_mask <= rob_uop_24_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1639)
      rob_uop_24_debug_fsrc <= 2'h3;
    else if (_GEN_176)
      rob_uop_24_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_178) begin
      rob_uop_25_uopc <= io_enq_uops_0_uopc;
      rob_uop_25_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_25_is_br <= io_enq_uops_0_is_br;
      rob_uop_25_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_25_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_25_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_25_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_25_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_25_pdst <= io_enq_uops_0_pdst;
      rob_uop_25_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_25_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_25_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_25_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_25_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_25_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_25_ldst <= io_enq_uops_0_ldst;
      rob_uop_25_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_25_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_25_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1608) | ~rob_val_25) begin
      if (_GEN_178)
        rob_uop_25_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_25_br_mask <= rob_uop_25_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1640)
      rob_uop_25_debug_fsrc <= 2'h3;
    else if (_GEN_178)
      rob_uop_25_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_180) begin
      rob_uop_26_uopc <= io_enq_uops_0_uopc;
      rob_uop_26_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_26_is_br <= io_enq_uops_0_is_br;
      rob_uop_26_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_26_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_26_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_26_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_26_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_26_pdst <= io_enq_uops_0_pdst;
      rob_uop_26_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_26_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_26_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_26_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_26_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_26_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_26_ldst <= io_enq_uops_0_ldst;
      rob_uop_26_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_26_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_26_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1609) | ~rob_val_26) begin
      if (_GEN_180)
        rob_uop_26_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_26_br_mask <= rob_uop_26_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1641)
      rob_uop_26_debug_fsrc <= 2'h3;
    else if (_GEN_180)
      rob_uop_26_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_182) begin
      rob_uop_27_uopc <= io_enq_uops_0_uopc;
      rob_uop_27_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_27_is_br <= io_enq_uops_0_is_br;
      rob_uop_27_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_27_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_27_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_27_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_27_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_27_pdst <= io_enq_uops_0_pdst;
      rob_uop_27_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_27_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_27_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_27_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_27_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_27_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_27_ldst <= io_enq_uops_0_ldst;
      rob_uop_27_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_27_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_27_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1610) | ~rob_val_27) begin
      if (_GEN_182)
        rob_uop_27_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_27_br_mask <= rob_uop_27_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1642)
      rob_uop_27_debug_fsrc <= 2'h3;
    else if (_GEN_182)
      rob_uop_27_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_184) begin
      rob_uop_28_uopc <= io_enq_uops_0_uopc;
      rob_uop_28_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_28_is_br <= io_enq_uops_0_is_br;
      rob_uop_28_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_28_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_28_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_28_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_28_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_28_pdst <= io_enq_uops_0_pdst;
      rob_uop_28_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_28_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_28_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_28_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_28_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_28_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_28_ldst <= io_enq_uops_0_ldst;
      rob_uop_28_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_28_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_28_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1611) | ~rob_val_28) begin
      if (_GEN_184)
        rob_uop_28_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_28_br_mask <= rob_uop_28_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1643)
      rob_uop_28_debug_fsrc <= 2'h3;
    else if (_GEN_184)
      rob_uop_28_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_186) begin
      rob_uop_29_uopc <= io_enq_uops_0_uopc;
      rob_uop_29_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_29_is_br <= io_enq_uops_0_is_br;
      rob_uop_29_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_29_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_29_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_29_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_29_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_29_pdst <= io_enq_uops_0_pdst;
      rob_uop_29_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_29_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_29_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_29_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_29_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_29_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_29_ldst <= io_enq_uops_0_ldst;
      rob_uop_29_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_29_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_29_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1612) | ~rob_val_29) begin
      if (_GEN_186)
        rob_uop_29_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_29_br_mask <= rob_uop_29_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1644)
      rob_uop_29_debug_fsrc <= 2'h3;
    else if (_GEN_186)
      rob_uop_29_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_188) begin
      rob_uop_30_uopc <= io_enq_uops_0_uopc;
      rob_uop_30_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_30_is_br <= io_enq_uops_0_is_br;
      rob_uop_30_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_30_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_30_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_30_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_30_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_30_pdst <= io_enq_uops_0_pdst;
      rob_uop_30_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_30_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_30_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_30_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_30_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_30_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_30_ldst <= io_enq_uops_0_ldst;
      rob_uop_30_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_30_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_30_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1613) | ~rob_val_30) begin
      if (_GEN_188)
        rob_uop_30_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_30_br_mask <= rob_uop_30_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & _GEN_1645)
      rob_uop_30_debug_fsrc <= 2'h3;
    else if (_GEN_188)
      rob_uop_30_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    if (_GEN_189) begin
      rob_uop_31_uopc <= io_enq_uops_0_uopc;
      rob_uop_31_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop_31_is_br <= io_enq_uops_0_is_br;
      rob_uop_31_is_jalr <= io_enq_uops_0_is_jalr;
      rob_uop_31_is_jal <= io_enq_uops_0_is_jal;
      rob_uop_31_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop_31_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop_31_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop_31_pdst <= io_enq_uops_0_pdst;
      rob_uop_31_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop_31_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop_31_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop_31_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop_31_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop_31_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop_31_ldst <= io_enq_uops_0_ldst;
      rob_uop_31_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop_31_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop_31_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_1614) | ~rob_val_31) begin
      if (_GEN_189)
        rob_uop_31_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop_31_br_mask <= rob_uop_31_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_15 & (&(io_brupdate_b2_uop_rob_idx[6:2])))
      rob_uop_31_debug_fsrc <= 2'h3;
    else if (_GEN_189)
      rob_uop_31_debug_fsrc <= io_enq_uops_0_debug_fsrc;
    rob_exception_0 <= ~_GEN_1521 & (_GEN_12 & _GEN_1489 | (_GEN_128 ? io_enq_uops_0_exception : rob_exception_0));
    rob_exception_1 <= ~_GEN_1523 & (_GEN_12 & _GEN_1490 | (_GEN_130 ? io_enq_uops_0_exception : rob_exception_1));
    rob_exception_2 <= ~_GEN_1525 & (_GEN_12 & _GEN_1491 | (_GEN_132 ? io_enq_uops_0_exception : rob_exception_2));
    rob_exception_3 <= ~_GEN_1527 & (_GEN_12 & _GEN_1492 | (_GEN_134 ? io_enq_uops_0_exception : rob_exception_3));
    rob_exception_4 <= ~_GEN_1529 & (_GEN_12 & _GEN_1493 | (_GEN_136 ? io_enq_uops_0_exception : rob_exception_4));
    rob_exception_5 <= ~_GEN_1531 & (_GEN_12 & _GEN_1494 | (_GEN_138 ? io_enq_uops_0_exception : rob_exception_5));
    rob_exception_6 <= ~_GEN_1533 & (_GEN_12 & _GEN_1495 | (_GEN_140 ? io_enq_uops_0_exception : rob_exception_6));
    rob_exception_7 <= ~_GEN_1535 & (_GEN_12 & _GEN_1496 | (_GEN_142 ? io_enq_uops_0_exception : rob_exception_7));
    rob_exception_8 <= ~_GEN_1537 & (_GEN_12 & _GEN_1497 | (_GEN_144 ? io_enq_uops_0_exception : rob_exception_8));
    rob_exception_9 <= ~_GEN_1539 & (_GEN_12 & _GEN_1498 | (_GEN_146 ? io_enq_uops_0_exception : rob_exception_9));
    rob_exception_10 <= ~_GEN_1541 & (_GEN_12 & _GEN_1499 | (_GEN_148 ? io_enq_uops_0_exception : rob_exception_10));
    rob_exception_11 <= ~_GEN_1543 & (_GEN_12 & _GEN_1500 | (_GEN_150 ? io_enq_uops_0_exception : rob_exception_11));
    rob_exception_12 <= ~_GEN_1545 & (_GEN_12 & _GEN_1501 | (_GEN_152 ? io_enq_uops_0_exception : rob_exception_12));
    rob_exception_13 <= ~_GEN_1547 & (_GEN_12 & _GEN_1502 | (_GEN_154 ? io_enq_uops_0_exception : rob_exception_13));
    rob_exception_14 <= ~_GEN_1549 & (_GEN_12 & _GEN_1503 | (_GEN_156 ? io_enq_uops_0_exception : rob_exception_14));
    rob_exception_15 <= ~_GEN_1551 & (_GEN_12 & _GEN_1504 | (_GEN_158 ? io_enq_uops_0_exception : rob_exception_15));
    rob_exception_16 <= ~_GEN_1553 & (_GEN_12 & _GEN_1505 | (_GEN_160 ? io_enq_uops_0_exception : rob_exception_16));
    rob_exception_17 <= ~_GEN_1555 & (_GEN_12 & _GEN_1506 | (_GEN_162 ? io_enq_uops_0_exception : rob_exception_17));
    rob_exception_18 <= ~_GEN_1557 & (_GEN_12 & _GEN_1507 | (_GEN_164 ? io_enq_uops_0_exception : rob_exception_18));
    rob_exception_19 <= ~_GEN_1559 & (_GEN_12 & _GEN_1508 | (_GEN_166 ? io_enq_uops_0_exception : rob_exception_19));
    rob_exception_20 <= ~_GEN_1561 & (_GEN_12 & _GEN_1509 | (_GEN_168 ? io_enq_uops_0_exception : rob_exception_20));
    rob_exception_21 <= ~_GEN_1563 & (_GEN_12 & _GEN_1510 | (_GEN_170 ? io_enq_uops_0_exception : rob_exception_21));
    rob_exception_22 <= ~_GEN_1565 & (_GEN_12 & _GEN_1511 | (_GEN_172 ? io_enq_uops_0_exception : rob_exception_22));
    rob_exception_23 <= ~_GEN_1567 & (_GEN_12 & _GEN_1512 | (_GEN_174 ? io_enq_uops_0_exception : rob_exception_23));
    rob_exception_24 <= ~_GEN_1569 & (_GEN_12 & _GEN_1513 | (_GEN_176 ? io_enq_uops_0_exception : rob_exception_24));
    rob_exception_25 <= ~_GEN_1571 & (_GEN_12 & _GEN_1514 | (_GEN_178 ? io_enq_uops_0_exception : rob_exception_25));
    rob_exception_26 <= ~_GEN_1573 & (_GEN_12 & _GEN_1515 | (_GEN_180 ? io_enq_uops_0_exception : rob_exception_26));
    rob_exception_27 <= ~_GEN_1575 & (_GEN_12 & _GEN_1516 | (_GEN_182 ? io_enq_uops_0_exception : rob_exception_27));
    rob_exception_28 <= ~_GEN_1577 & (_GEN_12 & _GEN_1517 | (_GEN_184 ? io_enq_uops_0_exception : rob_exception_28));
    rob_exception_29 <= ~_GEN_1579 & (_GEN_12 & _GEN_1518 | (_GEN_186 ? io_enq_uops_0_exception : rob_exception_29));
    rob_exception_30 <= ~_GEN_1581 & (_GEN_12 & _GEN_1519 | (_GEN_188 ? io_enq_uops_0_exception : rob_exception_30));
    rob_exception_31 <= ~_GEN_1582 & (_GEN_12 & (&(io_lxcpt_bits_uop_rob_idx[6:2])) | (_GEN_189 ? io_enq_uops_0_exception : rob_exception_31));
    rob_predicated_0 <= ~(_GEN_8 & _GEN_1077 | _GEN_1015 | _GEN_6 & _GEN_887) & (_GEN_825 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_697 | _GEN_635 | _GEN_2 & _GEN_507 | _GEN_445 | _GEN_0 & _GEN_317) & (_GEN_255 ? io_wb_resps_0_bits_predicated : ~_GEN_128 & rob_predicated_0));
    rob_predicated_1 <= ~(_GEN_8 & _GEN_1080 | _GEN_1017 | _GEN_6 & _GEN_890) & (_GEN_827 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_700 | _GEN_637 | _GEN_2 & _GEN_510 | _GEN_447 | _GEN_0 & _GEN_320) & (_GEN_257 ? io_wb_resps_0_bits_predicated : ~_GEN_130 & rob_predicated_1));
    rob_predicated_2 <= ~(_GEN_8 & _GEN_1083 | _GEN_1019 | _GEN_6 & _GEN_893) & (_GEN_829 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_703 | _GEN_639 | _GEN_2 & _GEN_513 | _GEN_449 | _GEN_0 & _GEN_323) & (_GEN_259 ? io_wb_resps_0_bits_predicated : ~_GEN_132 & rob_predicated_2));
    rob_predicated_3 <= ~(_GEN_8 & _GEN_1086 | _GEN_1021 | _GEN_6 & _GEN_896) & (_GEN_831 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_706 | _GEN_641 | _GEN_2 & _GEN_516 | _GEN_451 | _GEN_0 & _GEN_326) & (_GEN_261 ? io_wb_resps_0_bits_predicated : ~_GEN_134 & rob_predicated_3));
    rob_predicated_4 <= ~(_GEN_8 & _GEN_1089 | _GEN_1023 | _GEN_6 & _GEN_899) & (_GEN_833 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_709 | _GEN_643 | _GEN_2 & _GEN_519 | _GEN_453 | _GEN_0 & _GEN_329) & (_GEN_263 ? io_wb_resps_0_bits_predicated : ~_GEN_136 & rob_predicated_4));
    rob_predicated_5 <= ~(_GEN_8 & _GEN_1092 | _GEN_1025 | _GEN_6 & _GEN_902) & (_GEN_835 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_712 | _GEN_645 | _GEN_2 & _GEN_522 | _GEN_455 | _GEN_0 & _GEN_332) & (_GEN_265 ? io_wb_resps_0_bits_predicated : ~_GEN_138 & rob_predicated_5));
    rob_predicated_6 <= ~(_GEN_8 & _GEN_1095 | _GEN_1027 | _GEN_6 & _GEN_905) & (_GEN_837 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_715 | _GEN_647 | _GEN_2 & _GEN_525 | _GEN_457 | _GEN_0 & _GEN_335) & (_GEN_267 ? io_wb_resps_0_bits_predicated : ~_GEN_140 & rob_predicated_6));
    rob_predicated_7 <= ~(_GEN_8 & _GEN_1098 | _GEN_1029 | _GEN_6 & _GEN_908) & (_GEN_839 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_718 | _GEN_649 | _GEN_2 & _GEN_528 | _GEN_459 | _GEN_0 & _GEN_338) & (_GEN_269 ? io_wb_resps_0_bits_predicated : ~_GEN_142 & rob_predicated_7));
    rob_predicated_8 <= ~(_GEN_8 & _GEN_1101 | _GEN_1031 | _GEN_6 & _GEN_911) & (_GEN_841 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_721 | _GEN_651 | _GEN_2 & _GEN_531 | _GEN_461 | _GEN_0 & _GEN_341) & (_GEN_271 ? io_wb_resps_0_bits_predicated : ~_GEN_144 & rob_predicated_8));
    rob_predicated_9 <= ~(_GEN_8 & _GEN_1104 | _GEN_1033 | _GEN_6 & _GEN_914) & (_GEN_843 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_724 | _GEN_653 | _GEN_2 & _GEN_534 | _GEN_463 | _GEN_0 & _GEN_344) & (_GEN_273 ? io_wb_resps_0_bits_predicated : ~_GEN_146 & rob_predicated_9));
    rob_predicated_10 <= ~(_GEN_8 & _GEN_1107 | _GEN_1035 | _GEN_6 & _GEN_917) & (_GEN_845 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_727 | _GEN_655 | _GEN_2 & _GEN_537 | _GEN_465 | _GEN_0 & _GEN_347) & (_GEN_275 ? io_wb_resps_0_bits_predicated : ~_GEN_148 & rob_predicated_10));
    rob_predicated_11 <= ~(_GEN_8 & _GEN_1110 | _GEN_1037 | _GEN_6 & _GEN_920) & (_GEN_847 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_730 | _GEN_657 | _GEN_2 & _GEN_540 | _GEN_467 | _GEN_0 & _GEN_350) & (_GEN_277 ? io_wb_resps_0_bits_predicated : ~_GEN_150 & rob_predicated_11));
    rob_predicated_12 <= ~(_GEN_8 & _GEN_1113 | _GEN_1039 | _GEN_6 & _GEN_923) & (_GEN_849 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_733 | _GEN_659 | _GEN_2 & _GEN_543 | _GEN_469 | _GEN_0 & _GEN_353) & (_GEN_279 ? io_wb_resps_0_bits_predicated : ~_GEN_152 & rob_predicated_12));
    rob_predicated_13 <= ~(_GEN_8 & _GEN_1116 | _GEN_1041 | _GEN_6 & _GEN_926) & (_GEN_851 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_736 | _GEN_661 | _GEN_2 & _GEN_546 | _GEN_471 | _GEN_0 & _GEN_356) & (_GEN_281 ? io_wb_resps_0_bits_predicated : ~_GEN_154 & rob_predicated_13));
    rob_predicated_14 <= ~(_GEN_8 & _GEN_1119 | _GEN_1043 | _GEN_6 & _GEN_929) & (_GEN_853 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_739 | _GEN_663 | _GEN_2 & _GEN_549 | _GEN_473 | _GEN_0 & _GEN_359) & (_GEN_283 ? io_wb_resps_0_bits_predicated : ~_GEN_156 & rob_predicated_14));
    rob_predicated_15 <= ~(_GEN_8 & _GEN_1122 | _GEN_1045 | _GEN_6 & _GEN_932) & (_GEN_855 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_742 | _GEN_665 | _GEN_2 & _GEN_552 | _GEN_475 | _GEN_0 & _GEN_362) & (_GEN_285 ? io_wb_resps_0_bits_predicated : ~_GEN_158 & rob_predicated_15));
    rob_predicated_16 <= ~(_GEN_8 & _GEN_1125 | _GEN_1047 | _GEN_6 & _GEN_935) & (_GEN_857 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_745 | _GEN_667 | _GEN_2 & _GEN_555 | _GEN_477 | _GEN_0 & _GEN_365) & (_GEN_287 ? io_wb_resps_0_bits_predicated : ~_GEN_160 & rob_predicated_16));
    rob_predicated_17 <= ~(_GEN_8 & _GEN_1128 | _GEN_1049 | _GEN_6 & _GEN_938) & (_GEN_859 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_748 | _GEN_669 | _GEN_2 & _GEN_558 | _GEN_479 | _GEN_0 & _GEN_368) & (_GEN_289 ? io_wb_resps_0_bits_predicated : ~_GEN_162 & rob_predicated_17));
    rob_predicated_18 <= ~(_GEN_8 & _GEN_1131 | _GEN_1051 | _GEN_6 & _GEN_941) & (_GEN_861 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_751 | _GEN_671 | _GEN_2 & _GEN_561 | _GEN_481 | _GEN_0 & _GEN_371) & (_GEN_291 ? io_wb_resps_0_bits_predicated : ~_GEN_164 & rob_predicated_18));
    rob_predicated_19 <= ~(_GEN_8 & _GEN_1134 | _GEN_1053 | _GEN_6 & _GEN_944) & (_GEN_863 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_754 | _GEN_673 | _GEN_2 & _GEN_564 | _GEN_483 | _GEN_0 & _GEN_374) & (_GEN_293 ? io_wb_resps_0_bits_predicated : ~_GEN_166 & rob_predicated_19));
    rob_predicated_20 <= ~(_GEN_8 & _GEN_1137 | _GEN_1055 | _GEN_6 & _GEN_947) & (_GEN_865 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_757 | _GEN_675 | _GEN_2 & _GEN_567 | _GEN_485 | _GEN_0 & _GEN_377) & (_GEN_295 ? io_wb_resps_0_bits_predicated : ~_GEN_168 & rob_predicated_20));
    rob_predicated_21 <= ~(_GEN_8 & _GEN_1140 | _GEN_1057 | _GEN_6 & _GEN_950) & (_GEN_867 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_760 | _GEN_677 | _GEN_2 & _GEN_570 | _GEN_487 | _GEN_0 & _GEN_380) & (_GEN_297 ? io_wb_resps_0_bits_predicated : ~_GEN_170 & rob_predicated_21));
    rob_predicated_22 <= ~(_GEN_8 & _GEN_1143 | _GEN_1059 | _GEN_6 & _GEN_953) & (_GEN_869 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_763 | _GEN_679 | _GEN_2 & _GEN_573 | _GEN_489 | _GEN_0 & _GEN_383) & (_GEN_299 ? io_wb_resps_0_bits_predicated : ~_GEN_172 & rob_predicated_22));
    rob_predicated_23 <= ~(_GEN_8 & _GEN_1146 | _GEN_1061 | _GEN_6 & _GEN_956) & (_GEN_871 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_766 | _GEN_681 | _GEN_2 & _GEN_576 | _GEN_491 | _GEN_0 & _GEN_386) & (_GEN_301 ? io_wb_resps_0_bits_predicated : ~_GEN_174 & rob_predicated_23));
    rob_predicated_24 <= ~(_GEN_8 & _GEN_1149 | _GEN_1063 | _GEN_6 & _GEN_959) & (_GEN_873 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_769 | _GEN_683 | _GEN_2 & _GEN_579 | _GEN_493 | _GEN_0 & _GEN_389) & (_GEN_303 ? io_wb_resps_0_bits_predicated : ~_GEN_176 & rob_predicated_24));
    rob_predicated_25 <= ~(_GEN_8 & _GEN_1152 | _GEN_1065 | _GEN_6 & _GEN_962) & (_GEN_875 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_772 | _GEN_685 | _GEN_2 & _GEN_582 | _GEN_495 | _GEN_0 & _GEN_392) & (_GEN_305 ? io_wb_resps_0_bits_predicated : ~_GEN_178 & rob_predicated_25));
    rob_predicated_26 <= ~(_GEN_8 & _GEN_1155 | _GEN_1067 | _GEN_6 & _GEN_965) & (_GEN_877 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_775 | _GEN_687 | _GEN_2 & _GEN_585 | _GEN_497 | _GEN_0 & _GEN_395) & (_GEN_307 ? io_wb_resps_0_bits_predicated : ~_GEN_180 & rob_predicated_26));
    rob_predicated_27 <= ~(_GEN_8 & _GEN_1158 | _GEN_1069 | _GEN_6 & _GEN_968) & (_GEN_879 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_778 | _GEN_689 | _GEN_2 & _GEN_588 | _GEN_499 | _GEN_0 & _GEN_398) & (_GEN_309 ? io_wb_resps_0_bits_predicated : ~_GEN_182 & rob_predicated_27));
    rob_predicated_28 <= ~(_GEN_8 & _GEN_1161 | _GEN_1071 | _GEN_6 & _GEN_971) & (_GEN_881 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_781 | _GEN_691 | _GEN_2 & _GEN_591 | _GEN_501 | _GEN_0 & _GEN_401) & (_GEN_311 ? io_wb_resps_0_bits_predicated : ~_GEN_184 & rob_predicated_28));
    rob_predicated_29 <= ~(_GEN_8 & _GEN_1164 | _GEN_1073 | _GEN_6 & _GEN_974) & (_GEN_883 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_784 | _GEN_693 | _GEN_2 & _GEN_594 | _GEN_503 | _GEN_0 & _GEN_404) & (_GEN_313 ? io_wb_resps_0_bits_predicated : ~_GEN_186 & rob_predicated_29));
    rob_predicated_30 <= ~(_GEN_8 & _GEN_1167 | _GEN_1075 | _GEN_6 & _GEN_977) & (_GEN_885 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & _GEN_787 | _GEN_695 | _GEN_2 & _GEN_597 | _GEN_505 | _GEN_0 & _GEN_407) & (_GEN_315 ? io_wb_resps_0_bits_predicated : ~_GEN_188 & rob_predicated_30));
    rob_predicated_31 <= ~(_GEN_8 & (&(io_wb_resps_9_bits_uop_rob_idx[6:2])) | _GEN_1076 | _GEN_6 & (&(io_wb_resps_7_bits_uop_rob_idx[6:2]))) & (_GEN_886 ? io_wb_resps_6_bits_predicated : ~(_GEN_4 & (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_696 | _GEN_2 & (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_506 | _GEN_0 & (&(io_wb_resps_1_bits_uop_rob_idx[6:2]))) & (_GEN_316 ? io_wb_resps_0_bits_predicated : ~_GEN_189 & rob_predicated_31));
    rob_bsy_1_0 <= ~_GEN_2446 & (_GEN_28 ? ~_GEN_2414 & _GEN_2287 : ~_GEN_2382 & _GEN_2287);
    rob_bsy_1_1 <= ~_GEN_2447 & (_GEN_28 ? ~_GEN_2415 & _GEN_2289 : ~_GEN_2383 & _GEN_2289);
    rob_bsy_1_2 <= ~_GEN_2448 & (_GEN_28 ? ~_GEN_2416 & _GEN_2291 : ~_GEN_2384 & _GEN_2291);
    rob_bsy_1_3 <= ~_GEN_2449 & (_GEN_28 ? ~_GEN_2417 & _GEN_2293 : ~_GEN_2385 & _GEN_2293);
    rob_bsy_1_4 <= ~_GEN_2450 & (_GEN_28 ? ~_GEN_2418 & _GEN_2295 : ~_GEN_2386 & _GEN_2295);
    rob_bsy_1_5 <= ~_GEN_2451 & (_GEN_28 ? ~_GEN_2419 & _GEN_2297 : ~_GEN_2387 & _GEN_2297);
    rob_bsy_1_6 <= ~_GEN_2452 & (_GEN_28 ? ~_GEN_2420 & _GEN_2299 : ~_GEN_2388 & _GEN_2299);
    rob_bsy_1_7 <= ~_GEN_2453 & (_GEN_28 ? ~_GEN_2421 & _GEN_2301 : ~_GEN_2389 & _GEN_2301);
    rob_bsy_1_8 <= ~_GEN_2454 & (_GEN_28 ? ~_GEN_2422 & _GEN_2303 : ~_GEN_2390 & _GEN_2303);
    rob_bsy_1_9 <= ~_GEN_2455 & (_GEN_28 ? ~_GEN_2423 & _GEN_2305 : ~_GEN_2391 & _GEN_2305);
    rob_bsy_1_10 <= ~_GEN_2456 & (_GEN_28 ? ~_GEN_2424 & _GEN_2307 : ~_GEN_2392 & _GEN_2307);
    rob_bsy_1_11 <= ~_GEN_2457 & (_GEN_28 ? ~_GEN_2425 & _GEN_2309 : ~_GEN_2393 & _GEN_2309);
    rob_bsy_1_12 <= ~_GEN_2458 & (_GEN_28 ? ~_GEN_2426 & _GEN_2311 : ~_GEN_2394 & _GEN_2311);
    rob_bsy_1_13 <= ~_GEN_2459 & (_GEN_28 ? ~_GEN_2427 & _GEN_2313 : ~_GEN_2395 & _GEN_2313);
    rob_bsy_1_14 <= ~_GEN_2460 & (_GEN_28 ? ~_GEN_2428 & _GEN_2315 : ~_GEN_2396 & _GEN_2315);
    rob_bsy_1_15 <= ~_GEN_2461 & (_GEN_28 ? ~_GEN_2429 & _GEN_2317 : ~_GEN_2397 & _GEN_2317);
    rob_bsy_1_16 <= ~_GEN_2462 & (_GEN_28 ? ~_GEN_2430 & _GEN_2319 : ~_GEN_2398 & _GEN_2319);
    rob_bsy_1_17 <= ~_GEN_2463 & (_GEN_28 ? ~_GEN_2431 & _GEN_2321 : ~_GEN_2399 & _GEN_2321);
    rob_bsy_1_18 <= ~_GEN_2464 & (_GEN_28 ? ~_GEN_2432 & _GEN_2323 : ~_GEN_2400 & _GEN_2323);
    rob_bsy_1_19 <= ~_GEN_2465 & (_GEN_28 ? ~_GEN_2433 & _GEN_2325 : ~_GEN_2401 & _GEN_2325);
    rob_bsy_1_20 <= ~_GEN_2466 & (_GEN_28 ? ~_GEN_2434 & _GEN_2327 : ~_GEN_2402 & _GEN_2327);
    rob_bsy_1_21 <= ~_GEN_2467 & (_GEN_28 ? ~_GEN_2435 & _GEN_2329 : ~_GEN_2403 & _GEN_2329);
    rob_bsy_1_22 <= ~_GEN_2468 & (_GEN_28 ? ~_GEN_2436 & _GEN_2331 : ~_GEN_2404 & _GEN_2331);
    rob_bsy_1_23 <= ~_GEN_2469 & (_GEN_28 ? ~_GEN_2437 & _GEN_2333 : ~_GEN_2405 & _GEN_2333);
    rob_bsy_1_24 <= ~_GEN_2470 & (_GEN_28 ? ~_GEN_2438 & _GEN_2335 : ~_GEN_2406 & _GEN_2335);
    rob_bsy_1_25 <= ~_GEN_2471 & (_GEN_28 ? ~_GEN_2439 & _GEN_2337 : ~_GEN_2407 & _GEN_2337);
    rob_bsy_1_26 <= ~_GEN_2472 & (_GEN_28 ? ~_GEN_2440 & _GEN_2339 : ~_GEN_2408 & _GEN_2339);
    rob_bsy_1_27 <= ~_GEN_2473 & (_GEN_28 ? ~_GEN_2441 & _GEN_2341 : ~_GEN_2409 & _GEN_2341);
    rob_bsy_1_28 <= ~_GEN_2474 & (_GEN_28 ? ~_GEN_2442 & _GEN_2343 : ~_GEN_2410 & _GEN_2343);
    rob_bsy_1_29 <= ~_GEN_2475 & (_GEN_28 ? ~_GEN_2443 & _GEN_2345 : ~_GEN_2411 & _GEN_2345);
    rob_bsy_1_30 <= ~_GEN_2476 & (_GEN_28 ? ~_GEN_2444 & _GEN_2347 : ~_GEN_2412 & _GEN_2347);
    rob_bsy_1_31 <= ~_GEN_2477 & (_GEN_28 ? ~_GEN_2445 & _GEN_2349 : ~_GEN_2413 & _GEN_2349);
    rob_unsafe_1_0 <= ~_GEN_2446 & (_GEN_28 ? ~_GEN_2414 & _GEN_2350 : ~_GEN_2382 & _GEN_2350);
    rob_unsafe_1_1 <= ~_GEN_2447 & (_GEN_28 ? ~_GEN_2415 & _GEN_2351 : ~_GEN_2383 & _GEN_2351);
    rob_unsafe_1_2 <= ~_GEN_2448 & (_GEN_28 ? ~_GEN_2416 & _GEN_2352 : ~_GEN_2384 & _GEN_2352);
    rob_unsafe_1_3 <= ~_GEN_2449 & (_GEN_28 ? ~_GEN_2417 & _GEN_2353 : ~_GEN_2385 & _GEN_2353);
    rob_unsafe_1_4 <= ~_GEN_2450 & (_GEN_28 ? ~_GEN_2418 & _GEN_2354 : ~_GEN_2386 & _GEN_2354);
    rob_unsafe_1_5 <= ~_GEN_2451 & (_GEN_28 ? ~_GEN_2419 & _GEN_2355 : ~_GEN_2387 & _GEN_2355);
    rob_unsafe_1_6 <= ~_GEN_2452 & (_GEN_28 ? ~_GEN_2420 & _GEN_2356 : ~_GEN_2388 & _GEN_2356);
    rob_unsafe_1_7 <= ~_GEN_2453 & (_GEN_28 ? ~_GEN_2421 & _GEN_2357 : ~_GEN_2389 & _GEN_2357);
    rob_unsafe_1_8 <= ~_GEN_2454 & (_GEN_28 ? ~_GEN_2422 & _GEN_2358 : ~_GEN_2390 & _GEN_2358);
    rob_unsafe_1_9 <= ~_GEN_2455 & (_GEN_28 ? ~_GEN_2423 & _GEN_2359 : ~_GEN_2391 & _GEN_2359);
    rob_unsafe_1_10 <= ~_GEN_2456 & (_GEN_28 ? ~_GEN_2424 & _GEN_2360 : ~_GEN_2392 & _GEN_2360);
    rob_unsafe_1_11 <= ~_GEN_2457 & (_GEN_28 ? ~_GEN_2425 & _GEN_2361 : ~_GEN_2393 & _GEN_2361);
    rob_unsafe_1_12 <= ~_GEN_2458 & (_GEN_28 ? ~_GEN_2426 & _GEN_2362 : ~_GEN_2394 & _GEN_2362);
    rob_unsafe_1_13 <= ~_GEN_2459 & (_GEN_28 ? ~_GEN_2427 & _GEN_2363 : ~_GEN_2395 & _GEN_2363);
    rob_unsafe_1_14 <= ~_GEN_2460 & (_GEN_28 ? ~_GEN_2428 & _GEN_2364 : ~_GEN_2396 & _GEN_2364);
    rob_unsafe_1_15 <= ~_GEN_2461 & (_GEN_28 ? ~_GEN_2429 & _GEN_2365 : ~_GEN_2397 & _GEN_2365);
    rob_unsafe_1_16 <= ~_GEN_2462 & (_GEN_28 ? ~_GEN_2430 & _GEN_2366 : ~_GEN_2398 & _GEN_2366);
    rob_unsafe_1_17 <= ~_GEN_2463 & (_GEN_28 ? ~_GEN_2431 & _GEN_2367 : ~_GEN_2399 & _GEN_2367);
    rob_unsafe_1_18 <= ~_GEN_2464 & (_GEN_28 ? ~_GEN_2432 & _GEN_2368 : ~_GEN_2400 & _GEN_2368);
    rob_unsafe_1_19 <= ~_GEN_2465 & (_GEN_28 ? ~_GEN_2433 & _GEN_2369 : ~_GEN_2401 & _GEN_2369);
    rob_unsafe_1_20 <= ~_GEN_2466 & (_GEN_28 ? ~_GEN_2434 & _GEN_2370 : ~_GEN_2402 & _GEN_2370);
    rob_unsafe_1_21 <= ~_GEN_2467 & (_GEN_28 ? ~_GEN_2435 & _GEN_2371 : ~_GEN_2403 & _GEN_2371);
    rob_unsafe_1_22 <= ~_GEN_2468 & (_GEN_28 ? ~_GEN_2436 & _GEN_2372 : ~_GEN_2404 & _GEN_2372);
    rob_unsafe_1_23 <= ~_GEN_2469 & (_GEN_28 ? ~_GEN_2437 & _GEN_2373 : ~_GEN_2405 & _GEN_2373);
    rob_unsafe_1_24 <= ~_GEN_2470 & (_GEN_28 ? ~_GEN_2438 & _GEN_2374 : ~_GEN_2406 & _GEN_2374);
    rob_unsafe_1_25 <= ~_GEN_2471 & (_GEN_28 ? ~_GEN_2439 & _GEN_2375 : ~_GEN_2407 & _GEN_2375);
    rob_unsafe_1_26 <= ~_GEN_2472 & (_GEN_28 ? ~_GEN_2440 & _GEN_2376 : ~_GEN_2408 & _GEN_2376);
    rob_unsafe_1_27 <= ~_GEN_2473 & (_GEN_28 ? ~_GEN_2441 & _GEN_2377 : ~_GEN_2409 & _GEN_2377);
    rob_unsafe_1_28 <= ~_GEN_2474 & (_GEN_28 ? ~_GEN_2442 & _GEN_2378 : ~_GEN_2410 & _GEN_2378);
    rob_unsafe_1_29 <= ~_GEN_2475 & (_GEN_28 ? ~_GEN_2443 & _GEN_2379 : ~_GEN_2411 & _GEN_2379);
    rob_unsafe_1_30 <= ~_GEN_2476 & (_GEN_28 ? ~_GEN_2444 & _GEN_2380 : ~_GEN_2412 & _GEN_2380);
    rob_unsafe_1_31 <= ~_GEN_2477 & (_GEN_28 ? ~_GEN_2445 & _GEN_2381 : ~_GEN_2413 & _GEN_2381);
    if (_GEN_1646) begin
      rob_uop_1_0_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_0_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_0_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_0_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_0_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_0_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_0_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_0_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_0_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_0_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_0_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_0_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_0_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_0_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_0_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_0_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_0_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_0_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_0_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2513) | ~rob_val_1_0) begin
      if (_GEN_1646)
        rob_uop_1_0_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_0_br_mask <= rob_uop_1_0_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1615)
      rob_uop_1_0_debug_fsrc <= 2'h3;
    else if (_GEN_1646)
      rob_uop_1_0_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1647) begin
      rob_uop_1_1_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_1_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_1_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_1_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_1_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_1_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_1_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_1_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_1_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_1_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_1_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_1_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_1_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_1_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_1_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_1_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_1_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_1_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_1_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2514) | ~rob_val_1_1) begin
      if (_GEN_1647)
        rob_uop_1_1_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_1_br_mask <= rob_uop_1_1_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1616)
      rob_uop_1_1_debug_fsrc <= 2'h3;
    else if (_GEN_1647)
      rob_uop_1_1_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1648) begin
      rob_uop_1_2_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_2_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_2_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_2_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_2_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_2_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_2_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_2_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_2_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_2_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_2_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_2_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_2_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_2_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_2_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_2_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_2_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_2_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_2_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2515) | ~rob_val_1_2) begin
      if (_GEN_1648)
        rob_uop_1_2_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_2_br_mask <= rob_uop_1_2_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1617)
      rob_uop_1_2_debug_fsrc <= 2'h3;
    else if (_GEN_1648)
      rob_uop_1_2_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1649) begin
      rob_uop_1_3_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_3_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_3_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_3_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_3_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_3_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_3_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_3_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_3_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_3_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_3_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_3_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_3_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_3_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_3_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_3_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_3_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_3_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_3_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2516) | ~rob_val_1_3) begin
      if (_GEN_1649)
        rob_uop_1_3_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_3_br_mask <= rob_uop_1_3_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1618)
      rob_uop_1_3_debug_fsrc <= 2'h3;
    else if (_GEN_1649)
      rob_uop_1_3_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1650) begin
      rob_uop_1_4_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_4_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_4_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_4_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_4_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_4_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_4_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_4_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_4_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_4_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_4_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_4_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_4_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_4_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_4_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_4_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_4_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_4_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_4_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2517) | ~rob_val_1_4) begin
      if (_GEN_1650)
        rob_uop_1_4_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_4_br_mask <= rob_uop_1_4_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1619)
      rob_uop_1_4_debug_fsrc <= 2'h3;
    else if (_GEN_1650)
      rob_uop_1_4_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1651) begin
      rob_uop_1_5_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_5_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_5_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_5_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_5_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_5_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_5_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_5_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_5_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_5_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_5_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_5_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_5_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_5_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_5_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_5_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_5_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_5_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_5_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2518) | ~rob_val_1_5) begin
      if (_GEN_1651)
        rob_uop_1_5_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_5_br_mask <= rob_uop_1_5_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1620)
      rob_uop_1_5_debug_fsrc <= 2'h3;
    else if (_GEN_1651)
      rob_uop_1_5_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1652) begin
      rob_uop_1_6_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_6_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_6_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_6_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_6_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_6_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_6_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_6_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_6_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_6_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_6_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_6_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_6_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_6_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_6_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_6_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_6_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_6_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_6_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2519) | ~rob_val_1_6) begin
      if (_GEN_1652)
        rob_uop_1_6_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_6_br_mask <= rob_uop_1_6_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1621)
      rob_uop_1_6_debug_fsrc <= 2'h3;
    else if (_GEN_1652)
      rob_uop_1_6_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1653) begin
      rob_uop_1_7_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_7_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_7_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_7_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_7_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_7_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_7_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_7_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_7_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_7_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_7_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_7_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_7_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_7_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_7_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_7_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_7_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_7_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_7_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2520) | ~rob_val_1_7) begin
      if (_GEN_1653)
        rob_uop_1_7_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_7_br_mask <= rob_uop_1_7_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1622)
      rob_uop_1_7_debug_fsrc <= 2'h3;
    else if (_GEN_1653)
      rob_uop_1_7_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1654) begin
      rob_uop_1_8_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_8_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_8_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_8_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_8_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_8_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_8_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_8_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_8_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_8_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_8_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_8_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_8_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_8_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_8_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_8_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_8_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_8_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_8_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2521) | ~rob_val_1_8) begin
      if (_GEN_1654)
        rob_uop_1_8_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_8_br_mask <= rob_uop_1_8_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1623)
      rob_uop_1_8_debug_fsrc <= 2'h3;
    else if (_GEN_1654)
      rob_uop_1_8_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1655) begin
      rob_uop_1_9_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_9_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_9_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_9_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_9_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_9_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_9_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_9_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_9_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_9_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_9_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_9_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_9_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_9_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_9_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_9_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_9_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_9_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_9_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2522) | ~rob_val_1_9) begin
      if (_GEN_1655)
        rob_uop_1_9_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_9_br_mask <= rob_uop_1_9_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1624)
      rob_uop_1_9_debug_fsrc <= 2'h3;
    else if (_GEN_1655)
      rob_uop_1_9_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1656) begin
      rob_uop_1_10_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_10_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_10_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_10_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_10_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_10_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_10_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_10_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_10_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_10_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_10_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_10_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_10_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_10_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_10_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_10_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_10_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_10_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_10_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2523) | ~rob_val_1_10) begin
      if (_GEN_1656)
        rob_uop_1_10_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_10_br_mask <= rob_uop_1_10_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1625)
      rob_uop_1_10_debug_fsrc <= 2'h3;
    else if (_GEN_1656)
      rob_uop_1_10_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1657) begin
      rob_uop_1_11_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_11_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_11_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_11_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_11_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_11_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_11_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_11_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_11_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_11_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_11_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_11_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_11_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_11_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_11_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_11_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_11_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_11_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_11_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2524) | ~rob_val_1_11) begin
      if (_GEN_1657)
        rob_uop_1_11_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_11_br_mask <= rob_uop_1_11_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1626)
      rob_uop_1_11_debug_fsrc <= 2'h3;
    else if (_GEN_1657)
      rob_uop_1_11_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1658) begin
      rob_uop_1_12_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_12_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_12_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_12_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_12_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_12_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_12_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_12_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_12_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_12_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_12_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_12_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_12_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_12_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_12_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_12_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_12_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_12_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_12_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2525) | ~rob_val_1_12) begin
      if (_GEN_1658)
        rob_uop_1_12_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_12_br_mask <= rob_uop_1_12_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1627)
      rob_uop_1_12_debug_fsrc <= 2'h3;
    else if (_GEN_1658)
      rob_uop_1_12_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1659) begin
      rob_uop_1_13_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_13_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_13_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_13_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_13_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_13_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_13_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_13_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_13_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_13_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_13_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_13_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_13_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_13_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_13_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_13_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_13_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_13_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_13_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2526) | ~rob_val_1_13) begin
      if (_GEN_1659)
        rob_uop_1_13_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_13_br_mask <= rob_uop_1_13_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1628)
      rob_uop_1_13_debug_fsrc <= 2'h3;
    else if (_GEN_1659)
      rob_uop_1_13_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1660) begin
      rob_uop_1_14_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_14_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_14_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_14_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_14_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_14_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_14_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_14_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_14_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_14_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_14_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_14_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_14_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_14_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_14_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_14_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_14_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_14_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_14_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2527) | ~rob_val_1_14) begin
      if (_GEN_1660)
        rob_uop_1_14_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_14_br_mask <= rob_uop_1_14_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1629)
      rob_uop_1_14_debug_fsrc <= 2'h3;
    else if (_GEN_1660)
      rob_uop_1_14_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1661) begin
      rob_uop_1_15_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_15_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_15_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_15_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_15_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_15_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_15_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_15_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_15_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_15_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_15_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_15_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_15_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_15_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_15_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_15_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_15_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_15_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_15_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2528) | ~rob_val_1_15) begin
      if (_GEN_1661)
        rob_uop_1_15_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_15_br_mask <= rob_uop_1_15_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1630)
      rob_uop_1_15_debug_fsrc <= 2'h3;
    else if (_GEN_1661)
      rob_uop_1_15_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1662) begin
      rob_uop_1_16_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_16_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_16_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_16_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_16_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_16_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_16_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_16_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_16_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_16_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_16_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_16_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_16_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_16_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_16_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_16_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_16_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_16_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_16_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2529) | ~rob_val_1_16) begin
      if (_GEN_1662)
        rob_uop_1_16_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_16_br_mask <= rob_uop_1_16_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1631)
      rob_uop_1_16_debug_fsrc <= 2'h3;
    else if (_GEN_1662)
      rob_uop_1_16_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1663) begin
      rob_uop_1_17_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_17_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_17_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_17_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_17_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_17_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_17_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_17_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_17_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_17_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_17_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_17_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_17_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_17_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_17_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_17_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_17_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_17_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_17_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2530) | ~rob_val_1_17) begin
      if (_GEN_1663)
        rob_uop_1_17_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_17_br_mask <= rob_uop_1_17_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1632)
      rob_uop_1_17_debug_fsrc <= 2'h3;
    else if (_GEN_1663)
      rob_uop_1_17_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1664) begin
      rob_uop_1_18_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_18_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_18_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_18_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_18_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_18_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_18_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_18_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_18_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_18_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_18_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_18_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_18_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_18_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_18_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_18_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_18_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_18_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_18_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2531) | ~rob_val_1_18) begin
      if (_GEN_1664)
        rob_uop_1_18_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_18_br_mask <= rob_uop_1_18_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1633)
      rob_uop_1_18_debug_fsrc <= 2'h3;
    else if (_GEN_1664)
      rob_uop_1_18_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1665) begin
      rob_uop_1_19_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_19_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_19_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_19_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_19_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_19_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_19_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_19_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_19_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_19_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_19_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_19_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_19_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_19_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_19_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_19_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_19_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_19_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_19_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2532) | ~rob_val_1_19) begin
      if (_GEN_1665)
        rob_uop_1_19_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_19_br_mask <= rob_uop_1_19_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1634)
      rob_uop_1_19_debug_fsrc <= 2'h3;
    else if (_GEN_1665)
      rob_uop_1_19_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1666) begin
      rob_uop_1_20_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_20_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_20_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_20_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_20_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_20_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_20_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_20_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_20_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_20_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_20_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_20_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_20_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_20_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_20_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_20_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_20_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_20_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_20_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2533) | ~rob_val_1_20) begin
      if (_GEN_1666)
        rob_uop_1_20_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_20_br_mask <= rob_uop_1_20_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1635)
      rob_uop_1_20_debug_fsrc <= 2'h3;
    else if (_GEN_1666)
      rob_uop_1_20_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1667) begin
      rob_uop_1_21_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_21_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_21_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_21_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_21_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_21_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_21_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_21_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_21_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_21_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_21_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_21_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_21_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_21_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_21_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_21_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_21_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_21_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_21_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2534) | ~rob_val_1_21) begin
      if (_GEN_1667)
        rob_uop_1_21_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_21_br_mask <= rob_uop_1_21_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1636)
      rob_uop_1_21_debug_fsrc <= 2'h3;
    else if (_GEN_1667)
      rob_uop_1_21_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1668) begin
      rob_uop_1_22_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_22_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_22_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_22_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_22_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_22_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_22_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_22_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_22_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_22_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_22_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_22_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_22_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_22_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_22_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_22_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_22_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_22_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_22_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2535) | ~rob_val_1_22) begin
      if (_GEN_1668)
        rob_uop_1_22_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_22_br_mask <= rob_uop_1_22_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1637)
      rob_uop_1_22_debug_fsrc <= 2'h3;
    else if (_GEN_1668)
      rob_uop_1_22_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1669) begin
      rob_uop_1_23_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_23_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_23_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_23_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_23_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_23_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_23_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_23_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_23_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_23_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_23_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_23_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_23_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_23_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_23_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_23_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_23_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_23_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_23_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2536) | ~rob_val_1_23) begin
      if (_GEN_1669)
        rob_uop_1_23_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_23_br_mask <= rob_uop_1_23_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1638)
      rob_uop_1_23_debug_fsrc <= 2'h3;
    else if (_GEN_1669)
      rob_uop_1_23_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1670) begin
      rob_uop_1_24_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_24_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_24_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_24_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_24_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_24_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_24_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_24_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_24_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_24_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_24_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_24_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_24_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_24_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_24_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_24_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_24_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_24_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_24_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2537) | ~rob_val_1_24) begin
      if (_GEN_1670)
        rob_uop_1_24_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_24_br_mask <= rob_uop_1_24_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1639)
      rob_uop_1_24_debug_fsrc <= 2'h3;
    else if (_GEN_1670)
      rob_uop_1_24_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1671) begin
      rob_uop_1_25_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_25_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_25_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_25_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_25_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_25_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_25_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_25_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_25_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_25_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_25_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_25_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_25_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_25_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_25_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_25_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_25_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_25_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_25_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2538) | ~rob_val_1_25) begin
      if (_GEN_1671)
        rob_uop_1_25_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_25_br_mask <= rob_uop_1_25_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1640)
      rob_uop_1_25_debug_fsrc <= 2'h3;
    else if (_GEN_1671)
      rob_uop_1_25_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1672) begin
      rob_uop_1_26_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_26_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_26_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_26_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_26_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_26_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_26_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_26_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_26_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_26_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_26_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_26_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_26_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_26_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_26_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_26_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_26_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_26_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_26_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2539) | ~rob_val_1_26) begin
      if (_GEN_1672)
        rob_uop_1_26_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_26_br_mask <= rob_uop_1_26_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1641)
      rob_uop_1_26_debug_fsrc <= 2'h3;
    else if (_GEN_1672)
      rob_uop_1_26_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1673) begin
      rob_uop_1_27_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_27_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_27_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_27_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_27_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_27_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_27_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_27_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_27_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_27_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_27_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_27_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_27_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_27_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_27_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_27_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_27_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_27_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_27_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2540) | ~rob_val_1_27) begin
      if (_GEN_1673)
        rob_uop_1_27_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_27_br_mask <= rob_uop_1_27_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1642)
      rob_uop_1_27_debug_fsrc <= 2'h3;
    else if (_GEN_1673)
      rob_uop_1_27_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1674) begin
      rob_uop_1_28_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_28_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_28_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_28_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_28_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_28_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_28_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_28_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_28_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_28_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_28_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_28_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_28_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_28_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_28_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_28_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_28_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_28_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_28_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2541) | ~rob_val_1_28) begin
      if (_GEN_1674)
        rob_uop_1_28_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_28_br_mask <= rob_uop_1_28_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1643)
      rob_uop_1_28_debug_fsrc <= 2'h3;
    else if (_GEN_1674)
      rob_uop_1_28_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1675) begin
      rob_uop_1_29_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_29_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_29_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_29_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_29_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_29_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_29_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_29_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_29_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_29_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_29_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_29_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_29_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_29_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_29_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_29_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_29_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_29_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_29_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2542) | ~rob_val_1_29) begin
      if (_GEN_1675)
        rob_uop_1_29_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_29_br_mask <= rob_uop_1_29_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1644)
      rob_uop_1_29_debug_fsrc <= 2'h3;
    else if (_GEN_1675)
      rob_uop_1_29_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1676) begin
      rob_uop_1_30_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_30_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_30_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_30_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_30_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_30_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_30_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_30_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_30_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_30_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_30_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_30_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_30_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_30_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_30_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_30_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_30_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_30_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_30_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2543) | ~rob_val_1_30) begin
      if (_GEN_1676)
        rob_uop_1_30_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_30_br_mask <= rob_uop_1_30_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & _GEN_1645)
      rob_uop_1_30_debug_fsrc <= 2'h3;
    else if (_GEN_1676)
      rob_uop_1_30_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    if (_GEN_1677) begin
      rob_uop_1_31_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_31_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_31_is_br <= io_enq_uops_1_is_br;
      rob_uop_1_31_is_jalr <= io_enq_uops_1_is_jalr;
      rob_uop_1_31_is_jal <= io_enq_uops_1_is_jal;
      rob_uop_1_31_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_31_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_31_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_31_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_31_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_31_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_31_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_31_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_31_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_31_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_31_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_31_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_31_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_31_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2544) | ~rob_val_1_31) begin
      if (_GEN_1677)
        rob_uop_1_31_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_31_br_mask <= rob_uop_1_31_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_32 & (&(io_brupdate_b2_uop_rob_idx[6:2])))
      rob_uop_1_31_debug_fsrc <= 2'h3;
    else if (_GEN_1677)
      rob_uop_1_31_debug_fsrc <= io_enq_uops_1_debug_fsrc;
    rob_exception_1_0 <= ~_GEN_2481 & (_GEN_30 & _GEN_1489 | (_GEN_1646 ? io_enq_uops_1_exception : rob_exception_1_0));
    rob_exception_1_1 <= ~_GEN_2482 & (_GEN_30 & _GEN_1490 | (_GEN_1647 ? io_enq_uops_1_exception : rob_exception_1_1));
    rob_exception_1_2 <= ~_GEN_2483 & (_GEN_30 & _GEN_1491 | (_GEN_1648 ? io_enq_uops_1_exception : rob_exception_1_2));
    rob_exception_1_3 <= ~_GEN_2484 & (_GEN_30 & _GEN_1492 | (_GEN_1649 ? io_enq_uops_1_exception : rob_exception_1_3));
    rob_exception_1_4 <= ~_GEN_2485 & (_GEN_30 & _GEN_1493 | (_GEN_1650 ? io_enq_uops_1_exception : rob_exception_1_4));
    rob_exception_1_5 <= ~_GEN_2486 & (_GEN_30 & _GEN_1494 | (_GEN_1651 ? io_enq_uops_1_exception : rob_exception_1_5));
    rob_exception_1_6 <= ~_GEN_2487 & (_GEN_30 & _GEN_1495 | (_GEN_1652 ? io_enq_uops_1_exception : rob_exception_1_6));
    rob_exception_1_7 <= ~_GEN_2488 & (_GEN_30 & _GEN_1496 | (_GEN_1653 ? io_enq_uops_1_exception : rob_exception_1_7));
    rob_exception_1_8 <= ~_GEN_2489 & (_GEN_30 & _GEN_1497 | (_GEN_1654 ? io_enq_uops_1_exception : rob_exception_1_8));
    rob_exception_1_9 <= ~_GEN_2490 & (_GEN_30 & _GEN_1498 | (_GEN_1655 ? io_enq_uops_1_exception : rob_exception_1_9));
    rob_exception_1_10 <= ~_GEN_2491 & (_GEN_30 & _GEN_1499 | (_GEN_1656 ? io_enq_uops_1_exception : rob_exception_1_10));
    rob_exception_1_11 <= ~_GEN_2492 & (_GEN_30 & _GEN_1500 | (_GEN_1657 ? io_enq_uops_1_exception : rob_exception_1_11));
    rob_exception_1_12 <= ~_GEN_2493 & (_GEN_30 & _GEN_1501 | (_GEN_1658 ? io_enq_uops_1_exception : rob_exception_1_12));
    rob_exception_1_13 <= ~_GEN_2494 & (_GEN_30 & _GEN_1502 | (_GEN_1659 ? io_enq_uops_1_exception : rob_exception_1_13));
    rob_exception_1_14 <= ~_GEN_2495 & (_GEN_30 & _GEN_1503 | (_GEN_1660 ? io_enq_uops_1_exception : rob_exception_1_14));
    rob_exception_1_15 <= ~_GEN_2496 & (_GEN_30 & _GEN_1504 | (_GEN_1661 ? io_enq_uops_1_exception : rob_exception_1_15));
    rob_exception_1_16 <= ~_GEN_2497 & (_GEN_30 & _GEN_1505 | (_GEN_1662 ? io_enq_uops_1_exception : rob_exception_1_16));
    rob_exception_1_17 <= ~_GEN_2498 & (_GEN_30 & _GEN_1506 | (_GEN_1663 ? io_enq_uops_1_exception : rob_exception_1_17));
    rob_exception_1_18 <= ~_GEN_2499 & (_GEN_30 & _GEN_1507 | (_GEN_1664 ? io_enq_uops_1_exception : rob_exception_1_18));
    rob_exception_1_19 <= ~_GEN_2500 & (_GEN_30 & _GEN_1508 | (_GEN_1665 ? io_enq_uops_1_exception : rob_exception_1_19));
    rob_exception_1_20 <= ~_GEN_2501 & (_GEN_30 & _GEN_1509 | (_GEN_1666 ? io_enq_uops_1_exception : rob_exception_1_20));
    rob_exception_1_21 <= ~_GEN_2502 & (_GEN_30 & _GEN_1510 | (_GEN_1667 ? io_enq_uops_1_exception : rob_exception_1_21));
    rob_exception_1_22 <= ~_GEN_2503 & (_GEN_30 & _GEN_1511 | (_GEN_1668 ? io_enq_uops_1_exception : rob_exception_1_22));
    rob_exception_1_23 <= ~_GEN_2504 & (_GEN_30 & _GEN_1512 | (_GEN_1669 ? io_enq_uops_1_exception : rob_exception_1_23));
    rob_exception_1_24 <= ~_GEN_2505 & (_GEN_30 & _GEN_1513 | (_GEN_1670 ? io_enq_uops_1_exception : rob_exception_1_24));
    rob_exception_1_25 <= ~_GEN_2506 & (_GEN_30 & _GEN_1514 | (_GEN_1671 ? io_enq_uops_1_exception : rob_exception_1_25));
    rob_exception_1_26 <= ~_GEN_2507 & (_GEN_30 & _GEN_1515 | (_GEN_1672 ? io_enq_uops_1_exception : rob_exception_1_26));
    rob_exception_1_27 <= ~_GEN_2508 & (_GEN_30 & _GEN_1516 | (_GEN_1673 ? io_enq_uops_1_exception : rob_exception_1_27));
    rob_exception_1_28 <= ~_GEN_2509 & (_GEN_30 & _GEN_1517 | (_GEN_1674 ? io_enq_uops_1_exception : rob_exception_1_28));
    rob_exception_1_29 <= ~_GEN_2510 & (_GEN_30 & _GEN_1518 | (_GEN_1675 ? io_enq_uops_1_exception : rob_exception_1_29));
    rob_exception_1_30 <= ~_GEN_2511 & (_GEN_30 & _GEN_1519 | (_GEN_1676 ? io_enq_uops_1_exception : rob_exception_1_30));
    rob_exception_1_31 <= ~_GEN_2512 & (_GEN_30 & (&(io_lxcpt_bits_uop_rob_idx[6:2])) | (_GEN_1677 ? io_enq_uops_1_exception : rob_exception_1_31));
    rob_predicated_1_0 <= ~(_GEN_26 & _GEN_1077 | _GEN_2254 | _GEN_24 & _GEN_887) & (_GEN_2126 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_697 | _GEN_1998 | _GEN_20 & _GEN_507 | _GEN_1870 | _GEN_18 & _GEN_317) & (_GEN_1742 ? io_wb_resps_0_bits_predicated : ~_GEN_1646 & rob_predicated_1_0));
    rob_predicated_1_1 <= ~(_GEN_26 & _GEN_1080 | _GEN_2255 | _GEN_24 & _GEN_890) & (_GEN_2127 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_700 | _GEN_1999 | _GEN_20 & _GEN_510 | _GEN_1871 | _GEN_18 & _GEN_320) & (_GEN_1743 ? io_wb_resps_0_bits_predicated : ~_GEN_1647 & rob_predicated_1_1));
    rob_predicated_1_2 <= ~(_GEN_26 & _GEN_1083 | _GEN_2256 | _GEN_24 & _GEN_893) & (_GEN_2128 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_703 | _GEN_2000 | _GEN_20 & _GEN_513 | _GEN_1872 | _GEN_18 & _GEN_323) & (_GEN_1744 ? io_wb_resps_0_bits_predicated : ~_GEN_1648 & rob_predicated_1_2));
    rob_predicated_1_3 <= ~(_GEN_26 & _GEN_1086 | _GEN_2257 | _GEN_24 & _GEN_896) & (_GEN_2129 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_706 | _GEN_2001 | _GEN_20 & _GEN_516 | _GEN_1873 | _GEN_18 & _GEN_326) & (_GEN_1745 ? io_wb_resps_0_bits_predicated : ~_GEN_1649 & rob_predicated_1_3));
    rob_predicated_1_4 <= ~(_GEN_26 & _GEN_1089 | _GEN_2258 | _GEN_24 & _GEN_899) & (_GEN_2130 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_709 | _GEN_2002 | _GEN_20 & _GEN_519 | _GEN_1874 | _GEN_18 & _GEN_329) & (_GEN_1746 ? io_wb_resps_0_bits_predicated : ~_GEN_1650 & rob_predicated_1_4));
    rob_predicated_1_5 <= ~(_GEN_26 & _GEN_1092 | _GEN_2259 | _GEN_24 & _GEN_902) & (_GEN_2131 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_712 | _GEN_2003 | _GEN_20 & _GEN_522 | _GEN_1875 | _GEN_18 & _GEN_332) & (_GEN_1747 ? io_wb_resps_0_bits_predicated : ~_GEN_1651 & rob_predicated_1_5));
    rob_predicated_1_6 <= ~(_GEN_26 & _GEN_1095 | _GEN_2260 | _GEN_24 & _GEN_905) & (_GEN_2132 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_715 | _GEN_2004 | _GEN_20 & _GEN_525 | _GEN_1876 | _GEN_18 & _GEN_335) & (_GEN_1748 ? io_wb_resps_0_bits_predicated : ~_GEN_1652 & rob_predicated_1_6));
    rob_predicated_1_7 <= ~(_GEN_26 & _GEN_1098 | _GEN_2261 | _GEN_24 & _GEN_908) & (_GEN_2133 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_718 | _GEN_2005 | _GEN_20 & _GEN_528 | _GEN_1877 | _GEN_18 & _GEN_338) & (_GEN_1749 ? io_wb_resps_0_bits_predicated : ~_GEN_1653 & rob_predicated_1_7));
    rob_predicated_1_8 <= ~(_GEN_26 & _GEN_1101 | _GEN_2262 | _GEN_24 & _GEN_911) & (_GEN_2134 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_721 | _GEN_2006 | _GEN_20 & _GEN_531 | _GEN_1878 | _GEN_18 & _GEN_341) & (_GEN_1750 ? io_wb_resps_0_bits_predicated : ~_GEN_1654 & rob_predicated_1_8));
    rob_predicated_1_9 <= ~(_GEN_26 & _GEN_1104 | _GEN_2263 | _GEN_24 & _GEN_914) & (_GEN_2135 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_724 | _GEN_2007 | _GEN_20 & _GEN_534 | _GEN_1879 | _GEN_18 & _GEN_344) & (_GEN_1751 ? io_wb_resps_0_bits_predicated : ~_GEN_1655 & rob_predicated_1_9));
    rob_predicated_1_10 <= ~(_GEN_26 & _GEN_1107 | _GEN_2264 | _GEN_24 & _GEN_917) & (_GEN_2136 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_727 | _GEN_2008 | _GEN_20 & _GEN_537 | _GEN_1880 | _GEN_18 & _GEN_347) & (_GEN_1752 ? io_wb_resps_0_bits_predicated : ~_GEN_1656 & rob_predicated_1_10));
    rob_predicated_1_11 <= ~(_GEN_26 & _GEN_1110 | _GEN_2265 | _GEN_24 & _GEN_920) & (_GEN_2137 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_730 | _GEN_2009 | _GEN_20 & _GEN_540 | _GEN_1881 | _GEN_18 & _GEN_350) & (_GEN_1753 ? io_wb_resps_0_bits_predicated : ~_GEN_1657 & rob_predicated_1_11));
    rob_predicated_1_12 <= ~(_GEN_26 & _GEN_1113 | _GEN_2266 | _GEN_24 & _GEN_923) & (_GEN_2138 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_733 | _GEN_2010 | _GEN_20 & _GEN_543 | _GEN_1882 | _GEN_18 & _GEN_353) & (_GEN_1754 ? io_wb_resps_0_bits_predicated : ~_GEN_1658 & rob_predicated_1_12));
    rob_predicated_1_13 <= ~(_GEN_26 & _GEN_1116 | _GEN_2267 | _GEN_24 & _GEN_926) & (_GEN_2139 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_736 | _GEN_2011 | _GEN_20 & _GEN_546 | _GEN_1883 | _GEN_18 & _GEN_356) & (_GEN_1755 ? io_wb_resps_0_bits_predicated : ~_GEN_1659 & rob_predicated_1_13));
    rob_predicated_1_14 <= ~(_GEN_26 & _GEN_1119 | _GEN_2268 | _GEN_24 & _GEN_929) & (_GEN_2140 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_739 | _GEN_2012 | _GEN_20 & _GEN_549 | _GEN_1884 | _GEN_18 & _GEN_359) & (_GEN_1756 ? io_wb_resps_0_bits_predicated : ~_GEN_1660 & rob_predicated_1_14));
    rob_predicated_1_15 <= ~(_GEN_26 & _GEN_1122 | _GEN_2269 | _GEN_24 & _GEN_932) & (_GEN_2141 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_742 | _GEN_2013 | _GEN_20 & _GEN_552 | _GEN_1885 | _GEN_18 & _GEN_362) & (_GEN_1757 ? io_wb_resps_0_bits_predicated : ~_GEN_1661 & rob_predicated_1_15));
    rob_predicated_1_16 <= ~(_GEN_26 & _GEN_1125 | _GEN_2270 | _GEN_24 & _GEN_935) & (_GEN_2142 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_745 | _GEN_2014 | _GEN_20 & _GEN_555 | _GEN_1886 | _GEN_18 & _GEN_365) & (_GEN_1758 ? io_wb_resps_0_bits_predicated : ~_GEN_1662 & rob_predicated_1_16));
    rob_predicated_1_17 <= ~(_GEN_26 & _GEN_1128 | _GEN_2271 | _GEN_24 & _GEN_938) & (_GEN_2143 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_748 | _GEN_2015 | _GEN_20 & _GEN_558 | _GEN_1887 | _GEN_18 & _GEN_368) & (_GEN_1759 ? io_wb_resps_0_bits_predicated : ~_GEN_1663 & rob_predicated_1_17));
    rob_predicated_1_18 <= ~(_GEN_26 & _GEN_1131 | _GEN_2272 | _GEN_24 & _GEN_941) & (_GEN_2144 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_751 | _GEN_2016 | _GEN_20 & _GEN_561 | _GEN_1888 | _GEN_18 & _GEN_371) & (_GEN_1760 ? io_wb_resps_0_bits_predicated : ~_GEN_1664 & rob_predicated_1_18));
    rob_predicated_1_19 <= ~(_GEN_26 & _GEN_1134 | _GEN_2273 | _GEN_24 & _GEN_944) & (_GEN_2145 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_754 | _GEN_2017 | _GEN_20 & _GEN_564 | _GEN_1889 | _GEN_18 & _GEN_374) & (_GEN_1761 ? io_wb_resps_0_bits_predicated : ~_GEN_1665 & rob_predicated_1_19));
    rob_predicated_1_20 <= ~(_GEN_26 & _GEN_1137 | _GEN_2274 | _GEN_24 & _GEN_947) & (_GEN_2146 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_757 | _GEN_2018 | _GEN_20 & _GEN_567 | _GEN_1890 | _GEN_18 & _GEN_377) & (_GEN_1762 ? io_wb_resps_0_bits_predicated : ~_GEN_1666 & rob_predicated_1_20));
    rob_predicated_1_21 <= ~(_GEN_26 & _GEN_1140 | _GEN_2275 | _GEN_24 & _GEN_950) & (_GEN_2147 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_760 | _GEN_2019 | _GEN_20 & _GEN_570 | _GEN_1891 | _GEN_18 & _GEN_380) & (_GEN_1763 ? io_wb_resps_0_bits_predicated : ~_GEN_1667 & rob_predicated_1_21));
    rob_predicated_1_22 <= ~(_GEN_26 & _GEN_1143 | _GEN_2276 | _GEN_24 & _GEN_953) & (_GEN_2148 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_763 | _GEN_2020 | _GEN_20 & _GEN_573 | _GEN_1892 | _GEN_18 & _GEN_383) & (_GEN_1764 ? io_wb_resps_0_bits_predicated : ~_GEN_1668 & rob_predicated_1_22));
    rob_predicated_1_23 <= ~(_GEN_26 & _GEN_1146 | _GEN_2277 | _GEN_24 & _GEN_956) & (_GEN_2149 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_766 | _GEN_2021 | _GEN_20 & _GEN_576 | _GEN_1893 | _GEN_18 & _GEN_386) & (_GEN_1765 ? io_wb_resps_0_bits_predicated : ~_GEN_1669 & rob_predicated_1_23));
    rob_predicated_1_24 <= ~(_GEN_26 & _GEN_1149 | _GEN_2278 | _GEN_24 & _GEN_959) & (_GEN_2150 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_769 | _GEN_2022 | _GEN_20 & _GEN_579 | _GEN_1894 | _GEN_18 & _GEN_389) & (_GEN_1766 ? io_wb_resps_0_bits_predicated : ~_GEN_1670 & rob_predicated_1_24));
    rob_predicated_1_25 <= ~(_GEN_26 & _GEN_1152 | _GEN_2279 | _GEN_24 & _GEN_962) & (_GEN_2151 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_772 | _GEN_2023 | _GEN_20 & _GEN_582 | _GEN_1895 | _GEN_18 & _GEN_392) & (_GEN_1767 ? io_wb_resps_0_bits_predicated : ~_GEN_1671 & rob_predicated_1_25));
    rob_predicated_1_26 <= ~(_GEN_26 & _GEN_1155 | _GEN_2280 | _GEN_24 & _GEN_965) & (_GEN_2152 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_775 | _GEN_2024 | _GEN_20 & _GEN_585 | _GEN_1896 | _GEN_18 & _GEN_395) & (_GEN_1768 ? io_wb_resps_0_bits_predicated : ~_GEN_1672 & rob_predicated_1_26));
    rob_predicated_1_27 <= ~(_GEN_26 & _GEN_1158 | _GEN_2281 | _GEN_24 & _GEN_968) & (_GEN_2153 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_778 | _GEN_2025 | _GEN_20 & _GEN_588 | _GEN_1897 | _GEN_18 & _GEN_398) & (_GEN_1769 ? io_wb_resps_0_bits_predicated : ~_GEN_1673 & rob_predicated_1_27));
    rob_predicated_1_28 <= ~(_GEN_26 & _GEN_1161 | _GEN_2282 | _GEN_24 & _GEN_971) & (_GEN_2154 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_781 | _GEN_2026 | _GEN_20 & _GEN_591 | _GEN_1898 | _GEN_18 & _GEN_401) & (_GEN_1770 ? io_wb_resps_0_bits_predicated : ~_GEN_1674 & rob_predicated_1_28));
    rob_predicated_1_29 <= ~(_GEN_26 & _GEN_1164 | _GEN_2283 | _GEN_24 & _GEN_974) & (_GEN_2155 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_784 | _GEN_2027 | _GEN_20 & _GEN_594 | _GEN_1899 | _GEN_18 & _GEN_404) & (_GEN_1771 ? io_wb_resps_0_bits_predicated : ~_GEN_1675 & rob_predicated_1_29));
    rob_predicated_1_30 <= ~(_GEN_26 & _GEN_1167 | _GEN_2284 | _GEN_24 & _GEN_977) & (_GEN_2156 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & _GEN_787 | _GEN_2028 | _GEN_20 & _GEN_597 | _GEN_1900 | _GEN_18 & _GEN_407) & (_GEN_1772 ? io_wb_resps_0_bits_predicated : ~_GEN_1676 & rob_predicated_1_30));
    rob_predicated_1_31 <= ~(_GEN_26 & (&(io_wb_resps_9_bits_uop_rob_idx[6:2])) | _GEN_2285 | _GEN_24 & (&(io_wb_resps_7_bits_uop_rob_idx[6:2]))) & (_GEN_2157 ? io_wb_resps_6_bits_predicated : ~(_GEN_22 & (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_2029 | _GEN_20 & (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_1901 | _GEN_18 & (&(io_wb_resps_1_bits_uop_rob_idx[6:2]))) & (_GEN_1773 ? io_wb_resps_0_bits_predicated : ~_GEN_1677 & rob_predicated_1_31));
    rob_bsy_2_0 <= ~_GEN_3345 & (_GEN_44 ? ~_GEN_3313 & _GEN_3186 : ~_GEN_3281 & _GEN_3186);
    rob_bsy_2_1 <= ~_GEN_3346 & (_GEN_44 ? ~_GEN_3314 & _GEN_3188 : ~_GEN_3282 & _GEN_3188);
    rob_bsy_2_2 <= ~_GEN_3347 & (_GEN_44 ? ~_GEN_3315 & _GEN_3190 : ~_GEN_3283 & _GEN_3190);
    rob_bsy_2_3 <= ~_GEN_3348 & (_GEN_44 ? ~_GEN_3316 & _GEN_3192 : ~_GEN_3284 & _GEN_3192);
    rob_bsy_2_4 <= ~_GEN_3349 & (_GEN_44 ? ~_GEN_3317 & _GEN_3194 : ~_GEN_3285 & _GEN_3194);
    rob_bsy_2_5 <= ~_GEN_3350 & (_GEN_44 ? ~_GEN_3318 & _GEN_3196 : ~_GEN_3286 & _GEN_3196);
    rob_bsy_2_6 <= ~_GEN_3351 & (_GEN_44 ? ~_GEN_3319 & _GEN_3198 : ~_GEN_3287 & _GEN_3198);
    rob_bsy_2_7 <= ~_GEN_3352 & (_GEN_44 ? ~_GEN_3320 & _GEN_3200 : ~_GEN_3288 & _GEN_3200);
    rob_bsy_2_8 <= ~_GEN_3353 & (_GEN_44 ? ~_GEN_3321 & _GEN_3202 : ~_GEN_3289 & _GEN_3202);
    rob_bsy_2_9 <= ~_GEN_3354 & (_GEN_44 ? ~_GEN_3322 & _GEN_3204 : ~_GEN_3290 & _GEN_3204);
    rob_bsy_2_10 <= ~_GEN_3355 & (_GEN_44 ? ~_GEN_3323 & _GEN_3206 : ~_GEN_3291 & _GEN_3206);
    rob_bsy_2_11 <= ~_GEN_3356 & (_GEN_44 ? ~_GEN_3324 & _GEN_3208 : ~_GEN_3292 & _GEN_3208);
    rob_bsy_2_12 <= ~_GEN_3357 & (_GEN_44 ? ~_GEN_3325 & _GEN_3210 : ~_GEN_3293 & _GEN_3210);
    rob_bsy_2_13 <= ~_GEN_3358 & (_GEN_44 ? ~_GEN_3326 & _GEN_3212 : ~_GEN_3294 & _GEN_3212);
    rob_bsy_2_14 <= ~_GEN_3359 & (_GEN_44 ? ~_GEN_3327 & _GEN_3214 : ~_GEN_3295 & _GEN_3214);
    rob_bsy_2_15 <= ~_GEN_3360 & (_GEN_44 ? ~_GEN_3328 & _GEN_3216 : ~_GEN_3296 & _GEN_3216);
    rob_bsy_2_16 <= ~_GEN_3361 & (_GEN_44 ? ~_GEN_3329 & _GEN_3218 : ~_GEN_3297 & _GEN_3218);
    rob_bsy_2_17 <= ~_GEN_3362 & (_GEN_44 ? ~_GEN_3330 & _GEN_3220 : ~_GEN_3298 & _GEN_3220);
    rob_bsy_2_18 <= ~_GEN_3363 & (_GEN_44 ? ~_GEN_3331 & _GEN_3222 : ~_GEN_3299 & _GEN_3222);
    rob_bsy_2_19 <= ~_GEN_3364 & (_GEN_44 ? ~_GEN_3332 & _GEN_3224 : ~_GEN_3300 & _GEN_3224);
    rob_bsy_2_20 <= ~_GEN_3365 & (_GEN_44 ? ~_GEN_3333 & _GEN_3226 : ~_GEN_3301 & _GEN_3226);
    rob_bsy_2_21 <= ~_GEN_3366 & (_GEN_44 ? ~_GEN_3334 & _GEN_3228 : ~_GEN_3302 & _GEN_3228);
    rob_bsy_2_22 <= ~_GEN_3367 & (_GEN_44 ? ~_GEN_3335 & _GEN_3230 : ~_GEN_3303 & _GEN_3230);
    rob_bsy_2_23 <= ~_GEN_3368 & (_GEN_44 ? ~_GEN_3336 & _GEN_3232 : ~_GEN_3304 & _GEN_3232);
    rob_bsy_2_24 <= ~_GEN_3369 & (_GEN_44 ? ~_GEN_3337 & _GEN_3234 : ~_GEN_3305 & _GEN_3234);
    rob_bsy_2_25 <= ~_GEN_3370 & (_GEN_44 ? ~_GEN_3338 & _GEN_3236 : ~_GEN_3306 & _GEN_3236);
    rob_bsy_2_26 <= ~_GEN_3371 & (_GEN_44 ? ~_GEN_3339 & _GEN_3238 : ~_GEN_3307 & _GEN_3238);
    rob_bsy_2_27 <= ~_GEN_3372 & (_GEN_44 ? ~_GEN_3340 & _GEN_3240 : ~_GEN_3308 & _GEN_3240);
    rob_bsy_2_28 <= ~_GEN_3373 & (_GEN_44 ? ~_GEN_3341 & _GEN_3242 : ~_GEN_3309 & _GEN_3242);
    rob_bsy_2_29 <= ~_GEN_3374 & (_GEN_44 ? ~_GEN_3342 & _GEN_3244 : ~_GEN_3310 & _GEN_3244);
    rob_bsy_2_30 <= ~_GEN_3375 & (_GEN_44 ? ~_GEN_3343 & _GEN_3246 : ~_GEN_3311 & _GEN_3246);
    rob_bsy_2_31 <= ~_GEN_3376 & (_GEN_44 ? ~_GEN_3344 & _GEN_3248 : ~_GEN_3312 & _GEN_3248);
    rob_unsafe_2_0 <= ~_GEN_3345 & (_GEN_44 ? ~_GEN_3313 & _GEN_3249 : ~_GEN_3281 & _GEN_3249);
    rob_unsafe_2_1 <= ~_GEN_3346 & (_GEN_44 ? ~_GEN_3314 & _GEN_3250 : ~_GEN_3282 & _GEN_3250);
    rob_unsafe_2_2 <= ~_GEN_3347 & (_GEN_44 ? ~_GEN_3315 & _GEN_3251 : ~_GEN_3283 & _GEN_3251);
    rob_unsafe_2_3 <= ~_GEN_3348 & (_GEN_44 ? ~_GEN_3316 & _GEN_3252 : ~_GEN_3284 & _GEN_3252);
    rob_unsafe_2_4 <= ~_GEN_3349 & (_GEN_44 ? ~_GEN_3317 & _GEN_3253 : ~_GEN_3285 & _GEN_3253);
    rob_unsafe_2_5 <= ~_GEN_3350 & (_GEN_44 ? ~_GEN_3318 & _GEN_3254 : ~_GEN_3286 & _GEN_3254);
    rob_unsafe_2_6 <= ~_GEN_3351 & (_GEN_44 ? ~_GEN_3319 & _GEN_3255 : ~_GEN_3287 & _GEN_3255);
    rob_unsafe_2_7 <= ~_GEN_3352 & (_GEN_44 ? ~_GEN_3320 & _GEN_3256 : ~_GEN_3288 & _GEN_3256);
    rob_unsafe_2_8 <= ~_GEN_3353 & (_GEN_44 ? ~_GEN_3321 & _GEN_3257 : ~_GEN_3289 & _GEN_3257);
    rob_unsafe_2_9 <= ~_GEN_3354 & (_GEN_44 ? ~_GEN_3322 & _GEN_3258 : ~_GEN_3290 & _GEN_3258);
    rob_unsafe_2_10 <= ~_GEN_3355 & (_GEN_44 ? ~_GEN_3323 & _GEN_3259 : ~_GEN_3291 & _GEN_3259);
    rob_unsafe_2_11 <= ~_GEN_3356 & (_GEN_44 ? ~_GEN_3324 & _GEN_3260 : ~_GEN_3292 & _GEN_3260);
    rob_unsafe_2_12 <= ~_GEN_3357 & (_GEN_44 ? ~_GEN_3325 & _GEN_3261 : ~_GEN_3293 & _GEN_3261);
    rob_unsafe_2_13 <= ~_GEN_3358 & (_GEN_44 ? ~_GEN_3326 & _GEN_3262 : ~_GEN_3294 & _GEN_3262);
    rob_unsafe_2_14 <= ~_GEN_3359 & (_GEN_44 ? ~_GEN_3327 & _GEN_3263 : ~_GEN_3295 & _GEN_3263);
    rob_unsafe_2_15 <= ~_GEN_3360 & (_GEN_44 ? ~_GEN_3328 & _GEN_3264 : ~_GEN_3296 & _GEN_3264);
    rob_unsafe_2_16 <= ~_GEN_3361 & (_GEN_44 ? ~_GEN_3329 & _GEN_3265 : ~_GEN_3297 & _GEN_3265);
    rob_unsafe_2_17 <= ~_GEN_3362 & (_GEN_44 ? ~_GEN_3330 & _GEN_3266 : ~_GEN_3298 & _GEN_3266);
    rob_unsafe_2_18 <= ~_GEN_3363 & (_GEN_44 ? ~_GEN_3331 & _GEN_3267 : ~_GEN_3299 & _GEN_3267);
    rob_unsafe_2_19 <= ~_GEN_3364 & (_GEN_44 ? ~_GEN_3332 & _GEN_3268 : ~_GEN_3300 & _GEN_3268);
    rob_unsafe_2_20 <= ~_GEN_3365 & (_GEN_44 ? ~_GEN_3333 & _GEN_3269 : ~_GEN_3301 & _GEN_3269);
    rob_unsafe_2_21 <= ~_GEN_3366 & (_GEN_44 ? ~_GEN_3334 & _GEN_3270 : ~_GEN_3302 & _GEN_3270);
    rob_unsafe_2_22 <= ~_GEN_3367 & (_GEN_44 ? ~_GEN_3335 & _GEN_3271 : ~_GEN_3303 & _GEN_3271);
    rob_unsafe_2_23 <= ~_GEN_3368 & (_GEN_44 ? ~_GEN_3336 & _GEN_3272 : ~_GEN_3304 & _GEN_3272);
    rob_unsafe_2_24 <= ~_GEN_3369 & (_GEN_44 ? ~_GEN_3337 & _GEN_3273 : ~_GEN_3305 & _GEN_3273);
    rob_unsafe_2_25 <= ~_GEN_3370 & (_GEN_44 ? ~_GEN_3338 & _GEN_3274 : ~_GEN_3306 & _GEN_3274);
    rob_unsafe_2_26 <= ~_GEN_3371 & (_GEN_44 ? ~_GEN_3339 & _GEN_3275 : ~_GEN_3307 & _GEN_3275);
    rob_unsafe_2_27 <= ~_GEN_3372 & (_GEN_44 ? ~_GEN_3340 & _GEN_3276 : ~_GEN_3308 & _GEN_3276);
    rob_unsafe_2_28 <= ~_GEN_3373 & (_GEN_44 ? ~_GEN_3341 & _GEN_3277 : ~_GEN_3309 & _GEN_3277);
    rob_unsafe_2_29 <= ~_GEN_3374 & (_GEN_44 ? ~_GEN_3342 & _GEN_3278 : ~_GEN_3310 & _GEN_3278);
    rob_unsafe_2_30 <= ~_GEN_3375 & (_GEN_44 ? ~_GEN_3343 & _GEN_3279 : ~_GEN_3311 & _GEN_3279);
    rob_unsafe_2_31 <= ~_GEN_3376 & (_GEN_44 ? ~_GEN_3344 & _GEN_3280 : ~_GEN_3312 & _GEN_3280);
    if (_GEN_2545) begin
      rob_uop_2_0_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_0_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_0_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_0_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_0_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_0_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_0_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_0_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_0_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_0_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_0_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_0_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_0_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_0_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_0_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_0_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_0_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_0_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_0_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3412) | ~rob_val_2_0) begin
      if (_GEN_2545)
        rob_uop_2_0_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_0_br_mask <= rob_uop_2_0_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1615)
      rob_uop_2_0_debug_fsrc <= 2'h3;
    else if (_GEN_2545)
      rob_uop_2_0_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2546) begin
      rob_uop_2_1_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_1_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_1_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_1_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_1_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_1_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_1_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_1_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_1_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_1_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_1_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_1_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_1_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_1_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_1_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_1_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_1_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_1_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_1_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3413) | ~rob_val_2_1) begin
      if (_GEN_2546)
        rob_uop_2_1_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_1_br_mask <= rob_uop_2_1_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1616)
      rob_uop_2_1_debug_fsrc <= 2'h3;
    else if (_GEN_2546)
      rob_uop_2_1_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2547) begin
      rob_uop_2_2_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_2_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_2_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_2_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_2_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_2_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_2_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_2_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_2_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_2_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_2_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_2_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_2_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_2_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_2_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_2_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_2_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_2_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_2_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3414) | ~rob_val_2_2) begin
      if (_GEN_2547)
        rob_uop_2_2_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_2_br_mask <= rob_uop_2_2_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1617)
      rob_uop_2_2_debug_fsrc <= 2'h3;
    else if (_GEN_2547)
      rob_uop_2_2_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2548) begin
      rob_uop_2_3_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_3_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_3_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_3_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_3_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_3_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_3_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_3_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_3_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_3_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_3_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_3_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_3_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_3_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_3_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_3_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_3_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_3_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_3_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3415) | ~rob_val_2_3) begin
      if (_GEN_2548)
        rob_uop_2_3_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_3_br_mask <= rob_uop_2_3_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1618)
      rob_uop_2_3_debug_fsrc <= 2'h3;
    else if (_GEN_2548)
      rob_uop_2_3_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2549) begin
      rob_uop_2_4_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_4_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_4_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_4_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_4_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_4_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_4_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_4_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_4_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_4_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_4_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_4_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_4_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_4_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_4_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_4_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_4_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_4_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_4_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3416) | ~rob_val_2_4) begin
      if (_GEN_2549)
        rob_uop_2_4_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_4_br_mask <= rob_uop_2_4_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1619)
      rob_uop_2_4_debug_fsrc <= 2'h3;
    else if (_GEN_2549)
      rob_uop_2_4_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2550) begin
      rob_uop_2_5_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_5_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_5_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_5_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_5_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_5_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_5_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_5_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_5_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_5_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_5_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_5_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_5_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_5_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_5_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_5_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_5_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_5_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_5_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3417) | ~rob_val_2_5) begin
      if (_GEN_2550)
        rob_uop_2_5_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_5_br_mask <= rob_uop_2_5_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1620)
      rob_uop_2_5_debug_fsrc <= 2'h3;
    else if (_GEN_2550)
      rob_uop_2_5_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2551) begin
      rob_uop_2_6_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_6_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_6_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_6_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_6_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_6_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_6_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_6_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_6_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_6_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_6_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_6_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_6_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_6_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_6_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_6_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_6_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_6_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_6_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3418) | ~rob_val_2_6) begin
      if (_GEN_2551)
        rob_uop_2_6_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_6_br_mask <= rob_uop_2_6_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1621)
      rob_uop_2_6_debug_fsrc <= 2'h3;
    else if (_GEN_2551)
      rob_uop_2_6_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2552) begin
      rob_uop_2_7_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_7_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_7_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_7_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_7_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_7_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_7_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_7_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_7_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_7_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_7_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_7_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_7_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_7_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_7_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_7_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_7_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_7_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_7_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3419) | ~rob_val_2_7) begin
      if (_GEN_2552)
        rob_uop_2_7_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_7_br_mask <= rob_uop_2_7_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1622)
      rob_uop_2_7_debug_fsrc <= 2'h3;
    else if (_GEN_2552)
      rob_uop_2_7_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2553) begin
      rob_uop_2_8_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_8_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_8_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_8_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_8_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_8_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_8_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_8_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_8_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_8_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_8_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_8_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_8_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_8_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_8_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_8_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_8_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_8_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_8_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3420) | ~rob_val_2_8) begin
      if (_GEN_2553)
        rob_uop_2_8_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_8_br_mask <= rob_uop_2_8_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1623)
      rob_uop_2_8_debug_fsrc <= 2'h3;
    else if (_GEN_2553)
      rob_uop_2_8_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2554) begin
      rob_uop_2_9_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_9_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_9_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_9_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_9_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_9_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_9_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_9_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_9_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_9_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_9_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_9_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_9_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_9_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_9_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_9_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_9_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_9_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_9_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3421) | ~rob_val_2_9) begin
      if (_GEN_2554)
        rob_uop_2_9_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_9_br_mask <= rob_uop_2_9_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1624)
      rob_uop_2_9_debug_fsrc <= 2'h3;
    else if (_GEN_2554)
      rob_uop_2_9_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2555) begin
      rob_uop_2_10_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_10_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_10_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_10_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_10_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_10_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_10_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_10_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_10_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_10_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_10_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_10_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_10_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_10_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_10_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_10_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_10_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_10_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_10_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3422) | ~rob_val_2_10) begin
      if (_GEN_2555)
        rob_uop_2_10_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_10_br_mask <= rob_uop_2_10_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1625)
      rob_uop_2_10_debug_fsrc <= 2'h3;
    else if (_GEN_2555)
      rob_uop_2_10_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2556) begin
      rob_uop_2_11_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_11_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_11_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_11_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_11_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_11_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_11_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_11_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_11_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_11_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_11_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_11_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_11_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_11_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_11_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_11_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_11_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_11_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_11_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3423) | ~rob_val_2_11) begin
      if (_GEN_2556)
        rob_uop_2_11_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_11_br_mask <= rob_uop_2_11_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1626)
      rob_uop_2_11_debug_fsrc <= 2'h3;
    else if (_GEN_2556)
      rob_uop_2_11_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2557) begin
      rob_uop_2_12_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_12_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_12_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_12_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_12_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_12_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_12_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_12_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_12_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_12_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_12_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_12_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_12_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_12_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_12_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_12_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_12_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_12_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_12_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3424) | ~rob_val_2_12) begin
      if (_GEN_2557)
        rob_uop_2_12_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_12_br_mask <= rob_uop_2_12_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1627)
      rob_uop_2_12_debug_fsrc <= 2'h3;
    else if (_GEN_2557)
      rob_uop_2_12_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2558) begin
      rob_uop_2_13_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_13_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_13_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_13_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_13_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_13_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_13_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_13_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_13_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_13_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_13_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_13_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_13_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_13_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_13_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_13_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_13_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_13_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_13_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3425) | ~rob_val_2_13) begin
      if (_GEN_2558)
        rob_uop_2_13_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_13_br_mask <= rob_uop_2_13_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1628)
      rob_uop_2_13_debug_fsrc <= 2'h3;
    else if (_GEN_2558)
      rob_uop_2_13_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2559) begin
      rob_uop_2_14_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_14_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_14_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_14_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_14_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_14_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_14_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_14_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_14_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_14_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_14_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_14_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_14_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_14_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_14_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_14_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_14_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_14_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_14_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3426) | ~rob_val_2_14) begin
      if (_GEN_2559)
        rob_uop_2_14_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_14_br_mask <= rob_uop_2_14_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1629)
      rob_uop_2_14_debug_fsrc <= 2'h3;
    else if (_GEN_2559)
      rob_uop_2_14_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2560) begin
      rob_uop_2_15_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_15_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_15_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_15_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_15_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_15_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_15_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_15_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_15_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_15_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_15_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_15_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_15_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_15_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_15_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_15_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_15_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_15_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_15_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3427) | ~rob_val_2_15) begin
      if (_GEN_2560)
        rob_uop_2_15_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_15_br_mask <= rob_uop_2_15_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1630)
      rob_uop_2_15_debug_fsrc <= 2'h3;
    else if (_GEN_2560)
      rob_uop_2_15_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2561) begin
      rob_uop_2_16_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_16_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_16_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_16_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_16_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_16_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_16_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_16_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_16_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_16_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_16_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_16_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_16_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_16_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_16_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_16_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_16_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_16_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_16_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3428) | ~rob_val_2_16) begin
      if (_GEN_2561)
        rob_uop_2_16_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_16_br_mask <= rob_uop_2_16_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1631)
      rob_uop_2_16_debug_fsrc <= 2'h3;
    else if (_GEN_2561)
      rob_uop_2_16_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2562) begin
      rob_uop_2_17_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_17_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_17_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_17_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_17_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_17_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_17_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_17_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_17_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_17_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_17_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_17_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_17_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_17_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_17_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_17_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_17_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_17_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_17_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3429) | ~rob_val_2_17) begin
      if (_GEN_2562)
        rob_uop_2_17_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_17_br_mask <= rob_uop_2_17_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1632)
      rob_uop_2_17_debug_fsrc <= 2'h3;
    else if (_GEN_2562)
      rob_uop_2_17_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2563) begin
      rob_uop_2_18_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_18_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_18_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_18_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_18_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_18_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_18_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_18_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_18_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_18_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_18_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_18_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_18_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_18_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_18_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_18_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_18_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_18_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_18_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3430) | ~rob_val_2_18) begin
      if (_GEN_2563)
        rob_uop_2_18_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_18_br_mask <= rob_uop_2_18_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1633)
      rob_uop_2_18_debug_fsrc <= 2'h3;
    else if (_GEN_2563)
      rob_uop_2_18_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2564) begin
      rob_uop_2_19_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_19_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_19_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_19_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_19_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_19_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_19_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_19_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_19_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_19_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_19_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_19_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_19_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_19_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_19_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_19_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_19_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_19_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_19_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3431) | ~rob_val_2_19) begin
      if (_GEN_2564)
        rob_uop_2_19_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_19_br_mask <= rob_uop_2_19_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1634)
      rob_uop_2_19_debug_fsrc <= 2'h3;
    else if (_GEN_2564)
      rob_uop_2_19_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2565) begin
      rob_uop_2_20_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_20_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_20_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_20_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_20_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_20_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_20_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_20_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_20_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_20_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_20_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_20_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_20_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_20_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_20_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_20_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_20_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_20_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_20_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3432) | ~rob_val_2_20) begin
      if (_GEN_2565)
        rob_uop_2_20_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_20_br_mask <= rob_uop_2_20_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1635)
      rob_uop_2_20_debug_fsrc <= 2'h3;
    else if (_GEN_2565)
      rob_uop_2_20_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2566) begin
      rob_uop_2_21_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_21_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_21_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_21_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_21_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_21_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_21_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_21_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_21_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_21_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_21_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_21_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_21_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_21_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_21_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_21_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_21_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_21_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_21_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3433) | ~rob_val_2_21) begin
      if (_GEN_2566)
        rob_uop_2_21_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_21_br_mask <= rob_uop_2_21_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1636)
      rob_uop_2_21_debug_fsrc <= 2'h3;
    else if (_GEN_2566)
      rob_uop_2_21_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2567) begin
      rob_uop_2_22_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_22_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_22_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_22_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_22_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_22_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_22_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_22_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_22_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_22_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_22_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_22_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_22_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_22_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_22_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_22_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_22_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_22_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_22_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3434) | ~rob_val_2_22) begin
      if (_GEN_2567)
        rob_uop_2_22_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_22_br_mask <= rob_uop_2_22_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1637)
      rob_uop_2_22_debug_fsrc <= 2'h3;
    else if (_GEN_2567)
      rob_uop_2_22_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2568) begin
      rob_uop_2_23_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_23_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_23_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_23_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_23_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_23_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_23_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_23_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_23_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_23_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_23_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_23_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_23_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_23_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_23_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_23_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_23_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_23_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_23_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3435) | ~rob_val_2_23) begin
      if (_GEN_2568)
        rob_uop_2_23_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_23_br_mask <= rob_uop_2_23_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1638)
      rob_uop_2_23_debug_fsrc <= 2'h3;
    else if (_GEN_2568)
      rob_uop_2_23_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2569) begin
      rob_uop_2_24_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_24_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_24_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_24_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_24_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_24_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_24_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_24_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_24_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_24_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_24_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_24_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_24_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_24_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_24_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_24_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_24_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_24_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_24_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3436) | ~rob_val_2_24) begin
      if (_GEN_2569)
        rob_uop_2_24_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_24_br_mask <= rob_uop_2_24_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1639)
      rob_uop_2_24_debug_fsrc <= 2'h3;
    else if (_GEN_2569)
      rob_uop_2_24_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2570) begin
      rob_uop_2_25_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_25_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_25_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_25_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_25_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_25_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_25_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_25_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_25_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_25_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_25_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_25_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_25_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_25_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_25_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_25_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_25_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_25_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_25_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3437) | ~rob_val_2_25) begin
      if (_GEN_2570)
        rob_uop_2_25_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_25_br_mask <= rob_uop_2_25_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1640)
      rob_uop_2_25_debug_fsrc <= 2'h3;
    else if (_GEN_2570)
      rob_uop_2_25_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2571) begin
      rob_uop_2_26_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_26_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_26_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_26_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_26_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_26_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_26_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_26_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_26_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_26_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_26_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_26_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_26_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_26_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_26_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_26_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_26_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_26_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_26_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3438) | ~rob_val_2_26) begin
      if (_GEN_2571)
        rob_uop_2_26_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_26_br_mask <= rob_uop_2_26_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1641)
      rob_uop_2_26_debug_fsrc <= 2'h3;
    else if (_GEN_2571)
      rob_uop_2_26_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2572) begin
      rob_uop_2_27_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_27_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_27_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_27_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_27_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_27_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_27_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_27_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_27_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_27_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_27_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_27_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_27_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_27_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_27_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_27_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_27_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_27_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_27_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3439) | ~rob_val_2_27) begin
      if (_GEN_2572)
        rob_uop_2_27_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_27_br_mask <= rob_uop_2_27_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1642)
      rob_uop_2_27_debug_fsrc <= 2'h3;
    else if (_GEN_2572)
      rob_uop_2_27_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2573) begin
      rob_uop_2_28_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_28_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_28_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_28_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_28_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_28_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_28_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_28_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_28_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_28_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_28_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_28_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_28_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_28_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_28_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_28_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_28_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_28_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_28_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3440) | ~rob_val_2_28) begin
      if (_GEN_2573)
        rob_uop_2_28_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_28_br_mask <= rob_uop_2_28_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1643)
      rob_uop_2_28_debug_fsrc <= 2'h3;
    else if (_GEN_2573)
      rob_uop_2_28_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2574) begin
      rob_uop_2_29_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_29_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_29_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_29_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_29_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_29_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_29_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_29_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_29_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_29_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_29_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_29_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_29_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_29_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_29_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_29_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_29_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_29_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_29_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3441) | ~rob_val_2_29) begin
      if (_GEN_2574)
        rob_uop_2_29_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_29_br_mask <= rob_uop_2_29_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1644)
      rob_uop_2_29_debug_fsrc <= 2'h3;
    else if (_GEN_2574)
      rob_uop_2_29_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2575) begin
      rob_uop_2_30_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_30_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_30_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_30_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_30_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_30_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_30_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_30_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_30_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_30_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_30_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_30_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_30_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_30_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_30_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_30_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_30_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_30_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_30_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3442) | ~rob_val_2_30) begin
      if (_GEN_2575)
        rob_uop_2_30_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_30_br_mask <= rob_uop_2_30_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & _GEN_1645)
      rob_uop_2_30_debug_fsrc <= 2'h3;
    else if (_GEN_2575)
      rob_uop_2_30_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    if (_GEN_2576) begin
      rob_uop_2_31_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_31_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_31_is_br <= io_enq_uops_2_is_br;
      rob_uop_2_31_is_jalr <= io_enq_uops_2_is_jalr;
      rob_uop_2_31_is_jal <= io_enq_uops_2_is_jal;
      rob_uop_2_31_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_31_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_31_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_31_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_31_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_31_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_31_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_31_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_31_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_31_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_31_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_31_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_31_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_31_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_3443) | ~rob_val_2_31) begin
      if (_GEN_2576)
        rob_uop_2_31_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_31_br_mask <= rob_uop_2_31_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48 & (&(io_brupdate_b2_uop_rob_idx[6:2])))
      rob_uop_2_31_debug_fsrc <= 2'h3;
    else if (_GEN_2576)
      rob_uop_2_31_debug_fsrc <= io_enq_uops_2_debug_fsrc;
    rob_exception_2_0 <= ~_GEN_3380 & (_GEN_46 & _GEN_1489 | (_GEN_2545 ? io_enq_uops_2_exception : rob_exception_2_0));
    rob_exception_2_1 <= ~_GEN_3381 & (_GEN_46 & _GEN_1490 | (_GEN_2546 ? io_enq_uops_2_exception : rob_exception_2_1));
    rob_exception_2_2 <= ~_GEN_3382 & (_GEN_46 & _GEN_1491 | (_GEN_2547 ? io_enq_uops_2_exception : rob_exception_2_2));
    rob_exception_2_3 <= ~_GEN_3383 & (_GEN_46 & _GEN_1492 | (_GEN_2548 ? io_enq_uops_2_exception : rob_exception_2_3));
    rob_exception_2_4 <= ~_GEN_3384 & (_GEN_46 & _GEN_1493 | (_GEN_2549 ? io_enq_uops_2_exception : rob_exception_2_4));
    rob_exception_2_5 <= ~_GEN_3385 & (_GEN_46 & _GEN_1494 | (_GEN_2550 ? io_enq_uops_2_exception : rob_exception_2_5));
    rob_exception_2_6 <= ~_GEN_3386 & (_GEN_46 & _GEN_1495 | (_GEN_2551 ? io_enq_uops_2_exception : rob_exception_2_6));
    rob_exception_2_7 <= ~_GEN_3387 & (_GEN_46 & _GEN_1496 | (_GEN_2552 ? io_enq_uops_2_exception : rob_exception_2_7));
    rob_exception_2_8 <= ~_GEN_3388 & (_GEN_46 & _GEN_1497 | (_GEN_2553 ? io_enq_uops_2_exception : rob_exception_2_8));
    rob_exception_2_9 <= ~_GEN_3389 & (_GEN_46 & _GEN_1498 | (_GEN_2554 ? io_enq_uops_2_exception : rob_exception_2_9));
    rob_exception_2_10 <= ~_GEN_3390 & (_GEN_46 & _GEN_1499 | (_GEN_2555 ? io_enq_uops_2_exception : rob_exception_2_10));
    rob_exception_2_11 <= ~_GEN_3391 & (_GEN_46 & _GEN_1500 | (_GEN_2556 ? io_enq_uops_2_exception : rob_exception_2_11));
    rob_exception_2_12 <= ~_GEN_3392 & (_GEN_46 & _GEN_1501 | (_GEN_2557 ? io_enq_uops_2_exception : rob_exception_2_12));
    rob_exception_2_13 <= ~_GEN_3393 & (_GEN_46 & _GEN_1502 | (_GEN_2558 ? io_enq_uops_2_exception : rob_exception_2_13));
    rob_exception_2_14 <= ~_GEN_3394 & (_GEN_46 & _GEN_1503 | (_GEN_2559 ? io_enq_uops_2_exception : rob_exception_2_14));
    rob_exception_2_15 <= ~_GEN_3395 & (_GEN_46 & _GEN_1504 | (_GEN_2560 ? io_enq_uops_2_exception : rob_exception_2_15));
    rob_exception_2_16 <= ~_GEN_3396 & (_GEN_46 & _GEN_1505 | (_GEN_2561 ? io_enq_uops_2_exception : rob_exception_2_16));
    rob_exception_2_17 <= ~_GEN_3397 & (_GEN_46 & _GEN_1506 | (_GEN_2562 ? io_enq_uops_2_exception : rob_exception_2_17));
    rob_exception_2_18 <= ~_GEN_3398 & (_GEN_46 & _GEN_1507 | (_GEN_2563 ? io_enq_uops_2_exception : rob_exception_2_18));
    rob_exception_2_19 <= ~_GEN_3399 & (_GEN_46 & _GEN_1508 | (_GEN_2564 ? io_enq_uops_2_exception : rob_exception_2_19));
    rob_exception_2_20 <= ~_GEN_3400 & (_GEN_46 & _GEN_1509 | (_GEN_2565 ? io_enq_uops_2_exception : rob_exception_2_20));
    rob_exception_2_21 <= ~_GEN_3401 & (_GEN_46 & _GEN_1510 | (_GEN_2566 ? io_enq_uops_2_exception : rob_exception_2_21));
    rob_exception_2_22 <= ~_GEN_3402 & (_GEN_46 & _GEN_1511 | (_GEN_2567 ? io_enq_uops_2_exception : rob_exception_2_22));
    rob_exception_2_23 <= ~_GEN_3403 & (_GEN_46 & _GEN_1512 | (_GEN_2568 ? io_enq_uops_2_exception : rob_exception_2_23));
    rob_exception_2_24 <= ~_GEN_3404 & (_GEN_46 & _GEN_1513 | (_GEN_2569 ? io_enq_uops_2_exception : rob_exception_2_24));
    rob_exception_2_25 <= ~_GEN_3405 & (_GEN_46 & _GEN_1514 | (_GEN_2570 ? io_enq_uops_2_exception : rob_exception_2_25));
    rob_exception_2_26 <= ~_GEN_3406 & (_GEN_46 & _GEN_1515 | (_GEN_2571 ? io_enq_uops_2_exception : rob_exception_2_26));
    rob_exception_2_27 <= ~_GEN_3407 & (_GEN_46 & _GEN_1516 | (_GEN_2572 ? io_enq_uops_2_exception : rob_exception_2_27));
    rob_exception_2_28 <= ~_GEN_3408 & (_GEN_46 & _GEN_1517 | (_GEN_2573 ? io_enq_uops_2_exception : rob_exception_2_28));
    rob_exception_2_29 <= ~_GEN_3409 & (_GEN_46 & _GEN_1518 | (_GEN_2574 ? io_enq_uops_2_exception : rob_exception_2_29));
    rob_exception_2_30 <= ~_GEN_3410 & (_GEN_46 & _GEN_1519 | (_GEN_2575 ? io_enq_uops_2_exception : rob_exception_2_30));
    rob_exception_2_31 <= ~_GEN_3411 & (_GEN_46 & (&(io_lxcpt_bits_uop_rob_idx[6:2])) | (_GEN_2576 ? io_enq_uops_2_exception : rob_exception_2_31));
    rob_predicated_2_0 <= ~(_GEN_42 & _GEN_1077 | _GEN_3153 | _GEN_40 & _GEN_887) & (_GEN_3025 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_697 | _GEN_2897 | _GEN_36 & _GEN_507 | _GEN_2769 | _GEN_34 & _GEN_317) & (_GEN_2641 ? io_wb_resps_0_bits_predicated : ~_GEN_2545 & rob_predicated_2_0));
    rob_predicated_2_1 <= ~(_GEN_42 & _GEN_1080 | _GEN_3154 | _GEN_40 & _GEN_890) & (_GEN_3026 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_700 | _GEN_2898 | _GEN_36 & _GEN_510 | _GEN_2770 | _GEN_34 & _GEN_320) & (_GEN_2642 ? io_wb_resps_0_bits_predicated : ~_GEN_2546 & rob_predicated_2_1));
    rob_predicated_2_2 <= ~(_GEN_42 & _GEN_1083 | _GEN_3155 | _GEN_40 & _GEN_893) & (_GEN_3027 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_703 | _GEN_2899 | _GEN_36 & _GEN_513 | _GEN_2771 | _GEN_34 & _GEN_323) & (_GEN_2643 ? io_wb_resps_0_bits_predicated : ~_GEN_2547 & rob_predicated_2_2));
    rob_predicated_2_3 <= ~(_GEN_42 & _GEN_1086 | _GEN_3156 | _GEN_40 & _GEN_896) & (_GEN_3028 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_706 | _GEN_2900 | _GEN_36 & _GEN_516 | _GEN_2772 | _GEN_34 & _GEN_326) & (_GEN_2644 ? io_wb_resps_0_bits_predicated : ~_GEN_2548 & rob_predicated_2_3));
    rob_predicated_2_4 <= ~(_GEN_42 & _GEN_1089 | _GEN_3157 | _GEN_40 & _GEN_899) & (_GEN_3029 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_709 | _GEN_2901 | _GEN_36 & _GEN_519 | _GEN_2773 | _GEN_34 & _GEN_329) & (_GEN_2645 ? io_wb_resps_0_bits_predicated : ~_GEN_2549 & rob_predicated_2_4));
    rob_predicated_2_5 <= ~(_GEN_42 & _GEN_1092 | _GEN_3158 | _GEN_40 & _GEN_902) & (_GEN_3030 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_712 | _GEN_2902 | _GEN_36 & _GEN_522 | _GEN_2774 | _GEN_34 & _GEN_332) & (_GEN_2646 ? io_wb_resps_0_bits_predicated : ~_GEN_2550 & rob_predicated_2_5));
    rob_predicated_2_6 <= ~(_GEN_42 & _GEN_1095 | _GEN_3159 | _GEN_40 & _GEN_905) & (_GEN_3031 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_715 | _GEN_2903 | _GEN_36 & _GEN_525 | _GEN_2775 | _GEN_34 & _GEN_335) & (_GEN_2647 ? io_wb_resps_0_bits_predicated : ~_GEN_2551 & rob_predicated_2_6));
    rob_predicated_2_7 <= ~(_GEN_42 & _GEN_1098 | _GEN_3160 | _GEN_40 & _GEN_908) & (_GEN_3032 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_718 | _GEN_2904 | _GEN_36 & _GEN_528 | _GEN_2776 | _GEN_34 & _GEN_338) & (_GEN_2648 ? io_wb_resps_0_bits_predicated : ~_GEN_2552 & rob_predicated_2_7));
    rob_predicated_2_8 <= ~(_GEN_42 & _GEN_1101 | _GEN_3161 | _GEN_40 & _GEN_911) & (_GEN_3033 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_721 | _GEN_2905 | _GEN_36 & _GEN_531 | _GEN_2777 | _GEN_34 & _GEN_341) & (_GEN_2649 ? io_wb_resps_0_bits_predicated : ~_GEN_2553 & rob_predicated_2_8));
    rob_predicated_2_9 <= ~(_GEN_42 & _GEN_1104 | _GEN_3162 | _GEN_40 & _GEN_914) & (_GEN_3034 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_724 | _GEN_2906 | _GEN_36 & _GEN_534 | _GEN_2778 | _GEN_34 & _GEN_344) & (_GEN_2650 ? io_wb_resps_0_bits_predicated : ~_GEN_2554 & rob_predicated_2_9));
    rob_predicated_2_10 <= ~(_GEN_42 & _GEN_1107 | _GEN_3163 | _GEN_40 & _GEN_917) & (_GEN_3035 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_727 | _GEN_2907 | _GEN_36 & _GEN_537 | _GEN_2779 | _GEN_34 & _GEN_347) & (_GEN_2651 ? io_wb_resps_0_bits_predicated : ~_GEN_2555 & rob_predicated_2_10));
    rob_predicated_2_11 <= ~(_GEN_42 & _GEN_1110 | _GEN_3164 | _GEN_40 & _GEN_920) & (_GEN_3036 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_730 | _GEN_2908 | _GEN_36 & _GEN_540 | _GEN_2780 | _GEN_34 & _GEN_350) & (_GEN_2652 ? io_wb_resps_0_bits_predicated : ~_GEN_2556 & rob_predicated_2_11));
    rob_predicated_2_12 <= ~(_GEN_42 & _GEN_1113 | _GEN_3165 | _GEN_40 & _GEN_923) & (_GEN_3037 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_733 | _GEN_2909 | _GEN_36 & _GEN_543 | _GEN_2781 | _GEN_34 & _GEN_353) & (_GEN_2653 ? io_wb_resps_0_bits_predicated : ~_GEN_2557 & rob_predicated_2_12));
    rob_predicated_2_13 <= ~(_GEN_42 & _GEN_1116 | _GEN_3166 | _GEN_40 & _GEN_926) & (_GEN_3038 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_736 | _GEN_2910 | _GEN_36 & _GEN_546 | _GEN_2782 | _GEN_34 & _GEN_356) & (_GEN_2654 ? io_wb_resps_0_bits_predicated : ~_GEN_2558 & rob_predicated_2_13));
    rob_predicated_2_14 <= ~(_GEN_42 & _GEN_1119 | _GEN_3167 | _GEN_40 & _GEN_929) & (_GEN_3039 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_739 | _GEN_2911 | _GEN_36 & _GEN_549 | _GEN_2783 | _GEN_34 & _GEN_359) & (_GEN_2655 ? io_wb_resps_0_bits_predicated : ~_GEN_2559 & rob_predicated_2_14));
    rob_predicated_2_15 <= ~(_GEN_42 & _GEN_1122 | _GEN_3168 | _GEN_40 & _GEN_932) & (_GEN_3040 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_742 | _GEN_2912 | _GEN_36 & _GEN_552 | _GEN_2784 | _GEN_34 & _GEN_362) & (_GEN_2656 ? io_wb_resps_0_bits_predicated : ~_GEN_2560 & rob_predicated_2_15));
    rob_predicated_2_16 <= ~(_GEN_42 & _GEN_1125 | _GEN_3169 | _GEN_40 & _GEN_935) & (_GEN_3041 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_745 | _GEN_2913 | _GEN_36 & _GEN_555 | _GEN_2785 | _GEN_34 & _GEN_365) & (_GEN_2657 ? io_wb_resps_0_bits_predicated : ~_GEN_2561 & rob_predicated_2_16));
    rob_predicated_2_17 <= ~(_GEN_42 & _GEN_1128 | _GEN_3170 | _GEN_40 & _GEN_938) & (_GEN_3042 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_748 | _GEN_2914 | _GEN_36 & _GEN_558 | _GEN_2786 | _GEN_34 & _GEN_368) & (_GEN_2658 ? io_wb_resps_0_bits_predicated : ~_GEN_2562 & rob_predicated_2_17));
    rob_predicated_2_18 <= ~(_GEN_42 & _GEN_1131 | _GEN_3171 | _GEN_40 & _GEN_941) & (_GEN_3043 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_751 | _GEN_2915 | _GEN_36 & _GEN_561 | _GEN_2787 | _GEN_34 & _GEN_371) & (_GEN_2659 ? io_wb_resps_0_bits_predicated : ~_GEN_2563 & rob_predicated_2_18));
    rob_predicated_2_19 <= ~(_GEN_42 & _GEN_1134 | _GEN_3172 | _GEN_40 & _GEN_944) & (_GEN_3044 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_754 | _GEN_2916 | _GEN_36 & _GEN_564 | _GEN_2788 | _GEN_34 & _GEN_374) & (_GEN_2660 ? io_wb_resps_0_bits_predicated : ~_GEN_2564 & rob_predicated_2_19));
    rob_predicated_2_20 <= ~(_GEN_42 & _GEN_1137 | _GEN_3173 | _GEN_40 & _GEN_947) & (_GEN_3045 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_757 | _GEN_2917 | _GEN_36 & _GEN_567 | _GEN_2789 | _GEN_34 & _GEN_377) & (_GEN_2661 ? io_wb_resps_0_bits_predicated : ~_GEN_2565 & rob_predicated_2_20));
    rob_predicated_2_21 <= ~(_GEN_42 & _GEN_1140 | _GEN_3174 | _GEN_40 & _GEN_950) & (_GEN_3046 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_760 | _GEN_2918 | _GEN_36 & _GEN_570 | _GEN_2790 | _GEN_34 & _GEN_380) & (_GEN_2662 ? io_wb_resps_0_bits_predicated : ~_GEN_2566 & rob_predicated_2_21));
    rob_predicated_2_22 <= ~(_GEN_42 & _GEN_1143 | _GEN_3175 | _GEN_40 & _GEN_953) & (_GEN_3047 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_763 | _GEN_2919 | _GEN_36 & _GEN_573 | _GEN_2791 | _GEN_34 & _GEN_383) & (_GEN_2663 ? io_wb_resps_0_bits_predicated : ~_GEN_2567 & rob_predicated_2_22));
    rob_predicated_2_23 <= ~(_GEN_42 & _GEN_1146 | _GEN_3176 | _GEN_40 & _GEN_956) & (_GEN_3048 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_766 | _GEN_2920 | _GEN_36 & _GEN_576 | _GEN_2792 | _GEN_34 & _GEN_386) & (_GEN_2664 ? io_wb_resps_0_bits_predicated : ~_GEN_2568 & rob_predicated_2_23));
    rob_predicated_2_24 <= ~(_GEN_42 & _GEN_1149 | _GEN_3177 | _GEN_40 & _GEN_959) & (_GEN_3049 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_769 | _GEN_2921 | _GEN_36 & _GEN_579 | _GEN_2793 | _GEN_34 & _GEN_389) & (_GEN_2665 ? io_wb_resps_0_bits_predicated : ~_GEN_2569 & rob_predicated_2_24));
    rob_predicated_2_25 <= ~(_GEN_42 & _GEN_1152 | _GEN_3178 | _GEN_40 & _GEN_962) & (_GEN_3050 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_772 | _GEN_2922 | _GEN_36 & _GEN_582 | _GEN_2794 | _GEN_34 & _GEN_392) & (_GEN_2666 ? io_wb_resps_0_bits_predicated : ~_GEN_2570 & rob_predicated_2_25));
    rob_predicated_2_26 <= ~(_GEN_42 & _GEN_1155 | _GEN_3179 | _GEN_40 & _GEN_965) & (_GEN_3051 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_775 | _GEN_2923 | _GEN_36 & _GEN_585 | _GEN_2795 | _GEN_34 & _GEN_395) & (_GEN_2667 ? io_wb_resps_0_bits_predicated : ~_GEN_2571 & rob_predicated_2_26));
    rob_predicated_2_27 <= ~(_GEN_42 & _GEN_1158 | _GEN_3180 | _GEN_40 & _GEN_968) & (_GEN_3052 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_778 | _GEN_2924 | _GEN_36 & _GEN_588 | _GEN_2796 | _GEN_34 & _GEN_398) & (_GEN_2668 ? io_wb_resps_0_bits_predicated : ~_GEN_2572 & rob_predicated_2_27));
    rob_predicated_2_28 <= ~(_GEN_42 & _GEN_1161 | _GEN_3181 | _GEN_40 & _GEN_971) & (_GEN_3053 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_781 | _GEN_2925 | _GEN_36 & _GEN_591 | _GEN_2797 | _GEN_34 & _GEN_401) & (_GEN_2669 ? io_wb_resps_0_bits_predicated : ~_GEN_2573 & rob_predicated_2_28));
    rob_predicated_2_29 <= ~(_GEN_42 & _GEN_1164 | _GEN_3182 | _GEN_40 & _GEN_974) & (_GEN_3054 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_784 | _GEN_2926 | _GEN_36 & _GEN_594 | _GEN_2798 | _GEN_34 & _GEN_404) & (_GEN_2670 ? io_wb_resps_0_bits_predicated : ~_GEN_2574 & rob_predicated_2_29));
    rob_predicated_2_30 <= ~(_GEN_42 & _GEN_1167 | _GEN_3183 | _GEN_40 & _GEN_977) & (_GEN_3055 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & _GEN_787 | _GEN_2927 | _GEN_36 & _GEN_597 | _GEN_2799 | _GEN_34 & _GEN_407) & (_GEN_2671 ? io_wb_resps_0_bits_predicated : ~_GEN_2575 & rob_predicated_2_30));
    rob_predicated_2_31 <= ~(_GEN_42 & (&(io_wb_resps_9_bits_uop_rob_idx[6:2])) | _GEN_3184 | _GEN_40 & (&(io_wb_resps_7_bits_uop_rob_idx[6:2]))) & (_GEN_3056 ? io_wb_resps_6_bits_predicated : ~(_GEN_38 & (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_2928 | _GEN_36 & (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_2800 | _GEN_34 & (&(io_wb_resps_1_bits_uop_rob_idx[6:2]))) & (_GEN_2672 ? io_wb_resps_0_bits_predicated : ~_GEN_2576 & rob_predicated_2_31));
    rob_bsy_3_0 <= ~_GEN_4244 & (_GEN_60 ? ~_GEN_4212 & _GEN_4085 : ~_GEN_4180 & _GEN_4085);
    rob_bsy_3_1 <= ~_GEN_4245 & (_GEN_60 ? ~_GEN_4213 & _GEN_4087 : ~_GEN_4181 & _GEN_4087);
    rob_bsy_3_2 <= ~_GEN_4246 & (_GEN_60 ? ~_GEN_4214 & _GEN_4089 : ~_GEN_4182 & _GEN_4089);
    rob_bsy_3_3 <= ~_GEN_4247 & (_GEN_60 ? ~_GEN_4215 & _GEN_4091 : ~_GEN_4183 & _GEN_4091);
    rob_bsy_3_4 <= ~_GEN_4248 & (_GEN_60 ? ~_GEN_4216 & _GEN_4093 : ~_GEN_4184 & _GEN_4093);
    rob_bsy_3_5 <= ~_GEN_4249 & (_GEN_60 ? ~_GEN_4217 & _GEN_4095 : ~_GEN_4185 & _GEN_4095);
    rob_bsy_3_6 <= ~_GEN_4250 & (_GEN_60 ? ~_GEN_4218 & _GEN_4097 : ~_GEN_4186 & _GEN_4097);
    rob_bsy_3_7 <= ~_GEN_4251 & (_GEN_60 ? ~_GEN_4219 & _GEN_4099 : ~_GEN_4187 & _GEN_4099);
    rob_bsy_3_8 <= ~_GEN_4252 & (_GEN_60 ? ~_GEN_4220 & _GEN_4101 : ~_GEN_4188 & _GEN_4101);
    rob_bsy_3_9 <= ~_GEN_4253 & (_GEN_60 ? ~_GEN_4221 & _GEN_4103 : ~_GEN_4189 & _GEN_4103);
    rob_bsy_3_10 <= ~_GEN_4254 & (_GEN_60 ? ~_GEN_4222 & _GEN_4105 : ~_GEN_4190 & _GEN_4105);
    rob_bsy_3_11 <= ~_GEN_4255 & (_GEN_60 ? ~_GEN_4223 & _GEN_4107 : ~_GEN_4191 & _GEN_4107);
    rob_bsy_3_12 <= ~_GEN_4256 & (_GEN_60 ? ~_GEN_4224 & _GEN_4109 : ~_GEN_4192 & _GEN_4109);
    rob_bsy_3_13 <= ~_GEN_4257 & (_GEN_60 ? ~_GEN_4225 & _GEN_4111 : ~_GEN_4193 & _GEN_4111);
    rob_bsy_3_14 <= ~_GEN_4258 & (_GEN_60 ? ~_GEN_4226 & _GEN_4113 : ~_GEN_4194 & _GEN_4113);
    rob_bsy_3_15 <= ~_GEN_4259 & (_GEN_60 ? ~_GEN_4227 & _GEN_4115 : ~_GEN_4195 & _GEN_4115);
    rob_bsy_3_16 <= ~_GEN_4260 & (_GEN_60 ? ~_GEN_4228 & _GEN_4117 : ~_GEN_4196 & _GEN_4117);
    rob_bsy_3_17 <= ~_GEN_4261 & (_GEN_60 ? ~_GEN_4229 & _GEN_4119 : ~_GEN_4197 & _GEN_4119);
    rob_bsy_3_18 <= ~_GEN_4262 & (_GEN_60 ? ~_GEN_4230 & _GEN_4121 : ~_GEN_4198 & _GEN_4121);
    rob_bsy_3_19 <= ~_GEN_4263 & (_GEN_60 ? ~_GEN_4231 & _GEN_4123 : ~_GEN_4199 & _GEN_4123);
    rob_bsy_3_20 <= ~_GEN_4264 & (_GEN_60 ? ~_GEN_4232 & _GEN_4125 : ~_GEN_4200 & _GEN_4125);
    rob_bsy_3_21 <= ~_GEN_4265 & (_GEN_60 ? ~_GEN_4233 & _GEN_4127 : ~_GEN_4201 & _GEN_4127);
    rob_bsy_3_22 <= ~_GEN_4266 & (_GEN_60 ? ~_GEN_4234 & _GEN_4129 : ~_GEN_4202 & _GEN_4129);
    rob_bsy_3_23 <= ~_GEN_4267 & (_GEN_60 ? ~_GEN_4235 & _GEN_4131 : ~_GEN_4203 & _GEN_4131);
    rob_bsy_3_24 <= ~_GEN_4268 & (_GEN_60 ? ~_GEN_4236 & _GEN_4133 : ~_GEN_4204 & _GEN_4133);
    rob_bsy_3_25 <= ~_GEN_4269 & (_GEN_60 ? ~_GEN_4237 & _GEN_4135 : ~_GEN_4205 & _GEN_4135);
    rob_bsy_3_26 <= ~_GEN_4270 & (_GEN_60 ? ~_GEN_4238 & _GEN_4137 : ~_GEN_4206 & _GEN_4137);
    rob_bsy_3_27 <= ~_GEN_4271 & (_GEN_60 ? ~_GEN_4239 & _GEN_4139 : ~_GEN_4207 & _GEN_4139);
    rob_bsy_3_28 <= ~_GEN_4272 & (_GEN_60 ? ~_GEN_4240 & _GEN_4141 : ~_GEN_4208 & _GEN_4141);
    rob_bsy_3_29 <= ~_GEN_4273 & (_GEN_60 ? ~_GEN_4241 & _GEN_4143 : ~_GEN_4209 & _GEN_4143);
    rob_bsy_3_30 <= ~_GEN_4274 & (_GEN_60 ? ~_GEN_4242 & _GEN_4145 : ~_GEN_4210 & _GEN_4145);
    rob_bsy_3_31 <= ~_GEN_4275 & (_GEN_60 ? ~_GEN_4243 & _GEN_4147 : ~_GEN_4211 & _GEN_4147);
    rob_unsafe_3_0 <= ~_GEN_4244 & (_GEN_60 ? ~_GEN_4212 & _GEN_4148 : ~_GEN_4180 & _GEN_4148);
    rob_unsafe_3_1 <= ~_GEN_4245 & (_GEN_60 ? ~_GEN_4213 & _GEN_4149 : ~_GEN_4181 & _GEN_4149);
    rob_unsafe_3_2 <= ~_GEN_4246 & (_GEN_60 ? ~_GEN_4214 & _GEN_4150 : ~_GEN_4182 & _GEN_4150);
    rob_unsafe_3_3 <= ~_GEN_4247 & (_GEN_60 ? ~_GEN_4215 & _GEN_4151 : ~_GEN_4183 & _GEN_4151);
    rob_unsafe_3_4 <= ~_GEN_4248 & (_GEN_60 ? ~_GEN_4216 & _GEN_4152 : ~_GEN_4184 & _GEN_4152);
    rob_unsafe_3_5 <= ~_GEN_4249 & (_GEN_60 ? ~_GEN_4217 & _GEN_4153 : ~_GEN_4185 & _GEN_4153);
    rob_unsafe_3_6 <= ~_GEN_4250 & (_GEN_60 ? ~_GEN_4218 & _GEN_4154 : ~_GEN_4186 & _GEN_4154);
    rob_unsafe_3_7 <= ~_GEN_4251 & (_GEN_60 ? ~_GEN_4219 & _GEN_4155 : ~_GEN_4187 & _GEN_4155);
    rob_unsafe_3_8 <= ~_GEN_4252 & (_GEN_60 ? ~_GEN_4220 & _GEN_4156 : ~_GEN_4188 & _GEN_4156);
    rob_unsafe_3_9 <= ~_GEN_4253 & (_GEN_60 ? ~_GEN_4221 & _GEN_4157 : ~_GEN_4189 & _GEN_4157);
    rob_unsafe_3_10 <= ~_GEN_4254 & (_GEN_60 ? ~_GEN_4222 & _GEN_4158 : ~_GEN_4190 & _GEN_4158);
    rob_unsafe_3_11 <= ~_GEN_4255 & (_GEN_60 ? ~_GEN_4223 & _GEN_4159 : ~_GEN_4191 & _GEN_4159);
    rob_unsafe_3_12 <= ~_GEN_4256 & (_GEN_60 ? ~_GEN_4224 & _GEN_4160 : ~_GEN_4192 & _GEN_4160);
    rob_unsafe_3_13 <= ~_GEN_4257 & (_GEN_60 ? ~_GEN_4225 & _GEN_4161 : ~_GEN_4193 & _GEN_4161);
    rob_unsafe_3_14 <= ~_GEN_4258 & (_GEN_60 ? ~_GEN_4226 & _GEN_4162 : ~_GEN_4194 & _GEN_4162);
    rob_unsafe_3_15 <= ~_GEN_4259 & (_GEN_60 ? ~_GEN_4227 & _GEN_4163 : ~_GEN_4195 & _GEN_4163);
    rob_unsafe_3_16 <= ~_GEN_4260 & (_GEN_60 ? ~_GEN_4228 & _GEN_4164 : ~_GEN_4196 & _GEN_4164);
    rob_unsafe_3_17 <= ~_GEN_4261 & (_GEN_60 ? ~_GEN_4229 & _GEN_4165 : ~_GEN_4197 & _GEN_4165);
    rob_unsafe_3_18 <= ~_GEN_4262 & (_GEN_60 ? ~_GEN_4230 & _GEN_4166 : ~_GEN_4198 & _GEN_4166);
    rob_unsafe_3_19 <= ~_GEN_4263 & (_GEN_60 ? ~_GEN_4231 & _GEN_4167 : ~_GEN_4199 & _GEN_4167);
    rob_unsafe_3_20 <= ~_GEN_4264 & (_GEN_60 ? ~_GEN_4232 & _GEN_4168 : ~_GEN_4200 & _GEN_4168);
    rob_unsafe_3_21 <= ~_GEN_4265 & (_GEN_60 ? ~_GEN_4233 & _GEN_4169 : ~_GEN_4201 & _GEN_4169);
    rob_unsafe_3_22 <= ~_GEN_4266 & (_GEN_60 ? ~_GEN_4234 & _GEN_4170 : ~_GEN_4202 & _GEN_4170);
    rob_unsafe_3_23 <= ~_GEN_4267 & (_GEN_60 ? ~_GEN_4235 & _GEN_4171 : ~_GEN_4203 & _GEN_4171);
    rob_unsafe_3_24 <= ~_GEN_4268 & (_GEN_60 ? ~_GEN_4236 & _GEN_4172 : ~_GEN_4204 & _GEN_4172);
    rob_unsafe_3_25 <= ~_GEN_4269 & (_GEN_60 ? ~_GEN_4237 & _GEN_4173 : ~_GEN_4205 & _GEN_4173);
    rob_unsafe_3_26 <= ~_GEN_4270 & (_GEN_60 ? ~_GEN_4238 & _GEN_4174 : ~_GEN_4206 & _GEN_4174);
    rob_unsafe_3_27 <= ~_GEN_4271 & (_GEN_60 ? ~_GEN_4239 & _GEN_4175 : ~_GEN_4207 & _GEN_4175);
    rob_unsafe_3_28 <= ~_GEN_4272 & (_GEN_60 ? ~_GEN_4240 & _GEN_4176 : ~_GEN_4208 & _GEN_4176);
    rob_unsafe_3_29 <= ~_GEN_4273 & (_GEN_60 ? ~_GEN_4241 & _GEN_4177 : ~_GEN_4209 & _GEN_4177);
    rob_unsafe_3_30 <= ~_GEN_4274 & (_GEN_60 ? ~_GEN_4242 & _GEN_4178 : ~_GEN_4210 & _GEN_4178);
    rob_unsafe_3_31 <= ~_GEN_4275 & (_GEN_60 ? ~_GEN_4243 & _GEN_4179 : ~_GEN_4211 & _GEN_4179);
    if (_GEN_3444) begin
      rob_uop_3_0_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_0_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_0_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_0_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_0_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_0_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_0_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_0_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_0_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_0_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_0_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_0_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_0_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_0_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_0_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_0_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_0_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_0_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_0_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4311) | ~rob_val_3_0) begin
      if (_GEN_3444)
        rob_uop_3_0_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_0_br_mask <= rob_uop_3_0_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1615)
      rob_uop_3_0_debug_fsrc <= 2'h3;
    else if (_GEN_3444)
      rob_uop_3_0_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3445) begin
      rob_uop_3_1_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_1_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_1_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_1_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_1_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_1_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_1_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_1_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_1_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_1_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_1_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_1_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_1_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_1_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_1_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_1_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_1_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_1_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_1_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4312) | ~rob_val_3_1) begin
      if (_GEN_3445)
        rob_uop_3_1_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_1_br_mask <= rob_uop_3_1_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1616)
      rob_uop_3_1_debug_fsrc <= 2'h3;
    else if (_GEN_3445)
      rob_uop_3_1_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3446) begin
      rob_uop_3_2_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_2_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_2_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_2_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_2_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_2_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_2_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_2_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_2_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_2_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_2_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_2_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_2_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_2_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_2_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_2_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_2_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_2_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_2_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4313) | ~rob_val_3_2) begin
      if (_GEN_3446)
        rob_uop_3_2_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_2_br_mask <= rob_uop_3_2_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1617)
      rob_uop_3_2_debug_fsrc <= 2'h3;
    else if (_GEN_3446)
      rob_uop_3_2_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3447) begin
      rob_uop_3_3_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_3_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_3_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_3_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_3_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_3_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_3_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_3_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_3_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_3_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_3_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_3_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_3_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_3_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_3_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_3_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_3_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_3_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_3_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4314) | ~rob_val_3_3) begin
      if (_GEN_3447)
        rob_uop_3_3_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_3_br_mask <= rob_uop_3_3_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1618)
      rob_uop_3_3_debug_fsrc <= 2'h3;
    else if (_GEN_3447)
      rob_uop_3_3_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3448) begin
      rob_uop_3_4_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_4_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_4_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_4_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_4_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_4_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_4_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_4_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_4_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_4_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_4_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_4_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_4_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_4_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_4_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_4_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_4_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_4_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_4_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4315) | ~rob_val_3_4) begin
      if (_GEN_3448)
        rob_uop_3_4_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_4_br_mask <= rob_uop_3_4_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1619)
      rob_uop_3_4_debug_fsrc <= 2'h3;
    else if (_GEN_3448)
      rob_uop_3_4_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3449) begin
      rob_uop_3_5_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_5_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_5_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_5_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_5_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_5_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_5_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_5_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_5_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_5_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_5_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_5_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_5_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_5_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_5_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_5_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_5_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_5_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_5_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4316) | ~rob_val_3_5) begin
      if (_GEN_3449)
        rob_uop_3_5_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_5_br_mask <= rob_uop_3_5_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1620)
      rob_uop_3_5_debug_fsrc <= 2'h3;
    else if (_GEN_3449)
      rob_uop_3_5_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3450) begin
      rob_uop_3_6_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_6_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_6_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_6_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_6_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_6_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_6_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_6_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_6_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_6_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_6_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_6_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_6_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_6_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_6_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_6_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_6_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_6_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_6_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4317) | ~rob_val_3_6) begin
      if (_GEN_3450)
        rob_uop_3_6_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_6_br_mask <= rob_uop_3_6_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1621)
      rob_uop_3_6_debug_fsrc <= 2'h3;
    else if (_GEN_3450)
      rob_uop_3_6_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3451) begin
      rob_uop_3_7_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_7_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_7_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_7_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_7_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_7_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_7_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_7_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_7_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_7_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_7_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_7_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_7_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_7_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_7_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_7_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_7_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_7_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_7_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4318) | ~rob_val_3_7) begin
      if (_GEN_3451)
        rob_uop_3_7_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_7_br_mask <= rob_uop_3_7_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1622)
      rob_uop_3_7_debug_fsrc <= 2'h3;
    else if (_GEN_3451)
      rob_uop_3_7_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3452) begin
      rob_uop_3_8_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_8_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_8_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_8_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_8_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_8_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_8_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_8_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_8_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_8_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_8_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_8_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_8_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_8_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_8_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_8_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_8_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_8_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_8_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4319) | ~rob_val_3_8) begin
      if (_GEN_3452)
        rob_uop_3_8_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_8_br_mask <= rob_uop_3_8_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1623)
      rob_uop_3_8_debug_fsrc <= 2'h3;
    else if (_GEN_3452)
      rob_uop_3_8_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3453) begin
      rob_uop_3_9_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_9_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_9_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_9_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_9_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_9_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_9_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_9_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_9_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_9_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_9_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_9_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_9_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_9_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_9_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_9_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_9_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_9_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_9_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4320) | ~rob_val_3_9) begin
      if (_GEN_3453)
        rob_uop_3_9_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_9_br_mask <= rob_uop_3_9_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1624)
      rob_uop_3_9_debug_fsrc <= 2'h3;
    else if (_GEN_3453)
      rob_uop_3_9_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3454) begin
      rob_uop_3_10_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_10_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_10_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_10_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_10_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_10_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_10_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_10_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_10_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_10_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_10_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_10_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_10_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_10_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_10_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_10_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_10_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_10_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_10_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4321) | ~rob_val_3_10) begin
      if (_GEN_3454)
        rob_uop_3_10_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_10_br_mask <= rob_uop_3_10_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1625)
      rob_uop_3_10_debug_fsrc <= 2'h3;
    else if (_GEN_3454)
      rob_uop_3_10_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3455) begin
      rob_uop_3_11_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_11_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_11_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_11_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_11_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_11_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_11_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_11_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_11_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_11_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_11_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_11_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_11_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_11_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_11_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_11_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_11_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_11_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_11_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4322) | ~rob_val_3_11) begin
      if (_GEN_3455)
        rob_uop_3_11_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_11_br_mask <= rob_uop_3_11_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1626)
      rob_uop_3_11_debug_fsrc <= 2'h3;
    else if (_GEN_3455)
      rob_uop_3_11_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3456) begin
      rob_uop_3_12_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_12_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_12_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_12_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_12_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_12_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_12_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_12_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_12_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_12_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_12_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_12_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_12_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_12_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_12_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_12_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_12_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_12_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_12_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4323) | ~rob_val_3_12) begin
      if (_GEN_3456)
        rob_uop_3_12_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_12_br_mask <= rob_uop_3_12_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1627)
      rob_uop_3_12_debug_fsrc <= 2'h3;
    else if (_GEN_3456)
      rob_uop_3_12_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3457) begin
      rob_uop_3_13_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_13_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_13_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_13_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_13_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_13_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_13_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_13_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_13_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_13_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_13_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_13_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_13_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_13_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_13_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_13_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_13_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_13_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_13_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4324) | ~rob_val_3_13) begin
      if (_GEN_3457)
        rob_uop_3_13_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_13_br_mask <= rob_uop_3_13_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1628)
      rob_uop_3_13_debug_fsrc <= 2'h3;
    else if (_GEN_3457)
      rob_uop_3_13_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3458) begin
      rob_uop_3_14_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_14_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_14_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_14_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_14_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_14_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_14_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_14_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_14_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_14_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_14_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_14_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_14_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_14_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_14_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_14_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_14_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_14_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_14_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4325) | ~rob_val_3_14) begin
      if (_GEN_3458)
        rob_uop_3_14_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_14_br_mask <= rob_uop_3_14_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1629)
      rob_uop_3_14_debug_fsrc <= 2'h3;
    else if (_GEN_3458)
      rob_uop_3_14_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3459) begin
      rob_uop_3_15_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_15_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_15_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_15_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_15_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_15_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_15_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_15_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_15_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_15_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_15_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_15_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_15_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_15_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_15_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_15_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_15_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_15_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_15_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4326) | ~rob_val_3_15) begin
      if (_GEN_3459)
        rob_uop_3_15_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_15_br_mask <= rob_uop_3_15_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1630)
      rob_uop_3_15_debug_fsrc <= 2'h3;
    else if (_GEN_3459)
      rob_uop_3_15_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3460) begin
      rob_uop_3_16_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_16_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_16_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_16_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_16_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_16_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_16_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_16_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_16_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_16_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_16_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_16_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_16_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_16_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_16_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_16_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_16_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_16_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_16_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4327) | ~rob_val_3_16) begin
      if (_GEN_3460)
        rob_uop_3_16_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_16_br_mask <= rob_uop_3_16_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1631)
      rob_uop_3_16_debug_fsrc <= 2'h3;
    else if (_GEN_3460)
      rob_uop_3_16_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3461) begin
      rob_uop_3_17_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_17_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_17_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_17_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_17_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_17_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_17_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_17_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_17_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_17_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_17_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_17_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_17_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_17_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_17_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_17_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_17_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_17_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_17_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4328) | ~rob_val_3_17) begin
      if (_GEN_3461)
        rob_uop_3_17_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_17_br_mask <= rob_uop_3_17_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1632)
      rob_uop_3_17_debug_fsrc <= 2'h3;
    else if (_GEN_3461)
      rob_uop_3_17_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3462) begin
      rob_uop_3_18_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_18_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_18_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_18_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_18_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_18_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_18_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_18_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_18_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_18_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_18_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_18_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_18_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_18_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_18_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_18_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_18_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_18_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_18_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4329) | ~rob_val_3_18) begin
      if (_GEN_3462)
        rob_uop_3_18_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_18_br_mask <= rob_uop_3_18_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1633)
      rob_uop_3_18_debug_fsrc <= 2'h3;
    else if (_GEN_3462)
      rob_uop_3_18_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3463) begin
      rob_uop_3_19_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_19_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_19_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_19_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_19_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_19_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_19_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_19_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_19_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_19_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_19_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_19_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_19_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_19_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_19_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_19_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_19_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_19_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_19_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4330) | ~rob_val_3_19) begin
      if (_GEN_3463)
        rob_uop_3_19_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_19_br_mask <= rob_uop_3_19_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1634)
      rob_uop_3_19_debug_fsrc <= 2'h3;
    else if (_GEN_3463)
      rob_uop_3_19_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3464) begin
      rob_uop_3_20_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_20_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_20_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_20_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_20_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_20_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_20_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_20_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_20_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_20_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_20_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_20_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_20_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_20_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_20_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_20_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_20_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_20_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_20_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4331) | ~rob_val_3_20) begin
      if (_GEN_3464)
        rob_uop_3_20_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_20_br_mask <= rob_uop_3_20_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1635)
      rob_uop_3_20_debug_fsrc <= 2'h3;
    else if (_GEN_3464)
      rob_uop_3_20_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3465) begin
      rob_uop_3_21_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_21_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_21_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_21_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_21_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_21_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_21_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_21_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_21_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_21_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_21_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_21_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_21_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_21_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_21_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_21_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_21_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_21_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_21_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4332) | ~rob_val_3_21) begin
      if (_GEN_3465)
        rob_uop_3_21_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_21_br_mask <= rob_uop_3_21_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1636)
      rob_uop_3_21_debug_fsrc <= 2'h3;
    else if (_GEN_3465)
      rob_uop_3_21_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3466) begin
      rob_uop_3_22_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_22_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_22_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_22_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_22_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_22_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_22_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_22_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_22_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_22_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_22_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_22_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_22_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_22_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_22_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_22_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_22_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_22_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_22_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4333) | ~rob_val_3_22) begin
      if (_GEN_3466)
        rob_uop_3_22_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_22_br_mask <= rob_uop_3_22_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1637)
      rob_uop_3_22_debug_fsrc <= 2'h3;
    else if (_GEN_3466)
      rob_uop_3_22_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3467) begin
      rob_uop_3_23_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_23_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_23_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_23_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_23_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_23_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_23_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_23_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_23_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_23_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_23_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_23_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_23_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_23_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_23_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_23_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_23_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_23_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_23_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4334) | ~rob_val_3_23) begin
      if (_GEN_3467)
        rob_uop_3_23_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_23_br_mask <= rob_uop_3_23_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1638)
      rob_uop_3_23_debug_fsrc <= 2'h3;
    else if (_GEN_3467)
      rob_uop_3_23_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3468) begin
      rob_uop_3_24_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_24_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_24_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_24_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_24_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_24_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_24_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_24_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_24_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_24_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_24_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_24_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_24_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_24_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_24_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_24_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_24_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_24_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_24_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4335) | ~rob_val_3_24) begin
      if (_GEN_3468)
        rob_uop_3_24_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_24_br_mask <= rob_uop_3_24_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1639)
      rob_uop_3_24_debug_fsrc <= 2'h3;
    else if (_GEN_3468)
      rob_uop_3_24_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3469) begin
      rob_uop_3_25_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_25_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_25_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_25_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_25_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_25_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_25_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_25_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_25_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_25_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_25_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_25_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_25_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_25_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_25_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_25_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_25_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_25_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_25_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4336) | ~rob_val_3_25) begin
      if (_GEN_3469)
        rob_uop_3_25_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_25_br_mask <= rob_uop_3_25_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1640)
      rob_uop_3_25_debug_fsrc <= 2'h3;
    else if (_GEN_3469)
      rob_uop_3_25_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3470) begin
      rob_uop_3_26_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_26_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_26_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_26_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_26_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_26_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_26_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_26_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_26_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_26_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_26_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_26_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_26_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_26_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_26_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_26_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_26_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_26_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_26_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4337) | ~rob_val_3_26) begin
      if (_GEN_3470)
        rob_uop_3_26_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_26_br_mask <= rob_uop_3_26_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1641)
      rob_uop_3_26_debug_fsrc <= 2'h3;
    else if (_GEN_3470)
      rob_uop_3_26_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3471) begin
      rob_uop_3_27_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_27_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_27_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_27_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_27_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_27_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_27_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_27_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_27_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_27_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_27_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_27_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_27_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_27_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_27_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_27_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_27_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_27_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_27_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4338) | ~rob_val_3_27) begin
      if (_GEN_3471)
        rob_uop_3_27_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_27_br_mask <= rob_uop_3_27_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1642)
      rob_uop_3_27_debug_fsrc <= 2'h3;
    else if (_GEN_3471)
      rob_uop_3_27_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3472) begin
      rob_uop_3_28_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_28_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_28_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_28_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_28_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_28_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_28_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_28_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_28_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_28_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_28_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_28_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_28_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_28_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_28_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_28_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_28_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_28_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_28_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4339) | ~rob_val_3_28) begin
      if (_GEN_3472)
        rob_uop_3_28_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_28_br_mask <= rob_uop_3_28_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1643)
      rob_uop_3_28_debug_fsrc <= 2'h3;
    else if (_GEN_3472)
      rob_uop_3_28_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3473) begin
      rob_uop_3_29_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_29_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_29_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_29_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_29_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_29_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_29_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_29_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_29_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_29_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_29_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_29_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_29_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_29_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_29_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_29_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_29_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_29_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_29_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4340) | ~rob_val_3_29) begin
      if (_GEN_3473)
        rob_uop_3_29_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_29_br_mask <= rob_uop_3_29_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1644)
      rob_uop_3_29_debug_fsrc <= 2'h3;
    else if (_GEN_3473)
      rob_uop_3_29_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3474) begin
      rob_uop_3_30_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_30_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_30_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_30_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_30_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_30_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_30_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_30_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_30_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_30_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_30_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_30_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_30_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_30_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_30_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_30_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_30_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_30_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_30_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4341) | ~rob_val_3_30) begin
      if (_GEN_3474)
        rob_uop_3_30_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_30_br_mask <= rob_uop_3_30_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & _GEN_1645)
      rob_uop_3_30_debug_fsrc <= 2'h3;
    else if (_GEN_3474)
      rob_uop_3_30_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    if (_GEN_3475) begin
      rob_uop_3_31_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_31_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_31_is_br <= io_enq_uops_3_is_br;
      rob_uop_3_31_is_jalr <= io_enq_uops_3_is_jalr;
      rob_uop_3_31_is_jal <= io_enq_uops_3_is_jal;
      rob_uop_3_31_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_31_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_31_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_31_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_31_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_31_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_31_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_31_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_31_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_31_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_31_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_31_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_31_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_31_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_4342) | ~rob_val_3_31) begin
      if (_GEN_3475)
        rob_uop_3_31_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_31_br_mask <= rob_uop_3_31_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64 & (&(io_brupdate_b2_uop_rob_idx[6:2])))
      rob_uop_3_31_debug_fsrc <= 2'h3;
    else if (_GEN_3475)
      rob_uop_3_31_debug_fsrc <= io_enq_uops_3_debug_fsrc;
    rob_exception_3_0 <= ~_GEN_4279 & (_GEN_62 & _GEN_1489 | (_GEN_3444 ? io_enq_uops_3_exception : rob_exception_3_0));
    rob_exception_3_1 <= ~_GEN_4280 & (_GEN_62 & _GEN_1490 | (_GEN_3445 ? io_enq_uops_3_exception : rob_exception_3_1));
    rob_exception_3_2 <= ~_GEN_4281 & (_GEN_62 & _GEN_1491 | (_GEN_3446 ? io_enq_uops_3_exception : rob_exception_3_2));
    rob_exception_3_3 <= ~_GEN_4282 & (_GEN_62 & _GEN_1492 | (_GEN_3447 ? io_enq_uops_3_exception : rob_exception_3_3));
    rob_exception_3_4 <= ~_GEN_4283 & (_GEN_62 & _GEN_1493 | (_GEN_3448 ? io_enq_uops_3_exception : rob_exception_3_4));
    rob_exception_3_5 <= ~_GEN_4284 & (_GEN_62 & _GEN_1494 | (_GEN_3449 ? io_enq_uops_3_exception : rob_exception_3_5));
    rob_exception_3_6 <= ~_GEN_4285 & (_GEN_62 & _GEN_1495 | (_GEN_3450 ? io_enq_uops_3_exception : rob_exception_3_6));
    rob_exception_3_7 <= ~_GEN_4286 & (_GEN_62 & _GEN_1496 | (_GEN_3451 ? io_enq_uops_3_exception : rob_exception_3_7));
    rob_exception_3_8 <= ~_GEN_4287 & (_GEN_62 & _GEN_1497 | (_GEN_3452 ? io_enq_uops_3_exception : rob_exception_3_8));
    rob_exception_3_9 <= ~_GEN_4288 & (_GEN_62 & _GEN_1498 | (_GEN_3453 ? io_enq_uops_3_exception : rob_exception_3_9));
    rob_exception_3_10 <= ~_GEN_4289 & (_GEN_62 & _GEN_1499 | (_GEN_3454 ? io_enq_uops_3_exception : rob_exception_3_10));
    rob_exception_3_11 <= ~_GEN_4290 & (_GEN_62 & _GEN_1500 | (_GEN_3455 ? io_enq_uops_3_exception : rob_exception_3_11));
    rob_exception_3_12 <= ~_GEN_4291 & (_GEN_62 & _GEN_1501 | (_GEN_3456 ? io_enq_uops_3_exception : rob_exception_3_12));
    rob_exception_3_13 <= ~_GEN_4292 & (_GEN_62 & _GEN_1502 | (_GEN_3457 ? io_enq_uops_3_exception : rob_exception_3_13));
    rob_exception_3_14 <= ~_GEN_4293 & (_GEN_62 & _GEN_1503 | (_GEN_3458 ? io_enq_uops_3_exception : rob_exception_3_14));
    rob_exception_3_15 <= ~_GEN_4294 & (_GEN_62 & _GEN_1504 | (_GEN_3459 ? io_enq_uops_3_exception : rob_exception_3_15));
    rob_exception_3_16 <= ~_GEN_4295 & (_GEN_62 & _GEN_1505 | (_GEN_3460 ? io_enq_uops_3_exception : rob_exception_3_16));
    rob_exception_3_17 <= ~_GEN_4296 & (_GEN_62 & _GEN_1506 | (_GEN_3461 ? io_enq_uops_3_exception : rob_exception_3_17));
    rob_exception_3_18 <= ~_GEN_4297 & (_GEN_62 & _GEN_1507 | (_GEN_3462 ? io_enq_uops_3_exception : rob_exception_3_18));
    rob_exception_3_19 <= ~_GEN_4298 & (_GEN_62 & _GEN_1508 | (_GEN_3463 ? io_enq_uops_3_exception : rob_exception_3_19));
    rob_exception_3_20 <= ~_GEN_4299 & (_GEN_62 & _GEN_1509 | (_GEN_3464 ? io_enq_uops_3_exception : rob_exception_3_20));
    rob_exception_3_21 <= ~_GEN_4300 & (_GEN_62 & _GEN_1510 | (_GEN_3465 ? io_enq_uops_3_exception : rob_exception_3_21));
    rob_exception_3_22 <= ~_GEN_4301 & (_GEN_62 & _GEN_1511 | (_GEN_3466 ? io_enq_uops_3_exception : rob_exception_3_22));
    rob_exception_3_23 <= ~_GEN_4302 & (_GEN_62 & _GEN_1512 | (_GEN_3467 ? io_enq_uops_3_exception : rob_exception_3_23));
    rob_exception_3_24 <= ~_GEN_4303 & (_GEN_62 & _GEN_1513 | (_GEN_3468 ? io_enq_uops_3_exception : rob_exception_3_24));
    rob_exception_3_25 <= ~_GEN_4304 & (_GEN_62 & _GEN_1514 | (_GEN_3469 ? io_enq_uops_3_exception : rob_exception_3_25));
    rob_exception_3_26 <= ~_GEN_4305 & (_GEN_62 & _GEN_1515 | (_GEN_3470 ? io_enq_uops_3_exception : rob_exception_3_26));
    rob_exception_3_27 <= ~_GEN_4306 & (_GEN_62 & _GEN_1516 | (_GEN_3471 ? io_enq_uops_3_exception : rob_exception_3_27));
    rob_exception_3_28 <= ~_GEN_4307 & (_GEN_62 & _GEN_1517 | (_GEN_3472 ? io_enq_uops_3_exception : rob_exception_3_28));
    rob_exception_3_29 <= ~_GEN_4308 & (_GEN_62 & _GEN_1518 | (_GEN_3473 ? io_enq_uops_3_exception : rob_exception_3_29));
    rob_exception_3_30 <= ~_GEN_4309 & (_GEN_62 & _GEN_1519 | (_GEN_3474 ? io_enq_uops_3_exception : rob_exception_3_30));
    rob_exception_3_31 <= ~_GEN_4310 & (_GEN_62 & (&(io_lxcpt_bits_uop_rob_idx[6:2])) | (_GEN_3475 ? io_enq_uops_3_exception : rob_exception_3_31));
    rob_predicated_3_0 <= ~(_GEN_58 & _GEN_1077 | _GEN_4052 | _GEN_56 & _GEN_887) & (_GEN_3924 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_697 | _GEN_3796 | _GEN_52 & _GEN_507 | _GEN_3668 | _GEN_50 & _GEN_317) & (_GEN_3540 ? io_wb_resps_0_bits_predicated : ~_GEN_3444 & rob_predicated_3_0));
    rob_predicated_3_1 <= ~(_GEN_58 & _GEN_1080 | _GEN_4053 | _GEN_56 & _GEN_890) & (_GEN_3925 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_700 | _GEN_3797 | _GEN_52 & _GEN_510 | _GEN_3669 | _GEN_50 & _GEN_320) & (_GEN_3541 ? io_wb_resps_0_bits_predicated : ~_GEN_3445 & rob_predicated_3_1));
    rob_predicated_3_2 <= ~(_GEN_58 & _GEN_1083 | _GEN_4054 | _GEN_56 & _GEN_893) & (_GEN_3926 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_703 | _GEN_3798 | _GEN_52 & _GEN_513 | _GEN_3670 | _GEN_50 & _GEN_323) & (_GEN_3542 ? io_wb_resps_0_bits_predicated : ~_GEN_3446 & rob_predicated_3_2));
    rob_predicated_3_3 <= ~(_GEN_58 & _GEN_1086 | _GEN_4055 | _GEN_56 & _GEN_896) & (_GEN_3927 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_706 | _GEN_3799 | _GEN_52 & _GEN_516 | _GEN_3671 | _GEN_50 & _GEN_326) & (_GEN_3543 ? io_wb_resps_0_bits_predicated : ~_GEN_3447 & rob_predicated_3_3));
    rob_predicated_3_4 <= ~(_GEN_58 & _GEN_1089 | _GEN_4056 | _GEN_56 & _GEN_899) & (_GEN_3928 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_709 | _GEN_3800 | _GEN_52 & _GEN_519 | _GEN_3672 | _GEN_50 & _GEN_329) & (_GEN_3544 ? io_wb_resps_0_bits_predicated : ~_GEN_3448 & rob_predicated_3_4));
    rob_predicated_3_5 <= ~(_GEN_58 & _GEN_1092 | _GEN_4057 | _GEN_56 & _GEN_902) & (_GEN_3929 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_712 | _GEN_3801 | _GEN_52 & _GEN_522 | _GEN_3673 | _GEN_50 & _GEN_332) & (_GEN_3545 ? io_wb_resps_0_bits_predicated : ~_GEN_3449 & rob_predicated_3_5));
    rob_predicated_3_6 <= ~(_GEN_58 & _GEN_1095 | _GEN_4058 | _GEN_56 & _GEN_905) & (_GEN_3930 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_715 | _GEN_3802 | _GEN_52 & _GEN_525 | _GEN_3674 | _GEN_50 & _GEN_335) & (_GEN_3546 ? io_wb_resps_0_bits_predicated : ~_GEN_3450 & rob_predicated_3_6));
    rob_predicated_3_7 <= ~(_GEN_58 & _GEN_1098 | _GEN_4059 | _GEN_56 & _GEN_908) & (_GEN_3931 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_718 | _GEN_3803 | _GEN_52 & _GEN_528 | _GEN_3675 | _GEN_50 & _GEN_338) & (_GEN_3547 ? io_wb_resps_0_bits_predicated : ~_GEN_3451 & rob_predicated_3_7));
    rob_predicated_3_8 <= ~(_GEN_58 & _GEN_1101 | _GEN_4060 | _GEN_56 & _GEN_911) & (_GEN_3932 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_721 | _GEN_3804 | _GEN_52 & _GEN_531 | _GEN_3676 | _GEN_50 & _GEN_341) & (_GEN_3548 ? io_wb_resps_0_bits_predicated : ~_GEN_3452 & rob_predicated_3_8));
    rob_predicated_3_9 <= ~(_GEN_58 & _GEN_1104 | _GEN_4061 | _GEN_56 & _GEN_914) & (_GEN_3933 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_724 | _GEN_3805 | _GEN_52 & _GEN_534 | _GEN_3677 | _GEN_50 & _GEN_344) & (_GEN_3549 ? io_wb_resps_0_bits_predicated : ~_GEN_3453 & rob_predicated_3_9));
    rob_predicated_3_10 <= ~(_GEN_58 & _GEN_1107 | _GEN_4062 | _GEN_56 & _GEN_917) & (_GEN_3934 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_727 | _GEN_3806 | _GEN_52 & _GEN_537 | _GEN_3678 | _GEN_50 & _GEN_347) & (_GEN_3550 ? io_wb_resps_0_bits_predicated : ~_GEN_3454 & rob_predicated_3_10));
    rob_predicated_3_11 <= ~(_GEN_58 & _GEN_1110 | _GEN_4063 | _GEN_56 & _GEN_920) & (_GEN_3935 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_730 | _GEN_3807 | _GEN_52 & _GEN_540 | _GEN_3679 | _GEN_50 & _GEN_350) & (_GEN_3551 ? io_wb_resps_0_bits_predicated : ~_GEN_3455 & rob_predicated_3_11));
    rob_predicated_3_12 <= ~(_GEN_58 & _GEN_1113 | _GEN_4064 | _GEN_56 & _GEN_923) & (_GEN_3936 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_733 | _GEN_3808 | _GEN_52 & _GEN_543 | _GEN_3680 | _GEN_50 & _GEN_353) & (_GEN_3552 ? io_wb_resps_0_bits_predicated : ~_GEN_3456 & rob_predicated_3_12));
    rob_predicated_3_13 <= ~(_GEN_58 & _GEN_1116 | _GEN_4065 | _GEN_56 & _GEN_926) & (_GEN_3937 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_736 | _GEN_3809 | _GEN_52 & _GEN_546 | _GEN_3681 | _GEN_50 & _GEN_356) & (_GEN_3553 ? io_wb_resps_0_bits_predicated : ~_GEN_3457 & rob_predicated_3_13));
    rob_predicated_3_14 <= ~(_GEN_58 & _GEN_1119 | _GEN_4066 | _GEN_56 & _GEN_929) & (_GEN_3938 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_739 | _GEN_3810 | _GEN_52 & _GEN_549 | _GEN_3682 | _GEN_50 & _GEN_359) & (_GEN_3554 ? io_wb_resps_0_bits_predicated : ~_GEN_3458 & rob_predicated_3_14));
    rob_predicated_3_15 <= ~(_GEN_58 & _GEN_1122 | _GEN_4067 | _GEN_56 & _GEN_932) & (_GEN_3939 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_742 | _GEN_3811 | _GEN_52 & _GEN_552 | _GEN_3683 | _GEN_50 & _GEN_362) & (_GEN_3555 ? io_wb_resps_0_bits_predicated : ~_GEN_3459 & rob_predicated_3_15));
    rob_predicated_3_16 <= ~(_GEN_58 & _GEN_1125 | _GEN_4068 | _GEN_56 & _GEN_935) & (_GEN_3940 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_745 | _GEN_3812 | _GEN_52 & _GEN_555 | _GEN_3684 | _GEN_50 & _GEN_365) & (_GEN_3556 ? io_wb_resps_0_bits_predicated : ~_GEN_3460 & rob_predicated_3_16));
    rob_predicated_3_17 <= ~(_GEN_58 & _GEN_1128 | _GEN_4069 | _GEN_56 & _GEN_938) & (_GEN_3941 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_748 | _GEN_3813 | _GEN_52 & _GEN_558 | _GEN_3685 | _GEN_50 & _GEN_368) & (_GEN_3557 ? io_wb_resps_0_bits_predicated : ~_GEN_3461 & rob_predicated_3_17));
    rob_predicated_3_18 <= ~(_GEN_58 & _GEN_1131 | _GEN_4070 | _GEN_56 & _GEN_941) & (_GEN_3942 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_751 | _GEN_3814 | _GEN_52 & _GEN_561 | _GEN_3686 | _GEN_50 & _GEN_371) & (_GEN_3558 ? io_wb_resps_0_bits_predicated : ~_GEN_3462 & rob_predicated_3_18));
    rob_predicated_3_19 <= ~(_GEN_58 & _GEN_1134 | _GEN_4071 | _GEN_56 & _GEN_944) & (_GEN_3943 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_754 | _GEN_3815 | _GEN_52 & _GEN_564 | _GEN_3687 | _GEN_50 & _GEN_374) & (_GEN_3559 ? io_wb_resps_0_bits_predicated : ~_GEN_3463 & rob_predicated_3_19));
    rob_predicated_3_20 <= ~(_GEN_58 & _GEN_1137 | _GEN_4072 | _GEN_56 & _GEN_947) & (_GEN_3944 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_757 | _GEN_3816 | _GEN_52 & _GEN_567 | _GEN_3688 | _GEN_50 & _GEN_377) & (_GEN_3560 ? io_wb_resps_0_bits_predicated : ~_GEN_3464 & rob_predicated_3_20));
    rob_predicated_3_21 <= ~(_GEN_58 & _GEN_1140 | _GEN_4073 | _GEN_56 & _GEN_950) & (_GEN_3945 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_760 | _GEN_3817 | _GEN_52 & _GEN_570 | _GEN_3689 | _GEN_50 & _GEN_380) & (_GEN_3561 ? io_wb_resps_0_bits_predicated : ~_GEN_3465 & rob_predicated_3_21));
    rob_predicated_3_22 <= ~(_GEN_58 & _GEN_1143 | _GEN_4074 | _GEN_56 & _GEN_953) & (_GEN_3946 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_763 | _GEN_3818 | _GEN_52 & _GEN_573 | _GEN_3690 | _GEN_50 & _GEN_383) & (_GEN_3562 ? io_wb_resps_0_bits_predicated : ~_GEN_3466 & rob_predicated_3_22));
    rob_predicated_3_23 <= ~(_GEN_58 & _GEN_1146 | _GEN_4075 | _GEN_56 & _GEN_956) & (_GEN_3947 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_766 | _GEN_3819 | _GEN_52 & _GEN_576 | _GEN_3691 | _GEN_50 & _GEN_386) & (_GEN_3563 ? io_wb_resps_0_bits_predicated : ~_GEN_3467 & rob_predicated_3_23));
    rob_predicated_3_24 <= ~(_GEN_58 & _GEN_1149 | _GEN_4076 | _GEN_56 & _GEN_959) & (_GEN_3948 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_769 | _GEN_3820 | _GEN_52 & _GEN_579 | _GEN_3692 | _GEN_50 & _GEN_389) & (_GEN_3564 ? io_wb_resps_0_bits_predicated : ~_GEN_3468 & rob_predicated_3_24));
    rob_predicated_3_25 <= ~(_GEN_58 & _GEN_1152 | _GEN_4077 | _GEN_56 & _GEN_962) & (_GEN_3949 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_772 | _GEN_3821 | _GEN_52 & _GEN_582 | _GEN_3693 | _GEN_50 & _GEN_392) & (_GEN_3565 ? io_wb_resps_0_bits_predicated : ~_GEN_3469 & rob_predicated_3_25));
    rob_predicated_3_26 <= ~(_GEN_58 & _GEN_1155 | _GEN_4078 | _GEN_56 & _GEN_965) & (_GEN_3950 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_775 | _GEN_3822 | _GEN_52 & _GEN_585 | _GEN_3694 | _GEN_50 & _GEN_395) & (_GEN_3566 ? io_wb_resps_0_bits_predicated : ~_GEN_3470 & rob_predicated_3_26));
    rob_predicated_3_27 <= ~(_GEN_58 & _GEN_1158 | _GEN_4079 | _GEN_56 & _GEN_968) & (_GEN_3951 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_778 | _GEN_3823 | _GEN_52 & _GEN_588 | _GEN_3695 | _GEN_50 & _GEN_398) & (_GEN_3567 ? io_wb_resps_0_bits_predicated : ~_GEN_3471 & rob_predicated_3_27));
    rob_predicated_3_28 <= ~(_GEN_58 & _GEN_1161 | _GEN_4080 | _GEN_56 & _GEN_971) & (_GEN_3952 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_781 | _GEN_3824 | _GEN_52 & _GEN_591 | _GEN_3696 | _GEN_50 & _GEN_401) & (_GEN_3568 ? io_wb_resps_0_bits_predicated : ~_GEN_3472 & rob_predicated_3_28));
    rob_predicated_3_29 <= ~(_GEN_58 & _GEN_1164 | _GEN_4081 | _GEN_56 & _GEN_974) & (_GEN_3953 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_784 | _GEN_3825 | _GEN_52 & _GEN_594 | _GEN_3697 | _GEN_50 & _GEN_404) & (_GEN_3569 ? io_wb_resps_0_bits_predicated : ~_GEN_3473 & rob_predicated_3_29));
    rob_predicated_3_30 <= ~(_GEN_58 & _GEN_1167 | _GEN_4082 | _GEN_56 & _GEN_977) & (_GEN_3954 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & _GEN_787 | _GEN_3826 | _GEN_52 & _GEN_597 | _GEN_3698 | _GEN_50 & _GEN_407) & (_GEN_3570 ? io_wb_resps_0_bits_predicated : ~_GEN_3474 & rob_predicated_3_30));
    rob_predicated_3_31 <= ~(_GEN_58 & (&(io_wb_resps_9_bits_uop_rob_idx[6:2])) | _GEN_4083 | _GEN_56 & (&(io_wb_resps_7_bits_uop_rob_idx[6:2]))) & (_GEN_3955 ? io_wb_resps_6_bits_predicated : ~(_GEN_54 & (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_3827 | _GEN_52 & (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_3699 | _GEN_50 & (&(io_wb_resps_1_bits_uop_rob_idx[6:2]))) & (_GEN_3571 ? io_wb_resps_0_bits_predicated : ~_GEN_3475 & rob_predicated_3_31));
    block_commit_REG <= exception_thrown;
    block_commit_REG_1 <= exception_thrown;
    block_commit_REG_2 <= block_commit_REG_1;
    REG <= exception_thrown;
    REG_1 <= REG;
    REG_2 <= exception_thrown;
    io_com_load_is_at_rob_head_REG <= casez_tmp_316 & ~(will_commit_0 | will_commit_1 | will_commit_2 | will_commit_3);
  end // always @(posedge)
  assign io_rob_tail_idx = rob_tail_idx;
  assign io_rob_head_idx = rob_head_idx;
  assign io_commit_valids_0 = will_commit_0;
  assign io_commit_valids_1 = will_commit_1;
  assign io_commit_valids_2 = will_commit_2;
  assign io_commit_valids_3 = will_commit_3;
  assign io_commit_arch_valids_0 = will_commit_0 & ~casez_tmp_10;
  assign io_commit_arch_valids_1 = will_commit_1 & ~casez_tmp_88;
  assign io_commit_arch_valids_2 = will_commit_2 & ~casez_tmp_166;
  assign io_commit_arch_valids_3 = will_commit_3 & ~casez_tmp_244;
  assign io_commit_uops_0_is_br = casez_tmp_13;
  assign io_commit_uops_0_is_jalr = casez_tmp_14;
  assign io_commit_uops_0_is_jal = casez_tmp_15;
  assign io_commit_uops_0_ftq_idx = casez_tmp_16;
  assign io_commit_uops_0_pdst = casez_tmp_19;
  assign io_commit_uops_0_stale_pdst = casez_tmp_20;
  assign io_commit_uops_0_is_fencei = casez_tmp_21;
  assign io_commit_uops_0_uses_ldq = casez_tmp_22;
  assign io_commit_uops_0_uses_stq = casez_tmp_23;
  assign io_commit_uops_0_ldst = casez_tmp_26;
  assign io_commit_uops_0_ldst_val = casez_tmp_27;
  assign io_commit_uops_0_dst_rtype = casez_tmp_28;
  assign io_commit_uops_0_debug_fsrc = _GEN_15 & _GEN_16 ? 2'h3 : casez_tmp_30;
  assign io_commit_uops_1_is_br = casez_tmp_91;
  assign io_commit_uops_1_is_jalr = casez_tmp_92;
  assign io_commit_uops_1_is_jal = casez_tmp_93;
  assign io_commit_uops_1_ftq_idx = casez_tmp_94;
  assign io_commit_uops_1_pdst = casez_tmp_97;
  assign io_commit_uops_1_stale_pdst = casez_tmp_98;
  assign io_commit_uops_1_is_fencei = casez_tmp_99;
  assign io_commit_uops_1_uses_ldq = casez_tmp_100;
  assign io_commit_uops_1_uses_stq = casez_tmp_101;
  assign io_commit_uops_1_ldst = casez_tmp_104;
  assign io_commit_uops_1_ldst_val = casez_tmp_105;
  assign io_commit_uops_1_dst_rtype = casez_tmp_106;
  assign io_commit_uops_1_debug_fsrc = _GEN_32 & _GEN_16 ? 2'h3 : casez_tmp_108;
  assign io_commit_uops_2_is_br = casez_tmp_169;
  assign io_commit_uops_2_is_jalr = casez_tmp_170;
  assign io_commit_uops_2_is_jal = casez_tmp_171;
  assign io_commit_uops_2_ftq_idx = casez_tmp_172;
  assign io_commit_uops_2_pdst = casez_tmp_175;
  assign io_commit_uops_2_stale_pdst = casez_tmp_176;
  assign io_commit_uops_2_is_fencei = casez_tmp_177;
  assign io_commit_uops_2_uses_ldq = casez_tmp_178;
  assign io_commit_uops_2_uses_stq = casez_tmp_179;
  assign io_commit_uops_2_ldst = casez_tmp_182;
  assign io_commit_uops_2_ldst_val = casez_tmp_183;
  assign io_commit_uops_2_dst_rtype = casez_tmp_184;
  assign io_commit_uops_2_debug_fsrc = _GEN_48 & _GEN_16 ? 2'h3 : casez_tmp_186;
  assign io_commit_uops_3_is_br = casez_tmp_247;
  assign io_commit_uops_3_is_jalr = casez_tmp_248;
  assign io_commit_uops_3_is_jal = casez_tmp_249;
  assign io_commit_uops_3_ftq_idx = casez_tmp_250;
  assign io_commit_uops_3_pdst = casez_tmp_253;
  assign io_commit_uops_3_stale_pdst = casez_tmp_254;
  assign io_commit_uops_3_is_fencei = casez_tmp_255;
  assign io_commit_uops_3_uses_ldq = casez_tmp_256;
  assign io_commit_uops_3_uses_stq = casez_tmp_257;
  assign io_commit_uops_3_ldst = casez_tmp_260;
  assign io_commit_uops_3_ldst_val = casez_tmp_261;
  assign io_commit_uops_3_dst_rtype = casez_tmp_262;
  assign io_commit_uops_3_debug_fsrc = _GEN_64 & _GEN_16 ? 2'h3 : casez_tmp_264;
  assign io_commit_fflags_valid = fflags_val_0 | fflags_val_1 | fflags_val_2 | fflags_val_3;
  assign io_commit_fflags_bits = (fflags_val_0 ? casez_tmp_32 : 5'h0) | (fflags_val_1 ? casez_tmp_110 : 5'h0) | (fflags_val_2 ? casez_tmp_188 : 5'h0) | (fflags_val_3 ? casez_tmp_266 : 5'h0);
  assign io_commit_rbk_valids_0 = _io_commit_rbk_valids_0_output;
  assign io_commit_rbk_valids_1 = _io_commit_rbk_valids_1_output;
  assign io_commit_rbk_valids_2 = _io_commit_rbk_valids_2_output;
  assign io_commit_rbk_valids_3 = _io_commit_rbk_valids_3_output;
  assign io_commit_rollback = _io_commit_rollback_T_3;
  assign io_com_load_is_at_rob_head = io_com_load_is_at_rob_head_REG;
  assign io_com_xcpt_valid = exception_thrown & ~is_mini_exception;
  assign io_com_xcpt_bits_ftq_idx = com_xcpt_uop_ftq_idx;
  assign io_com_xcpt_bits_edge_inst = com_xcpt_uop_edge_inst;
  assign io_com_xcpt_bits_pc_lob = com_xcpt_uop_pc_lob;
  assign io_com_xcpt_bits_cause = r_xcpt_uop_exc_cause;
  assign io_com_xcpt_bits_badvaddr = {{24{r_xcpt_badvaddr[39]}}, r_xcpt_badvaddr};
  assign io_flush_valid = _io_flush_valid_output;
  assign io_flush_bits_ftq_idx = exception_thrown ? com_xcpt_uop_ftq_idx : (flush_commit_mask_0 ? casez_tmp_16 : 6'h0) | (flush_commit_mask_1 ? casez_tmp_94 : 6'h0) | (flush_commit_mask_2 ? casez_tmp_172 : 6'h0) | (flush_commit_mask_3 ? casez_tmp_250 : 6'h0);
  assign io_flush_bits_edge_inst = exception_thrown ? com_xcpt_uop_edge_inst : flush_commit_mask_0 & casez_tmp_17 | flush_commit_mask_1 & casez_tmp_95 | flush_commit_mask_2 & casez_tmp_173 | flush_commit_mask_3 & casez_tmp_251;
  assign io_flush_bits_is_rvc = exception_thrown ? (casez_tmp_7 ? casez_tmp_12 : casez_tmp_85 ? casez_tmp_90 : casez_tmp_163 ? casez_tmp_168 : casez_tmp_246) : flush_commit_mask_0 & casez_tmp_12 | flush_commit_mask_1 & casez_tmp_90 | flush_commit_mask_2 & casez_tmp_168 | flush_commit_mask_3 & casez_tmp_246;
  assign io_flush_bits_pc_lob = exception_thrown ? com_xcpt_uop_pc_lob : (flush_commit_mask_0 ? casez_tmp_18 : 6'h0) | (flush_commit_mask_1 ? casez_tmp_96 : 6'h0) | (flush_commit_mask_2 ? casez_tmp_174 : 6'h0) | (flush_commit_mask_3 ? casez_tmp_252 : 6'h0);
  assign io_flush_bits_flush_typ = _io_flush_valid_output ? (flush_commit & (exception_thrown ? (casez_tmp_7 ? casez_tmp_11 : casez_tmp_85 ? casez_tmp_89 : casez_tmp_163 ? casez_tmp_167 : casez_tmp_245) : (flush_commit_mask_0 ? casez_tmp_11 : 7'h0) | (flush_commit_mask_1 ? casez_tmp_89 : 7'h0) | (flush_commit_mask_2 ? casez_tmp_167 : 7'h0) | (flush_commit_mask_3 ? casez_tmp_245 : 7'h0)) == 7'h6A ? 3'h3 : exception_thrown & ~is_mini_exception ? 3'h1 : exception_thrown | (casez_tmp_7 | casez_tmp_85 | casez_tmp_163 | casez_tmp_241) & (casez_tmp_7 ? casez_tmp_24 : casez_tmp_85 ? casez_tmp_102 : casez_tmp_163 ? casez_tmp_180 : casez_tmp_258) ? 3'h2 : 3'h4) : 3'h0;
  assign io_empty = empty;
  assign io_ready = _io_ready_T & ~full & ~r_xcpt_val;
  assign io_flush_frontend = r_xcpt_val;
endmodule

