VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS
MACRO memMod_dist_0
  FOREIGN memMod_dist_0 0 0 ;
  CLASS BLOCK ;
  SIZE 84.39 BY 67.91 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal7 ;
        RECT  2.9 42.7 59.38 44.1 ;
        RECT  2.9 2.7 59.38 4.1 ;
      LAYER metal4 ;
        RECT  58.9 1.315 59.38 65.885 ;
        RECT  2.9 1.315 3.38 65.885 ;
      LAYER metal1 ;
        RECT  1.14 65.715 83.22 65.885 ;
        RECT  1.14 62.915 83.22 63.085 ;
        RECT  1.14 60.115 83.22 60.285 ;
        RECT  1.14 57.315 83.22 57.485 ;
        RECT  1.14 54.515 83.22 54.685 ;
        RECT  1.14 51.715 83.22 51.885 ;
        RECT  1.14 48.915 83.22 49.085 ;
        RECT  1.14 46.115 83.22 46.285 ;
        RECT  1.14 43.315 83.22 43.485 ;
        RECT  1.14 40.515 83.22 40.685 ;
        RECT  1.14 37.715 83.22 37.885 ;
        RECT  1.14 34.915 83.22 35.085 ;
        RECT  1.14 32.115 83.22 32.285 ;
        RECT  1.14 29.315 83.22 29.485 ;
        RECT  1.14 26.515 83.22 26.685 ;
        RECT  1.14 23.715 83.22 23.885 ;
        RECT  1.14 20.915 83.22 21.085 ;
        RECT  1.14 18.115 83.22 18.285 ;
        RECT  1.14 15.315 83.22 15.485 ;
        RECT  1.14 12.515 83.22 12.685 ;
        RECT  1.14 9.715 83.22 9.885 ;
        RECT  1.14 6.915 83.22 7.085 ;
        RECT  1.14 4.115 83.22 4.285 ;
        RECT  1.14 1.315 83.22 1.485 ;
      VIA 59.14 43.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 43.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 43.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 59.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 59.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 43.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 43.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 43.4 via4_5_960_2800_5_2_600_600 ;
      VIA 3.14 3.4 via6_7_960_2800_4_1_600_600 ;
      VIA 3.14 3.4 via5_6_960_2800_5_2_600_600 ;
      VIA 3.14 3.4 via4_5_960_2800_5_2_600_600 ;
      VIA 59.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 59.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 59.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 59.14 1.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 65.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 65.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 65.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 63 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 63 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 63 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 60.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 60.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 60.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 57.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 57.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 57.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 54.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 54.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 54.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 51.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 51.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 51.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 49 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 49 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 49 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 46.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 46.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 46.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 43.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 43.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 43.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 40.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 40.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 40.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 37.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 37.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 37.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 35 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 35 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 35 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 32.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 32.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 32.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 29.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 29.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 29.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 26.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 26.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 26.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 23.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 23.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 23.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 21 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 21 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 21 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 18.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 18.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 18.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 15.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 15.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 15.4 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 12.6 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 12.6 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 12.6 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 9.8 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 9.8 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 9.8 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 7 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 7 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 7 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 4.2 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 4.2 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 4.2 via1_2_960_340_1_3_300_300 ;
      VIA 3.14 1.4 via3_4_960_340_1_3_320_320 ;
      VIA 3.14 1.4 via2_3_960_340_1_3_320_320 ;
      VIA 3.14 1.4 via1_2_960_340_1_3_300_300 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  30.9 2.715 31.38 64.485 ;
      LAYER metal1 ;
        RECT  1.14 64.315 83.22 64.485 ;
        RECT  1.14 61.515 83.22 61.685 ;
        RECT  1.14 58.715 83.22 58.885 ;
        RECT  1.14 55.915 83.22 56.085 ;
        RECT  1.14 53.115 83.22 53.285 ;
        RECT  1.14 50.315 83.22 50.485 ;
        RECT  1.14 47.515 83.22 47.685 ;
        RECT  1.14 44.715 83.22 44.885 ;
        RECT  1.14 41.915 83.22 42.085 ;
        RECT  1.14 39.115 83.22 39.285 ;
        RECT  1.14 36.315 83.22 36.485 ;
        RECT  1.14 33.515 83.22 33.685 ;
        RECT  1.14 30.715 83.22 30.885 ;
        RECT  1.14 27.915 83.22 28.085 ;
        RECT  1.14 25.115 83.22 25.285 ;
        RECT  1.14 22.315 83.22 22.485 ;
        RECT  1.14 19.515 83.22 19.685 ;
        RECT  1.14 16.715 83.22 16.885 ;
        RECT  1.14 13.915 83.22 14.085 ;
        RECT  1.14 11.115 83.22 11.285 ;
        RECT  1.14 8.315 83.22 8.485 ;
        RECT  1.14 5.515 83.22 5.685 ;
        RECT  1.14 2.715 83.22 2.885 ;
      VIA 31.14 64.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 64.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 64.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 61.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 61.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 61.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 58.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 58.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 58.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 56 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 56 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 56 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 53.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 53.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 53.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 50.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 50.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 50.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 47.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 47.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 47.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 44.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 44.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 44.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 42 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 42 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 42 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 39.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 39.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 39.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 36.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 36.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 36.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 33.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 33.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 33.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 30.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 30.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 30.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 28 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 28 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 28 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 25.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 25.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 25.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 22.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 22.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 22.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 19.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 19.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 19.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 16.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 16.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 16.8 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 14 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 14 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 14 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 11.2 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 11.2 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 11.2 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 8.4 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 8.4 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 8.4 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 5.6 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 5.6 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 5.6 via1_2_960_340_1_3_300_300 ;
      VIA 31.14 2.8 via3_4_960_340_1_3_320_320 ;
      VIA 31.14 2.8 via2_3_960_340_1_3_320_320 ;
      VIA 31.14 2.8 via1_2_960_340_1_3_300_300 ;
    END
  END VDD
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  3.385 0 3.525 0.14 ;
    END
  END clk
  PIN inAddr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  49.865 67.77 50.005 67.91 ;
    END
  END inAddr[0]
  PIN inAddr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  48.745 67.77 48.885 67.91 ;
    END
  END inAddr[1]
  PIN inAddr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  44.265 67.77 44.405 67.91 ;
    END
  END inAddr[2]
  PIN inAddr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  44.825 67.77 44.965 67.91 ;
    END
  END inAddr[3]
  PIN in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  19.625 0 19.765 0.14 ;
    END
  END in[0]
  PIN in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  84.25 12.88 84.39 13.02 ;
    END
  END in[10]
  PIN in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 63.84 0.14 63.98 ;
    END
  END in[11]
  PIN in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  59.945 67.77 60.085 67.91 ;
    END
  END in[12]
  PIN in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  36.425 0 36.565 0.14 ;
    END
  END in[13]
  PIN in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 11.2 0.14 11.34 ;
    END
  END in[14]
  PIN in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 37.52 0.14 37.66 ;
    END
  END in[15]
  PIN in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  49.865 0 50.005 0.14 ;
    END
  END in[16]
  PIN in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  43.145 0 43.285 0.14 ;
    END
  END in[17]
  PIN in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  84.25 35.84 84.39 35.98 ;
    END
  END in[18]
  PIN in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  84.25 50.96 84.39 51.1 ;
    END
  END in[19]
  PIN in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  35.865 0 36.005 0.14 ;
    END
  END in[1]
  PIN in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  84.25 28 84.39 28.14 ;
    END
  END in[20]
  PIN in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 53.76 0.14 53.9 ;
    END
  END in[21]
  PIN in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  73.385 67.77 73.525 67.91 ;
    END
  END in[22]
  PIN in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  26.345 67.77 26.485 67.91 ;
    END
  END in[23]
  PIN in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  38.105 67.77 38.245 67.91 ;
    END
  END in[24]
  PIN in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  84.25 20.72 84.39 20.86 ;
    END
  END in[25]
  PIN in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  84.25 29.68 84.39 29.82 ;
    END
  END in[26]
  PIN in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 19.04 0.14 19.18 ;
    END
  END in[27]
  PIN in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  47.065 67.77 47.205 67.91 ;
    END
  END in[28]
  PIN in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  47.625 67.77 47.765 67.91 ;
    END
  END in[29]
  PIN in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 49.28 0.14 49.42 ;
    END
  END in[2]
  PIN in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  31.385 0 31.525 0.14 ;
    END
  END in[30]
  PIN in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  53.785 0 53.925 0.14 ;
    END
  END in[31]
  PIN in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  58.825 67.77 58.965 67.91 ;
    END
  END in[3]
  PIN in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  65.545 0 65.685 0.14 ;
    END
  END in[4]
  PIN in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 43.68 0.14 43.82 ;
    END
  END in[5]
  PIN in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  84.25 43.68 84.39 43.82 ;
    END
  END in[6]
  PIN in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 35.28 0.14 35.42 ;
    END
  END in[7]
  PIN in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 26.88 0.14 27.02 ;
    END
  END in[8]
  PIN in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  24.105 0 24.245 0.14 ;
    END
  END in[9]
  PIN outAddr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  4.505 0 4.645 0.14 ;
    END
  END outAddr[0]
  PIN outAddr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  5.065 0 5.205 0.14 ;
    END
  END outAddr[1]
  PIN outAddr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  8.425 0 8.565 0.14 ;
    END
  END outAddr[2]
  PIN outAddr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  10.665 0 10.805 0.14 ;
    END
  END outAddr[3]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  26.905 0 27.045 0.14 ;
    END
  END out[0]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  84.25 16.8 84.39 16.94 ;
    END
  END out[10]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  17.385 67.77 17.525 67.91 ;
    END
  END out[11]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  59.385 67.77 59.525 67.91 ;
    END
  END out[12]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  43.705 0 43.845 0.14 ;
    END
  END out[13]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  12.905 0 13.045 0.14 ;
    END
  END out[14]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 34.16 0.14 34.3 ;
    END
  END out[15]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  56.585 0 56.725 0.14 ;
    END
  END out[16]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  49.305 0 49.445 0.14 ;
    END
  END out[17]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  84.25 39.76 84.39 39.9 ;
    END
  END out[18]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  84.25 54.88 84.39 55.02 ;
    END
  END out[19]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  42.585 0 42.725 0.14 ;
    END
  END out[1]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  84.25 31.36 84.39 31.5 ;
    END
  END out[20]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 49.84 0.14 49.98 ;
    END
  END out[21]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  72.265 67.77 72.405 67.91 ;
    END
  END out[22]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  26.905 67.77 27.045 67.91 ;
    END
  END out[23]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  36.985 67.77 37.125 67.91 ;
    END
  END out[24]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  84.25 21.84 84.39 21.98 ;
    END
  END out[25]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  84.25 33.6 84.39 33.74 ;
    END
  END out[26]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 16.8 0.14 16.94 ;
    END
  END out[27]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  41.465 67.77 41.605 67.91 ;
    END
  END out[28]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  48.185 67.77 48.325 67.91 ;
    END
  END out[29]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  28.585 67.77 28.725 67.91 ;
    END
  END out[2]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  40.345 0 40.485 0.14 ;
    END
  END out[30]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  59.945 0 60.085 0.14 ;
    END
  END out[31]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  84.25 44.24 84.39 44.38 ;
    END
  END out[3]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  84.25 6.72 84.39 6.86 ;
    END
  END out[4]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 41.44 0.14 41.58 ;
    END
  END out[5]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  84.25 44.8 84.39 44.94 ;
    END
  END out[6]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 33.6 0.14 33.74 ;
    END
  END out[7]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 25.76 0.14 25.9 ;
    END
  END out[8]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  29.705 0 29.845 0.14 ;
    END
  END out[9]
  PIN writeSel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  49.305 67.77 49.445 67.91 ;
    END
  END writeSel
  OBS
    LAYER metal1 ;
     RECT  0 0 84.39 67.91 ;
    LAYER metal2 ;
     RECT  0 0 84.39 67.91 ;
    LAYER metal3 ;
     RECT  0 0 84.39 67.91 ;
    LAYER metal4 ;
     RECT  0 0 84.39 67.91 ;
    LAYER metal5 ;
     RECT  0 0 84.39 67.91 ;
    LAYER metal6 ;
     RECT  0 0 84.39 67.91 ;
    LAYER metal7 ;
     RECT  0 0 84.39 67.91 ;
  END
END memMod_dist_0
END LIBRARY
