../../nangate45/lef/fakeram45_1024x32.lef