module MuxTest_width_64_inputs_16_outputs_16_pipeline_5( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [3:0]  io_selects_0_0, // @[:@6.4]
  input  [3:0]  io_selects_0_1, // @[:@6.4]
  input  [3:0]  io_selects_1_0, // @[:@6.4]
  input  [3:0]  io_selects_1_1, // @[:@6.4]
  input  [3:0]  io_selects_2_0, // @[:@6.4]
  input  [3:0]  io_selects_2_1, // @[:@6.4]
  input  [3:0]  io_selects_3_0, // @[:@6.4]
  input  [3:0]  io_selects_3_1, // @[:@6.4]
  input  [3:0]  io_selects_4_0, // @[:@6.4]
  input  [3:0]  io_selects_4_1, // @[:@6.4]
  input  [3:0]  io_selects_5_0, // @[:@6.4]
  input  [3:0]  io_selects_5_1, // @[:@6.4]
  input  [3:0]  io_selects_6_0, // @[:@6.4]
  input  [3:0]  io_selects_6_1, // @[:@6.4]
  input  [3:0]  io_selects_7_0, // @[:@6.4]
  input  [3:0]  io_selects_7_1, // @[:@6.4]
  input  [3:0]  io_selects_8_0, // @[:@6.4]
  input  [3:0]  io_selects_8_1, // @[:@6.4]
  input  [3:0]  io_selects_9_0, // @[:@6.4]
  input  [3:0]  io_selects_9_1, // @[:@6.4]
  input  [3:0]  io_selects_10_0, // @[:@6.4]
  input  [3:0]  io_selects_10_1, // @[:@6.4]
  input  [3:0]  io_selects_11_0, // @[:@6.4]
  input  [3:0]  io_selects_11_1, // @[:@6.4]
  input  [3:0]  io_selects_12_0, // @[:@6.4]
  input  [3:0]  io_selects_12_1, // @[:@6.4]
  input  [3:0]  io_selects_13_0, // @[:@6.4]
  input  [3:0]  io_selects_13_1, // @[:@6.4]
  input  [3:0]  io_selects_14_0, // @[:@6.4]
  input  [3:0]  io_selects_14_1, // @[:@6.4]
  input  [3:0]  io_selects_15_0, // @[:@6.4]
  input  [3:0]  io_selects_15_1, // @[:@6.4]
  input  [2:0]  io_operation_0, // @[:@6.4]
  input  [2:0]  io_operation_1, // @[:@6.4]
  input  [2:0]  io_operation_2, // @[:@6.4]
  input  [2:0]  io_operation_3, // @[:@6.4]
  input  [2:0]  io_operation_4, // @[:@6.4]
  input  [2:0]  io_operation_5, // @[:@6.4]
  input  [2:0]  io_operation_6, // @[:@6.4]
  input  [2:0]  io_operation_7, // @[:@6.4]
  input  [2:0]  io_operation_8, // @[:@6.4]
  input  [2:0]  io_operation_9, // @[:@6.4]
  input  [2:0]  io_operation_10, // @[:@6.4]
  input  [2:0]  io_operation_11, // @[:@6.4]
  input  [2:0]  io_operation_12, // @[:@6.4]
  input  [2:0]  io_operation_13, // @[:@6.4]
  input  [2:0]  io_operation_14, // @[:@6.4]
  input  [2:0]  io_operation_15, // @[:@6.4]
  input  [63:0] io_inputs_0, // @[:@6.4]
  input  [63:0] io_inputs_1, // @[:@6.4]
  input  [63:0] io_inputs_2, // @[:@6.4]
  input  [63:0] io_inputs_3, // @[:@6.4]
  input  [63:0] io_inputs_4, // @[:@6.4]
  input  [63:0] io_inputs_5, // @[:@6.4]
  input  [63:0] io_inputs_6, // @[:@6.4]
  input  [63:0] io_inputs_7, // @[:@6.4]
  input  [63:0] io_inputs_8, // @[:@6.4]
  input  [63:0] io_inputs_9, // @[:@6.4]
  input  [63:0] io_inputs_10, // @[:@6.4]
  input  [63:0] io_inputs_11, // @[:@6.4]
  input  [63:0] io_inputs_12, // @[:@6.4]
  input  [63:0] io_inputs_13, // @[:@6.4]
  input  [63:0] io_inputs_14, // @[:@6.4]
  input  [63:0] io_inputs_15, // @[:@6.4]
  output [63:0] io_outputs_0, // @[:@6.4]
  output [63:0] io_outputs_1, // @[:@6.4]
  output [63:0] io_outputs_2, // @[:@6.4]
  output [63:0] io_outputs_3, // @[:@6.4]
  output [63:0] io_outputs_4, // @[:@6.4]
  output [63:0] io_outputs_5, // @[:@6.4]
  output [63:0] io_outputs_6, // @[:@6.4]
  output [63:0] io_outputs_7, // @[:@6.4]
  output [63:0] io_outputs_8, // @[:@6.4]
  output [63:0] io_outputs_9, // @[:@6.4]
  output [63:0] io_outputs_10, // @[:@6.4]
  output [63:0] io_outputs_11, // @[:@6.4]
  output [63:0] io_outputs_12, // @[:@6.4]
  output [63:0] io_outputs_13, // @[:@6.4]
  output [63:0] io_outputs_14, // @[:@6.4]
  output [63:0] io_outputs_15 // @[:@6.4]
);
  wire [63:0] _GEN_1; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_2; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_3; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_4; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_5; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_6; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_7; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_8; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_9; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_10; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_11; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_12; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_13; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_14; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_15; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_17; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_18; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_19; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_20; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_21; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_22; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_23; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_24; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_25; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_26; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_27; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_28; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_29; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_30; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _GEN_31; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [64:0] _T_722; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [63:0] _T_723; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@9.4]
  wire [127:0] _T_725; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@10.4]
  wire [63:0] _T_727; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@11.4]
  wire  _T_728; // @[Mux.scala 46:19:@12.4]
  wire [63:0] _T_729; // @[Mux.scala 46:16:@13.4]
  wire  _T_730; // @[Mux.scala 46:19:@14.4]
  wire [127:0] _T_731; // @[Mux.scala 46:16:@15.4]
  wire  _T_732; // @[Mux.scala 46:19:@16.4]
  wire [127:0] _T_733; // @[Mux.scala 46:16:@17.4]
  wire  _T_734; // @[Mux.scala 46:19:@18.4]
  wire [63:0] _GEN_33; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_34; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_35; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_36; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_37; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_38; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_39; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_40; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_41; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_42; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_43; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_44; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_45; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_46; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_47; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_49; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_50; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_51; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_52; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_53; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_54; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_55; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_56; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_57; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_58; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_59; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_60; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_61; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_62; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _GEN_63; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [64:0] _T_739; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [63:0] _T_740; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@21.4]
  wire [127:0] _T_742; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@22.4]
  wire [63:0] _T_744; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@23.4]
  wire  _T_745; // @[Mux.scala 46:19:@24.4]
  wire [63:0] _T_746; // @[Mux.scala 46:16:@25.4]
  wire  _T_747; // @[Mux.scala 46:19:@26.4]
  wire [127:0] _T_748; // @[Mux.scala 46:16:@27.4]
  wire  _T_749; // @[Mux.scala 46:19:@28.4]
  wire [127:0] _T_750; // @[Mux.scala 46:16:@29.4]
  wire  _T_751; // @[Mux.scala 46:19:@30.4]
  wire [63:0] _GEN_65; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_66; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_67; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_68; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_69; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_70; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_71; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_72; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_73; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_74; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_75; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_76; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_77; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_78; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_79; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_81; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_82; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_83; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_84; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_85; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_86; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_87; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_88; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_89; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_90; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_91; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_92; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_93; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_94; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _GEN_95; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [64:0] _T_756; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [63:0] _T_757; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@33.4]
  wire [127:0] _T_759; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@34.4]
  wire [63:0] _T_761; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@35.4]
  wire  _T_762; // @[Mux.scala 46:19:@36.4]
  wire [63:0] _T_763; // @[Mux.scala 46:16:@37.4]
  wire  _T_764; // @[Mux.scala 46:19:@38.4]
  wire [127:0] _T_765; // @[Mux.scala 46:16:@39.4]
  wire  _T_766; // @[Mux.scala 46:19:@40.4]
  wire [127:0] _T_767; // @[Mux.scala 46:16:@41.4]
  wire  _T_768; // @[Mux.scala 46:19:@42.4]
  wire [63:0] _GEN_97; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_98; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_99; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_100; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_101; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_102; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_103; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_104; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_105; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_106; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_107; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_108; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_109; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_110; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_111; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_113; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_114; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_115; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_116; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_117; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_118; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_119; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_120; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_121; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_122; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_123; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_124; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_125; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_126; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _GEN_127; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [64:0] _T_773; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [63:0] _T_774; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@45.4]
  wire [127:0] _T_776; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@46.4]
  wire [63:0] _T_778; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@47.4]
  wire  _T_779; // @[Mux.scala 46:19:@48.4]
  wire [63:0] _T_780; // @[Mux.scala 46:16:@49.4]
  wire  _T_781; // @[Mux.scala 46:19:@50.4]
  wire [127:0] _T_782; // @[Mux.scala 46:16:@51.4]
  wire  _T_783; // @[Mux.scala 46:19:@52.4]
  wire [127:0] _T_784; // @[Mux.scala 46:16:@53.4]
  wire  _T_785; // @[Mux.scala 46:19:@54.4]
  wire [63:0] _GEN_129; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_130; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_131; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_132; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_133; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_134; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_135; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_136; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_137; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_138; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_139; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_140; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_141; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_142; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_143; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_145; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_146; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_147; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_148; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_149; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_150; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_151; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_152; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_153; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_154; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_155; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_156; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_157; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_158; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _GEN_159; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [64:0] _T_790; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [63:0] _T_791; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@57.4]
  wire [127:0] _T_793; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@58.4]
  wire [63:0] _T_795; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@59.4]
  wire  _T_796; // @[Mux.scala 46:19:@60.4]
  wire [63:0] _T_797; // @[Mux.scala 46:16:@61.4]
  wire  _T_798; // @[Mux.scala 46:19:@62.4]
  wire [127:0] _T_799; // @[Mux.scala 46:16:@63.4]
  wire  _T_800; // @[Mux.scala 46:19:@64.4]
  wire [127:0] _T_801; // @[Mux.scala 46:16:@65.4]
  wire  _T_802; // @[Mux.scala 46:19:@66.4]
  wire [63:0] _GEN_161; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_162; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_163; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_164; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_165; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_166; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_167; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_168; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_169; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_170; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_171; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_172; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_173; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_174; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_175; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_177; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_178; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_179; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_180; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_181; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_182; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_183; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_184; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_185; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_186; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_187; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_188; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_189; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_190; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _GEN_191; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [64:0] _T_807; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [63:0] _T_808; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@69.4]
  wire [127:0] _T_810; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@70.4]
  wire [63:0] _T_812; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@71.4]
  wire  _T_813; // @[Mux.scala 46:19:@72.4]
  wire [63:0] _T_814; // @[Mux.scala 46:16:@73.4]
  wire  _T_815; // @[Mux.scala 46:19:@74.4]
  wire [127:0] _T_816; // @[Mux.scala 46:16:@75.4]
  wire  _T_817; // @[Mux.scala 46:19:@76.4]
  wire [127:0] _T_818; // @[Mux.scala 46:16:@77.4]
  wire  _T_819; // @[Mux.scala 46:19:@78.4]
  wire [63:0] _GEN_193; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_194; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_195; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_196; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_197; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_198; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_199; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_200; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_201; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_202; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_203; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_204; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_205; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_206; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_207; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_209; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_210; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_211; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_212; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_213; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_214; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_215; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_216; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_217; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_218; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_219; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_220; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_221; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_222; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _GEN_223; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [64:0] _T_824; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [63:0] _T_825; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@81.4]
  wire [127:0] _T_827; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@82.4]
  wire [63:0] _T_829; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@83.4]
  wire  _T_830; // @[Mux.scala 46:19:@84.4]
  wire [63:0] _T_831; // @[Mux.scala 46:16:@85.4]
  wire  _T_832; // @[Mux.scala 46:19:@86.4]
  wire [127:0] _T_833; // @[Mux.scala 46:16:@87.4]
  wire  _T_834; // @[Mux.scala 46:19:@88.4]
  wire [127:0] _T_835; // @[Mux.scala 46:16:@89.4]
  wire  _T_836; // @[Mux.scala 46:19:@90.4]
  wire [63:0] _GEN_225; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_226; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_227; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_228; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_229; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_230; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_231; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_232; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_233; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_234; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_235; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_236; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_237; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_238; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_239; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_241; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_242; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_243; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_244; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_245; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_246; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_247; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_248; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_249; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_250; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_251; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_252; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_253; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_254; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _GEN_255; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [64:0] _T_841; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [63:0] _T_842; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@93.4]
  wire [127:0] _T_844; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@94.4]
  wire [63:0] _T_846; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@95.4]
  wire  _T_847; // @[Mux.scala 46:19:@96.4]
  wire [63:0] _T_848; // @[Mux.scala 46:16:@97.4]
  wire  _T_849; // @[Mux.scala 46:19:@98.4]
  wire [127:0] _T_850; // @[Mux.scala 46:16:@99.4]
  wire  _T_851; // @[Mux.scala 46:19:@100.4]
  wire [127:0] _T_852; // @[Mux.scala 46:16:@101.4]
  wire  _T_853; // @[Mux.scala 46:19:@102.4]
  wire [63:0] _GEN_257; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_258; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_259; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_260; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_261; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_262; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_263; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_264; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_265; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_266; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_267; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_268; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_269; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_270; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_271; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_273; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_274; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_275; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_276; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_277; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_278; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_279; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_280; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_281; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_282; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_283; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_284; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_285; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_286; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _GEN_287; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [64:0] _T_858; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [63:0] _T_859; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@105.4]
  wire [127:0] _T_861; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@106.4]
  wire [63:0] _T_863; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@107.4]
  wire  _T_864; // @[Mux.scala 46:19:@108.4]
  wire [63:0] _T_865; // @[Mux.scala 46:16:@109.4]
  wire  _T_866; // @[Mux.scala 46:19:@110.4]
  wire [127:0] _T_867; // @[Mux.scala 46:16:@111.4]
  wire  _T_868; // @[Mux.scala 46:19:@112.4]
  wire [127:0] _T_869; // @[Mux.scala 46:16:@113.4]
  wire  _T_870; // @[Mux.scala 46:19:@114.4]
  wire [63:0] _GEN_289; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_290; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_291; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_292; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_293; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_294; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_295; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_296; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_297; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_298; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_299; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_300; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_301; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_302; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_303; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_305; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_306; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_307; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_308; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_309; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_310; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_311; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_312; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_313; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_314; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_315; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_316; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_317; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_318; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _GEN_319; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [64:0] _T_875; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [63:0] _T_876; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@117.4]
  wire [127:0] _T_878; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@118.4]
  wire [63:0] _T_880; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@119.4]
  wire  _T_881; // @[Mux.scala 46:19:@120.4]
  wire [63:0] _T_882; // @[Mux.scala 46:16:@121.4]
  wire  _T_883; // @[Mux.scala 46:19:@122.4]
  wire [127:0] _T_884; // @[Mux.scala 46:16:@123.4]
  wire  _T_885; // @[Mux.scala 46:19:@124.4]
  wire [127:0] _T_886; // @[Mux.scala 46:16:@125.4]
  wire  _T_887; // @[Mux.scala 46:19:@126.4]
  wire [63:0] _GEN_321; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_322; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_323; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_324; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_325; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_326; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_327; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_328; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_329; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_330; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_331; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_332; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_333; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_334; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_335; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_337; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_338; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_339; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_340; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_341; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_342; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_343; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_344; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_345; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_346; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_347; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_348; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_349; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_350; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _GEN_351; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [64:0] _T_892; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [63:0] _T_893; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@129.4]
  wire [127:0] _T_895; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@130.4]
  wire [63:0] _T_897; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@131.4]
  wire  _T_898; // @[Mux.scala 46:19:@132.4]
  wire [63:0] _T_899; // @[Mux.scala 46:16:@133.4]
  wire  _T_900; // @[Mux.scala 46:19:@134.4]
  wire [127:0] _T_901; // @[Mux.scala 46:16:@135.4]
  wire  _T_902; // @[Mux.scala 46:19:@136.4]
  wire [127:0] _T_903; // @[Mux.scala 46:16:@137.4]
  wire  _T_904; // @[Mux.scala 46:19:@138.4]
  wire [63:0] _GEN_353; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_354; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_355; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_356; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_357; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_358; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_359; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_360; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_361; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_362; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_363; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_364; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_365; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_366; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_367; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_369; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_370; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_371; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_372; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_373; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_374; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_375; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_376; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_377; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_378; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_379; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_380; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_381; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_382; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _GEN_383; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [64:0] _T_909; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [63:0] _T_910; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@141.4]
  wire [127:0] _T_912; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@142.4]
  wire [63:0] _T_914; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@143.4]
  wire  _T_915; // @[Mux.scala 46:19:@144.4]
  wire [63:0] _T_916; // @[Mux.scala 46:16:@145.4]
  wire  _T_917; // @[Mux.scala 46:19:@146.4]
  wire [127:0] _T_918; // @[Mux.scala 46:16:@147.4]
  wire  _T_919; // @[Mux.scala 46:19:@148.4]
  wire [127:0] _T_920; // @[Mux.scala 46:16:@149.4]
  wire  _T_921; // @[Mux.scala 46:19:@150.4]
  wire [63:0] _GEN_385; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_386; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_387; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_388; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_389; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_390; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_391; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_392; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_393; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_394; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_395; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_396; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_397; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_398; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_399; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_401; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_402; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_403; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_404; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_405; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_406; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_407; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_408; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_409; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_410; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_411; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_412; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_413; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_414; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _GEN_415; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [64:0] _T_926; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [63:0] _T_927; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@153.4]
  wire [127:0] _T_929; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@154.4]
  wire [63:0] _T_931; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@155.4]
  wire  _T_932; // @[Mux.scala 46:19:@156.4]
  wire [63:0] _T_933; // @[Mux.scala 46:16:@157.4]
  wire  _T_934; // @[Mux.scala 46:19:@158.4]
  wire [127:0] _T_935; // @[Mux.scala 46:16:@159.4]
  wire  _T_936; // @[Mux.scala 46:19:@160.4]
  wire [127:0] _T_937; // @[Mux.scala 46:16:@161.4]
  wire  _T_938; // @[Mux.scala 46:19:@162.4]
  wire [63:0] _GEN_417; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_418; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_419; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_420; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_421; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_422; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_423; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_424; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_425; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_426; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_427; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_428; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_429; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_430; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_431; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_433; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_434; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_435; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_436; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_437; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_438; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_439; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_440; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_441; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_442; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_443; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_444; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_445; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_446; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _GEN_447; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [64:0] _T_943; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [63:0] _T_944; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@165.4]
  wire [127:0] _T_946; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@166.4]
  wire [63:0] _T_948; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@167.4]
  wire  _T_949; // @[Mux.scala 46:19:@168.4]
  wire [63:0] _T_950; // @[Mux.scala 46:16:@169.4]
  wire  _T_951; // @[Mux.scala 46:19:@170.4]
  wire [127:0] _T_952; // @[Mux.scala 46:16:@171.4]
  wire  _T_953; // @[Mux.scala 46:19:@172.4]
  wire [127:0] _T_954; // @[Mux.scala 46:16:@173.4]
  wire  _T_955; // @[Mux.scala 46:19:@174.4]
  wire [63:0] _GEN_449; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_450; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_451; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_452; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_453; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_454; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_455; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_456; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_457; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_458; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_459; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_460; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_461; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_462; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_463; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_465; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_466; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_467; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_468; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_469; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_470; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_471; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_472; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_473; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_474; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_475; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_476; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_477; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_478; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _GEN_479; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [64:0] _T_960; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [63:0] _T_961; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@177.4]
  wire [127:0] _T_963; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@178.4]
  wire [63:0] _T_965; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@179.4]
  wire  _T_966; // @[Mux.scala 46:19:@180.4]
  wire [63:0] _T_967; // @[Mux.scala 46:16:@181.4]
  wire  _T_968; // @[Mux.scala 46:19:@182.4]
  wire [127:0] _T_969; // @[Mux.scala 46:16:@183.4]
  wire  _T_970; // @[Mux.scala 46:19:@184.4]
  wire [127:0] _T_971; // @[Mux.scala 46:16:@185.4]
  wire  _T_972; // @[Mux.scala 46:19:@186.4]
  wire [63:0] _GEN_481; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_482; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_483; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_484; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_485; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_486; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_487; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_488; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_489; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_490; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_491; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_492; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_493; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_494; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_495; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_497; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_498; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_499; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_500; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_501; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_502; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_503; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_504; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_505; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_506; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_507; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_508; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_509; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_510; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _GEN_511; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [64:0] _T_977; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [63:0] _T_978; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@189.4]
  wire [127:0] _T_980; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@190.4]
  wire [63:0] _T_982; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@191.4]
  wire  _T_983; // @[Mux.scala 46:19:@192.4]
  wire [63:0] _T_984; // @[Mux.scala 46:16:@193.4]
  wire  _T_985; // @[Mux.scala 46:19:@194.4]
  wire [127:0] _T_986; // @[Mux.scala 46:16:@195.4]
  wire  _T_987; // @[Mux.scala 46:19:@196.4]
  wire [127:0] _T_988; // @[Mux.scala 46:16:@197.4]
  wire  _T_989; // @[Mux.scala 46:19:@198.4]
  reg [127:0] _T_993; // @[Reg.scala 11:16:@200.4]
  reg [127:0] _RAND_0;
  reg [127:0] _T_995; // @[Reg.scala 11:16:@204.4]
  reg [127:0] _RAND_1;
  reg [127:0] _T_997; // @[Reg.scala 11:16:@208.4]
  reg [127:0] _RAND_2;
  reg [127:0] _T_999; // @[Reg.scala 11:16:@212.4]
  reg [127:0] _RAND_3;
  reg [127:0] _T_1001; // @[Reg.scala 11:16:@216.4]
  reg [127:0] _RAND_4;
  reg [127:0] _T_1004; // @[Reg.scala 11:16:@220.4]
  reg [127:0] _RAND_5;
  reg [127:0] _T_1006; // @[Reg.scala 11:16:@224.4]
  reg [127:0] _RAND_6;
  reg [127:0] _T_1008; // @[Reg.scala 11:16:@228.4]
  reg [127:0] _RAND_7;
  reg [127:0] _T_1010; // @[Reg.scala 11:16:@232.4]
  reg [127:0] _RAND_8;
  reg [127:0] _T_1012; // @[Reg.scala 11:16:@236.4]
  reg [127:0] _RAND_9;
  reg [127:0] _T_1015; // @[Reg.scala 11:16:@240.4]
  reg [127:0] _RAND_10;
  reg [127:0] _T_1017; // @[Reg.scala 11:16:@244.4]
  reg [127:0] _RAND_11;
  reg [127:0] _T_1019; // @[Reg.scala 11:16:@248.4]
  reg [127:0] _RAND_12;
  reg [127:0] _T_1021; // @[Reg.scala 11:16:@252.4]
  reg [127:0] _RAND_13;
  reg [127:0] _T_1023; // @[Reg.scala 11:16:@256.4]
  reg [127:0] _RAND_14;
  reg [127:0] _T_1026; // @[Reg.scala 11:16:@260.4]
  reg [127:0] _RAND_15;
  reg [127:0] _T_1028; // @[Reg.scala 11:16:@264.4]
  reg [127:0] _RAND_16;
  reg [127:0] _T_1030; // @[Reg.scala 11:16:@268.4]
  reg [127:0] _RAND_17;
  reg [127:0] _T_1032; // @[Reg.scala 11:16:@272.4]
  reg [127:0] _RAND_18;
  reg [127:0] _T_1034; // @[Reg.scala 11:16:@276.4]
  reg [127:0] _RAND_19;
  reg [127:0] _T_1037; // @[Reg.scala 11:16:@280.4]
  reg [127:0] _RAND_20;
  reg [127:0] _T_1039; // @[Reg.scala 11:16:@284.4]
  reg [127:0] _RAND_21;
  reg [127:0] _T_1041; // @[Reg.scala 11:16:@288.4]
  reg [127:0] _RAND_22;
  reg [127:0] _T_1043; // @[Reg.scala 11:16:@292.4]
  reg [127:0] _RAND_23;
  reg [127:0] _T_1045; // @[Reg.scala 11:16:@296.4]
  reg [127:0] _RAND_24;
  reg [127:0] _T_1048; // @[Reg.scala 11:16:@300.4]
  reg [127:0] _RAND_25;
  reg [127:0] _T_1050; // @[Reg.scala 11:16:@304.4]
  reg [127:0] _RAND_26;
  reg [127:0] _T_1052; // @[Reg.scala 11:16:@308.4]
  reg [127:0] _RAND_27;
  reg [127:0] _T_1054; // @[Reg.scala 11:16:@312.4]
  reg [127:0] _RAND_28;
  reg [127:0] _T_1056; // @[Reg.scala 11:16:@316.4]
  reg [127:0] _RAND_29;
  reg [127:0] _T_1059; // @[Reg.scala 11:16:@320.4]
  reg [127:0] _RAND_30;
  reg [127:0] _T_1061; // @[Reg.scala 11:16:@324.4]
  reg [127:0] _RAND_31;
  reg [127:0] _T_1063; // @[Reg.scala 11:16:@328.4]
  reg [127:0] _RAND_32;
  reg [127:0] _T_1065; // @[Reg.scala 11:16:@332.4]
  reg [127:0] _RAND_33;
  reg [127:0] _T_1067; // @[Reg.scala 11:16:@336.4]
  reg [127:0] _RAND_34;
  reg [127:0] _T_1070; // @[Reg.scala 11:16:@340.4]
  reg [127:0] _RAND_35;
  reg [127:0] _T_1072; // @[Reg.scala 11:16:@344.4]
  reg [127:0] _RAND_36;
  reg [127:0] _T_1074; // @[Reg.scala 11:16:@348.4]
  reg [127:0] _RAND_37;
  reg [127:0] _T_1076; // @[Reg.scala 11:16:@352.4]
  reg [127:0] _RAND_38;
  reg [127:0] _T_1078; // @[Reg.scala 11:16:@356.4]
  reg [127:0] _RAND_39;
  reg [127:0] _T_1081; // @[Reg.scala 11:16:@360.4]
  reg [127:0] _RAND_40;
  reg [127:0] _T_1083; // @[Reg.scala 11:16:@364.4]
  reg [127:0] _RAND_41;
  reg [127:0] _T_1085; // @[Reg.scala 11:16:@368.4]
  reg [127:0] _RAND_42;
  reg [127:0] _T_1087; // @[Reg.scala 11:16:@372.4]
  reg [127:0] _RAND_43;
  reg [127:0] _T_1089; // @[Reg.scala 11:16:@376.4]
  reg [127:0] _RAND_44;
  reg [127:0] _T_1092; // @[Reg.scala 11:16:@380.4]
  reg [127:0] _RAND_45;
  reg [127:0] _T_1094; // @[Reg.scala 11:16:@384.4]
  reg [127:0] _RAND_46;
  reg [127:0] _T_1096; // @[Reg.scala 11:16:@388.4]
  reg [127:0] _RAND_47;
  reg [127:0] _T_1098; // @[Reg.scala 11:16:@392.4]
  reg [127:0] _RAND_48;
  reg [127:0] _T_1100; // @[Reg.scala 11:16:@396.4]
  reg [127:0] _RAND_49;
  reg [127:0] _T_1103; // @[Reg.scala 11:16:@400.4]
  reg [127:0] _RAND_50;
  reg [127:0] _T_1105; // @[Reg.scala 11:16:@404.4]
  reg [127:0] _RAND_51;
  reg [127:0] _T_1107; // @[Reg.scala 11:16:@408.4]
  reg [127:0] _RAND_52;
  reg [127:0] _T_1109; // @[Reg.scala 11:16:@412.4]
  reg [127:0] _RAND_53;
  reg [127:0] _T_1111; // @[Reg.scala 11:16:@416.4]
  reg [127:0] _RAND_54;
  reg [127:0] _T_1114; // @[Reg.scala 11:16:@420.4]
  reg [127:0] _RAND_55;
  reg [127:0] _T_1116; // @[Reg.scala 11:16:@424.4]
  reg [127:0] _RAND_56;
  reg [127:0] _T_1118; // @[Reg.scala 11:16:@428.4]
  reg [127:0] _RAND_57;
  reg [127:0] _T_1120; // @[Reg.scala 11:16:@432.4]
  reg [127:0] _RAND_58;
  reg [127:0] _T_1122; // @[Reg.scala 11:16:@436.4]
  reg [127:0] _RAND_59;
  reg [127:0] _T_1125; // @[Reg.scala 11:16:@440.4]
  reg [127:0] _RAND_60;
  reg [127:0] _T_1127; // @[Reg.scala 11:16:@444.4]
  reg [127:0] _RAND_61;
  reg [127:0] _T_1129; // @[Reg.scala 11:16:@448.4]
  reg [127:0] _RAND_62;
  reg [127:0] _T_1131; // @[Reg.scala 11:16:@452.4]
  reg [127:0] _RAND_63;
  reg [127:0] _T_1133; // @[Reg.scala 11:16:@456.4]
  reg [127:0] _RAND_64;
  reg [127:0] _T_1136; // @[Reg.scala 11:16:@460.4]
  reg [127:0] _RAND_65;
  reg [127:0] _T_1138; // @[Reg.scala 11:16:@464.4]
  reg [127:0] _RAND_66;
  reg [127:0] _T_1140; // @[Reg.scala 11:16:@468.4]
  reg [127:0] _RAND_67;
  reg [127:0] _T_1142; // @[Reg.scala 11:16:@472.4]
  reg [127:0] _RAND_68;
  reg [127:0] _T_1144; // @[Reg.scala 11:16:@476.4]
  reg [127:0] _RAND_69;
  reg [127:0] _T_1147; // @[Reg.scala 11:16:@480.4]
  reg [127:0] _RAND_70;
  reg [127:0] _T_1149; // @[Reg.scala 11:16:@484.4]
  reg [127:0] _RAND_71;
  reg [127:0] _T_1151; // @[Reg.scala 11:16:@488.4]
  reg [127:0] _RAND_72;
  reg [127:0] _T_1153; // @[Reg.scala 11:16:@492.4]
  reg [127:0] _RAND_73;
  reg [127:0] _T_1155; // @[Reg.scala 11:16:@496.4]
  reg [127:0] _RAND_74;
  reg [127:0] _T_1158; // @[Reg.scala 11:16:@500.4]
  reg [127:0] _RAND_75;
  reg [127:0] _T_1160; // @[Reg.scala 11:16:@504.4]
  reg [127:0] _RAND_76;
  reg [127:0] _T_1162; // @[Reg.scala 11:16:@508.4]
  reg [127:0] _RAND_77;
  reg [127:0] _T_1164; // @[Reg.scala 11:16:@512.4]
  reg [127:0] _RAND_78;
  reg [127:0] _T_1166; // @[Reg.scala 11:16:@516.4]
  reg [127:0] _RAND_79;
  assign _GEN_1 = 4'h1 == io_selects_0_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_2 = 4'h2 == io_selects_0_0 ? io_inputs_2 : _GEN_1; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_3 = 4'h3 == io_selects_0_0 ? io_inputs_3 : _GEN_2; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_4 = 4'h4 == io_selects_0_0 ? io_inputs_4 : _GEN_3; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_5 = 4'h5 == io_selects_0_0 ? io_inputs_5 : _GEN_4; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_6 = 4'h6 == io_selects_0_0 ? io_inputs_6 : _GEN_5; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_7 = 4'h7 == io_selects_0_0 ? io_inputs_7 : _GEN_6; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_8 = 4'h8 == io_selects_0_0 ? io_inputs_8 : _GEN_7; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_9 = 4'h9 == io_selects_0_0 ? io_inputs_9 : _GEN_8; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_10 = 4'ha == io_selects_0_0 ? io_inputs_10 : _GEN_9; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_11 = 4'hb == io_selects_0_0 ? io_inputs_11 : _GEN_10; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_12 = 4'hc == io_selects_0_0 ? io_inputs_12 : _GEN_11; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_13 = 4'hd == io_selects_0_0 ? io_inputs_13 : _GEN_12; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_14 = 4'he == io_selects_0_0 ? io_inputs_14 : _GEN_13; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_15 = 4'hf == io_selects_0_0 ? io_inputs_15 : _GEN_14; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_17 = 4'h1 == io_selects_0_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_18 = 4'h2 == io_selects_0_1 ? io_inputs_2 : _GEN_17; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_19 = 4'h3 == io_selects_0_1 ? io_inputs_3 : _GEN_18; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_20 = 4'h4 == io_selects_0_1 ? io_inputs_4 : _GEN_19; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_21 = 4'h5 == io_selects_0_1 ? io_inputs_5 : _GEN_20; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_22 = 4'h6 == io_selects_0_1 ? io_inputs_6 : _GEN_21; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_23 = 4'h7 == io_selects_0_1 ? io_inputs_7 : _GEN_22; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_24 = 4'h8 == io_selects_0_1 ? io_inputs_8 : _GEN_23; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_25 = 4'h9 == io_selects_0_1 ? io_inputs_9 : _GEN_24; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_26 = 4'ha == io_selects_0_1 ? io_inputs_10 : _GEN_25; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_27 = 4'hb == io_selects_0_1 ? io_inputs_11 : _GEN_26; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_28 = 4'hc == io_selects_0_1 ? io_inputs_12 : _GEN_27; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_29 = 4'hd == io_selects_0_1 ? io_inputs_13 : _GEN_28; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_30 = 4'he == io_selects_0_1 ? io_inputs_14 : _GEN_29; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_31 = 4'hf == io_selects_0_1 ? io_inputs_15 : _GEN_30; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _T_722 = _GEN_15 + _GEN_31; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _T_723 = _GEN_15 + _GEN_31; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@9.4]
  assign _T_725 = _GEN_15 * _GEN_31; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@10.4]
  assign _T_727 = _GEN_15 / _GEN_31; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@11.4]
  assign _T_728 = 3'h3 == io_operation_0; // @[Mux.scala 46:19:@12.4]
  assign _T_729 = _T_728 ? _T_727 : 64'h0; // @[Mux.scala 46:16:@13.4]
  assign _T_730 = 3'h2 == io_operation_0; // @[Mux.scala 46:19:@14.4]
  assign _T_731 = _T_730 ? _T_725 : {{64'd0}, _T_729}; // @[Mux.scala 46:16:@15.4]
  assign _T_732 = 3'h1 == io_operation_0; // @[Mux.scala 46:19:@16.4]
  assign _T_733 = _T_732 ? {{64'd0}, _T_723} : _T_731; // @[Mux.scala 46:16:@17.4]
  assign _T_734 = 3'h0 == io_operation_0; // @[Mux.scala 46:19:@18.4]
  assign _GEN_33 = 4'h1 == io_selects_1_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_34 = 4'h2 == io_selects_1_0 ? io_inputs_2 : _GEN_33; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_35 = 4'h3 == io_selects_1_0 ? io_inputs_3 : _GEN_34; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_36 = 4'h4 == io_selects_1_0 ? io_inputs_4 : _GEN_35; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_37 = 4'h5 == io_selects_1_0 ? io_inputs_5 : _GEN_36; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_38 = 4'h6 == io_selects_1_0 ? io_inputs_6 : _GEN_37; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_39 = 4'h7 == io_selects_1_0 ? io_inputs_7 : _GEN_38; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_40 = 4'h8 == io_selects_1_0 ? io_inputs_8 : _GEN_39; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_41 = 4'h9 == io_selects_1_0 ? io_inputs_9 : _GEN_40; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_42 = 4'ha == io_selects_1_0 ? io_inputs_10 : _GEN_41; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_43 = 4'hb == io_selects_1_0 ? io_inputs_11 : _GEN_42; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_44 = 4'hc == io_selects_1_0 ? io_inputs_12 : _GEN_43; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_45 = 4'hd == io_selects_1_0 ? io_inputs_13 : _GEN_44; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_46 = 4'he == io_selects_1_0 ? io_inputs_14 : _GEN_45; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_47 = 4'hf == io_selects_1_0 ? io_inputs_15 : _GEN_46; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_49 = 4'h1 == io_selects_1_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_50 = 4'h2 == io_selects_1_1 ? io_inputs_2 : _GEN_49; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_51 = 4'h3 == io_selects_1_1 ? io_inputs_3 : _GEN_50; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_52 = 4'h4 == io_selects_1_1 ? io_inputs_4 : _GEN_51; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_53 = 4'h5 == io_selects_1_1 ? io_inputs_5 : _GEN_52; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_54 = 4'h6 == io_selects_1_1 ? io_inputs_6 : _GEN_53; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_55 = 4'h7 == io_selects_1_1 ? io_inputs_7 : _GEN_54; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_56 = 4'h8 == io_selects_1_1 ? io_inputs_8 : _GEN_55; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_57 = 4'h9 == io_selects_1_1 ? io_inputs_9 : _GEN_56; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_58 = 4'ha == io_selects_1_1 ? io_inputs_10 : _GEN_57; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_59 = 4'hb == io_selects_1_1 ? io_inputs_11 : _GEN_58; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_60 = 4'hc == io_selects_1_1 ? io_inputs_12 : _GEN_59; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_61 = 4'hd == io_selects_1_1 ? io_inputs_13 : _GEN_60; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_62 = 4'he == io_selects_1_1 ? io_inputs_14 : _GEN_61; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_63 = 4'hf == io_selects_1_1 ? io_inputs_15 : _GEN_62; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _T_739 = _GEN_47 + _GEN_63; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _T_740 = _GEN_47 + _GEN_63; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@21.4]
  assign _T_742 = _GEN_47 * _GEN_63; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@22.4]
  assign _T_744 = _GEN_47 / _GEN_63; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@23.4]
  assign _T_745 = 3'h3 == io_operation_1; // @[Mux.scala 46:19:@24.4]
  assign _T_746 = _T_745 ? _T_744 : 64'h0; // @[Mux.scala 46:16:@25.4]
  assign _T_747 = 3'h2 == io_operation_1; // @[Mux.scala 46:19:@26.4]
  assign _T_748 = _T_747 ? _T_742 : {{64'd0}, _T_746}; // @[Mux.scala 46:16:@27.4]
  assign _T_749 = 3'h1 == io_operation_1; // @[Mux.scala 46:19:@28.4]
  assign _T_750 = _T_749 ? {{64'd0}, _T_740} : _T_748; // @[Mux.scala 46:16:@29.4]
  assign _T_751 = 3'h0 == io_operation_1; // @[Mux.scala 46:19:@30.4]
  assign _GEN_65 = 4'h1 == io_selects_2_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_66 = 4'h2 == io_selects_2_0 ? io_inputs_2 : _GEN_65; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_67 = 4'h3 == io_selects_2_0 ? io_inputs_3 : _GEN_66; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_68 = 4'h4 == io_selects_2_0 ? io_inputs_4 : _GEN_67; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_69 = 4'h5 == io_selects_2_0 ? io_inputs_5 : _GEN_68; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_70 = 4'h6 == io_selects_2_0 ? io_inputs_6 : _GEN_69; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_71 = 4'h7 == io_selects_2_0 ? io_inputs_7 : _GEN_70; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_72 = 4'h8 == io_selects_2_0 ? io_inputs_8 : _GEN_71; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_73 = 4'h9 == io_selects_2_0 ? io_inputs_9 : _GEN_72; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_74 = 4'ha == io_selects_2_0 ? io_inputs_10 : _GEN_73; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_75 = 4'hb == io_selects_2_0 ? io_inputs_11 : _GEN_74; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_76 = 4'hc == io_selects_2_0 ? io_inputs_12 : _GEN_75; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_77 = 4'hd == io_selects_2_0 ? io_inputs_13 : _GEN_76; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_78 = 4'he == io_selects_2_0 ? io_inputs_14 : _GEN_77; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_79 = 4'hf == io_selects_2_0 ? io_inputs_15 : _GEN_78; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_81 = 4'h1 == io_selects_2_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_82 = 4'h2 == io_selects_2_1 ? io_inputs_2 : _GEN_81; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_83 = 4'h3 == io_selects_2_1 ? io_inputs_3 : _GEN_82; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_84 = 4'h4 == io_selects_2_1 ? io_inputs_4 : _GEN_83; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_85 = 4'h5 == io_selects_2_1 ? io_inputs_5 : _GEN_84; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_86 = 4'h6 == io_selects_2_1 ? io_inputs_6 : _GEN_85; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_87 = 4'h7 == io_selects_2_1 ? io_inputs_7 : _GEN_86; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_88 = 4'h8 == io_selects_2_1 ? io_inputs_8 : _GEN_87; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_89 = 4'h9 == io_selects_2_1 ? io_inputs_9 : _GEN_88; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_90 = 4'ha == io_selects_2_1 ? io_inputs_10 : _GEN_89; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_91 = 4'hb == io_selects_2_1 ? io_inputs_11 : _GEN_90; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_92 = 4'hc == io_selects_2_1 ? io_inputs_12 : _GEN_91; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_93 = 4'hd == io_selects_2_1 ? io_inputs_13 : _GEN_92; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_94 = 4'he == io_selects_2_1 ? io_inputs_14 : _GEN_93; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_95 = 4'hf == io_selects_2_1 ? io_inputs_15 : _GEN_94; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _T_756 = _GEN_79 + _GEN_95; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _T_757 = _GEN_79 + _GEN_95; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@33.4]
  assign _T_759 = _GEN_79 * _GEN_95; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@34.4]
  assign _T_761 = _GEN_79 / _GEN_95; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@35.4]
  assign _T_762 = 3'h3 == io_operation_2; // @[Mux.scala 46:19:@36.4]
  assign _T_763 = _T_762 ? _T_761 : 64'h0; // @[Mux.scala 46:16:@37.4]
  assign _T_764 = 3'h2 == io_operation_2; // @[Mux.scala 46:19:@38.4]
  assign _T_765 = _T_764 ? _T_759 : {{64'd0}, _T_763}; // @[Mux.scala 46:16:@39.4]
  assign _T_766 = 3'h1 == io_operation_2; // @[Mux.scala 46:19:@40.4]
  assign _T_767 = _T_766 ? {{64'd0}, _T_757} : _T_765; // @[Mux.scala 46:16:@41.4]
  assign _T_768 = 3'h0 == io_operation_2; // @[Mux.scala 46:19:@42.4]
  assign _GEN_97 = 4'h1 == io_selects_3_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_98 = 4'h2 == io_selects_3_0 ? io_inputs_2 : _GEN_97; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_99 = 4'h3 == io_selects_3_0 ? io_inputs_3 : _GEN_98; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_100 = 4'h4 == io_selects_3_0 ? io_inputs_4 : _GEN_99; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_101 = 4'h5 == io_selects_3_0 ? io_inputs_5 : _GEN_100; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_102 = 4'h6 == io_selects_3_0 ? io_inputs_6 : _GEN_101; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_103 = 4'h7 == io_selects_3_0 ? io_inputs_7 : _GEN_102; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_104 = 4'h8 == io_selects_3_0 ? io_inputs_8 : _GEN_103; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_105 = 4'h9 == io_selects_3_0 ? io_inputs_9 : _GEN_104; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_106 = 4'ha == io_selects_3_0 ? io_inputs_10 : _GEN_105; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_107 = 4'hb == io_selects_3_0 ? io_inputs_11 : _GEN_106; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_108 = 4'hc == io_selects_3_0 ? io_inputs_12 : _GEN_107; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_109 = 4'hd == io_selects_3_0 ? io_inputs_13 : _GEN_108; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_110 = 4'he == io_selects_3_0 ? io_inputs_14 : _GEN_109; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_111 = 4'hf == io_selects_3_0 ? io_inputs_15 : _GEN_110; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_113 = 4'h1 == io_selects_3_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_114 = 4'h2 == io_selects_3_1 ? io_inputs_2 : _GEN_113; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_115 = 4'h3 == io_selects_3_1 ? io_inputs_3 : _GEN_114; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_116 = 4'h4 == io_selects_3_1 ? io_inputs_4 : _GEN_115; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_117 = 4'h5 == io_selects_3_1 ? io_inputs_5 : _GEN_116; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_118 = 4'h6 == io_selects_3_1 ? io_inputs_6 : _GEN_117; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_119 = 4'h7 == io_selects_3_1 ? io_inputs_7 : _GEN_118; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_120 = 4'h8 == io_selects_3_1 ? io_inputs_8 : _GEN_119; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_121 = 4'h9 == io_selects_3_1 ? io_inputs_9 : _GEN_120; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_122 = 4'ha == io_selects_3_1 ? io_inputs_10 : _GEN_121; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_123 = 4'hb == io_selects_3_1 ? io_inputs_11 : _GEN_122; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_124 = 4'hc == io_selects_3_1 ? io_inputs_12 : _GEN_123; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_125 = 4'hd == io_selects_3_1 ? io_inputs_13 : _GEN_124; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_126 = 4'he == io_selects_3_1 ? io_inputs_14 : _GEN_125; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_127 = 4'hf == io_selects_3_1 ? io_inputs_15 : _GEN_126; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _T_773 = _GEN_111 + _GEN_127; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _T_774 = _GEN_111 + _GEN_127; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@45.4]
  assign _T_776 = _GEN_111 * _GEN_127; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@46.4]
  assign _T_778 = _GEN_111 / _GEN_127; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@47.4]
  assign _T_779 = 3'h3 == io_operation_3; // @[Mux.scala 46:19:@48.4]
  assign _T_780 = _T_779 ? _T_778 : 64'h0; // @[Mux.scala 46:16:@49.4]
  assign _T_781 = 3'h2 == io_operation_3; // @[Mux.scala 46:19:@50.4]
  assign _T_782 = _T_781 ? _T_776 : {{64'd0}, _T_780}; // @[Mux.scala 46:16:@51.4]
  assign _T_783 = 3'h1 == io_operation_3; // @[Mux.scala 46:19:@52.4]
  assign _T_784 = _T_783 ? {{64'd0}, _T_774} : _T_782; // @[Mux.scala 46:16:@53.4]
  assign _T_785 = 3'h0 == io_operation_3; // @[Mux.scala 46:19:@54.4]
  assign _GEN_129 = 4'h1 == io_selects_4_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_130 = 4'h2 == io_selects_4_0 ? io_inputs_2 : _GEN_129; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_131 = 4'h3 == io_selects_4_0 ? io_inputs_3 : _GEN_130; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_132 = 4'h4 == io_selects_4_0 ? io_inputs_4 : _GEN_131; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_133 = 4'h5 == io_selects_4_0 ? io_inputs_5 : _GEN_132; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_134 = 4'h6 == io_selects_4_0 ? io_inputs_6 : _GEN_133; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_135 = 4'h7 == io_selects_4_0 ? io_inputs_7 : _GEN_134; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_136 = 4'h8 == io_selects_4_0 ? io_inputs_8 : _GEN_135; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_137 = 4'h9 == io_selects_4_0 ? io_inputs_9 : _GEN_136; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_138 = 4'ha == io_selects_4_0 ? io_inputs_10 : _GEN_137; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_139 = 4'hb == io_selects_4_0 ? io_inputs_11 : _GEN_138; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_140 = 4'hc == io_selects_4_0 ? io_inputs_12 : _GEN_139; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_141 = 4'hd == io_selects_4_0 ? io_inputs_13 : _GEN_140; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_142 = 4'he == io_selects_4_0 ? io_inputs_14 : _GEN_141; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_143 = 4'hf == io_selects_4_0 ? io_inputs_15 : _GEN_142; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_145 = 4'h1 == io_selects_4_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_146 = 4'h2 == io_selects_4_1 ? io_inputs_2 : _GEN_145; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_147 = 4'h3 == io_selects_4_1 ? io_inputs_3 : _GEN_146; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_148 = 4'h4 == io_selects_4_1 ? io_inputs_4 : _GEN_147; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_149 = 4'h5 == io_selects_4_1 ? io_inputs_5 : _GEN_148; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_150 = 4'h6 == io_selects_4_1 ? io_inputs_6 : _GEN_149; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_151 = 4'h7 == io_selects_4_1 ? io_inputs_7 : _GEN_150; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_152 = 4'h8 == io_selects_4_1 ? io_inputs_8 : _GEN_151; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_153 = 4'h9 == io_selects_4_1 ? io_inputs_9 : _GEN_152; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_154 = 4'ha == io_selects_4_1 ? io_inputs_10 : _GEN_153; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_155 = 4'hb == io_selects_4_1 ? io_inputs_11 : _GEN_154; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_156 = 4'hc == io_selects_4_1 ? io_inputs_12 : _GEN_155; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_157 = 4'hd == io_selects_4_1 ? io_inputs_13 : _GEN_156; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_158 = 4'he == io_selects_4_1 ? io_inputs_14 : _GEN_157; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_159 = 4'hf == io_selects_4_1 ? io_inputs_15 : _GEN_158; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _T_790 = _GEN_143 + _GEN_159; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _T_791 = _GEN_143 + _GEN_159; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@57.4]
  assign _T_793 = _GEN_143 * _GEN_159; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@58.4]
  assign _T_795 = _GEN_143 / _GEN_159; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@59.4]
  assign _T_796 = 3'h3 == io_operation_4; // @[Mux.scala 46:19:@60.4]
  assign _T_797 = _T_796 ? _T_795 : 64'h0; // @[Mux.scala 46:16:@61.4]
  assign _T_798 = 3'h2 == io_operation_4; // @[Mux.scala 46:19:@62.4]
  assign _T_799 = _T_798 ? _T_793 : {{64'd0}, _T_797}; // @[Mux.scala 46:16:@63.4]
  assign _T_800 = 3'h1 == io_operation_4; // @[Mux.scala 46:19:@64.4]
  assign _T_801 = _T_800 ? {{64'd0}, _T_791} : _T_799; // @[Mux.scala 46:16:@65.4]
  assign _T_802 = 3'h0 == io_operation_4; // @[Mux.scala 46:19:@66.4]
  assign _GEN_161 = 4'h1 == io_selects_5_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_162 = 4'h2 == io_selects_5_0 ? io_inputs_2 : _GEN_161; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_163 = 4'h3 == io_selects_5_0 ? io_inputs_3 : _GEN_162; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_164 = 4'h4 == io_selects_5_0 ? io_inputs_4 : _GEN_163; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_165 = 4'h5 == io_selects_5_0 ? io_inputs_5 : _GEN_164; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_166 = 4'h6 == io_selects_5_0 ? io_inputs_6 : _GEN_165; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_167 = 4'h7 == io_selects_5_0 ? io_inputs_7 : _GEN_166; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_168 = 4'h8 == io_selects_5_0 ? io_inputs_8 : _GEN_167; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_169 = 4'h9 == io_selects_5_0 ? io_inputs_9 : _GEN_168; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_170 = 4'ha == io_selects_5_0 ? io_inputs_10 : _GEN_169; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_171 = 4'hb == io_selects_5_0 ? io_inputs_11 : _GEN_170; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_172 = 4'hc == io_selects_5_0 ? io_inputs_12 : _GEN_171; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_173 = 4'hd == io_selects_5_0 ? io_inputs_13 : _GEN_172; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_174 = 4'he == io_selects_5_0 ? io_inputs_14 : _GEN_173; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_175 = 4'hf == io_selects_5_0 ? io_inputs_15 : _GEN_174; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_177 = 4'h1 == io_selects_5_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_178 = 4'h2 == io_selects_5_1 ? io_inputs_2 : _GEN_177; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_179 = 4'h3 == io_selects_5_1 ? io_inputs_3 : _GEN_178; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_180 = 4'h4 == io_selects_5_1 ? io_inputs_4 : _GEN_179; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_181 = 4'h5 == io_selects_5_1 ? io_inputs_5 : _GEN_180; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_182 = 4'h6 == io_selects_5_1 ? io_inputs_6 : _GEN_181; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_183 = 4'h7 == io_selects_5_1 ? io_inputs_7 : _GEN_182; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_184 = 4'h8 == io_selects_5_1 ? io_inputs_8 : _GEN_183; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_185 = 4'h9 == io_selects_5_1 ? io_inputs_9 : _GEN_184; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_186 = 4'ha == io_selects_5_1 ? io_inputs_10 : _GEN_185; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_187 = 4'hb == io_selects_5_1 ? io_inputs_11 : _GEN_186; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_188 = 4'hc == io_selects_5_1 ? io_inputs_12 : _GEN_187; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_189 = 4'hd == io_selects_5_1 ? io_inputs_13 : _GEN_188; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_190 = 4'he == io_selects_5_1 ? io_inputs_14 : _GEN_189; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_191 = 4'hf == io_selects_5_1 ? io_inputs_15 : _GEN_190; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _T_807 = _GEN_175 + _GEN_191; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _T_808 = _GEN_175 + _GEN_191; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@69.4]
  assign _T_810 = _GEN_175 * _GEN_191; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@70.4]
  assign _T_812 = _GEN_175 / _GEN_191; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@71.4]
  assign _T_813 = 3'h3 == io_operation_5; // @[Mux.scala 46:19:@72.4]
  assign _T_814 = _T_813 ? _T_812 : 64'h0; // @[Mux.scala 46:16:@73.4]
  assign _T_815 = 3'h2 == io_operation_5; // @[Mux.scala 46:19:@74.4]
  assign _T_816 = _T_815 ? _T_810 : {{64'd0}, _T_814}; // @[Mux.scala 46:16:@75.4]
  assign _T_817 = 3'h1 == io_operation_5; // @[Mux.scala 46:19:@76.4]
  assign _T_818 = _T_817 ? {{64'd0}, _T_808} : _T_816; // @[Mux.scala 46:16:@77.4]
  assign _T_819 = 3'h0 == io_operation_5; // @[Mux.scala 46:19:@78.4]
  assign _GEN_193 = 4'h1 == io_selects_6_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_194 = 4'h2 == io_selects_6_0 ? io_inputs_2 : _GEN_193; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_195 = 4'h3 == io_selects_6_0 ? io_inputs_3 : _GEN_194; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_196 = 4'h4 == io_selects_6_0 ? io_inputs_4 : _GEN_195; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_197 = 4'h5 == io_selects_6_0 ? io_inputs_5 : _GEN_196; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_198 = 4'h6 == io_selects_6_0 ? io_inputs_6 : _GEN_197; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_199 = 4'h7 == io_selects_6_0 ? io_inputs_7 : _GEN_198; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_200 = 4'h8 == io_selects_6_0 ? io_inputs_8 : _GEN_199; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_201 = 4'h9 == io_selects_6_0 ? io_inputs_9 : _GEN_200; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_202 = 4'ha == io_selects_6_0 ? io_inputs_10 : _GEN_201; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_203 = 4'hb == io_selects_6_0 ? io_inputs_11 : _GEN_202; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_204 = 4'hc == io_selects_6_0 ? io_inputs_12 : _GEN_203; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_205 = 4'hd == io_selects_6_0 ? io_inputs_13 : _GEN_204; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_206 = 4'he == io_selects_6_0 ? io_inputs_14 : _GEN_205; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_207 = 4'hf == io_selects_6_0 ? io_inputs_15 : _GEN_206; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_209 = 4'h1 == io_selects_6_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_210 = 4'h2 == io_selects_6_1 ? io_inputs_2 : _GEN_209; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_211 = 4'h3 == io_selects_6_1 ? io_inputs_3 : _GEN_210; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_212 = 4'h4 == io_selects_6_1 ? io_inputs_4 : _GEN_211; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_213 = 4'h5 == io_selects_6_1 ? io_inputs_5 : _GEN_212; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_214 = 4'h6 == io_selects_6_1 ? io_inputs_6 : _GEN_213; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_215 = 4'h7 == io_selects_6_1 ? io_inputs_7 : _GEN_214; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_216 = 4'h8 == io_selects_6_1 ? io_inputs_8 : _GEN_215; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_217 = 4'h9 == io_selects_6_1 ? io_inputs_9 : _GEN_216; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_218 = 4'ha == io_selects_6_1 ? io_inputs_10 : _GEN_217; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_219 = 4'hb == io_selects_6_1 ? io_inputs_11 : _GEN_218; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_220 = 4'hc == io_selects_6_1 ? io_inputs_12 : _GEN_219; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_221 = 4'hd == io_selects_6_1 ? io_inputs_13 : _GEN_220; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_222 = 4'he == io_selects_6_1 ? io_inputs_14 : _GEN_221; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_223 = 4'hf == io_selects_6_1 ? io_inputs_15 : _GEN_222; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _T_824 = _GEN_207 + _GEN_223; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _T_825 = _GEN_207 + _GEN_223; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@81.4]
  assign _T_827 = _GEN_207 * _GEN_223; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@82.4]
  assign _T_829 = _GEN_207 / _GEN_223; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@83.4]
  assign _T_830 = 3'h3 == io_operation_6; // @[Mux.scala 46:19:@84.4]
  assign _T_831 = _T_830 ? _T_829 : 64'h0; // @[Mux.scala 46:16:@85.4]
  assign _T_832 = 3'h2 == io_operation_6; // @[Mux.scala 46:19:@86.4]
  assign _T_833 = _T_832 ? _T_827 : {{64'd0}, _T_831}; // @[Mux.scala 46:16:@87.4]
  assign _T_834 = 3'h1 == io_operation_6; // @[Mux.scala 46:19:@88.4]
  assign _T_835 = _T_834 ? {{64'd0}, _T_825} : _T_833; // @[Mux.scala 46:16:@89.4]
  assign _T_836 = 3'h0 == io_operation_6; // @[Mux.scala 46:19:@90.4]
  assign _GEN_225 = 4'h1 == io_selects_7_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_226 = 4'h2 == io_selects_7_0 ? io_inputs_2 : _GEN_225; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_227 = 4'h3 == io_selects_7_0 ? io_inputs_3 : _GEN_226; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_228 = 4'h4 == io_selects_7_0 ? io_inputs_4 : _GEN_227; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_229 = 4'h5 == io_selects_7_0 ? io_inputs_5 : _GEN_228; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_230 = 4'h6 == io_selects_7_0 ? io_inputs_6 : _GEN_229; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_231 = 4'h7 == io_selects_7_0 ? io_inputs_7 : _GEN_230; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_232 = 4'h8 == io_selects_7_0 ? io_inputs_8 : _GEN_231; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_233 = 4'h9 == io_selects_7_0 ? io_inputs_9 : _GEN_232; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_234 = 4'ha == io_selects_7_0 ? io_inputs_10 : _GEN_233; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_235 = 4'hb == io_selects_7_0 ? io_inputs_11 : _GEN_234; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_236 = 4'hc == io_selects_7_0 ? io_inputs_12 : _GEN_235; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_237 = 4'hd == io_selects_7_0 ? io_inputs_13 : _GEN_236; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_238 = 4'he == io_selects_7_0 ? io_inputs_14 : _GEN_237; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_239 = 4'hf == io_selects_7_0 ? io_inputs_15 : _GEN_238; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_241 = 4'h1 == io_selects_7_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_242 = 4'h2 == io_selects_7_1 ? io_inputs_2 : _GEN_241; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_243 = 4'h3 == io_selects_7_1 ? io_inputs_3 : _GEN_242; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_244 = 4'h4 == io_selects_7_1 ? io_inputs_4 : _GEN_243; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_245 = 4'h5 == io_selects_7_1 ? io_inputs_5 : _GEN_244; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_246 = 4'h6 == io_selects_7_1 ? io_inputs_6 : _GEN_245; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_247 = 4'h7 == io_selects_7_1 ? io_inputs_7 : _GEN_246; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_248 = 4'h8 == io_selects_7_1 ? io_inputs_8 : _GEN_247; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_249 = 4'h9 == io_selects_7_1 ? io_inputs_9 : _GEN_248; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_250 = 4'ha == io_selects_7_1 ? io_inputs_10 : _GEN_249; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_251 = 4'hb == io_selects_7_1 ? io_inputs_11 : _GEN_250; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_252 = 4'hc == io_selects_7_1 ? io_inputs_12 : _GEN_251; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_253 = 4'hd == io_selects_7_1 ? io_inputs_13 : _GEN_252; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_254 = 4'he == io_selects_7_1 ? io_inputs_14 : _GEN_253; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_255 = 4'hf == io_selects_7_1 ? io_inputs_15 : _GEN_254; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _T_841 = _GEN_239 + _GEN_255; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _T_842 = _GEN_239 + _GEN_255; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@93.4]
  assign _T_844 = _GEN_239 * _GEN_255; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@94.4]
  assign _T_846 = _GEN_239 / _GEN_255; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@95.4]
  assign _T_847 = 3'h3 == io_operation_7; // @[Mux.scala 46:19:@96.4]
  assign _T_848 = _T_847 ? _T_846 : 64'h0; // @[Mux.scala 46:16:@97.4]
  assign _T_849 = 3'h2 == io_operation_7; // @[Mux.scala 46:19:@98.4]
  assign _T_850 = _T_849 ? _T_844 : {{64'd0}, _T_848}; // @[Mux.scala 46:16:@99.4]
  assign _T_851 = 3'h1 == io_operation_7; // @[Mux.scala 46:19:@100.4]
  assign _T_852 = _T_851 ? {{64'd0}, _T_842} : _T_850; // @[Mux.scala 46:16:@101.4]
  assign _T_853 = 3'h0 == io_operation_7; // @[Mux.scala 46:19:@102.4]
  assign _GEN_257 = 4'h1 == io_selects_8_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_258 = 4'h2 == io_selects_8_0 ? io_inputs_2 : _GEN_257; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_259 = 4'h3 == io_selects_8_0 ? io_inputs_3 : _GEN_258; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_260 = 4'h4 == io_selects_8_0 ? io_inputs_4 : _GEN_259; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_261 = 4'h5 == io_selects_8_0 ? io_inputs_5 : _GEN_260; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_262 = 4'h6 == io_selects_8_0 ? io_inputs_6 : _GEN_261; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_263 = 4'h7 == io_selects_8_0 ? io_inputs_7 : _GEN_262; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_264 = 4'h8 == io_selects_8_0 ? io_inputs_8 : _GEN_263; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_265 = 4'h9 == io_selects_8_0 ? io_inputs_9 : _GEN_264; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_266 = 4'ha == io_selects_8_0 ? io_inputs_10 : _GEN_265; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_267 = 4'hb == io_selects_8_0 ? io_inputs_11 : _GEN_266; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_268 = 4'hc == io_selects_8_0 ? io_inputs_12 : _GEN_267; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_269 = 4'hd == io_selects_8_0 ? io_inputs_13 : _GEN_268; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_270 = 4'he == io_selects_8_0 ? io_inputs_14 : _GEN_269; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_271 = 4'hf == io_selects_8_0 ? io_inputs_15 : _GEN_270; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_273 = 4'h1 == io_selects_8_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_274 = 4'h2 == io_selects_8_1 ? io_inputs_2 : _GEN_273; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_275 = 4'h3 == io_selects_8_1 ? io_inputs_3 : _GEN_274; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_276 = 4'h4 == io_selects_8_1 ? io_inputs_4 : _GEN_275; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_277 = 4'h5 == io_selects_8_1 ? io_inputs_5 : _GEN_276; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_278 = 4'h6 == io_selects_8_1 ? io_inputs_6 : _GEN_277; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_279 = 4'h7 == io_selects_8_1 ? io_inputs_7 : _GEN_278; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_280 = 4'h8 == io_selects_8_1 ? io_inputs_8 : _GEN_279; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_281 = 4'h9 == io_selects_8_1 ? io_inputs_9 : _GEN_280; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_282 = 4'ha == io_selects_8_1 ? io_inputs_10 : _GEN_281; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_283 = 4'hb == io_selects_8_1 ? io_inputs_11 : _GEN_282; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_284 = 4'hc == io_selects_8_1 ? io_inputs_12 : _GEN_283; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_285 = 4'hd == io_selects_8_1 ? io_inputs_13 : _GEN_284; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_286 = 4'he == io_selects_8_1 ? io_inputs_14 : _GEN_285; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_287 = 4'hf == io_selects_8_1 ? io_inputs_15 : _GEN_286; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _T_858 = _GEN_271 + _GEN_287; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _T_859 = _GEN_271 + _GEN_287; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@105.4]
  assign _T_861 = _GEN_271 * _GEN_287; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@106.4]
  assign _T_863 = _GEN_271 / _GEN_287; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@107.4]
  assign _T_864 = 3'h3 == io_operation_8; // @[Mux.scala 46:19:@108.4]
  assign _T_865 = _T_864 ? _T_863 : 64'h0; // @[Mux.scala 46:16:@109.4]
  assign _T_866 = 3'h2 == io_operation_8; // @[Mux.scala 46:19:@110.4]
  assign _T_867 = _T_866 ? _T_861 : {{64'd0}, _T_865}; // @[Mux.scala 46:16:@111.4]
  assign _T_868 = 3'h1 == io_operation_8; // @[Mux.scala 46:19:@112.4]
  assign _T_869 = _T_868 ? {{64'd0}, _T_859} : _T_867; // @[Mux.scala 46:16:@113.4]
  assign _T_870 = 3'h0 == io_operation_8; // @[Mux.scala 46:19:@114.4]
  assign _GEN_289 = 4'h1 == io_selects_9_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_290 = 4'h2 == io_selects_9_0 ? io_inputs_2 : _GEN_289; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_291 = 4'h3 == io_selects_9_0 ? io_inputs_3 : _GEN_290; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_292 = 4'h4 == io_selects_9_0 ? io_inputs_4 : _GEN_291; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_293 = 4'h5 == io_selects_9_0 ? io_inputs_5 : _GEN_292; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_294 = 4'h6 == io_selects_9_0 ? io_inputs_6 : _GEN_293; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_295 = 4'h7 == io_selects_9_0 ? io_inputs_7 : _GEN_294; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_296 = 4'h8 == io_selects_9_0 ? io_inputs_8 : _GEN_295; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_297 = 4'h9 == io_selects_9_0 ? io_inputs_9 : _GEN_296; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_298 = 4'ha == io_selects_9_0 ? io_inputs_10 : _GEN_297; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_299 = 4'hb == io_selects_9_0 ? io_inputs_11 : _GEN_298; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_300 = 4'hc == io_selects_9_0 ? io_inputs_12 : _GEN_299; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_301 = 4'hd == io_selects_9_0 ? io_inputs_13 : _GEN_300; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_302 = 4'he == io_selects_9_0 ? io_inputs_14 : _GEN_301; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_303 = 4'hf == io_selects_9_0 ? io_inputs_15 : _GEN_302; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_305 = 4'h1 == io_selects_9_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_306 = 4'h2 == io_selects_9_1 ? io_inputs_2 : _GEN_305; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_307 = 4'h3 == io_selects_9_1 ? io_inputs_3 : _GEN_306; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_308 = 4'h4 == io_selects_9_1 ? io_inputs_4 : _GEN_307; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_309 = 4'h5 == io_selects_9_1 ? io_inputs_5 : _GEN_308; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_310 = 4'h6 == io_selects_9_1 ? io_inputs_6 : _GEN_309; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_311 = 4'h7 == io_selects_9_1 ? io_inputs_7 : _GEN_310; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_312 = 4'h8 == io_selects_9_1 ? io_inputs_8 : _GEN_311; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_313 = 4'h9 == io_selects_9_1 ? io_inputs_9 : _GEN_312; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_314 = 4'ha == io_selects_9_1 ? io_inputs_10 : _GEN_313; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_315 = 4'hb == io_selects_9_1 ? io_inputs_11 : _GEN_314; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_316 = 4'hc == io_selects_9_1 ? io_inputs_12 : _GEN_315; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_317 = 4'hd == io_selects_9_1 ? io_inputs_13 : _GEN_316; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_318 = 4'he == io_selects_9_1 ? io_inputs_14 : _GEN_317; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_319 = 4'hf == io_selects_9_1 ? io_inputs_15 : _GEN_318; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _T_875 = _GEN_303 + _GEN_319; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _T_876 = _GEN_303 + _GEN_319; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@117.4]
  assign _T_878 = _GEN_303 * _GEN_319; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@118.4]
  assign _T_880 = _GEN_303 / _GEN_319; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@119.4]
  assign _T_881 = 3'h3 == io_operation_9; // @[Mux.scala 46:19:@120.4]
  assign _T_882 = _T_881 ? _T_880 : 64'h0; // @[Mux.scala 46:16:@121.4]
  assign _T_883 = 3'h2 == io_operation_9; // @[Mux.scala 46:19:@122.4]
  assign _T_884 = _T_883 ? _T_878 : {{64'd0}, _T_882}; // @[Mux.scala 46:16:@123.4]
  assign _T_885 = 3'h1 == io_operation_9; // @[Mux.scala 46:19:@124.4]
  assign _T_886 = _T_885 ? {{64'd0}, _T_876} : _T_884; // @[Mux.scala 46:16:@125.4]
  assign _T_887 = 3'h0 == io_operation_9; // @[Mux.scala 46:19:@126.4]
  assign _GEN_321 = 4'h1 == io_selects_10_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_322 = 4'h2 == io_selects_10_0 ? io_inputs_2 : _GEN_321; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_323 = 4'h3 == io_selects_10_0 ? io_inputs_3 : _GEN_322; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_324 = 4'h4 == io_selects_10_0 ? io_inputs_4 : _GEN_323; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_325 = 4'h5 == io_selects_10_0 ? io_inputs_5 : _GEN_324; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_326 = 4'h6 == io_selects_10_0 ? io_inputs_6 : _GEN_325; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_327 = 4'h7 == io_selects_10_0 ? io_inputs_7 : _GEN_326; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_328 = 4'h8 == io_selects_10_0 ? io_inputs_8 : _GEN_327; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_329 = 4'h9 == io_selects_10_0 ? io_inputs_9 : _GEN_328; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_330 = 4'ha == io_selects_10_0 ? io_inputs_10 : _GEN_329; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_331 = 4'hb == io_selects_10_0 ? io_inputs_11 : _GEN_330; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_332 = 4'hc == io_selects_10_0 ? io_inputs_12 : _GEN_331; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_333 = 4'hd == io_selects_10_0 ? io_inputs_13 : _GEN_332; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_334 = 4'he == io_selects_10_0 ? io_inputs_14 : _GEN_333; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_335 = 4'hf == io_selects_10_0 ? io_inputs_15 : _GEN_334; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_337 = 4'h1 == io_selects_10_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_338 = 4'h2 == io_selects_10_1 ? io_inputs_2 : _GEN_337; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_339 = 4'h3 == io_selects_10_1 ? io_inputs_3 : _GEN_338; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_340 = 4'h4 == io_selects_10_1 ? io_inputs_4 : _GEN_339; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_341 = 4'h5 == io_selects_10_1 ? io_inputs_5 : _GEN_340; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_342 = 4'h6 == io_selects_10_1 ? io_inputs_6 : _GEN_341; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_343 = 4'h7 == io_selects_10_1 ? io_inputs_7 : _GEN_342; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_344 = 4'h8 == io_selects_10_1 ? io_inputs_8 : _GEN_343; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_345 = 4'h9 == io_selects_10_1 ? io_inputs_9 : _GEN_344; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_346 = 4'ha == io_selects_10_1 ? io_inputs_10 : _GEN_345; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_347 = 4'hb == io_selects_10_1 ? io_inputs_11 : _GEN_346; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_348 = 4'hc == io_selects_10_1 ? io_inputs_12 : _GEN_347; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_349 = 4'hd == io_selects_10_1 ? io_inputs_13 : _GEN_348; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_350 = 4'he == io_selects_10_1 ? io_inputs_14 : _GEN_349; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_351 = 4'hf == io_selects_10_1 ? io_inputs_15 : _GEN_350; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _T_892 = _GEN_335 + _GEN_351; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _T_893 = _GEN_335 + _GEN_351; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@129.4]
  assign _T_895 = _GEN_335 * _GEN_351; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@130.4]
  assign _T_897 = _GEN_335 / _GEN_351; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@131.4]
  assign _T_898 = 3'h3 == io_operation_10; // @[Mux.scala 46:19:@132.4]
  assign _T_899 = _T_898 ? _T_897 : 64'h0; // @[Mux.scala 46:16:@133.4]
  assign _T_900 = 3'h2 == io_operation_10; // @[Mux.scala 46:19:@134.4]
  assign _T_901 = _T_900 ? _T_895 : {{64'd0}, _T_899}; // @[Mux.scala 46:16:@135.4]
  assign _T_902 = 3'h1 == io_operation_10; // @[Mux.scala 46:19:@136.4]
  assign _T_903 = _T_902 ? {{64'd0}, _T_893} : _T_901; // @[Mux.scala 46:16:@137.4]
  assign _T_904 = 3'h0 == io_operation_10; // @[Mux.scala 46:19:@138.4]
  assign _GEN_353 = 4'h1 == io_selects_11_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_354 = 4'h2 == io_selects_11_0 ? io_inputs_2 : _GEN_353; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_355 = 4'h3 == io_selects_11_0 ? io_inputs_3 : _GEN_354; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_356 = 4'h4 == io_selects_11_0 ? io_inputs_4 : _GEN_355; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_357 = 4'h5 == io_selects_11_0 ? io_inputs_5 : _GEN_356; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_358 = 4'h6 == io_selects_11_0 ? io_inputs_6 : _GEN_357; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_359 = 4'h7 == io_selects_11_0 ? io_inputs_7 : _GEN_358; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_360 = 4'h8 == io_selects_11_0 ? io_inputs_8 : _GEN_359; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_361 = 4'h9 == io_selects_11_0 ? io_inputs_9 : _GEN_360; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_362 = 4'ha == io_selects_11_0 ? io_inputs_10 : _GEN_361; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_363 = 4'hb == io_selects_11_0 ? io_inputs_11 : _GEN_362; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_364 = 4'hc == io_selects_11_0 ? io_inputs_12 : _GEN_363; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_365 = 4'hd == io_selects_11_0 ? io_inputs_13 : _GEN_364; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_366 = 4'he == io_selects_11_0 ? io_inputs_14 : _GEN_365; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_367 = 4'hf == io_selects_11_0 ? io_inputs_15 : _GEN_366; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_369 = 4'h1 == io_selects_11_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_370 = 4'h2 == io_selects_11_1 ? io_inputs_2 : _GEN_369; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_371 = 4'h3 == io_selects_11_1 ? io_inputs_3 : _GEN_370; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_372 = 4'h4 == io_selects_11_1 ? io_inputs_4 : _GEN_371; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_373 = 4'h5 == io_selects_11_1 ? io_inputs_5 : _GEN_372; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_374 = 4'h6 == io_selects_11_1 ? io_inputs_6 : _GEN_373; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_375 = 4'h7 == io_selects_11_1 ? io_inputs_7 : _GEN_374; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_376 = 4'h8 == io_selects_11_1 ? io_inputs_8 : _GEN_375; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_377 = 4'h9 == io_selects_11_1 ? io_inputs_9 : _GEN_376; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_378 = 4'ha == io_selects_11_1 ? io_inputs_10 : _GEN_377; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_379 = 4'hb == io_selects_11_1 ? io_inputs_11 : _GEN_378; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_380 = 4'hc == io_selects_11_1 ? io_inputs_12 : _GEN_379; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_381 = 4'hd == io_selects_11_1 ? io_inputs_13 : _GEN_380; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_382 = 4'he == io_selects_11_1 ? io_inputs_14 : _GEN_381; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_383 = 4'hf == io_selects_11_1 ? io_inputs_15 : _GEN_382; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _T_909 = _GEN_367 + _GEN_383; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _T_910 = _GEN_367 + _GEN_383; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@141.4]
  assign _T_912 = _GEN_367 * _GEN_383; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@142.4]
  assign _T_914 = _GEN_367 / _GEN_383; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@143.4]
  assign _T_915 = 3'h3 == io_operation_11; // @[Mux.scala 46:19:@144.4]
  assign _T_916 = _T_915 ? _T_914 : 64'h0; // @[Mux.scala 46:16:@145.4]
  assign _T_917 = 3'h2 == io_operation_11; // @[Mux.scala 46:19:@146.4]
  assign _T_918 = _T_917 ? _T_912 : {{64'd0}, _T_916}; // @[Mux.scala 46:16:@147.4]
  assign _T_919 = 3'h1 == io_operation_11; // @[Mux.scala 46:19:@148.4]
  assign _T_920 = _T_919 ? {{64'd0}, _T_910} : _T_918; // @[Mux.scala 46:16:@149.4]
  assign _T_921 = 3'h0 == io_operation_11; // @[Mux.scala 46:19:@150.4]
  assign _GEN_385 = 4'h1 == io_selects_12_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_386 = 4'h2 == io_selects_12_0 ? io_inputs_2 : _GEN_385; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_387 = 4'h3 == io_selects_12_0 ? io_inputs_3 : _GEN_386; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_388 = 4'h4 == io_selects_12_0 ? io_inputs_4 : _GEN_387; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_389 = 4'h5 == io_selects_12_0 ? io_inputs_5 : _GEN_388; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_390 = 4'h6 == io_selects_12_0 ? io_inputs_6 : _GEN_389; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_391 = 4'h7 == io_selects_12_0 ? io_inputs_7 : _GEN_390; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_392 = 4'h8 == io_selects_12_0 ? io_inputs_8 : _GEN_391; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_393 = 4'h9 == io_selects_12_0 ? io_inputs_9 : _GEN_392; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_394 = 4'ha == io_selects_12_0 ? io_inputs_10 : _GEN_393; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_395 = 4'hb == io_selects_12_0 ? io_inputs_11 : _GEN_394; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_396 = 4'hc == io_selects_12_0 ? io_inputs_12 : _GEN_395; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_397 = 4'hd == io_selects_12_0 ? io_inputs_13 : _GEN_396; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_398 = 4'he == io_selects_12_0 ? io_inputs_14 : _GEN_397; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_399 = 4'hf == io_selects_12_0 ? io_inputs_15 : _GEN_398; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_401 = 4'h1 == io_selects_12_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_402 = 4'h2 == io_selects_12_1 ? io_inputs_2 : _GEN_401; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_403 = 4'h3 == io_selects_12_1 ? io_inputs_3 : _GEN_402; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_404 = 4'h4 == io_selects_12_1 ? io_inputs_4 : _GEN_403; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_405 = 4'h5 == io_selects_12_1 ? io_inputs_5 : _GEN_404; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_406 = 4'h6 == io_selects_12_1 ? io_inputs_6 : _GEN_405; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_407 = 4'h7 == io_selects_12_1 ? io_inputs_7 : _GEN_406; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_408 = 4'h8 == io_selects_12_1 ? io_inputs_8 : _GEN_407; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_409 = 4'h9 == io_selects_12_1 ? io_inputs_9 : _GEN_408; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_410 = 4'ha == io_selects_12_1 ? io_inputs_10 : _GEN_409; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_411 = 4'hb == io_selects_12_1 ? io_inputs_11 : _GEN_410; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_412 = 4'hc == io_selects_12_1 ? io_inputs_12 : _GEN_411; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_413 = 4'hd == io_selects_12_1 ? io_inputs_13 : _GEN_412; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_414 = 4'he == io_selects_12_1 ? io_inputs_14 : _GEN_413; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_415 = 4'hf == io_selects_12_1 ? io_inputs_15 : _GEN_414; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _T_926 = _GEN_399 + _GEN_415; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _T_927 = _GEN_399 + _GEN_415; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@153.4]
  assign _T_929 = _GEN_399 * _GEN_415; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@154.4]
  assign _T_931 = _GEN_399 / _GEN_415; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@155.4]
  assign _T_932 = 3'h3 == io_operation_12; // @[Mux.scala 46:19:@156.4]
  assign _T_933 = _T_932 ? _T_931 : 64'h0; // @[Mux.scala 46:16:@157.4]
  assign _T_934 = 3'h2 == io_operation_12; // @[Mux.scala 46:19:@158.4]
  assign _T_935 = _T_934 ? _T_929 : {{64'd0}, _T_933}; // @[Mux.scala 46:16:@159.4]
  assign _T_936 = 3'h1 == io_operation_12; // @[Mux.scala 46:19:@160.4]
  assign _T_937 = _T_936 ? {{64'd0}, _T_927} : _T_935; // @[Mux.scala 46:16:@161.4]
  assign _T_938 = 3'h0 == io_operation_12; // @[Mux.scala 46:19:@162.4]
  assign _GEN_417 = 4'h1 == io_selects_13_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_418 = 4'h2 == io_selects_13_0 ? io_inputs_2 : _GEN_417; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_419 = 4'h3 == io_selects_13_0 ? io_inputs_3 : _GEN_418; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_420 = 4'h4 == io_selects_13_0 ? io_inputs_4 : _GEN_419; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_421 = 4'h5 == io_selects_13_0 ? io_inputs_5 : _GEN_420; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_422 = 4'h6 == io_selects_13_0 ? io_inputs_6 : _GEN_421; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_423 = 4'h7 == io_selects_13_0 ? io_inputs_7 : _GEN_422; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_424 = 4'h8 == io_selects_13_0 ? io_inputs_8 : _GEN_423; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_425 = 4'h9 == io_selects_13_0 ? io_inputs_9 : _GEN_424; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_426 = 4'ha == io_selects_13_0 ? io_inputs_10 : _GEN_425; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_427 = 4'hb == io_selects_13_0 ? io_inputs_11 : _GEN_426; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_428 = 4'hc == io_selects_13_0 ? io_inputs_12 : _GEN_427; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_429 = 4'hd == io_selects_13_0 ? io_inputs_13 : _GEN_428; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_430 = 4'he == io_selects_13_0 ? io_inputs_14 : _GEN_429; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_431 = 4'hf == io_selects_13_0 ? io_inputs_15 : _GEN_430; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_433 = 4'h1 == io_selects_13_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_434 = 4'h2 == io_selects_13_1 ? io_inputs_2 : _GEN_433; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_435 = 4'h3 == io_selects_13_1 ? io_inputs_3 : _GEN_434; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_436 = 4'h4 == io_selects_13_1 ? io_inputs_4 : _GEN_435; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_437 = 4'h5 == io_selects_13_1 ? io_inputs_5 : _GEN_436; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_438 = 4'h6 == io_selects_13_1 ? io_inputs_6 : _GEN_437; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_439 = 4'h7 == io_selects_13_1 ? io_inputs_7 : _GEN_438; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_440 = 4'h8 == io_selects_13_1 ? io_inputs_8 : _GEN_439; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_441 = 4'h9 == io_selects_13_1 ? io_inputs_9 : _GEN_440; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_442 = 4'ha == io_selects_13_1 ? io_inputs_10 : _GEN_441; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_443 = 4'hb == io_selects_13_1 ? io_inputs_11 : _GEN_442; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_444 = 4'hc == io_selects_13_1 ? io_inputs_12 : _GEN_443; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_445 = 4'hd == io_selects_13_1 ? io_inputs_13 : _GEN_444; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_446 = 4'he == io_selects_13_1 ? io_inputs_14 : _GEN_445; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_447 = 4'hf == io_selects_13_1 ? io_inputs_15 : _GEN_446; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _T_943 = _GEN_431 + _GEN_447; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _T_944 = _GEN_431 + _GEN_447; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@165.4]
  assign _T_946 = _GEN_431 * _GEN_447; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@166.4]
  assign _T_948 = _GEN_431 / _GEN_447; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@167.4]
  assign _T_949 = 3'h3 == io_operation_13; // @[Mux.scala 46:19:@168.4]
  assign _T_950 = _T_949 ? _T_948 : 64'h0; // @[Mux.scala 46:16:@169.4]
  assign _T_951 = 3'h2 == io_operation_13; // @[Mux.scala 46:19:@170.4]
  assign _T_952 = _T_951 ? _T_946 : {{64'd0}, _T_950}; // @[Mux.scala 46:16:@171.4]
  assign _T_953 = 3'h1 == io_operation_13; // @[Mux.scala 46:19:@172.4]
  assign _T_954 = _T_953 ? {{64'd0}, _T_944} : _T_952; // @[Mux.scala 46:16:@173.4]
  assign _T_955 = 3'h0 == io_operation_13; // @[Mux.scala 46:19:@174.4]
  assign _GEN_449 = 4'h1 == io_selects_14_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_450 = 4'h2 == io_selects_14_0 ? io_inputs_2 : _GEN_449; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_451 = 4'h3 == io_selects_14_0 ? io_inputs_3 : _GEN_450; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_452 = 4'h4 == io_selects_14_0 ? io_inputs_4 : _GEN_451; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_453 = 4'h5 == io_selects_14_0 ? io_inputs_5 : _GEN_452; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_454 = 4'h6 == io_selects_14_0 ? io_inputs_6 : _GEN_453; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_455 = 4'h7 == io_selects_14_0 ? io_inputs_7 : _GEN_454; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_456 = 4'h8 == io_selects_14_0 ? io_inputs_8 : _GEN_455; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_457 = 4'h9 == io_selects_14_0 ? io_inputs_9 : _GEN_456; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_458 = 4'ha == io_selects_14_0 ? io_inputs_10 : _GEN_457; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_459 = 4'hb == io_selects_14_0 ? io_inputs_11 : _GEN_458; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_460 = 4'hc == io_selects_14_0 ? io_inputs_12 : _GEN_459; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_461 = 4'hd == io_selects_14_0 ? io_inputs_13 : _GEN_460; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_462 = 4'he == io_selects_14_0 ? io_inputs_14 : _GEN_461; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_463 = 4'hf == io_selects_14_0 ? io_inputs_15 : _GEN_462; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_465 = 4'h1 == io_selects_14_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_466 = 4'h2 == io_selects_14_1 ? io_inputs_2 : _GEN_465; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_467 = 4'h3 == io_selects_14_1 ? io_inputs_3 : _GEN_466; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_468 = 4'h4 == io_selects_14_1 ? io_inputs_4 : _GEN_467; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_469 = 4'h5 == io_selects_14_1 ? io_inputs_5 : _GEN_468; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_470 = 4'h6 == io_selects_14_1 ? io_inputs_6 : _GEN_469; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_471 = 4'h7 == io_selects_14_1 ? io_inputs_7 : _GEN_470; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_472 = 4'h8 == io_selects_14_1 ? io_inputs_8 : _GEN_471; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_473 = 4'h9 == io_selects_14_1 ? io_inputs_9 : _GEN_472; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_474 = 4'ha == io_selects_14_1 ? io_inputs_10 : _GEN_473; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_475 = 4'hb == io_selects_14_1 ? io_inputs_11 : _GEN_474; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_476 = 4'hc == io_selects_14_1 ? io_inputs_12 : _GEN_475; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_477 = 4'hd == io_selects_14_1 ? io_inputs_13 : _GEN_476; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_478 = 4'he == io_selects_14_1 ? io_inputs_14 : _GEN_477; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_479 = 4'hf == io_selects_14_1 ? io_inputs_15 : _GEN_478; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _T_960 = _GEN_463 + _GEN_479; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _T_961 = _GEN_463 + _GEN_479; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@177.4]
  assign _T_963 = _GEN_463 * _GEN_479; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@178.4]
  assign _T_965 = _GEN_463 / _GEN_479; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@179.4]
  assign _T_966 = 3'h3 == io_operation_14; // @[Mux.scala 46:19:@180.4]
  assign _T_967 = _T_966 ? _T_965 : 64'h0; // @[Mux.scala 46:16:@181.4]
  assign _T_968 = 3'h2 == io_operation_14; // @[Mux.scala 46:19:@182.4]
  assign _T_969 = _T_968 ? _T_963 : {{64'd0}, _T_967}; // @[Mux.scala 46:16:@183.4]
  assign _T_970 = 3'h1 == io_operation_14; // @[Mux.scala 46:19:@184.4]
  assign _T_971 = _T_970 ? {{64'd0}, _T_961} : _T_969; // @[Mux.scala 46:16:@185.4]
  assign _T_972 = 3'h0 == io_operation_14; // @[Mux.scala 46:19:@186.4]
  assign _GEN_481 = 4'h1 == io_selects_15_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_482 = 4'h2 == io_selects_15_0 ? io_inputs_2 : _GEN_481; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_483 = 4'h3 == io_selects_15_0 ? io_inputs_3 : _GEN_482; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_484 = 4'h4 == io_selects_15_0 ? io_inputs_4 : _GEN_483; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_485 = 4'h5 == io_selects_15_0 ? io_inputs_5 : _GEN_484; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_486 = 4'h6 == io_selects_15_0 ? io_inputs_6 : _GEN_485; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_487 = 4'h7 == io_selects_15_0 ? io_inputs_7 : _GEN_486; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_488 = 4'h8 == io_selects_15_0 ? io_inputs_8 : _GEN_487; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_489 = 4'h9 == io_selects_15_0 ? io_inputs_9 : _GEN_488; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_490 = 4'ha == io_selects_15_0 ? io_inputs_10 : _GEN_489; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_491 = 4'hb == io_selects_15_0 ? io_inputs_11 : _GEN_490; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_492 = 4'hc == io_selects_15_0 ? io_inputs_12 : _GEN_491; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_493 = 4'hd == io_selects_15_0 ? io_inputs_13 : _GEN_492; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_494 = 4'he == io_selects_15_0 ? io_inputs_14 : _GEN_493; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_495 = 4'hf == io_selects_15_0 ? io_inputs_15 : _GEN_494; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_497 = 4'h1 == io_selects_15_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_498 = 4'h2 == io_selects_15_1 ? io_inputs_2 : _GEN_497; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_499 = 4'h3 == io_selects_15_1 ? io_inputs_3 : _GEN_498; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_500 = 4'h4 == io_selects_15_1 ? io_inputs_4 : _GEN_499; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_501 = 4'h5 == io_selects_15_1 ? io_inputs_5 : _GEN_500; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_502 = 4'h6 == io_selects_15_1 ? io_inputs_6 : _GEN_501; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_503 = 4'h7 == io_selects_15_1 ? io_inputs_7 : _GEN_502; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_504 = 4'h8 == io_selects_15_1 ? io_inputs_8 : _GEN_503; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_505 = 4'h9 == io_selects_15_1 ? io_inputs_9 : _GEN_504; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_506 = 4'ha == io_selects_15_1 ? io_inputs_10 : _GEN_505; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_507 = 4'hb == io_selects_15_1 ? io_inputs_11 : _GEN_506; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_508 = 4'hc == io_selects_15_1 ? io_inputs_12 : _GEN_507; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_509 = 4'hd == io_selects_15_1 ? io_inputs_13 : _GEN_508; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_510 = 4'he == io_selects_15_1 ? io_inputs_14 : _GEN_509; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_511 = 4'hf == io_selects_15_1 ? io_inputs_15 : _GEN_510; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _T_977 = _GEN_495 + _GEN_511; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _T_978 = _GEN_495 + _GEN_511; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 32:53:@189.4]
  assign _T_980 = _GEN_495 * _GEN_511; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 33:58:@190.4]
  assign _T_982 = _GEN_495 / _GEN_511; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 34:56:@191.4]
  assign _T_983 = 3'h3 == io_operation_15; // @[Mux.scala 46:19:@192.4]
  assign _T_984 = _T_983 ? _T_982 : 64'h0; // @[Mux.scala 46:16:@193.4]
  assign _T_985 = 3'h2 == io_operation_15; // @[Mux.scala 46:19:@194.4]
  assign _T_986 = _T_985 ? _T_980 : {{64'd0}, _T_984}; // @[Mux.scala 46:16:@195.4]
  assign _T_987 = 3'h1 == io_operation_15; // @[Mux.scala 46:19:@196.4]
  assign _T_988 = _T_987 ? {{64'd0}, _T_978} : _T_986; // @[Mux.scala 46:16:@197.4]
  assign _T_989 = 3'h0 == io_operation_15; // @[Mux.scala 46:19:@198.4]
  assign io_outputs_0 = _T_1001[63:0]; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 23:14:@520.4]
  assign io_outputs_1 = _T_1012[63:0]; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 23:14:@521.4]
  assign io_outputs_2 = _T_1023[63:0]; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 23:14:@522.4]
  assign io_outputs_3 = _T_1034[63:0]; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 23:14:@523.4]
  assign io_outputs_4 = _T_1045[63:0]; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 23:14:@524.4]
  assign io_outputs_5 = _T_1056[63:0]; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 23:14:@525.4]
  assign io_outputs_6 = _T_1067[63:0]; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 23:14:@526.4]
  assign io_outputs_7 = _T_1078[63:0]; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 23:14:@527.4]
  assign io_outputs_8 = _T_1089[63:0]; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 23:14:@528.4]
  assign io_outputs_9 = _T_1100[63:0]; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 23:14:@529.4]
  assign io_outputs_10 = _T_1111[63:0]; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 23:14:@530.4]
  assign io_outputs_11 = _T_1122[63:0]; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 23:14:@531.4]
  assign io_outputs_12 = _T_1133[63:0]; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 23:14:@532.4]
  assign io_outputs_13 = _T_1144[63:0]; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 23:14:@533.4]
  assign io_outputs_14 = _T_1155[63:0]; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 23:14:@534.4]
  assign io_outputs_15 = _T_1166[63:0]; // @[MuxTest_width_64_inputs_16_outputs_16_pipeline_5s.scala 23:14:@535.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  _T_993 = _RAND_0[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {4{`RANDOM}};
  _T_995 = _RAND_1[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {4{`RANDOM}};
  _T_997 = _RAND_2[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {4{`RANDOM}};
  _T_999 = _RAND_3[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {4{`RANDOM}};
  _T_1001 = _RAND_4[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {4{`RANDOM}};
  _T_1004 = _RAND_5[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {4{`RANDOM}};
  _T_1006 = _RAND_6[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {4{`RANDOM}};
  _T_1008 = _RAND_7[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {4{`RANDOM}};
  _T_1010 = _RAND_8[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {4{`RANDOM}};
  _T_1012 = _RAND_9[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {4{`RANDOM}};
  _T_1015 = _RAND_10[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {4{`RANDOM}};
  _T_1017 = _RAND_11[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {4{`RANDOM}};
  _T_1019 = _RAND_12[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {4{`RANDOM}};
  _T_1021 = _RAND_13[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {4{`RANDOM}};
  _T_1023 = _RAND_14[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {4{`RANDOM}};
  _T_1026 = _RAND_15[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {4{`RANDOM}};
  _T_1028 = _RAND_16[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {4{`RANDOM}};
  _T_1030 = _RAND_17[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {4{`RANDOM}};
  _T_1032 = _RAND_18[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {4{`RANDOM}};
  _T_1034 = _RAND_19[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {4{`RANDOM}};
  _T_1037 = _RAND_20[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {4{`RANDOM}};
  _T_1039 = _RAND_21[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {4{`RANDOM}};
  _T_1041 = _RAND_22[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {4{`RANDOM}};
  _T_1043 = _RAND_23[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {4{`RANDOM}};
  _T_1045 = _RAND_24[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {4{`RANDOM}};
  _T_1048 = _RAND_25[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {4{`RANDOM}};
  _T_1050 = _RAND_26[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {4{`RANDOM}};
  _T_1052 = _RAND_27[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {4{`RANDOM}};
  _T_1054 = _RAND_28[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {4{`RANDOM}};
  _T_1056 = _RAND_29[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {4{`RANDOM}};
  _T_1059 = _RAND_30[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {4{`RANDOM}};
  _T_1061 = _RAND_31[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {4{`RANDOM}};
  _T_1063 = _RAND_32[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {4{`RANDOM}};
  _T_1065 = _RAND_33[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {4{`RANDOM}};
  _T_1067 = _RAND_34[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {4{`RANDOM}};
  _T_1070 = _RAND_35[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {4{`RANDOM}};
  _T_1072 = _RAND_36[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {4{`RANDOM}};
  _T_1074 = _RAND_37[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {4{`RANDOM}};
  _T_1076 = _RAND_38[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {4{`RANDOM}};
  _T_1078 = _RAND_39[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {4{`RANDOM}};
  _T_1081 = _RAND_40[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {4{`RANDOM}};
  _T_1083 = _RAND_41[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {4{`RANDOM}};
  _T_1085 = _RAND_42[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {4{`RANDOM}};
  _T_1087 = _RAND_43[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {4{`RANDOM}};
  _T_1089 = _RAND_44[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {4{`RANDOM}};
  _T_1092 = _RAND_45[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {4{`RANDOM}};
  _T_1094 = _RAND_46[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {4{`RANDOM}};
  _T_1096 = _RAND_47[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {4{`RANDOM}};
  _T_1098 = _RAND_48[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {4{`RANDOM}};
  _T_1100 = _RAND_49[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {4{`RANDOM}};
  _T_1103 = _RAND_50[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {4{`RANDOM}};
  _T_1105 = _RAND_51[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {4{`RANDOM}};
  _T_1107 = _RAND_52[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {4{`RANDOM}};
  _T_1109 = _RAND_53[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {4{`RANDOM}};
  _T_1111 = _RAND_54[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {4{`RANDOM}};
  _T_1114 = _RAND_55[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {4{`RANDOM}};
  _T_1116 = _RAND_56[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {4{`RANDOM}};
  _T_1118 = _RAND_57[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {4{`RANDOM}};
  _T_1120 = _RAND_58[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {4{`RANDOM}};
  _T_1122 = _RAND_59[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {4{`RANDOM}};
  _T_1125 = _RAND_60[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {4{`RANDOM}};
  _T_1127 = _RAND_61[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {4{`RANDOM}};
  _T_1129 = _RAND_62[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {4{`RANDOM}};
  _T_1131 = _RAND_63[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {4{`RANDOM}};
  _T_1133 = _RAND_64[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {4{`RANDOM}};
  _T_1136 = _RAND_65[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {4{`RANDOM}};
  _T_1138 = _RAND_66[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {4{`RANDOM}};
  _T_1140 = _RAND_67[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {4{`RANDOM}};
  _T_1142 = _RAND_68[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {4{`RANDOM}};
  _T_1144 = _RAND_69[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {4{`RANDOM}};
  _T_1147 = _RAND_70[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {4{`RANDOM}};
  _T_1149 = _RAND_71[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {4{`RANDOM}};
  _T_1151 = _RAND_72[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {4{`RANDOM}};
  _T_1153 = _RAND_73[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {4{`RANDOM}};
  _T_1155 = _RAND_74[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {4{`RANDOM}};
  _T_1158 = _RAND_75[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {4{`RANDOM}};
  _T_1160 = _RAND_76[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {4{`RANDOM}};
  _T_1162 = _RAND_77[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {4{`RANDOM}};
  _T_1164 = _RAND_78[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {4{`RANDOM}};
  _T_1166 = _RAND_79[127:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_734) begin
      _T_993 <= {{64'd0}, _GEN_15};
    end else begin
      _T_993 <= _T_733;
    end
    _T_995 <= _T_993;
    _T_997 <= _T_995;
    _T_999 <= _T_997;
    _T_1001 <= _T_999;
    if (_T_751) begin
      _T_1004 <= {{64'd0}, _GEN_47};
    end else begin
      _T_1004 <= _T_750;
    end
    _T_1006 <= _T_1004;
    _T_1008 <= _T_1006;
    _T_1010 <= _T_1008;
    _T_1012 <= _T_1010;
    if (_T_768) begin
      _T_1015 <= {{64'd0}, _GEN_79};
    end else begin
      _T_1015 <= _T_767;
    end
    _T_1017 <= _T_1015;
    _T_1019 <= _T_1017;
    _T_1021 <= _T_1019;
    _T_1023 <= _T_1021;
    if (_T_785) begin
      _T_1026 <= {{64'd0}, _GEN_111};
    end else begin
      _T_1026 <= _T_784;
    end
    _T_1028 <= _T_1026;
    _T_1030 <= _T_1028;
    _T_1032 <= _T_1030;
    _T_1034 <= _T_1032;
    if (_T_802) begin
      _T_1037 <= {{64'd0}, _GEN_143};
    end else begin
      _T_1037 <= _T_801;
    end
    _T_1039 <= _T_1037;
    _T_1041 <= _T_1039;
    _T_1043 <= _T_1041;
    _T_1045 <= _T_1043;
    if (_T_819) begin
      _T_1048 <= {{64'd0}, _GEN_175};
    end else begin
      _T_1048 <= _T_818;
    end
    _T_1050 <= _T_1048;
    _T_1052 <= _T_1050;
    _T_1054 <= _T_1052;
    _T_1056 <= _T_1054;
    if (_T_836) begin
      _T_1059 <= {{64'd0}, _GEN_207};
    end else begin
      _T_1059 <= _T_835;
    end
    _T_1061 <= _T_1059;
    _T_1063 <= _T_1061;
    _T_1065 <= _T_1063;
    _T_1067 <= _T_1065;
    if (_T_853) begin
      _T_1070 <= {{64'd0}, _GEN_239};
    end else begin
      _T_1070 <= _T_852;
    end
    _T_1072 <= _T_1070;
    _T_1074 <= _T_1072;
    _T_1076 <= _T_1074;
    _T_1078 <= _T_1076;
    if (_T_870) begin
      _T_1081 <= {{64'd0}, _GEN_271};
    end else begin
      _T_1081 <= _T_869;
    end
    _T_1083 <= _T_1081;
    _T_1085 <= _T_1083;
    _T_1087 <= _T_1085;
    _T_1089 <= _T_1087;
    if (_T_887) begin
      _T_1092 <= {{64'd0}, _GEN_303};
    end else begin
      _T_1092 <= _T_886;
    end
    _T_1094 <= _T_1092;
    _T_1096 <= _T_1094;
    _T_1098 <= _T_1096;
    _T_1100 <= _T_1098;
    if (_T_904) begin
      _T_1103 <= {{64'd0}, _GEN_335};
    end else begin
      _T_1103 <= _T_903;
    end
    _T_1105 <= _T_1103;
    _T_1107 <= _T_1105;
    _T_1109 <= _T_1107;
    _T_1111 <= _T_1109;
    if (_T_921) begin
      _T_1114 <= {{64'd0}, _GEN_367};
    end else begin
      _T_1114 <= _T_920;
    end
    _T_1116 <= _T_1114;
    _T_1118 <= _T_1116;
    _T_1120 <= _T_1118;
    _T_1122 <= _T_1120;
    if (_T_938) begin
      _T_1125 <= {{64'd0}, _GEN_399};
    end else begin
      _T_1125 <= _T_937;
    end
    _T_1127 <= _T_1125;
    _T_1129 <= _T_1127;
    _T_1131 <= _T_1129;
    _T_1133 <= _T_1131;
    if (_T_955) begin
      _T_1136 <= {{64'd0}, _GEN_431};
    end else begin
      _T_1136 <= _T_954;
    end
    _T_1138 <= _T_1136;
    _T_1140 <= _T_1138;
    _T_1142 <= _T_1140;
    _T_1144 <= _T_1142;
    if (_T_972) begin
      _T_1147 <= {{64'd0}, _GEN_463};
    end else begin
      _T_1147 <= _T_971;
    end
    _T_1149 <= _T_1147;
    _T_1151 <= _T_1149;
    _T_1153 <= _T_1151;
    _T_1155 <= _T_1153;
    if (_T_989) begin
      _T_1158 <= {{64'd0}, _GEN_495};
    end else begin
      _T_1158 <= _T_988;
    end
    _T_1160 <= _T_1158;
    _T_1162 <= _T_1160;
    _T_1164 <= _T_1162;
    _T_1166 <= _T_1164;
  end
endmodule
