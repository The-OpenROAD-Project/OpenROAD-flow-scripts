(* blackbox *) module A2O1A1Ixp33_ASAP7_75t_L (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module A2O1A1O1Ixp25_ASAP7_75t_L (Y, A1, A2, B, C, D);
	output Y;
	input A1, A2, B, C, D;
endmodule
(* blackbox *) module AO211x2_ASAP7_75t_L (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module AO21x1_ASAP7_75t_L (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AO21x2_ASAP7_75t_L (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AO221x1_ASAP7_75t_L (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module AO221x2_ASAP7_75t_L (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module AO222x2_ASAP7_75t_L (Y, A1, A2, B1, B2, C1, C2);
	output Y;
	input A1, A2, B1, B2, C1, C2;
endmodule
(* blackbox *) module AO22x1_ASAP7_75t_L (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AO22x2_ASAP7_75t_L (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AO31x2_ASAP7_75t_L (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module AO322x2_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, C1, C2;
endmodule
(* blackbox *) module AO32x1_ASAP7_75t_L (Y, A1, A2, A3, B1, B2);
	output Y;
	input A1, A2, A3, B1, B2;
endmodule
(* blackbox *) module AO32x2_ASAP7_75t_L (Y, A1, A2, A3, B1, B2);
	output Y;
	input A1, A2, A3, B1, B2;
endmodule
(* blackbox *) module AO331x1_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C);
	output Y;
	input A1, A2, A3, B1, B2, B3, C;
endmodule
(* blackbox *) module AO331x2_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C);
	output Y;
	input A1, A2, A3, B1, B2, B3, C;
endmodule
(* blackbox *) module AO332x1_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module AO332x2_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module AO333x1_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module AO333x2_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module AO33x2_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3);
	output Y;
	input A1, A2, A3, B1, B2, B3;
endmodule
(* blackbox *) module AOI211x1_ASAP7_75t_L (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module AOI211xp5_ASAP7_75t_L (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module AOI21x1_ASAP7_75t_L (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AOI21xp33_ASAP7_75t_L (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AOI21xp5_ASAP7_75t_L (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AOI221x1_ASAP7_75t_L (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module AOI221xp5_ASAP7_75t_L (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module AOI222xp33_ASAP7_75t_L (Y, A1, A2, B1, B2, C1, C2);
	output Y;
	input A1, A2, B1, B2, C1, C2;
endmodule
(* blackbox *) module AOI22x1_ASAP7_75t_L (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AOI22xp33_ASAP7_75t_L (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AOI22xp5_ASAP7_75t_L (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AOI311xp33_ASAP7_75t_L (Y, A1, A2, A3, B, C);
	output Y;
	input A1, A2, A3, B, C;
endmodule
(* blackbox *) module AOI31xp33_ASAP7_75t_L (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module AOI31xp67_ASAP7_75t_L (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module AOI321xp33_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, C);
	output Y;
	input A1, A2, A3, B1, B2, C;
endmodule
(* blackbox *) module AOI322xp5_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, C1, C2;
endmodule
(* blackbox *) module AOI32xp33_ASAP7_75t_L (Y, A1, A2, A3, B1, B2);
	output Y;
	input A1, A2, A3, B1, B2;
endmodule
(* blackbox *) module AOI331xp33_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C1);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1;
endmodule
(* blackbox *) module AOI332xp33_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module AOI333xp33_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module AOI33xp33_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3);
	output Y;
	input A1, A2, A3, B1, B2, B3;
endmodule
(* blackbox *) module A2O1A1Ixp33_ASAP7_75t_R (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module A2O1A1O1Ixp25_ASAP7_75t_R (Y, A1, A2, B, C, D);
	output Y;
	input A1, A2, B, C, D;
endmodule
(* blackbox *) module AO211x2_ASAP7_75t_R (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module AO21x1_ASAP7_75t_R (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AO21x2_ASAP7_75t_R (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AO221x1_ASAP7_75t_R (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module AO221x2_ASAP7_75t_R (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module AO222x2_ASAP7_75t_R (Y, A1, A2, B1, B2, C1, C2);
	output Y;
	input A1, A2, B1, B2, C1, C2;
endmodule
(* blackbox *) module AO22x1_ASAP7_75t_R (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AO22x2_ASAP7_75t_R (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AO31x2_ASAP7_75t_R (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module AO322x2_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, C1, C2;
endmodule
(* blackbox *) module AO32x1_ASAP7_75t_R (Y, A1, A2, A3, B1, B2);
	output Y;
	input A1, A2, A3, B1, B2;
endmodule
(* blackbox *) module AO32x2_ASAP7_75t_R (Y, A1, A2, A3, B1, B2);
	output Y;
	input A1, A2, A3, B1, B2;
endmodule
(* blackbox *) module AO331x1_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, B3, C);
	output Y;
	input A1, A2, A3, B1, B2, B3, C;
endmodule
(* blackbox *) module AO331x2_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, B3, C);
	output Y;
	input A1, A2, A3, B1, B2, B3, C;
endmodule
(* blackbox *) module AO332x1_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module AO332x2_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module AO333x1_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module AO333x2_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module AO33x2_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, B3);
	output Y;
	input A1, A2, A3, B1, B2, B3;
endmodule
(* blackbox *) module AOI211x1_ASAP7_75t_R (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module AOI211xp5_ASAP7_75t_R (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module AOI21x1_ASAP7_75t_R (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AOI21xp33_ASAP7_75t_R (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AOI21xp5_ASAP7_75t_R (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AOI221x1_ASAP7_75t_R (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module AOI221xp5_ASAP7_75t_R (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module AOI222xp33_ASAP7_75t_R (Y, A1, A2, B1, B2, C1, C2);
	output Y;
	input A1, A2, B1, B2, C1, C2;
endmodule
(* blackbox *) module AOI22x1_ASAP7_75t_R (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AOI22xp33_ASAP7_75t_R (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AOI22xp5_ASAP7_75t_R (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AOI311xp33_ASAP7_75t_R (Y, A1, A2, A3, B, C);
	output Y;
	input A1, A2, A3, B, C;
endmodule
(* blackbox *) module AOI31xp33_ASAP7_75t_R (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module AOI31xp67_ASAP7_75t_R (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module AOI321xp33_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, C);
	output Y;
	input A1, A2, A3, B1, B2, C;
endmodule
(* blackbox *) module AOI322xp5_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, C1, C2;
endmodule
(* blackbox *) module AOI32xp33_ASAP7_75t_R (Y, A1, A2, A3, B1, B2);
	output Y;
	input A1, A2, A3, B1, B2;
endmodule
(* blackbox *) module AOI331xp33_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, B3, C1);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1;
endmodule
(* blackbox *) module AOI332xp33_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module AOI333xp33_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module AOI33xp33_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, B3);
	output Y;
	input A1, A2, A3, B1, B2, B3;
endmodule
(* blackbox *) module A2O1A1Ixp33_ASAP7_75t_SL (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module A2O1A1O1Ixp25_ASAP7_75t_SL (Y, A1, A2, B, C, D);
	output Y;
	input A1, A2, B, C, D;
endmodule
(* blackbox *) module AO211x2_ASAP7_75t_SL (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module AO21x1_ASAP7_75t_SL (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AO21x2_ASAP7_75t_SL (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AO221x1_ASAP7_75t_SL (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module AO221x2_ASAP7_75t_SL (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module AO222x2_ASAP7_75t_SL (Y, A1, A2, B1, B2, C1, C2);
	output Y;
	input A1, A2, B1, B2, C1, C2;
endmodule
(* blackbox *) module AO22x1_ASAP7_75t_SL (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AO22x2_ASAP7_75t_SL (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AO31x2_ASAP7_75t_SL (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module AO322x2_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, C1, C2;
endmodule
(* blackbox *) module AO32x1_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2);
	output Y;
	input A1, A2, A3, B1, B2;
endmodule
(* blackbox *) module AO32x2_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2);
	output Y;
	input A1, A2, A3, B1, B2;
endmodule
(* blackbox *) module AO331x1_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C);
	output Y;
	input A1, A2, A3, B1, B2, B3, C;
endmodule
(* blackbox *) module AO331x2_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C);
	output Y;
	input A1, A2, A3, B1, B2, B3, C;
endmodule
(* blackbox *) module AO332x1_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module AO332x2_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module AO333x1_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module AO333x2_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module AO33x2_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3);
	output Y;
	input A1, A2, A3, B1, B2, B3;
endmodule
(* blackbox *) module AOI211x1_ASAP7_75t_SL (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module AOI211xp5_ASAP7_75t_SL (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module AOI21x1_ASAP7_75t_SL (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AOI21xp33_ASAP7_75t_SL (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AOI21xp5_ASAP7_75t_SL (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AOI221x1_ASAP7_75t_SL (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module AOI221xp5_ASAP7_75t_SL (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module AOI222xp33_ASAP7_75t_SL (Y, A1, A2, B1, B2, C1, C2);
	output Y;
	input A1, A2, B1, B2, C1, C2;
endmodule
(* blackbox *) module AOI22x1_ASAP7_75t_SL (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AOI22xp33_ASAP7_75t_SL (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AOI22xp5_ASAP7_75t_SL (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AOI311xp33_ASAP7_75t_SL (Y, A1, A2, A3, B, C);
	output Y;
	input A1, A2, A3, B, C;
endmodule
(* blackbox *) module AOI31xp33_ASAP7_75t_SL (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module AOI31xp67_ASAP7_75t_SL (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module AOI321xp33_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, C);
	output Y;
	input A1, A2, A3, B1, B2, C;
endmodule
(* blackbox *) module AOI322xp5_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, C1, C2;
endmodule
(* blackbox *) module AOI32xp33_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2);
	output Y;
	input A1, A2, A3, B1, B2;
endmodule
(* blackbox *) module AOI331xp33_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1;
endmodule
(* blackbox *) module AOI332xp33_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module AOI333xp33_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module AOI33xp33_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3);
	output Y;
	input A1, A2, A3, B1, B2, B3;
endmodule
(* blackbox *) module A2O1A1Ixp33_ASAP7_75t_SRAM (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module A2O1A1O1Ixp25_ASAP7_75t_SRAM (Y, A1, A2, B, C, D);
	output Y;
	input A1, A2, B, C, D;
endmodule
(* blackbox *) module AO211x2_ASAP7_75t_SRAM (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module AO21x1_ASAP7_75t_SRAM (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AO21x2_ASAP7_75t_SRAM (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AO221x1_ASAP7_75t_SRAM (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module AO221x2_ASAP7_75t_SRAM (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module AO222x2_ASAP7_75t_SRAM (Y, A1, A2, B1, B2, C1, C2);
	output Y;
	input A1, A2, B1, B2, C1, C2;
endmodule
(* blackbox *) module AO22x1_ASAP7_75t_SRAM (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AO22x2_ASAP7_75t_SRAM (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AO31x2_ASAP7_75t_SRAM (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module AO322x2_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, C1, C2;
endmodule
(* blackbox *) module AO32x1_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2);
	output Y;
	input A1, A2, A3, B1, B2;
endmodule
(* blackbox *) module AO32x2_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2);
	output Y;
	input A1, A2, A3, B1, B2;
endmodule
(* blackbox *) module AO331x1_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, B3, C);
	output Y;
	input A1, A2, A3, B1, B2, B3, C;
endmodule
(* blackbox *) module AO331x2_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, B3, C);
	output Y;
	input A1, A2, A3, B1, B2, B3, C;
endmodule
(* blackbox *) module AO332x1_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module AO332x2_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module AO333x1_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module AO333x2_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module AO33x2_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, B3);
	output Y;
	input A1, A2, A3, B1, B2, B3;
endmodule
(* blackbox *) module AOI211x1_ASAP7_75t_SRAM (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module AOI211xp5_ASAP7_75t_SRAM (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module AOI21x1_ASAP7_75t_SRAM (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AOI21xp33_ASAP7_75t_SRAM (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AOI21xp5_ASAP7_75t_SRAM (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module AOI221x1_ASAP7_75t_SRAM (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module AOI221xp5_ASAP7_75t_SRAM (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module AOI222xp33_ASAP7_75t_SRAM (Y, A1, A2, B1, B2, C1, C2);
	output Y;
	input A1, A2, B1, B2, C1, C2;
endmodule
(* blackbox *) module AOI22x1_ASAP7_75t_SRAM (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AOI22xp33_ASAP7_75t_SRAM (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AOI22xp5_ASAP7_75t_SRAM (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module AOI311xp33_ASAP7_75t_SRAM (Y, A1, A2, A3, B, C);
	output Y;
	input A1, A2, A3, B, C;
endmodule
(* blackbox *) module AOI31xp33_ASAP7_75t_SRAM (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module AOI31xp67_ASAP7_75t_SRAM (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module AOI321xp33_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, C);
	output Y;
	input A1, A2, A3, B1, B2, C;
endmodule
(* blackbox *) module AOI322xp5_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, C1, C2;
endmodule
(* blackbox *) module AOI32xp33_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2);
	output Y;
	input A1, A2, A3, B1, B2;
endmodule
(* blackbox *) module AOI331xp33_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, B3, C1);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1;
endmodule
(* blackbox *) module AOI332xp33_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module AOI333xp33_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module AOI33xp33_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, B3);
	output Y;
	input A1, A2, A3, B1, B2, B3;
endmodule
(* blackbox *) module BUFx10_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx12_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx12f_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx16f_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx24_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx2_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx3_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx4_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx4f_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx5_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx6f_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx8_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx10_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx11_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx12_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx14_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx16_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx20_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx5p33_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx6p67_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx8_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx9p33_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module HB1xp67_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module HB2xp67_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module HB3xp67_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module HB4xp67_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx11_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx13_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx1_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx2_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx3_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx4_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx5_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx6_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx8_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVxp33_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVxp67_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx10_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx12_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx12f_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx16f_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx24_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx2_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx3_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx4_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx4f_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx5_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx6f_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx8_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx10_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx11_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx12_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx14_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx16_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx20_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx5p33_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx6p67_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx8_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx9p33_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module HB1xp67_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module HB2xp67_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module HB3xp67_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module HB4xp67_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx11_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx13_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx1_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx2_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx3_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx4_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx5_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx6_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx8_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVxp33_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVxp67_ASAP7_75t_R (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx10_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx12_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx12f_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx16f_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx24_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx2_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx3_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx4_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx4f_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx5_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx6f_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx8_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx10_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx11_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx12_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx14_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx16_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx20_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx5p33_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx6p67_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx8_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx9p33_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module HB1xp67_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module HB2xp67_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module HB3xp67_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module HB4xp67_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx11_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx13_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx1_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx2_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx3_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx4_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx5_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx6_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx8_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVxp33_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVxp67_ASAP7_75t_SL (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx10_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx12_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx12f_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx16f_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx24_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx2_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx3_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx4_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx4f_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx5_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx6f_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx8_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx10_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx11_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx12_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx14_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx16_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx20_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx5p33_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx6p67_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx8_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx9p33_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module HB1xp67_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module HB2xp67_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module HB3xp67_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module HB4xp67_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx11_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx13_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx1_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx2_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx3_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx4_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx5_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx6_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx8_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVxp33_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVxp67_ASAP7_75t_SRAM (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module O2A1O1Ixp33_ASAP7_75t_L (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module O2A1O1Ixp5_ASAP7_75t_L (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module OA211x2_ASAP7_75t_L (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module OA21x2_ASAP7_75t_L (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module OA221x2_ASAP7_75t_L (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module OA222x2_ASAP7_75t_L (Y, A1, A2, B1, B2, C1, C2);
	output Y;
	input A1, A2, B1, B2, C1, C2;
endmodule
(* blackbox *) module OA22x2_ASAP7_75t_L (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module OA31x2_ASAP7_75t_L (Y, A1, A2, A3, B1);
	output Y;
	input A1, A2, A3, B1;
endmodule
(* blackbox *) module OA331x1_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C1);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1;
endmodule
(* blackbox *) module OA331x2_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C1);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1;
endmodule
(* blackbox *) module OA332x1_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module OA332x2_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module OA333x1_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module OA333x2_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module OA33x2_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3);
	output Y;
	input A1, A2, A3, B1, B2, B3;
endmodule
(* blackbox *) module OAI211xp5_ASAP7_75t_L (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module OAI21x1_ASAP7_75t_L (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module OAI21xp33_ASAP7_75t_L (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module OAI21xp5_ASAP7_75t_L (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module OAI221xp5_ASAP7_75t_L (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module OAI222xp33_ASAP7_75t_L (Y, A1, A2, B1, B2, C1, C2);
	output Y;
	input A1, A2, B1, B2, C1, C2;
endmodule
(* blackbox *) module OAI22x1_ASAP7_75t_L (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module OAI22xp33_ASAP7_75t_L (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module OAI22xp5_ASAP7_75t_L (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module OAI311xp33_ASAP7_75t_L (Y, A1, A2, A3, B1, C1);
	output Y;
	input A1, A2, A3, B1, C1;
endmodule
(* blackbox *) module OAI31xp33_ASAP7_75t_L (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module OAI31xp67_ASAP7_75t_L (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module OAI321xp33_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, C);
	output Y;
	input A1, A2, A3, B1, B2, C;
endmodule
(* blackbox *) module OAI322xp33_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, C1, C2;
endmodule
(* blackbox *) module OAI32xp33_ASAP7_75t_L (Y, A1, A2, A3, B1, B2);
	output Y;
	input A1, A2, A3, B1, B2;
endmodule
(* blackbox *) module OAI331xp33_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C1);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1;
endmodule
(* blackbox *) module OAI332xp33_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module OAI333xp33_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module OAI33xp33_ASAP7_75t_L (Y, A1, A2, A3, B1, B2, B3);
	output Y;
	input A1, A2, A3, B1, B2, B3;
endmodule
(* blackbox *) module O2A1O1Ixp33_ASAP7_75t_R (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module O2A1O1Ixp5_ASAP7_75t_R (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module OA211x2_ASAP7_75t_R (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module OA21x2_ASAP7_75t_R (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module OA221x2_ASAP7_75t_R (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module OA222x2_ASAP7_75t_R (Y, A1, A2, B1, B2, C1, C2);
	output Y;
	input A1, A2, B1, B2, C1, C2;
endmodule
(* blackbox *) module OA22x2_ASAP7_75t_R (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module OA31x2_ASAP7_75t_R (Y, A1, A2, A3, B1);
	output Y;
	input A1, A2, A3, B1;
endmodule
(* blackbox *) module OA331x1_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, B3, C1);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1;
endmodule
(* blackbox *) module OA331x2_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, B3, C1);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1;
endmodule
(* blackbox *) module OA332x1_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module OA332x2_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module OA333x1_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module OA333x2_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module OA33x2_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, B3);
	output Y;
	input A1, A2, A3, B1, B2, B3;
endmodule
(* blackbox *) module OAI211xp5_ASAP7_75t_R (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module OAI21x1_ASAP7_75t_R (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module OAI21xp33_ASAP7_75t_R (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module OAI21xp5_ASAP7_75t_R (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module OAI221xp5_ASAP7_75t_R (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module OAI222xp33_ASAP7_75t_R (Y, A1, A2, B1, B2, C1, C2);
	output Y;
	input A1, A2, B1, B2, C1, C2;
endmodule
(* blackbox *) module OAI22x1_ASAP7_75t_R (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module OAI22xp33_ASAP7_75t_R (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module OAI22xp5_ASAP7_75t_R (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module OAI311xp33_ASAP7_75t_R (Y, A1, A2, A3, B1, C1);
	output Y;
	input A1, A2, A3, B1, C1;
endmodule
(* blackbox *) module OAI31xp33_ASAP7_75t_R (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module OAI31xp67_ASAP7_75t_R (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module OAI321xp33_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, C);
	output Y;
	input A1, A2, A3, B1, B2, C;
endmodule
(* blackbox *) module OAI322xp33_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, C1, C2;
endmodule
(* blackbox *) module OAI32xp33_ASAP7_75t_R (Y, A1, A2, A3, B1, B2);
	output Y;
	input A1, A2, A3, B1, B2;
endmodule
(* blackbox *) module OAI331xp33_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, B3, C1);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1;
endmodule
(* blackbox *) module OAI332xp33_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module OAI333xp33_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module OAI33xp33_ASAP7_75t_R (Y, A1, A2, A3, B1, B2, B3);
	output Y;
	input A1, A2, A3, B1, B2, B3;
endmodule
(* blackbox *) module O2A1O1Ixp33_ASAP7_75t_SL (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module O2A1O1Ixp5_ASAP7_75t_SL (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module OA211x2_ASAP7_75t_SL (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module OA21x2_ASAP7_75t_SL (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module OA221x2_ASAP7_75t_SL (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module OA222x2_ASAP7_75t_SL (Y, A1, A2, B1, B2, C1, C2);
	output Y;
	input A1, A2, B1, B2, C1, C2;
endmodule
(* blackbox *) module OA22x2_ASAP7_75t_SL (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module OA31x2_ASAP7_75t_SL (Y, A1, A2, A3, B1);
	output Y;
	input A1, A2, A3, B1;
endmodule
(* blackbox *) module OA331x1_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1;
endmodule
(* blackbox *) module OA331x2_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1;
endmodule
(* blackbox *) module OA332x1_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module OA332x2_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module OA333x1_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module OA333x2_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module OA33x2_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3);
	output Y;
	input A1, A2, A3, B1, B2, B3;
endmodule
(* blackbox *) module OAI211xp5_ASAP7_75t_SL (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module OAI21x1_ASAP7_75t_SL (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module OAI21xp33_ASAP7_75t_SL (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module OAI21xp5_ASAP7_75t_SL (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module OAI221xp5_ASAP7_75t_SL (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module OAI222xp33_ASAP7_75t_SL (Y, A1, A2, B1, B2, C1, C2);
	output Y;
	input A1, A2, B1, B2, C1, C2;
endmodule
(* blackbox *) module OAI22x1_ASAP7_75t_SL (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module OAI22xp33_ASAP7_75t_SL (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module OAI22xp5_ASAP7_75t_SL (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module OAI311xp33_ASAP7_75t_SL (Y, A1, A2, A3, B1, C1);
	output Y;
	input A1, A2, A3, B1, C1;
endmodule
(* blackbox *) module OAI31xp33_ASAP7_75t_SL (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module OAI31xp67_ASAP7_75t_SL (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module OAI321xp33_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, C);
	output Y;
	input A1, A2, A3, B1, B2, C;
endmodule
(* blackbox *) module OAI322xp33_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, C1, C2;
endmodule
(* blackbox *) module OAI32xp33_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2);
	output Y;
	input A1, A2, A3, B1, B2;
endmodule
(* blackbox *) module OAI331xp33_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1;
endmodule
(* blackbox *) module OAI332xp33_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module OAI333xp33_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module OAI33xp33_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3);
	output Y;
	input A1, A2, A3, B1, B2, B3;
endmodule
(* blackbox *) module O2A1O1Ixp33_ASAP7_75t_SRAM (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module O2A1O1Ixp5_ASAP7_75t_SRAM (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module OA211x2_ASAP7_75t_SRAM (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module OA21x2_ASAP7_75t_SRAM (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module OA221x2_ASAP7_75t_SRAM (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module OA222x2_ASAP7_75t_SRAM (Y, A1, A2, B1, B2, C1, C2);
	output Y;
	input A1, A2, B1, B2, C1, C2;
endmodule
(* blackbox *) module OA22x2_ASAP7_75t_SRAM (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module OA31x2_ASAP7_75t_SRAM (Y, A1, A2, A3, B1);
	output Y;
	input A1, A2, A3, B1;
endmodule
(* blackbox *) module OA331x1_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, B3, C1);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1;
endmodule
(* blackbox *) module OA331x2_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, B3, C1);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1;
endmodule
(* blackbox *) module OA332x1_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module OA332x2_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module OA333x1_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module OA333x2_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module OA33x2_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, B3);
	output Y;
	input A1, A2, A3, B1, B2, B3;
endmodule
(* blackbox *) module OAI211xp5_ASAP7_75t_SRAM (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module OAI21x1_ASAP7_75t_SRAM (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module OAI21xp33_ASAP7_75t_SRAM (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module OAI21xp5_ASAP7_75t_SRAM (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module OAI221xp5_ASAP7_75t_SRAM (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module OAI222xp33_ASAP7_75t_SRAM (Y, A1, A2, B1, B2, C1, C2);
	output Y;
	input A1, A2, B1, B2, C1, C2;
endmodule
(* blackbox *) module OAI22x1_ASAP7_75t_SRAM (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module OAI22xp33_ASAP7_75t_SRAM (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module OAI22xp5_ASAP7_75t_SRAM (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module OAI311xp33_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, C1);
	output Y;
	input A1, A2, A3, B1, C1;
endmodule
(* blackbox *) module OAI31xp33_ASAP7_75t_SRAM (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module OAI31xp67_ASAP7_75t_SRAM (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module OAI321xp33_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, C);
	output Y;
	input A1, A2, A3, B1, B2, C;
endmodule
(* blackbox *) module OAI322xp33_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, C1, C2;
endmodule
(* blackbox *) module OAI32xp33_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2);
	output Y;
	input A1, A2, A3, B1, B2;
endmodule
(* blackbox *) module OAI331xp33_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, B3, C1);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1;
endmodule
(* blackbox *) module OAI332xp33_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module OAI333xp33_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module OAI33xp33_ASAP7_75t_SRAM (Y, A1, A2, A3, B1, B2, B3);
	output Y;
	input A1, A2, A3, B1, B2, B3;
endmodule
(* blackbox *) module ASYNC_DFFHx1_ASAP7_75t_L (QN, D, RESET, SET, CLK);
	output QN;
	input D, RESET, SET, CLK;
endmodule
(* blackbox *) module DFFHQNx1_ASAP7_75t_L (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFHQNx2_ASAP7_75t_L (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFHQNx3_ASAP7_75t_L (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFHQx4_ASAP7_75t_L (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DFFLQNx1_ASAP7_75t_L (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFLQNx2_ASAP7_75t_L (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFLQNx3_ASAP7_75t_L (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFLQx4_ASAP7_75t_L (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DHLx1_ASAP7_75t_L (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DHLx2_ASAP7_75t_L (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DHLx3_ASAP7_75t_L (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DLLx1_ASAP7_75t_L (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DLLx2_ASAP7_75t_L (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DLLx3_ASAP7_75t_L (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module ICGx1_ASAP7_75t_L (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx2_ASAP7_75t_L (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx2p67DC_ASAP7_75t_L (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx3_ASAP7_75t_L (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx4DC_ASAP7_75t_L (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx4_ASAP7_75t_L (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx5_ASAP7_75t_L (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx5p33DC_ASAP7_75t_L (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx6p67DC_ASAP7_75t_L (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx8DC_ASAP7_75t_L (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module SDFHx1_ASAP7_75t_L (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFHx2_ASAP7_75t_L (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFHx3_ASAP7_75t_L (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFHx4_ASAP7_75t_L (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFLx1_ASAP7_75t_L (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFLx2_ASAP7_75t_L (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFLx3_ASAP7_75t_L (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFLx4_ASAP7_75t_L (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module ASYNC_DFFHx1_ASAP7_75t_R (QN, D, RESET, SET, CLK);
	output QN;
	input D, RESET, SET, CLK;
endmodule
(* blackbox *) module DFFHQNx1_ASAP7_75t_R (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFHQNx2_ASAP7_75t_R (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFHQNx3_ASAP7_75t_R (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFHQx4_ASAP7_75t_R (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DFFLQNx1_ASAP7_75t_R (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFLQNx2_ASAP7_75t_R (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFLQNx3_ASAP7_75t_R (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFLQx4_ASAP7_75t_R (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DHLx1_ASAP7_75t_R (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DHLx2_ASAP7_75t_R (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DHLx3_ASAP7_75t_R (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DLLx1_ASAP7_75t_R (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DLLx2_ASAP7_75t_R (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DLLx3_ASAP7_75t_R (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module ICGx1_ASAP7_75t_R (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx2_ASAP7_75t_R (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx2p67DC_ASAP7_75t_R (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx3_ASAP7_75t_R (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx4DC_ASAP7_75t_R (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx4_ASAP7_75t_R (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx5_ASAP7_75t_R (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx5p33DC_ASAP7_75t_R (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx6p67DC_ASAP7_75t_R (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx8DC_ASAP7_75t_R (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module SDFHx1_ASAP7_75t_R (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFHx2_ASAP7_75t_R (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFHx3_ASAP7_75t_R (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFHx4_ASAP7_75t_R (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFLx1_ASAP7_75t_R (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFLx2_ASAP7_75t_R (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFLx3_ASAP7_75t_R (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFLx4_ASAP7_75t_R (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module ASYNC_DFFHx1_ASAP7_75t_SL (QN, D, RESET, SET, CLK);
	output QN;
	input D, RESET, SET, CLK;
endmodule
(* blackbox *) module DFFHQNx1_ASAP7_75t_SL (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFHQNx2_ASAP7_75t_SL (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFHQNx3_ASAP7_75t_SL (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFHQx4_ASAP7_75t_SL (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DFFLQNx1_ASAP7_75t_SL (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFLQNx2_ASAP7_75t_SL (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFLQNx3_ASAP7_75t_SL (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFLQx4_ASAP7_75t_SL (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DHLx1_ASAP7_75t_SL (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DHLx2_ASAP7_75t_SL (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DHLx3_ASAP7_75t_SL (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DLLx1_ASAP7_75t_SL (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DLLx2_ASAP7_75t_SL (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DLLx3_ASAP7_75t_SL (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module ICGx1_ASAP7_75t_SL (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx2_ASAP7_75t_SL (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx2p67DC_ASAP7_75t_SL (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx3_ASAP7_75t_SL (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx4DC_ASAP7_75t_SL (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx4_ASAP7_75t_SL (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx5_ASAP7_75t_SL (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx5p33DC_ASAP7_75t_SL (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx6p67DC_ASAP7_75t_SL (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx8DC_ASAP7_75t_SL (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module SDFHx1_ASAP7_75t_SL (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFHx2_ASAP7_75t_SL (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFHx3_ASAP7_75t_SL (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFHx4_ASAP7_75t_SL (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFLx1_ASAP7_75t_SL (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFLx2_ASAP7_75t_SL (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFLx3_ASAP7_75t_SL (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFLx4_ASAP7_75t_SL (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module ASYNC_DFFHx1_ASAP7_75t_SRAM (QN, D, RESET, SET, CLK);
	output QN;
	input D, RESET, SET, CLK;
endmodule
(* blackbox *) module DFFHQNx1_ASAP7_75t_SRAM (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFHQNx2_ASAP7_75t_SRAM (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFHQNx3_ASAP7_75t_SRAM (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFHQx4_ASAP7_75t_SRAM (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DFFLQNx1_ASAP7_75t_SRAM (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFLQNx2_ASAP7_75t_SRAM (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFLQNx3_ASAP7_75t_SRAM (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFLQx4_ASAP7_75t_SRAM (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DHLx1_ASAP7_75t_SRAM (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DHLx2_ASAP7_75t_SRAM (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DHLx3_ASAP7_75t_SRAM (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DLLx1_ASAP7_75t_SRAM (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DLLx2_ASAP7_75t_SRAM (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DLLx3_ASAP7_75t_SRAM (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module ICGx1_ASAP7_75t_SRAM (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx2_ASAP7_75t_SRAM (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx2p67DC_ASAP7_75t_SRAM (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx3_ASAP7_75t_SRAM (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx4DC_ASAP7_75t_SRAM (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx4_ASAP7_75t_SRAM (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx5_ASAP7_75t_SRAM (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx5p33DC_ASAP7_75t_SRAM (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx6p67DC_ASAP7_75t_SRAM (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx8DC_ASAP7_75t_SRAM (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module SDFHx1_ASAP7_75t_SRAM (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFHx2_ASAP7_75t_SRAM (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFHx3_ASAP7_75t_SRAM (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFHx4_ASAP7_75t_SRAM (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFLx1_ASAP7_75t_SRAM (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFLx2_ASAP7_75t_SRAM (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFLx3_ASAP7_75t_SRAM (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFLx4_ASAP7_75t_SRAM (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module AND2x2_ASAP7_75t_L (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module AND2x4_ASAP7_75t_L (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module AND2x6_ASAP7_75t_L (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module AND3x1_ASAP7_75t_L (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module AND3x2_ASAP7_75t_L (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module AND3x4_ASAP7_75t_L (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module AND4x1_ASAP7_75t_L (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module AND4x2_ASAP7_75t_L (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module AND5x1_ASAP7_75t_L (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module AND5x2_ASAP7_75t_L (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module FAx1_ASAP7_75t_L (CON, SN, A, B, CI);
	output CON, SN;
	input A, B, CI;
endmodule
(* blackbox *) module HAxp5_ASAP7_75t_L (CON, SN, A, B);
	output CON, SN;
	input A, B;
endmodule
(* blackbox *) module MAJIxp5_ASAP7_75t_L (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module MAJx2_ASAP7_75t_L (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module MAJx3_ASAP7_75t_L (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NAND2x1_ASAP7_75t_L (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2x1p5_ASAP7_75t_L (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2x2_ASAP7_75t_L (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2xp33_ASAP7_75t_L (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2xp5_ASAP7_75t_L (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2xp67_ASAP7_75t_L (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND3x1_ASAP7_75t_L (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NAND3x2_ASAP7_75t_L (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NAND3xp33_ASAP7_75t_L (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NAND4xp25_ASAP7_75t_L (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module NAND4xp75_ASAP7_75t_L (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module NAND5xp2_ASAP7_75t_L (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module NOR2x1_ASAP7_75t_L (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR2x1p5_ASAP7_75t_L (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR2x2_ASAP7_75t_L (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR2xp33_ASAP7_75t_L (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR2xp67_ASAP7_75t_L (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR3x1_ASAP7_75t_L (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NOR3x2_ASAP7_75t_L (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NOR3xp33_ASAP7_75t_L (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NOR4xp25_ASAP7_75t_L (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module NOR4xp75_ASAP7_75t_L (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module NOR5xp2_ASAP7_75t_L (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module OR2x2_ASAP7_75t_L (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module OR2x4_ASAP7_75t_L (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module OR2x6_ASAP7_75t_L (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module OR3x1_ASAP7_75t_L (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module OR3x2_ASAP7_75t_L (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module OR3x4_ASAP7_75t_L (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module OR4x1_ASAP7_75t_L (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module OR4x2_ASAP7_75t_L (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module OR5x1_ASAP7_75t_L (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module OR5x2_ASAP7_75t_L (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module TIEHIx1_ASAP7_75t_L (H);
	output H;
endmodule
(* blackbox *) module TIELOx1_ASAP7_75t_L (L);
	output L;
endmodule
(* blackbox *) module XNOR2x1_ASAP7_75t_L (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XNOR2x2_ASAP7_75t_L (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XNOR2xp5_ASAP7_75t_L (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XOR2x1_ASAP7_75t_L (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XOR2x2_ASAP7_75t_L (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XOR2xp5_ASAP7_75t_L (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module AND2x2_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module AND2x4_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module AND2x6_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module AND3x1_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module AND3x2_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module AND3x4_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module AND4x1_ASAP7_75t_R (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module AND4x2_ASAP7_75t_R (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module AND5x1_ASAP7_75t_R (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module AND5x2_ASAP7_75t_R (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module FAx1_ASAP7_75t_R (CON, SN, A, B, CI);
	output CON, SN;
	input A, B, CI;
endmodule
(* blackbox *) module HAxp5_ASAP7_75t_R (CON, SN, A, B);
	output CON, SN;
	input A, B;
endmodule
(* blackbox *) module MAJIxp5_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module MAJx2_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module MAJx3_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NAND2x1_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2x1p5_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2x2_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2xp33_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2xp5_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2xp67_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND3x1_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NAND3x2_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NAND3xp33_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NAND4xp25_ASAP7_75t_R (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module NAND4xp75_ASAP7_75t_R (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module NAND5xp2_ASAP7_75t_R (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module NOR2x1_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR2x1p5_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR2x2_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR2xp33_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR2xp67_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR3x1_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NOR3x2_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NOR3xp33_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NOR4xp25_ASAP7_75t_R (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module NOR4xp75_ASAP7_75t_R (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module NOR5xp2_ASAP7_75t_R (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module OR2x2_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module OR2x4_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module OR2x6_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module OR3x1_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module OR3x2_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module OR3x4_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module OR4x1_ASAP7_75t_R (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module OR4x2_ASAP7_75t_R (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module OR5x1_ASAP7_75t_R (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module OR5x2_ASAP7_75t_R (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module TIEHIx1_ASAP7_75t_R (H);
	output H;
endmodule
(* blackbox *) module TIELOx1_ASAP7_75t_R (L);
	output L;
endmodule
(* blackbox *) module XNOR2x1_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XNOR2x2_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XNOR2xp5_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XOR2x1_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XOR2x2_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XOR2xp5_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module AND2x2_ASAP7_75t_SL (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module AND2x4_ASAP7_75t_SL (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module AND2x6_ASAP7_75t_SL (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module AND3x1_ASAP7_75t_SL (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module AND3x2_ASAP7_75t_SL (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module AND3x4_ASAP7_75t_SL (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module AND4x1_ASAP7_75t_SL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module AND4x2_ASAP7_75t_SL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module AND5x1_ASAP7_75t_SL (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module AND5x2_ASAP7_75t_SL (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module FAx1_ASAP7_75t_SL (CON, SN, A, B, CI);
	output CON, SN;
	input A, B, CI;
endmodule
(* blackbox *) module HAxp5_ASAP7_75t_SL (CON, SN, A, B);
	output CON, SN;
	input A, B;
endmodule
(* blackbox *) module MAJIxp5_ASAP7_75t_SL (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module MAJx2_ASAP7_75t_SL (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module MAJx3_ASAP7_75t_SL (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NAND2x1_ASAP7_75t_SL (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2x1p5_ASAP7_75t_SL (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2x2_ASAP7_75t_SL (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2xp33_ASAP7_75t_SL (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2xp5_ASAP7_75t_SL (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2xp67_ASAP7_75t_SL (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND3x1_ASAP7_75t_SL (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NAND3x2_ASAP7_75t_SL (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NAND3xp33_ASAP7_75t_SL (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NAND4xp25_ASAP7_75t_SL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module NAND4xp75_ASAP7_75t_SL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module NAND5xp2_ASAP7_75t_SL (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module NOR2x1_ASAP7_75t_SL (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR2x1p5_ASAP7_75t_SL (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR2x2_ASAP7_75t_SL (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR2xp33_ASAP7_75t_SL (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR2xp67_ASAP7_75t_SL (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR3x1_ASAP7_75t_SL (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NOR3x2_ASAP7_75t_SL (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NOR3xp33_ASAP7_75t_SL (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NOR4xp25_ASAP7_75t_SL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module NOR4xp75_ASAP7_75t_SL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module NOR5xp2_ASAP7_75t_SL (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module OR2x2_ASAP7_75t_SL (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module OR2x4_ASAP7_75t_SL (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module OR2x6_ASAP7_75t_SL (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module OR3x1_ASAP7_75t_SL (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module OR3x2_ASAP7_75t_SL (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module OR3x4_ASAP7_75t_SL (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module OR4x1_ASAP7_75t_SL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module OR4x2_ASAP7_75t_SL (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module OR5x1_ASAP7_75t_SL (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module OR5x2_ASAP7_75t_SL (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module TIEHIx1_ASAP7_75t_SL (H);
	output H;
endmodule
(* blackbox *) module TIELOx1_ASAP7_75t_SL (L);
	output L;
endmodule
(* blackbox *) module XNOR2x1_ASAP7_75t_SL (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XNOR2x2_ASAP7_75t_SL (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XNOR2xp5_ASAP7_75t_SL (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XOR2x1_ASAP7_75t_SL (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XOR2x2_ASAP7_75t_SL (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XOR2xp5_ASAP7_75t_SL (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module AND2x2_ASAP7_75t_SRAM (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module AND2x4_ASAP7_75t_SRAM (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module AND2x6_ASAP7_75t_SRAM (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module AND3x1_ASAP7_75t_SRAM (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module AND3x2_ASAP7_75t_SRAM (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module AND3x4_ASAP7_75t_SRAM (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module AND4x1_ASAP7_75t_SRAM (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module AND4x2_ASAP7_75t_SRAM (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module AND5x1_ASAP7_75t_SRAM (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module AND5x2_ASAP7_75t_SRAM (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module FAx1_ASAP7_75t_SRAM (CON, SN, A, B, CI);
	output CON, SN;
	input A, B, CI;
endmodule
(* blackbox *) module HAxp5_ASAP7_75t_SRAM (CON, SN, A, B);
	output CON, SN;
	input A, B;
endmodule
(* blackbox *) module MAJIxp5_ASAP7_75t_SRAM (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module MAJx2_ASAP7_75t_SRAM (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module MAJx3_ASAP7_75t_SRAM (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NAND2x1_ASAP7_75t_SRAM (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2x1p5_ASAP7_75t_SRAM (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2x2_ASAP7_75t_SRAM (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2xp33_ASAP7_75t_SRAM (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2xp5_ASAP7_75t_SRAM (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2xp67_ASAP7_75t_SRAM (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND3x1_ASAP7_75t_SRAM (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NAND3x2_ASAP7_75t_SRAM (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NAND3xp33_ASAP7_75t_SRAM (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NAND4xp25_ASAP7_75t_SRAM (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module NAND4xp75_ASAP7_75t_SRAM (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module NAND5xp2_ASAP7_75t_SRAM (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module NOR2x1_ASAP7_75t_SRAM (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR2x1p5_ASAP7_75t_SRAM (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR2x2_ASAP7_75t_SRAM (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR2xp33_ASAP7_75t_SRAM (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR2xp67_ASAP7_75t_SRAM (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR3x1_ASAP7_75t_SRAM (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NOR3x2_ASAP7_75t_SRAM (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NOR3xp33_ASAP7_75t_SRAM (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NOR4xp25_ASAP7_75t_SRAM (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module NOR4xp75_ASAP7_75t_SRAM (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module NOR5xp2_ASAP7_75t_SRAM (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module OR2x2_ASAP7_75t_SRAM (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module OR2x4_ASAP7_75t_SRAM (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module OR2x6_ASAP7_75t_SRAM (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module OR3x1_ASAP7_75t_SRAM (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module OR3x2_ASAP7_75t_SRAM (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module OR3x4_ASAP7_75t_SRAM (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module OR4x1_ASAP7_75t_SRAM (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module OR4x2_ASAP7_75t_SRAM (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module OR5x1_ASAP7_75t_SRAM (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module OR5x2_ASAP7_75t_SRAM (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module TIEHIx1_ASAP7_75t_SRAM (H);
	output H;
endmodule
(* blackbox *) module TIELOx1_ASAP7_75t_SRAM (L);
	output L;
endmodule
(* blackbox *) module XNOR2x1_ASAP7_75t_SRAM (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XNOR2x2_ASAP7_75t_SRAM (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XNOR2xp5_ASAP7_75t_SRAM (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XOR2x1_ASAP7_75t_SRAM (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XOR2x2_ASAP7_75t_SRAM (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XOR2xp5_ASAP7_75t_SRAM (Y, A, B);
	output Y;
	input A, B;
endmodule
