module MockArray(
  input         clock,
  input         reset,
  input  [63:0] io_ins_down_0,
  input  [63:0] io_ins_down_1,
  input  [63:0] io_ins_down_2,
  input  [63:0] io_ins_down_3,
  input  [63:0] io_ins_down_4,
  input  [63:0] io_ins_down_5,
  input  [63:0] io_ins_down_6,
  input  [63:0] io_ins_down_7,
  input  [63:0] io_ins_up_0,
  input  [63:0] io_ins_up_1,
  input  [63:0] io_ins_up_2,
  input  [63:0] io_ins_up_3,
  input  [63:0] io_ins_up_4,
  input  [63:0] io_ins_up_5,
  input  [63:0] io_ins_up_6,
  input  [63:0] io_ins_up_7,
  input  [63:0] io_ins_right_0,
  input  [63:0] io_ins_right_1,
  input  [63:0] io_ins_right_2,
  input  [63:0] io_ins_right_3,
  input  [63:0] io_ins_right_4,
  input  [63:0] io_ins_right_5,
  input  [63:0] io_ins_right_6,
  input  [63:0] io_ins_right_7,
  input  [63:0] io_ins_left_0,
  input  [63:0] io_ins_left_1,
  input  [63:0] io_ins_left_2,
  input  [63:0] io_ins_left_3,
  input  [63:0] io_ins_left_4,
  input  [63:0] io_ins_left_5,
  input  [63:0] io_ins_left_6,
  input  [63:0] io_ins_left_7,
  output [63:0] io_outs_down_0,
  output [63:0] io_outs_down_1,
  output [63:0] io_outs_down_2,
  output [63:0] io_outs_down_3,
  output [63:0] io_outs_down_4,
  output [63:0] io_outs_down_5,
  output [63:0] io_outs_down_6,
  output [63:0] io_outs_down_7,
  output [63:0] io_outs_up_0,
  output [63:0] io_outs_up_1,
  output [63:0] io_outs_up_2,
  output [63:0] io_outs_up_3,
  output [63:0] io_outs_up_4,
  output [63:0] io_outs_up_5,
  output [63:0] io_outs_up_6,
  output [63:0] io_outs_up_7,
  output [63:0] io_outs_right_0,
  output [63:0] io_outs_right_1,
  output [63:0] io_outs_right_2,
  output [63:0] io_outs_right_3,
  output [63:0] io_outs_right_4,
  output [63:0] io_outs_right_5,
  output [63:0] io_outs_right_6,
  output [63:0] io_outs_right_7,
  output [63:0] io_outs_left_0,
  output [63:0] io_outs_left_1,
  output [63:0] io_outs_left_2,
  output [63:0] io_outs_left_3,
  output [63:0] io_outs_left_4,
  output [63:0] io_outs_left_5,
  output [63:0] io_outs_left_6,
  output [63:0] io_outs_left_7,
  output        io_lsbs_0,
  output        io_lsbs_1,
  output        io_lsbs_2,
  output        io_lsbs_3,
  output        io_lsbs_4,
  output        io_lsbs_5,
  output        io_lsbs_6,
  output        io_lsbs_7,
  output        io_lsbs_8,
  output        io_lsbs_9,
  output        io_lsbs_10,
  output        io_lsbs_11,
  output        io_lsbs_12,
  output        io_lsbs_13,
  output        io_lsbs_14,
  output        io_lsbs_15,
  output        io_lsbs_16,
  output        io_lsbs_17,
  output        io_lsbs_18,
  output        io_lsbs_19,
  output        io_lsbs_20,
  output        io_lsbs_21,
  output        io_lsbs_22,
  output        io_lsbs_23,
  output        io_lsbs_24,
  output        io_lsbs_25,
  output        io_lsbs_26,
  output        io_lsbs_27,
  output        io_lsbs_28,
  output        io_lsbs_29,
  output        io_lsbs_30,
  output        io_lsbs_31,
  output        io_lsbs_32,
  output        io_lsbs_33,
  output        io_lsbs_34,
  output        io_lsbs_35,
  output        io_lsbs_36,
  output        io_lsbs_37,
  output        io_lsbs_38,
  output        io_lsbs_39,
  output        io_lsbs_40,
  output        io_lsbs_41,
  output        io_lsbs_42,
  output        io_lsbs_43,
  output        io_lsbs_44,
  output        io_lsbs_45,
  output        io_lsbs_46,
  output        io_lsbs_47,
  output        io_lsbs_48,
  output        io_lsbs_49,
  output        io_lsbs_50,
  output        io_lsbs_51,
  output        io_lsbs_52,
  output        io_lsbs_53,
  output        io_lsbs_54,
  output        io_lsbs_55,
  output        io_lsbs_56,
  output        io_lsbs_57,
  output        io_lsbs_58,
  output        io_lsbs_59,
  output        io_lsbs_60,
  output        io_lsbs_61,
  output        io_lsbs_62,
  output        io_lsbs_63
);
  wire  ces_0_0_clock;
  wire  ces_0_0_io_clockOutRight;
  wire [63:0] ces_0_0_io_ins_down;
  wire [63:0] ces_0_0_io_ins_right;
  wire [63:0] ces_0_0_io_ins_up;
  wire [63:0] ces_0_0_io_ins_left;
  wire [63:0] ces_0_0_io_outs_down;
  wire [63:0] ces_0_0_io_outs_right;
  wire [63:0] ces_0_0_io_outs_up;
  wire [63:0] ces_0_0_io_outs_left;
  wire  ces_0_0_io_lsbIns_1;
  wire  ces_0_0_io_lsbIns_2;
  wire  ces_0_0_io_lsbIns_3;
  wire  ces_0_0_io_lsbIns_4;
  wire  ces_0_0_io_lsbIns_5;
  wire  ces_0_0_io_lsbIns_6;
  wire  ces_0_0_io_lsbIns_7;
  wire  ces_0_0_io_lsbOuts_0;
  wire  ces_0_0_io_lsbOuts_1;
  wire  ces_0_0_io_lsbOuts_2;
  wire  ces_0_0_io_lsbOuts_3;
  wire  ces_0_0_io_lsbOuts_4;
  wire  ces_0_0_io_lsbOuts_5;
  wire  ces_0_0_io_lsbOuts_6;
  wire  ces_0_0_io_lsbOuts_7;
  wire  ces_0_1_clock;
  wire  ces_0_1_io_clockOutRight;
  wire [63:0] ces_0_1_io_ins_down;
  wire [63:0] ces_0_1_io_ins_right;
  wire [63:0] ces_0_1_io_ins_up;
  wire [63:0] ces_0_1_io_ins_left;
  wire [63:0] ces_0_1_io_outs_down;
  wire [63:0] ces_0_1_io_outs_right;
  wire [63:0] ces_0_1_io_outs_up;
  wire [63:0] ces_0_1_io_outs_left;
  wire  ces_0_1_io_lsbIns_1;
  wire  ces_0_1_io_lsbIns_2;
  wire  ces_0_1_io_lsbIns_3;
  wire  ces_0_1_io_lsbIns_4;
  wire  ces_0_1_io_lsbIns_5;
  wire  ces_0_1_io_lsbIns_6;
  wire  ces_0_1_io_lsbIns_7;
  wire  ces_0_1_io_lsbOuts_0;
  wire  ces_0_1_io_lsbOuts_1;
  wire  ces_0_1_io_lsbOuts_2;
  wire  ces_0_1_io_lsbOuts_3;
  wire  ces_0_1_io_lsbOuts_4;
  wire  ces_0_1_io_lsbOuts_5;
  wire  ces_0_1_io_lsbOuts_6;
  wire  ces_0_1_io_lsbOuts_7;
  wire  ces_0_2_clock;
  wire  ces_0_2_io_clockOutRight;
  wire [63:0] ces_0_2_io_ins_down;
  wire [63:0] ces_0_2_io_ins_right;
  wire [63:0] ces_0_2_io_ins_up;
  wire [63:0] ces_0_2_io_ins_left;
  wire [63:0] ces_0_2_io_outs_down;
  wire [63:0] ces_0_2_io_outs_right;
  wire [63:0] ces_0_2_io_outs_up;
  wire [63:0] ces_0_2_io_outs_left;
  wire  ces_0_2_io_lsbIns_1;
  wire  ces_0_2_io_lsbIns_2;
  wire  ces_0_2_io_lsbIns_3;
  wire  ces_0_2_io_lsbIns_4;
  wire  ces_0_2_io_lsbIns_5;
  wire  ces_0_2_io_lsbIns_6;
  wire  ces_0_2_io_lsbIns_7;
  wire  ces_0_2_io_lsbOuts_0;
  wire  ces_0_2_io_lsbOuts_1;
  wire  ces_0_2_io_lsbOuts_2;
  wire  ces_0_2_io_lsbOuts_3;
  wire  ces_0_2_io_lsbOuts_4;
  wire  ces_0_2_io_lsbOuts_5;
  wire  ces_0_2_io_lsbOuts_6;
  wire  ces_0_2_io_lsbOuts_7;
  wire  ces_0_3_clock;
  wire  ces_0_3_io_clockOutRight;
  wire [63:0] ces_0_3_io_ins_down;
  wire [63:0] ces_0_3_io_ins_right;
  wire [63:0] ces_0_3_io_ins_up;
  wire [63:0] ces_0_3_io_ins_left;
  wire [63:0] ces_0_3_io_outs_down;
  wire [63:0] ces_0_3_io_outs_right;
  wire [63:0] ces_0_3_io_outs_up;
  wire [63:0] ces_0_3_io_outs_left;
  wire  ces_0_3_io_lsbIns_1;
  wire  ces_0_3_io_lsbIns_2;
  wire  ces_0_3_io_lsbIns_3;
  wire  ces_0_3_io_lsbIns_4;
  wire  ces_0_3_io_lsbIns_5;
  wire  ces_0_3_io_lsbIns_6;
  wire  ces_0_3_io_lsbIns_7;
  wire  ces_0_3_io_lsbOuts_0;
  wire  ces_0_3_io_lsbOuts_1;
  wire  ces_0_3_io_lsbOuts_2;
  wire  ces_0_3_io_lsbOuts_3;
  wire  ces_0_3_io_lsbOuts_4;
  wire  ces_0_3_io_lsbOuts_5;
  wire  ces_0_3_io_lsbOuts_6;
  wire  ces_0_3_io_lsbOuts_7;
  wire  ces_0_4_clock;
  wire  ces_0_4_io_clockOutRight;
  wire [63:0] ces_0_4_io_ins_down;
  wire [63:0] ces_0_4_io_ins_right;
  wire [63:0] ces_0_4_io_ins_up;
  wire [63:0] ces_0_4_io_ins_left;
  wire [63:0] ces_0_4_io_outs_down;
  wire [63:0] ces_0_4_io_outs_right;
  wire [63:0] ces_0_4_io_outs_up;
  wire [63:0] ces_0_4_io_outs_left;
  wire  ces_0_4_io_lsbIns_1;
  wire  ces_0_4_io_lsbIns_2;
  wire  ces_0_4_io_lsbIns_3;
  wire  ces_0_4_io_lsbIns_4;
  wire  ces_0_4_io_lsbIns_5;
  wire  ces_0_4_io_lsbIns_6;
  wire  ces_0_4_io_lsbIns_7;
  wire  ces_0_4_io_lsbOuts_0;
  wire  ces_0_4_io_lsbOuts_1;
  wire  ces_0_4_io_lsbOuts_2;
  wire  ces_0_4_io_lsbOuts_3;
  wire  ces_0_4_io_lsbOuts_4;
  wire  ces_0_4_io_lsbOuts_5;
  wire  ces_0_4_io_lsbOuts_6;
  wire  ces_0_4_io_lsbOuts_7;
  wire  ces_0_5_clock;
  wire  ces_0_5_io_clockOutRight;
  wire [63:0] ces_0_5_io_ins_down;
  wire [63:0] ces_0_5_io_ins_right;
  wire [63:0] ces_0_5_io_ins_up;
  wire [63:0] ces_0_5_io_ins_left;
  wire [63:0] ces_0_5_io_outs_down;
  wire [63:0] ces_0_5_io_outs_right;
  wire [63:0] ces_0_5_io_outs_up;
  wire [63:0] ces_0_5_io_outs_left;
  wire  ces_0_5_io_lsbIns_1;
  wire  ces_0_5_io_lsbIns_2;
  wire  ces_0_5_io_lsbIns_3;
  wire  ces_0_5_io_lsbIns_4;
  wire  ces_0_5_io_lsbIns_5;
  wire  ces_0_5_io_lsbIns_6;
  wire  ces_0_5_io_lsbIns_7;
  wire  ces_0_5_io_lsbOuts_0;
  wire  ces_0_5_io_lsbOuts_1;
  wire  ces_0_5_io_lsbOuts_2;
  wire  ces_0_5_io_lsbOuts_3;
  wire  ces_0_5_io_lsbOuts_4;
  wire  ces_0_5_io_lsbOuts_5;
  wire  ces_0_5_io_lsbOuts_6;
  wire  ces_0_5_io_lsbOuts_7;
  wire  ces_0_6_clock;
  wire  ces_0_6_io_clockOutRight;
  wire [63:0] ces_0_6_io_ins_down;
  wire [63:0] ces_0_6_io_ins_right;
  wire [63:0] ces_0_6_io_ins_up;
  wire [63:0] ces_0_6_io_ins_left;
  wire [63:0] ces_0_6_io_outs_down;
  wire [63:0] ces_0_6_io_outs_right;
  wire [63:0] ces_0_6_io_outs_up;
  wire [63:0] ces_0_6_io_outs_left;
  wire  ces_0_6_io_lsbIns_1;
  wire  ces_0_6_io_lsbIns_2;
  wire  ces_0_6_io_lsbIns_3;
  wire  ces_0_6_io_lsbIns_4;
  wire  ces_0_6_io_lsbIns_5;
  wire  ces_0_6_io_lsbIns_6;
  wire  ces_0_6_io_lsbIns_7;
  wire  ces_0_6_io_lsbOuts_0;
  wire  ces_0_6_io_lsbOuts_1;
  wire  ces_0_6_io_lsbOuts_2;
  wire  ces_0_6_io_lsbOuts_3;
  wire  ces_0_6_io_lsbOuts_4;
  wire  ces_0_6_io_lsbOuts_5;
  wire  ces_0_6_io_lsbOuts_6;
  wire  ces_0_6_io_lsbOuts_7;
  wire  ces_0_7_clock;
  wire  ces_0_7_io_clockOutRight;
  wire [63:0] ces_0_7_io_ins_down;
  wire [63:0] ces_0_7_io_ins_right;
  wire [63:0] ces_0_7_io_ins_up;
  wire [63:0] ces_0_7_io_ins_left;
  wire [63:0] ces_0_7_io_outs_down;
  wire [63:0] ces_0_7_io_outs_right;
  wire [63:0] ces_0_7_io_outs_up;
  wire [63:0] ces_0_7_io_outs_left;
  wire  ces_0_7_io_lsbIns_1;
  wire  ces_0_7_io_lsbIns_2;
  wire  ces_0_7_io_lsbIns_3;
  wire  ces_0_7_io_lsbIns_4;
  wire  ces_0_7_io_lsbIns_5;
  wire  ces_0_7_io_lsbIns_6;
  wire  ces_0_7_io_lsbIns_7;
  wire  ces_0_7_io_lsbOuts_0;
  wire  ces_0_7_io_lsbOuts_1;
  wire  ces_0_7_io_lsbOuts_2;
  wire  ces_0_7_io_lsbOuts_3;
  wire  ces_0_7_io_lsbOuts_4;
  wire  ces_0_7_io_lsbOuts_5;
  wire  ces_0_7_io_lsbOuts_6;
  wire  ces_0_7_io_lsbOuts_7;
  wire  ces_1_0_clock;
  wire  ces_1_0_io_clockOutRight;
  wire [63:0] ces_1_0_io_ins_down;
  wire [63:0] ces_1_0_io_ins_right;
  wire [63:0] ces_1_0_io_ins_up;
  wire [63:0] ces_1_0_io_ins_left;
  wire [63:0] ces_1_0_io_outs_down;
  wire [63:0] ces_1_0_io_outs_right;
  wire [63:0] ces_1_0_io_outs_up;
  wire [63:0] ces_1_0_io_outs_left;
  wire  ces_1_0_io_lsbIns_1;
  wire  ces_1_0_io_lsbIns_2;
  wire  ces_1_0_io_lsbIns_3;
  wire  ces_1_0_io_lsbIns_4;
  wire  ces_1_0_io_lsbIns_5;
  wire  ces_1_0_io_lsbIns_6;
  wire  ces_1_0_io_lsbIns_7;
  wire  ces_1_0_io_lsbOuts_0;
  wire  ces_1_0_io_lsbOuts_1;
  wire  ces_1_0_io_lsbOuts_2;
  wire  ces_1_0_io_lsbOuts_3;
  wire  ces_1_0_io_lsbOuts_4;
  wire  ces_1_0_io_lsbOuts_5;
  wire  ces_1_0_io_lsbOuts_6;
  wire  ces_1_0_io_lsbOuts_7;
  wire  ces_1_1_clock;
  wire  ces_1_1_io_clockOutRight;
  wire [63:0] ces_1_1_io_ins_down;
  wire [63:0] ces_1_1_io_ins_right;
  wire [63:0] ces_1_1_io_ins_up;
  wire [63:0] ces_1_1_io_ins_left;
  wire [63:0] ces_1_1_io_outs_down;
  wire [63:0] ces_1_1_io_outs_right;
  wire [63:0] ces_1_1_io_outs_up;
  wire [63:0] ces_1_1_io_outs_left;
  wire  ces_1_1_io_lsbIns_1;
  wire  ces_1_1_io_lsbIns_2;
  wire  ces_1_1_io_lsbIns_3;
  wire  ces_1_1_io_lsbIns_4;
  wire  ces_1_1_io_lsbIns_5;
  wire  ces_1_1_io_lsbIns_6;
  wire  ces_1_1_io_lsbIns_7;
  wire  ces_1_1_io_lsbOuts_0;
  wire  ces_1_1_io_lsbOuts_1;
  wire  ces_1_1_io_lsbOuts_2;
  wire  ces_1_1_io_lsbOuts_3;
  wire  ces_1_1_io_lsbOuts_4;
  wire  ces_1_1_io_lsbOuts_5;
  wire  ces_1_1_io_lsbOuts_6;
  wire  ces_1_1_io_lsbOuts_7;
  wire  ces_1_2_clock;
  wire  ces_1_2_io_clockOutRight;
  wire [63:0] ces_1_2_io_ins_down;
  wire [63:0] ces_1_2_io_ins_right;
  wire [63:0] ces_1_2_io_ins_up;
  wire [63:0] ces_1_2_io_ins_left;
  wire [63:0] ces_1_2_io_outs_down;
  wire [63:0] ces_1_2_io_outs_right;
  wire [63:0] ces_1_2_io_outs_up;
  wire [63:0] ces_1_2_io_outs_left;
  wire  ces_1_2_io_lsbIns_1;
  wire  ces_1_2_io_lsbIns_2;
  wire  ces_1_2_io_lsbIns_3;
  wire  ces_1_2_io_lsbIns_4;
  wire  ces_1_2_io_lsbIns_5;
  wire  ces_1_2_io_lsbIns_6;
  wire  ces_1_2_io_lsbIns_7;
  wire  ces_1_2_io_lsbOuts_0;
  wire  ces_1_2_io_lsbOuts_1;
  wire  ces_1_2_io_lsbOuts_2;
  wire  ces_1_2_io_lsbOuts_3;
  wire  ces_1_2_io_lsbOuts_4;
  wire  ces_1_2_io_lsbOuts_5;
  wire  ces_1_2_io_lsbOuts_6;
  wire  ces_1_2_io_lsbOuts_7;
  wire  ces_1_3_clock;
  wire  ces_1_3_io_clockOutRight;
  wire [63:0] ces_1_3_io_ins_down;
  wire [63:0] ces_1_3_io_ins_right;
  wire [63:0] ces_1_3_io_ins_up;
  wire [63:0] ces_1_3_io_ins_left;
  wire [63:0] ces_1_3_io_outs_down;
  wire [63:0] ces_1_3_io_outs_right;
  wire [63:0] ces_1_3_io_outs_up;
  wire [63:0] ces_1_3_io_outs_left;
  wire  ces_1_3_io_lsbIns_1;
  wire  ces_1_3_io_lsbIns_2;
  wire  ces_1_3_io_lsbIns_3;
  wire  ces_1_3_io_lsbIns_4;
  wire  ces_1_3_io_lsbIns_5;
  wire  ces_1_3_io_lsbIns_6;
  wire  ces_1_3_io_lsbIns_7;
  wire  ces_1_3_io_lsbOuts_0;
  wire  ces_1_3_io_lsbOuts_1;
  wire  ces_1_3_io_lsbOuts_2;
  wire  ces_1_3_io_lsbOuts_3;
  wire  ces_1_3_io_lsbOuts_4;
  wire  ces_1_3_io_lsbOuts_5;
  wire  ces_1_3_io_lsbOuts_6;
  wire  ces_1_3_io_lsbOuts_7;
  wire  ces_1_4_clock;
  wire  ces_1_4_io_clockOutRight;
  wire [63:0] ces_1_4_io_ins_down;
  wire [63:0] ces_1_4_io_ins_right;
  wire [63:0] ces_1_4_io_ins_up;
  wire [63:0] ces_1_4_io_ins_left;
  wire [63:0] ces_1_4_io_outs_down;
  wire [63:0] ces_1_4_io_outs_right;
  wire [63:0] ces_1_4_io_outs_up;
  wire [63:0] ces_1_4_io_outs_left;
  wire  ces_1_4_io_lsbIns_1;
  wire  ces_1_4_io_lsbIns_2;
  wire  ces_1_4_io_lsbIns_3;
  wire  ces_1_4_io_lsbIns_4;
  wire  ces_1_4_io_lsbIns_5;
  wire  ces_1_4_io_lsbIns_6;
  wire  ces_1_4_io_lsbIns_7;
  wire  ces_1_4_io_lsbOuts_0;
  wire  ces_1_4_io_lsbOuts_1;
  wire  ces_1_4_io_lsbOuts_2;
  wire  ces_1_4_io_lsbOuts_3;
  wire  ces_1_4_io_lsbOuts_4;
  wire  ces_1_4_io_lsbOuts_5;
  wire  ces_1_4_io_lsbOuts_6;
  wire  ces_1_4_io_lsbOuts_7;
  wire  ces_1_5_clock;
  wire  ces_1_5_io_clockOutRight;
  wire [63:0] ces_1_5_io_ins_down;
  wire [63:0] ces_1_5_io_ins_right;
  wire [63:0] ces_1_5_io_ins_up;
  wire [63:0] ces_1_5_io_ins_left;
  wire [63:0] ces_1_5_io_outs_down;
  wire [63:0] ces_1_5_io_outs_right;
  wire [63:0] ces_1_5_io_outs_up;
  wire [63:0] ces_1_5_io_outs_left;
  wire  ces_1_5_io_lsbIns_1;
  wire  ces_1_5_io_lsbIns_2;
  wire  ces_1_5_io_lsbIns_3;
  wire  ces_1_5_io_lsbIns_4;
  wire  ces_1_5_io_lsbIns_5;
  wire  ces_1_5_io_lsbIns_6;
  wire  ces_1_5_io_lsbIns_7;
  wire  ces_1_5_io_lsbOuts_0;
  wire  ces_1_5_io_lsbOuts_1;
  wire  ces_1_5_io_lsbOuts_2;
  wire  ces_1_5_io_lsbOuts_3;
  wire  ces_1_5_io_lsbOuts_4;
  wire  ces_1_5_io_lsbOuts_5;
  wire  ces_1_5_io_lsbOuts_6;
  wire  ces_1_5_io_lsbOuts_7;
  wire  ces_1_6_clock;
  wire  ces_1_6_io_clockOutRight;
  wire [63:0] ces_1_6_io_ins_down;
  wire [63:0] ces_1_6_io_ins_right;
  wire [63:0] ces_1_6_io_ins_up;
  wire [63:0] ces_1_6_io_ins_left;
  wire [63:0] ces_1_6_io_outs_down;
  wire [63:0] ces_1_6_io_outs_right;
  wire [63:0] ces_1_6_io_outs_up;
  wire [63:0] ces_1_6_io_outs_left;
  wire  ces_1_6_io_lsbIns_1;
  wire  ces_1_6_io_lsbIns_2;
  wire  ces_1_6_io_lsbIns_3;
  wire  ces_1_6_io_lsbIns_4;
  wire  ces_1_6_io_lsbIns_5;
  wire  ces_1_6_io_lsbIns_6;
  wire  ces_1_6_io_lsbIns_7;
  wire  ces_1_6_io_lsbOuts_0;
  wire  ces_1_6_io_lsbOuts_1;
  wire  ces_1_6_io_lsbOuts_2;
  wire  ces_1_6_io_lsbOuts_3;
  wire  ces_1_6_io_lsbOuts_4;
  wire  ces_1_6_io_lsbOuts_5;
  wire  ces_1_6_io_lsbOuts_6;
  wire  ces_1_6_io_lsbOuts_7;
  wire  ces_1_7_clock;
  wire  ces_1_7_io_clockOutRight;
  wire [63:0] ces_1_7_io_ins_down;
  wire [63:0] ces_1_7_io_ins_right;
  wire [63:0] ces_1_7_io_ins_up;
  wire [63:0] ces_1_7_io_ins_left;
  wire [63:0] ces_1_7_io_outs_down;
  wire [63:0] ces_1_7_io_outs_right;
  wire [63:0] ces_1_7_io_outs_up;
  wire [63:0] ces_1_7_io_outs_left;
  wire  ces_1_7_io_lsbIns_1;
  wire  ces_1_7_io_lsbIns_2;
  wire  ces_1_7_io_lsbIns_3;
  wire  ces_1_7_io_lsbIns_4;
  wire  ces_1_7_io_lsbIns_5;
  wire  ces_1_7_io_lsbIns_6;
  wire  ces_1_7_io_lsbIns_7;
  wire  ces_1_7_io_lsbOuts_0;
  wire  ces_1_7_io_lsbOuts_1;
  wire  ces_1_7_io_lsbOuts_2;
  wire  ces_1_7_io_lsbOuts_3;
  wire  ces_1_7_io_lsbOuts_4;
  wire  ces_1_7_io_lsbOuts_5;
  wire  ces_1_7_io_lsbOuts_6;
  wire  ces_1_7_io_lsbOuts_7;
  wire  ces_2_0_clock;
  wire  ces_2_0_io_clockOutRight;
  wire [63:0] ces_2_0_io_ins_down;
  wire [63:0] ces_2_0_io_ins_right;
  wire [63:0] ces_2_0_io_ins_up;
  wire [63:0] ces_2_0_io_ins_left;
  wire [63:0] ces_2_0_io_outs_down;
  wire [63:0] ces_2_0_io_outs_right;
  wire [63:0] ces_2_0_io_outs_up;
  wire [63:0] ces_2_0_io_outs_left;
  wire  ces_2_0_io_lsbIns_1;
  wire  ces_2_0_io_lsbIns_2;
  wire  ces_2_0_io_lsbIns_3;
  wire  ces_2_0_io_lsbIns_4;
  wire  ces_2_0_io_lsbIns_5;
  wire  ces_2_0_io_lsbIns_6;
  wire  ces_2_0_io_lsbIns_7;
  wire  ces_2_0_io_lsbOuts_0;
  wire  ces_2_0_io_lsbOuts_1;
  wire  ces_2_0_io_lsbOuts_2;
  wire  ces_2_0_io_lsbOuts_3;
  wire  ces_2_0_io_lsbOuts_4;
  wire  ces_2_0_io_lsbOuts_5;
  wire  ces_2_0_io_lsbOuts_6;
  wire  ces_2_0_io_lsbOuts_7;
  wire  ces_2_1_clock;
  wire  ces_2_1_io_clockOutRight;
  wire [63:0] ces_2_1_io_ins_down;
  wire [63:0] ces_2_1_io_ins_right;
  wire [63:0] ces_2_1_io_ins_up;
  wire [63:0] ces_2_1_io_ins_left;
  wire [63:0] ces_2_1_io_outs_down;
  wire [63:0] ces_2_1_io_outs_right;
  wire [63:0] ces_2_1_io_outs_up;
  wire [63:0] ces_2_1_io_outs_left;
  wire  ces_2_1_io_lsbIns_1;
  wire  ces_2_1_io_lsbIns_2;
  wire  ces_2_1_io_lsbIns_3;
  wire  ces_2_1_io_lsbIns_4;
  wire  ces_2_1_io_lsbIns_5;
  wire  ces_2_1_io_lsbIns_6;
  wire  ces_2_1_io_lsbIns_7;
  wire  ces_2_1_io_lsbOuts_0;
  wire  ces_2_1_io_lsbOuts_1;
  wire  ces_2_1_io_lsbOuts_2;
  wire  ces_2_1_io_lsbOuts_3;
  wire  ces_2_1_io_lsbOuts_4;
  wire  ces_2_1_io_lsbOuts_5;
  wire  ces_2_1_io_lsbOuts_6;
  wire  ces_2_1_io_lsbOuts_7;
  wire  ces_2_2_clock;
  wire  ces_2_2_io_clockOutRight;
  wire [63:0] ces_2_2_io_ins_down;
  wire [63:0] ces_2_2_io_ins_right;
  wire [63:0] ces_2_2_io_ins_up;
  wire [63:0] ces_2_2_io_ins_left;
  wire [63:0] ces_2_2_io_outs_down;
  wire [63:0] ces_2_2_io_outs_right;
  wire [63:0] ces_2_2_io_outs_up;
  wire [63:0] ces_2_2_io_outs_left;
  wire  ces_2_2_io_lsbIns_1;
  wire  ces_2_2_io_lsbIns_2;
  wire  ces_2_2_io_lsbIns_3;
  wire  ces_2_2_io_lsbIns_4;
  wire  ces_2_2_io_lsbIns_5;
  wire  ces_2_2_io_lsbIns_6;
  wire  ces_2_2_io_lsbIns_7;
  wire  ces_2_2_io_lsbOuts_0;
  wire  ces_2_2_io_lsbOuts_1;
  wire  ces_2_2_io_lsbOuts_2;
  wire  ces_2_2_io_lsbOuts_3;
  wire  ces_2_2_io_lsbOuts_4;
  wire  ces_2_2_io_lsbOuts_5;
  wire  ces_2_2_io_lsbOuts_6;
  wire  ces_2_2_io_lsbOuts_7;
  wire  ces_2_3_clock;
  wire  ces_2_3_io_clockOutRight;
  wire [63:0] ces_2_3_io_ins_down;
  wire [63:0] ces_2_3_io_ins_right;
  wire [63:0] ces_2_3_io_ins_up;
  wire [63:0] ces_2_3_io_ins_left;
  wire [63:0] ces_2_3_io_outs_down;
  wire [63:0] ces_2_3_io_outs_right;
  wire [63:0] ces_2_3_io_outs_up;
  wire [63:0] ces_2_3_io_outs_left;
  wire  ces_2_3_io_lsbIns_1;
  wire  ces_2_3_io_lsbIns_2;
  wire  ces_2_3_io_lsbIns_3;
  wire  ces_2_3_io_lsbIns_4;
  wire  ces_2_3_io_lsbIns_5;
  wire  ces_2_3_io_lsbIns_6;
  wire  ces_2_3_io_lsbIns_7;
  wire  ces_2_3_io_lsbOuts_0;
  wire  ces_2_3_io_lsbOuts_1;
  wire  ces_2_3_io_lsbOuts_2;
  wire  ces_2_3_io_lsbOuts_3;
  wire  ces_2_3_io_lsbOuts_4;
  wire  ces_2_3_io_lsbOuts_5;
  wire  ces_2_3_io_lsbOuts_6;
  wire  ces_2_3_io_lsbOuts_7;
  wire  ces_2_4_clock;
  wire  ces_2_4_io_clockOutRight;
  wire [63:0] ces_2_4_io_ins_down;
  wire [63:0] ces_2_4_io_ins_right;
  wire [63:0] ces_2_4_io_ins_up;
  wire [63:0] ces_2_4_io_ins_left;
  wire [63:0] ces_2_4_io_outs_down;
  wire [63:0] ces_2_4_io_outs_right;
  wire [63:0] ces_2_4_io_outs_up;
  wire [63:0] ces_2_4_io_outs_left;
  wire  ces_2_4_io_lsbIns_1;
  wire  ces_2_4_io_lsbIns_2;
  wire  ces_2_4_io_lsbIns_3;
  wire  ces_2_4_io_lsbIns_4;
  wire  ces_2_4_io_lsbIns_5;
  wire  ces_2_4_io_lsbIns_6;
  wire  ces_2_4_io_lsbIns_7;
  wire  ces_2_4_io_lsbOuts_0;
  wire  ces_2_4_io_lsbOuts_1;
  wire  ces_2_4_io_lsbOuts_2;
  wire  ces_2_4_io_lsbOuts_3;
  wire  ces_2_4_io_lsbOuts_4;
  wire  ces_2_4_io_lsbOuts_5;
  wire  ces_2_4_io_lsbOuts_6;
  wire  ces_2_4_io_lsbOuts_7;
  wire  ces_2_5_clock;
  wire  ces_2_5_io_clockOutRight;
  wire [63:0] ces_2_5_io_ins_down;
  wire [63:0] ces_2_5_io_ins_right;
  wire [63:0] ces_2_5_io_ins_up;
  wire [63:0] ces_2_5_io_ins_left;
  wire [63:0] ces_2_5_io_outs_down;
  wire [63:0] ces_2_5_io_outs_right;
  wire [63:0] ces_2_5_io_outs_up;
  wire [63:0] ces_2_5_io_outs_left;
  wire  ces_2_5_io_lsbIns_1;
  wire  ces_2_5_io_lsbIns_2;
  wire  ces_2_5_io_lsbIns_3;
  wire  ces_2_5_io_lsbIns_4;
  wire  ces_2_5_io_lsbIns_5;
  wire  ces_2_5_io_lsbIns_6;
  wire  ces_2_5_io_lsbIns_7;
  wire  ces_2_5_io_lsbOuts_0;
  wire  ces_2_5_io_lsbOuts_1;
  wire  ces_2_5_io_lsbOuts_2;
  wire  ces_2_5_io_lsbOuts_3;
  wire  ces_2_5_io_lsbOuts_4;
  wire  ces_2_5_io_lsbOuts_5;
  wire  ces_2_5_io_lsbOuts_6;
  wire  ces_2_5_io_lsbOuts_7;
  wire  ces_2_6_clock;
  wire  ces_2_6_io_clockOutRight;
  wire [63:0] ces_2_6_io_ins_down;
  wire [63:0] ces_2_6_io_ins_right;
  wire [63:0] ces_2_6_io_ins_up;
  wire [63:0] ces_2_6_io_ins_left;
  wire [63:0] ces_2_6_io_outs_down;
  wire [63:0] ces_2_6_io_outs_right;
  wire [63:0] ces_2_6_io_outs_up;
  wire [63:0] ces_2_6_io_outs_left;
  wire  ces_2_6_io_lsbIns_1;
  wire  ces_2_6_io_lsbIns_2;
  wire  ces_2_6_io_lsbIns_3;
  wire  ces_2_6_io_lsbIns_4;
  wire  ces_2_6_io_lsbIns_5;
  wire  ces_2_6_io_lsbIns_6;
  wire  ces_2_6_io_lsbIns_7;
  wire  ces_2_6_io_lsbOuts_0;
  wire  ces_2_6_io_lsbOuts_1;
  wire  ces_2_6_io_lsbOuts_2;
  wire  ces_2_6_io_lsbOuts_3;
  wire  ces_2_6_io_lsbOuts_4;
  wire  ces_2_6_io_lsbOuts_5;
  wire  ces_2_6_io_lsbOuts_6;
  wire  ces_2_6_io_lsbOuts_7;
  wire  ces_2_7_clock;
  wire  ces_2_7_io_clockOutRight;
  wire [63:0] ces_2_7_io_ins_down;
  wire [63:0] ces_2_7_io_ins_right;
  wire [63:0] ces_2_7_io_ins_up;
  wire [63:0] ces_2_7_io_ins_left;
  wire [63:0] ces_2_7_io_outs_down;
  wire [63:0] ces_2_7_io_outs_right;
  wire [63:0] ces_2_7_io_outs_up;
  wire [63:0] ces_2_7_io_outs_left;
  wire  ces_2_7_io_lsbIns_1;
  wire  ces_2_7_io_lsbIns_2;
  wire  ces_2_7_io_lsbIns_3;
  wire  ces_2_7_io_lsbIns_4;
  wire  ces_2_7_io_lsbIns_5;
  wire  ces_2_7_io_lsbIns_6;
  wire  ces_2_7_io_lsbIns_7;
  wire  ces_2_7_io_lsbOuts_0;
  wire  ces_2_7_io_lsbOuts_1;
  wire  ces_2_7_io_lsbOuts_2;
  wire  ces_2_7_io_lsbOuts_3;
  wire  ces_2_7_io_lsbOuts_4;
  wire  ces_2_7_io_lsbOuts_5;
  wire  ces_2_7_io_lsbOuts_6;
  wire  ces_2_7_io_lsbOuts_7;
  wire  ces_3_0_clock;
  wire  ces_3_0_io_clockOutRight;
  wire [63:0] ces_3_0_io_ins_down;
  wire [63:0] ces_3_0_io_ins_right;
  wire [63:0] ces_3_0_io_ins_up;
  wire [63:0] ces_3_0_io_ins_left;
  wire [63:0] ces_3_0_io_outs_down;
  wire [63:0] ces_3_0_io_outs_right;
  wire [63:0] ces_3_0_io_outs_up;
  wire [63:0] ces_3_0_io_outs_left;
  wire  ces_3_0_io_lsbIns_1;
  wire  ces_3_0_io_lsbIns_2;
  wire  ces_3_0_io_lsbIns_3;
  wire  ces_3_0_io_lsbIns_4;
  wire  ces_3_0_io_lsbIns_5;
  wire  ces_3_0_io_lsbIns_6;
  wire  ces_3_0_io_lsbIns_7;
  wire  ces_3_0_io_lsbOuts_0;
  wire  ces_3_0_io_lsbOuts_1;
  wire  ces_3_0_io_lsbOuts_2;
  wire  ces_3_0_io_lsbOuts_3;
  wire  ces_3_0_io_lsbOuts_4;
  wire  ces_3_0_io_lsbOuts_5;
  wire  ces_3_0_io_lsbOuts_6;
  wire  ces_3_0_io_lsbOuts_7;
  wire  ces_3_1_clock;
  wire  ces_3_1_io_clockOutRight;
  wire [63:0] ces_3_1_io_ins_down;
  wire [63:0] ces_3_1_io_ins_right;
  wire [63:0] ces_3_1_io_ins_up;
  wire [63:0] ces_3_1_io_ins_left;
  wire [63:0] ces_3_1_io_outs_down;
  wire [63:0] ces_3_1_io_outs_right;
  wire [63:0] ces_3_1_io_outs_up;
  wire [63:0] ces_3_1_io_outs_left;
  wire  ces_3_1_io_lsbIns_1;
  wire  ces_3_1_io_lsbIns_2;
  wire  ces_3_1_io_lsbIns_3;
  wire  ces_3_1_io_lsbIns_4;
  wire  ces_3_1_io_lsbIns_5;
  wire  ces_3_1_io_lsbIns_6;
  wire  ces_3_1_io_lsbIns_7;
  wire  ces_3_1_io_lsbOuts_0;
  wire  ces_3_1_io_lsbOuts_1;
  wire  ces_3_1_io_lsbOuts_2;
  wire  ces_3_1_io_lsbOuts_3;
  wire  ces_3_1_io_lsbOuts_4;
  wire  ces_3_1_io_lsbOuts_5;
  wire  ces_3_1_io_lsbOuts_6;
  wire  ces_3_1_io_lsbOuts_7;
  wire  ces_3_2_clock;
  wire  ces_3_2_io_clockOutRight;
  wire [63:0] ces_3_2_io_ins_down;
  wire [63:0] ces_3_2_io_ins_right;
  wire [63:0] ces_3_2_io_ins_up;
  wire [63:0] ces_3_2_io_ins_left;
  wire [63:0] ces_3_2_io_outs_down;
  wire [63:0] ces_3_2_io_outs_right;
  wire [63:0] ces_3_2_io_outs_up;
  wire [63:0] ces_3_2_io_outs_left;
  wire  ces_3_2_io_lsbIns_1;
  wire  ces_3_2_io_lsbIns_2;
  wire  ces_3_2_io_lsbIns_3;
  wire  ces_3_2_io_lsbIns_4;
  wire  ces_3_2_io_lsbIns_5;
  wire  ces_3_2_io_lsbIns_6;
  wire  ces_3_2_io_lsbIns_7;
  wire  ces_3_2_io_lsbOuts_0;
  wire  ces_3_2_io_lsbOuts_1;
  wire  ces_3_2_io_lsbOuts_2;
  wire  ces_3_2_io_lsbOuts_3;
  wire  ces_3_2_io_lsbOuts_4;
  wire  ces_3_2_io_lsbOuts_5;
  wire  ces_3_2_io_lsbOuts_6;
  wire  ces_3_2_io_lsbOuts_7;
  wire  ces_3_3_clock;
  wire  ces_3_3_io_clockOutRight;
  wire [63:0] ces_3_3_io_ins_down;
  wire [63:0] ces_3_3_io_ins_right;
  wire [63:0] ces_3_3_io_ins_up;
  wire [63:0] ces_3_3_io_ins_left;
  wire [63:0] ces_3_3_io_outs_down;
  wire [63:0] ces_3_3_io_outs_right;
  wire [63:0] ces_3_3_io_outs_up;
  wire [63:0] ces_3_3_io_outs_left;
  wire  ces_3_3_io_lsbIns_1;
  wire  ces_3_3_io_lsbIns_2;
  wire  ces_3_3_io_lsbIns_3;
  wire  ces_3_3_io_lsbIns_4;
  wire  ces_3_3_io_lsbIns_5;
  wire  ces_3_3_io_lsbIns_6;
  wire  ces_3_3_io_lsbIns_7;
  wire  ces_3_3_io_lsbOuts_0;
  wire  ces_3_3_io_lsbOuts_1;
  wire  ces_3_3_io_lsbOuts_2;
  wire  ces_3_3_io_lsbOuts_3;
  wire  ces_3_3_io_lsbOuts_4;
  wire  ces_3_3_io_lsbOuts_5;
  wire  ces_3_3_io_lsbOuts_6;
  wire  ces_3_3_io_lsbOuts_7;
  wire  ces_3_4_clock;
  wire  ces_3_4_io_clockOutRight;
  wire [63:0] ces_3_4_io_ins_down;
  wire [63:0] ces_3_4_io_ins_right;
  wire [63:0] ces_3_4_io_ins_up;
  wire [63:0] ces_3_4_io_ins_left;
  wire [63:0] ces_3_4_io_outs_down;
  wire [63:0] ces_3_4_io_outs_right;
  wire [63:0] ces_3_4_io_outs_up;
  wire [63:0] ces_3_4_io_outs_left;
  wire  ces_3_4_io_lsbIns_1;
  wire  ces_3_4_io_lsbIns_2;
  wire  ces_3_4_io_lsbIns_3;
  wire  ces_3_4_io_lsbIns_4;
  wire  ces_3_4_io_lsbIns_5;
  wire  ces_3_4_io_lsbIns_6;
  wire  ces_3_4_io_lsbIns_7;
  wire  ces_3_4_io_lsbOuts_0;
  wire  ces_3_4_io_lsbOuts_1;
  wire  ces_3_4_io_lsbOuts_2;
  wire  ces_3_4_io_lsbOuts_3;
  wire  ces_3_4_io_lsbOuts_4;
  wire  ces_3_4_io_lsbOuts_5;
  wire  ces_3_4_io_lsbOuts_6;
  wire  ces_3_4_io_lsbOuts_7;
  wire  ces_3_5_clock;
  wire  ces_3_5_io_clockOutRight;
  wire [63:0] ces_3_5_io_ins_down;
  wire [63:0] ces_3_5_io_ins_right;
  wire [63:0] ces_3_5_io_ins_up;
  wire [63:0] ces_3_5_io_ins_left;
  wire [63:0] ces_3_5_io_outs_down;
  wire [63:0] ces_3_5_io_outs_right;
  wire [63:0] ces_3_5_io_outs_up;
  wire [63:0] ces_3_5_io_outs_left;
  wire  ces_3_5_io_lsbIns_1;
  wire  ces_3_5_io_lsbIns_2;
  wire  ces_3_5_io_lsbIns_3;
  wire  ces_3_5_io_lsbIns_4;
  wire  ces_3_5_io_lsbIns_5;
  wire  ces_3_5_io_lsbIns_6;
  wire  ces_3_5_io_lsbIns_7;
  wire  ces_3_5_io_lsbOuts_0;
  wire  ces_3_5_io_lsbOuts_1;
  wire  ces_3_5_io_lsbOuts_2;
  wire  ces_3_5_io_lsbOuts_3;
  wire  ces_3_5_io_lsbOuts_4;
  wire  ces_3_5_io_lsbOuts_5;
  wire  ces_3_5_io_lsbOuts_6;
  wire  ces_3_5_io_lsbOuts_7;
  wire  ces_3_6_clock;
  wire  ces_3_6_io_clockOutRight;
  wire [63:0] ces_3_6_io_ins_down;
  wire [63:0] ces_3_6_io_ins_right;
  wire [63:0] ces_3_6_io_ins_up;
  wire [63:0] ces_3_6_io_ins_left;
  wire [63:0] ces_3_6_io_outs_down;
  wire [63:0] ces_3_6_io_outs_right;
  wire [63:0] ces_3_6_io_outs_up;
  wire [63:0] ces_3_6_io_outs_left;
  wire  ces_3_6_io_lsbIns_1;
  wire  ces_3_6_io_lsbIns_2;
  wire  ces_3_6_io_lsbIns_3;
  wire  ces_3_6_io_lsbIns_4;
  wire  ces_3_6_io_lsbIns_5;
  wire  ces_3_6_io_lsbIns_6;
  wire  ces_3_6_io_lsbIns_7;
  wire  ces_3_6_io_lsbOuts_0;
  wire  ces_3_6_io_lsbOuts_1;
  wire  ces_3_6_io_lsbOuts_2;
  wire  ces_3_6_io_lsbOuts_3;
  wire  ces_3_6_io_lsbOuts_4;
  wire  ces_3_6_io_lsbOuts_5;
  wire  ces_3_6_io_lsbOuts_6;
  wire  ces_3_6_io_lsbOuts_7;
  wire  ces_3_7_clock;
  wire  ces_3_7_io_clockOutRight;
  wire [63:0] ces_3_7_io_ins_down;
  wire [63:0] ces_3_7_io_ins_right;
  wire [63:0] ces_3_7_io_ins_up;
  wire [63:0] ces_3_7_io_ins_left;
  wire [63:0] ces_3_7_io_outs_down;
  wire [63:0] ces_3_7_io_outs_right;
  wire [63:0] ces_3_7_io_outs_up;
  wire [63:0] ces_3_7_io_outs_left;
  wire  ces_3_7_io_lsbIns_1;
  wire  ces_3_7_io_lsbIns_2;
  wire  ces_3_7_io_lsbIns_3;
  wire  ces_3_7_io_lsbIns_4;
  wire  ces_3_7_io_lsbIns_5;
  wire  ces_3_7_io_lsbIns_6;
  wire  ces_3_7_io_lsbIns_7;
  wire  ces_3_7_io_lsbOuts_0;
  wire  ces_3_7_io_lsbOuts_1;
  wire  ces_3_7_io_lsbOuts_2;
  wire  ces_3_7_io_lsbOuts_3;
  wire  ces_3_7_io_lsbOuts_4;
  wire  ces_3_7_io_lsbOuts_5;
  wire  ces_3_7_io_lsbOuts_6;
  wire  ces_3_7_io_lsbOuts_7;
  wire  ces_4_0_clock;
  wire  ces_4_0_io_clockOutRight;
  wire [63:0] ces_4_0_io_ins_down;
  wire [63:0] ces_4_0_io_ins_right;
  wire [63:0] ces_4_0_io_ins_up;
  wire [63:0] ces_4_0_io_ins_left;
  wire [63:0] ces_4_0_io_outs_down;
  wire [63:0] ces_4_0_io_outs_right;
  wire [63:0] ces_4_0_io_outs_up;
  wire [63:0] ces_4_0_io_outs_left;
  wire  ces_4_0_io_lsbIns_1;
  wire  ces_4_0_io_lsbIns_2;
  wire  ces_4_0_io_lsbIns_3;
  wire  ces_4_0_io_lsbIns_4;
  wire  ces_4_0_io_lsbIns_5;
  wire  ces_4_0_io_lsbIns_6;
  wire  ces_4_0_io_lsbIns_7;
  wire  ces_4_0_io_lsbOuts_0;
  wire  ces_4_0_io_lsbOuts_1;
  wire  ces_4_0_io_lsbOuts_2;
  wire  ces_4_0_io_lsbOuts_3;
  wire  ces_4_0_io_lsbOuts_4;
  wire  ces_4_0_io_lsbOuts_5;
  wire  ces_4_0_io_lsbOuts_6;
  wire  ces_4_0_io_lsbOuts_7;
  wire  ces_4_1_clock;
  wire  ces_4_1_io_clockOutRight;
  wire [63:0] ces_4_1_io_ins_down;
  wire [63:0] ces_4_1_io_ins_right;
  wire [63:0] ces_4_1_io_ins_up;
  wire [63:0] ces_4_1_io_ins_left;
  wire [63:0] ces_4_1_io_outs_down;
  wire [63:0] ces_4_1_io_outs_right;
  wire [63:0] ces_4_1_io_outs_up;
  wire [63:0] ces_4_1_io_outs_left;
  wire  ces_4_1_io_lsbIns_1;
  wire  ces_4_1_io_lsbIns_2;
  wire  ces_4_1_io_lsbIns_3;
  wire  ces_4_1_io_lsbIns_4;
  wire  ces_4_1_io_lsbIns_5;
  wire  ces_4_1_io_lsbIns_6;
  wire  ces_4_1_io_lsbIns_7;
  wire  ces_4_1_io_lsbOuts_0;
  wire  ces_4_1_io_lsbOuts_1;
  wire  ces_4_1_io_lsbOuts_2;
  wire  ces_4_1_io_lsbOuts_3;
  wire  ces_4_1_io_lsbOuts_4;
  wire  ces_4_1_io_lsbOuts_5;
  wire  ces_4_1_io_lsbOuts_6;
  wire  ces_4_1_io_lsbOuts_7;
  wire  ces_4_2_clock;
  wire  ces_4_2_io_clockOutRight;
  wire [63:0] ces_4_2_io_ins_down;
  wire [63:0] ces_4_2_io_ins_right;
  wire [63:0] ces_4_2_io_ins_up;
  wire [63:0] ces_4_2_io_ins_left;
  wire [63:0] ces_4_2_io_outs_down;
  wire [63:0] ces_4_2_io_outs_right;
  wire [63:0] ces_4_2_io_outs_up;
  wire [63:0] ces_4_2_io_outs_left;
  wire  ces_4_2_io_lsbIns_1;
  wire  ces_4_2_io_lsbIns_2;
  wire  ces_4_2_io_lsbIns_3;
  wire  ces_4_2_io_lsbIns_4;
  wire  ces_4_2_io_lsbIns_5;
  wire  ces_4_2_io_lsbIns_6;
  wire  ces_4_2_io_lsbIns_7;
  wire  ces_4_2_io_lsbOuts_0;
  wire  ces_4_2_io_lsbOuts_1;
  wire  ces_4_2_io_lsbOuts_2;
  wire  ces_4_2_io_lsbOuts_3;
  wire  ces_4_2_io_lsbOuts_4;
  wire  ces_4_2_io_lsbOuts_5;
  wire  ces_4_2_io_lsbOuts_6;
  wire  ces_4_2_io_lsbOuts_7;
  wire  ces_4_3_clock;
  wire  ces_4_3_io_clockOutRight;
  wire [63:0] ces_4_3_io_ins_down;
  wire [63:0] ces_4_3_io_ins_right;
  wire [63:0] ces_4_3_io_ins_up;
  wire [63:0] ces_4_3_io_ins_left;
  wire [63:0] ces_4_3_io_outs_down;
  wire [63:0] ces_4_3_io_outs_right;
  wire [63:0] ces_4_3_io_outs_up;
  wire [63:0] ces_4_3_io_outs_left;
  wire  ces_4_3_io_lsbIns_1;
  wire  ces_4_3_io_lsbIns_2;
  wire  ces_4_3_io_lsbIns_3;
  wire  ces_4_3_io_lsbIns_4;
  wire  ces_4_3_io_lsbIns_5;
  wire  ces_4_3_io_lsbIns_6;
  wire  ces_4_3_io_lsbIns_7;
  wire  ces_4_3_io_lsbOuts_0;
  wire  ces_4_3_io_lsbOuts_1;
  wire  ces_4_3_io_lsbOuts_2;
  wire  ces_4_3_io_lsbOuts_3;
  wire  ces_4_3_io_lsbOuts_4;
  wire  ces_4_3_io_lsbOuts_5;
  wire  ces_4_3_io_lsbOuts_6;
  wire  ces_4_3_io_lsbOuts_7;
  wire  ces_4_4_clock;
  wire  ces_4_4_io_clockOutRight;
  wire [63:0] ces_4_4_io_ins_down;
  wire [63:0] ces_4_4_io_ins_right;
  wire [63:0] ces_4_4_io_ins_up;
  wire [63:0] ces_4_4_io_ins_left;
  wire [63:0] ces_4_4_io_outs_down;
  wire [63:0] ces_4_4_io_outs_right;
  wire [63:0] ces_4_4_io_outs_up;
  wire [63:0] ces_4_4_io_outs_left;
  wire  ces_4_4_io_lsbIns_1;
  wire  ces_4_4_io_lsbIns_2;
  wire  ces_4_4_io_lsbIns_3;
  wire  ces_4_4_io_lsbIns_4;
  wire  ces_4_4_io_lsbIns_5;
  wire  ces_4_4_io_lsbIns_6;
  wire  ces_4_4_io_lsbIns_7;
  wire  ces_4_4_io_lsbOuts_0;
  wire  ces_4_4_io_lsbOuts_1;
  wire  ces_4_4_io_lsbOuts_2;
  wire  ces_4_4_io_lsbOuts_3;
  wire  ces_4_4_io_lsbOuts_4;
  wire  ces_4_4_io_lsbOuts_5;
  wire  ces_4_4_io_lsbOuts_6;
  wire  ces_4_4_io_lsbOuts_7;
  wire  ces_4_5_clock;
  wire  ces_4_5_io_clockOutRight;
  wire [63:0] ces_4_5_io_ins_down;
  wire [63:0] ces_4_5_io_ins_right;
  wire [63:0] ces_4_5_io_ins_up;
  wire [63:0] ces_4_5_io_ins_left;
  wire [63:0] ces_4_5_io_outs_down;
  wire [63:0] ces_4_5_io_outs_right;
  wire [63:0] ces_4_5_io_outs_up;
  wire [63:0] ces_4_5_io_outs_left;
  wire  ces_4_5_io_lsbIns_1;
  wire  ces_4_5_io_lsbIns_2;
  wire  ces_4_5_io_lsbIns_3;
  wire  ces_4_5_io_lsbIns_4;
  wire  ces_4_5_io_lsbIns_5;
  wire  ces_4_5_io_lsbIns_6;
  wire  ces_4_5_io_lsbIns_7;
  wire  ces_4_5_io_lsbOuts_0;
  wire  ces_4_5_io_lsbOuts_1;
  wire  ces_4_5_io_lsbOuts_2;
  wire  ces_4_5_io_lsbOuts_3;
  wire  ces_4_5_io_lsbOuts_4;
  wire  ces_4_5_io_lsbOuts_5;
  wire  ces_4_5_io_lsbOuts_6;
  wire  ces_4_5_io_lsbOuts_7;
  wire  ces_4_6_clock;
  wire  ces_4_6_io_clockOutRight;
  wire [63:0] ces_4_6_io_ins_down;
  wire [63:0] ces_4_6_io_ins_right;
  wire [63:0] ces_4_6_io_ins_up;
  wire [63:0] ces_4_6_io_ins_left;
  wire [63:0] ces_4_6_io_outs_down;
  wire [63:0] ces_4_6_io_outs_right;
  wire [63:0] ces_4_6_io_outs_up;
  wire [63:0] ces_4_6_io_outs_left;
  wire  ces_4_6_io_lsbIns_1;
  wire  ces_4_6_io_lsbIns_2;
  wire  ces_4_6_io_lsbIns_3;
  wire  ces_4_6_io_lsbIns_4;
  wire  ces_4_6_io_lsbIns_5;
  wire  ces_4_6_io_lsbIns_6;
  wire  ces_4_6_io_lsbIns_7;
  wire  ces_4_6_io_lsbOuts_0;
  wire  ces_4_6_io_lsbOuts_1;
  wire  ces_4_6_io_lsbOuts_2;
  wire  ces_4_6_io_lsbOuts_3;
  wire  ces_4_6_io_lsbOuts_4;
  wire  ces_4_6_io_lsbOuts_5;
  wire  ces_4_6_io_lsbOuts_6;
  wire  ces_4_6_io_lsbOuts_7;
  wire  ces_4_7_clock;
  wire  ces_4_7_io_clockOutRight;
  wire [63:0] ces_4_7_io_ins_down;
  wire [63:0] ces_4_7_io_ins_right;
  wire [63:0] ces_4_7_io_ins_up;
  wire [63:0] ces_4_7_io_ins_left;
  wire [63:0] ces_4_7_io_outs_down;
  wire [63:0] ces_4_7_io_outs_right;
  wire [63:0] ces_4_7_io_outs_up;
  wire [63:0] ces_4_7_io_outs_left;
  wire  ces_4_7_io_lsbIns_1;
  wire  ces_4_7_io_lsbIns_2;
  wire  ces_4_7_io_lsbIns_3;
  wire  ces_4_7_io_lsbIns_4;
  wire  ces_4_7_io_lsbIns_5;
  wire  ces_4_7_io_lsbIns_6;
  wire  ces_4_7_io_lsbIns_7;
  wire  ces_4_7_io_lsbOuts_0;
  wire  ces_4_7_io_lsbOuts_1;
  wire  ces_4_7_io_lsbOuts_2;
  wire  ces_4_7_io_lsbOuts_3;
  wire  ces_4_7_io_lsbOuts_4;
  wire  ces_4_7_io_lsbOuts_5;
  wire  ces_4_7_io_lsbOuts_6;
  wire  ces_4_7_io_lsbOuts_7;
  wire  ces_5_0_clock;
  wire  ces_5_0_io_clockOutRight;
  wire [63:0] ces_5_0_io_ins_down;
  wire [63:0] ces_5_0_io_ins_right;
  wire [63:0] ces_5_0_io_ins_up;
  wire [63:0] ces_5_0_io_ins_left;
  wire [63:0] ces_5_0_io_outs_down;
  wire [63:0] ces_5_0_io_outs_right;
  wire [63:0] ces_5_0_io_outs_up;
  wire [63:0] ces_5_0_io_outs_left;
  wire  ces_5_0_io_lsbIns_1;
  wire  ces_5_0_io_lsbIns_2;
  wire  ces_5_0_io_lsbIns_3;
  wire  ces_5_0_io_lsbIns_4;
  wire  ces_5_0_io_lsbIns_5;
  wire  ces_5_0_io_lsbIns_6;
  wire  ces_5_0_io_lsbIns_7;
  wire  ces_5_0_io_lsbOuts_0;
  wire  ces_5_0_io_lsbOuts_1;
  wire  ces_5_0_io_lsbOuts_2;
  wire  ces_5_0_io_lsbOuts_3;
  wire  ces_5_0_io_lsbOuts_4;
  wire  ces_5_0_io_lsbOuts_5;
  wire  ces_5_0_io_lsbOuts_6;
  wire  ces_5_0_io_lsbOuts_7;
  wire  ces_5_1_clock;
  wire  ces_5_1_io_clockOutRight;
  wire [63:0] ces_5_1_io_ins_down;
  wire [63:0] ces_5_1_io_ins_right;
  wire [63:0] ces_5_1_io_ins_up;
  wire [63:0] ces_5_1_io_ins_left;
  wire [63:0] ces_5_1_io_outs_down;
  wire [63:0] ces_5_1_io_outs_right;
  wire [63:0] ces_5_1_io_outs_up;
  wire [63:0] ces_5_1_io_outs_left;
  wire  ces_5_1_io_lsbIns_1;
  wire  ces_5_1_io_lsbIns_2;
  wire  ces_5_1_io_lsbIns_3;
  wire  ces_5_1_io_lsbIns_4;
  wire  ces_5_1_io_lsbIns_5;
  wire  ces_5_1_io_lsbIns_6;
  wire  ces_5_1_io_lsbIns_7;
  wire  ces_5_1_io_lsbOuts_0;
  wire  ces_5_1_io_lsbOuts_1;
  wire  ces_5_1_io_lsbOuts_2;
  wire  ces_5_1_io_lsbOuts_3;
  wire  ces_5_1_io_lsbOuts_4;
  wire  ces_5_1_io_lsbOuts_5;
  wire  ces_5_1_io_lsbOuts_6;
  wire  ces_5_1_io_lsbOuts_7;
  wire  ces_5_2_clock;
  wire  ces_5_2_io_clockOutRight;
  wire [63:0] ces_5_2_io_ins_down;
  wire [63:0] ces_5_2_io_ins_right;
  wire [63:0] ces_5_2_io_ins_up;
  wire [63:0] ces_5_2_io_ins_left;
  wire [63:0] ces_5_2_io_outs_down;
  wire [63:0] ces_5_2_io_outs_right;
  wire [63:0] ces_5_2_io_outs_up;
  wire [63:0] ces_5_2_io_outs_left;
  wire  ces_5_2_io_lsbIns_1;
  wire  ces_5_2_io_lsbIns_2;
  wire  ces_5_2_io_lsbIns_3;
  wire  ces_5_2_io_lsbIns_4;
  wire  ces_5_2_io_lsbIns_5;
  wire  ces_5_2_io_lsbIns_6;
  wire  ces_5_2_io_lsbIns_7;
  wire  ces_5_2_io_lsbOuts_0;
  wire  ces_5_2_io_lsbOuts_1;
  wire  ces_5_2_io_lsbOuts_2;
  wire  ces_5_2_io_lsbOuts_3;
  wire  ces_5_2_io_lsbOuts_4;
  wire  ces_5_2_io_lsbOuts_5;
  wire  ces_5_2_io_lsbOuts_6;
  wire  ces_5_2_io_lsbOuts_7;
  wire  ces_5_3_clock;
  wire  ces_5_3_io_clockOutRight;
  wire [63:0] ces_5_3_io_ins_down;
  wire [63:0] ces_5_3_io_ins_right;
  wire [63:0] ces_5_3_io_ins_up;
  wire [63:0] ces_5_3_io_ins_left;
  wire [63:0] ces_5_3_io_outs_down;
  wire [63:0] ces_5_3_io_outs_right;
  wire [63:0] ces_5_3_io_outs_up;
  wire [63:0] ces_5_3_io_outs_left;
  wire  ces_5_3_io_lsbIns_1;
  wire  ces_5_3_io_lsbIns_2;
  wire  ces_5_3_io_lsbIns_3;
  wire  ces_5_3_io_lsbIns_4;
  wire  ces_5_3_io_lsbIns_5;
  wire  ces_5_3_io_lsbIns_6;
  wire  ces_5_3_io_lsbIns_7;
  wire  ces_5_3_io_lsbOuts_0;
  wire  ces_5_3_io_lsbOuts_1;
  wire  ces_5_3_io_lsbOuts_2;
  wire  ces_5_3_io_lsbOuts_3;
  wire  ces_5_3_io_lsbOuts_4;
  wire  ces_5_3_io_lsbOuts_5;
  wire  ces_5_3_io_lsbOuts_6;
  wire  ces_5_3_io_lsbOuts_7;
  wire  ces_5_4_clock;
  wire  ces_5_4_io_clockOutRight;
  wire [63:0] ces_5_4_io_ins_down;
  wire [63:0] ces_5_4_io_ins_right;
  wire [63:0] ces_5_4_io_ins_up;
  wire [63:0] ces_5_4_io_ins_left;
  wire [63:0] ces_5_4_io_outs_down;
  wire [63:0] ces_5_4_io_outs_right;
  wire [63:0] ces_5_4_io_outs_up;
  wire [63:0] ces_5_4_io_outs_left;
  wire  ces_5_4_io_lsbIns_1;
  wire  ces_5_4_io_lsbIns_2;
  wire  ces_5_4_io_lsbIns_3;
  wire  ces_5_4_io_lsbIns_4;
  wire  ces_5_4_io_lsbIns_5;
  wire  ces_5_4_io_lsbIns_6;
  wire  ces_5_4_io_lsbIns_7;
  wire  ces_5_4_io_lsbOuts_0;
  wire  ces_5_4_io_lsbOuts_1;
  wire  ces_5_4_io_lsbOuts_2;
  wire  ces_5_4_io_lsbOuts_3;
  wire  ces_5_4_io_lsbOuts_4;
  wire  ces_5_4_io_lsbOuts_5;
  wire  ces_5_4_io_lsbOuts_6;
  wire  ces_5_4_io_lsbOuts_7;
  wire  ces_5_5_clock;
  wire  ces_5_5_io_clockOutRight;
  wire [63:0] ces_5_5_io_ins_down;
  wire [63:0] ces_5_5_io_ins_right;
  wire [63:0] ces_5_5_io_ins_up;
  wire [63:0] ces_5_5_io_ins_left;
  wire [63:0] ces_5_5_io_outs_down;
  wire [63:0] ces_5_5_io_outs_right;
  wire [63:0] ces_5_5_io_outs_up;
  wire [63:0] ces_5_5_io_outs_left;
  wire  ces_5_5_io_lsbIns_1;
  wire  ces_5_5_io_lsbIns_2;
  wire  ces_5_5_io_lsbIns_3;
  wire  ces_5_5_io_lsbIns_4;
  wire  ces_5_5_io_lsbIns_5;
  wire  ces_5_5_io_lsbIns_6;
  wire  ces_5_5_io_lsbIns_7;
  wire  ces_5_5_io_lsbOuts_0;
  wire  ces_5_5_io_lsbOuts_1;
  wire  ces_5_5_io_lsbOuts_2;
  wire  ces_5_5_io_lsbOuts_3;
  wire  ces_5_5_io_lsbOuts_4;
  wire  ces_5_5_io_lsbOuts_5;
  wire  ces_5_5_io_lsbOuts_6;
  wire  ces_5_5_io_lsbOuts_7;
  wire  ces_5_6_clock;
  wire  ces_5_6_io_clockOutRight;
  wire [63:0] ces_5_6_io_ins_down;
  wire [63:0] ces_5_6_io_ins_right;
  wire [63:0] ces_5_6_io_ins_up;
  wire [63:0] ces_5_6_io_ins_left;
  wire [63:0] ces_5_6_io_outs_down;
  wire [63:0] ces_5_6_io_outs_right;
  wire [63:0] ces_5_6_io_outs_up;
  wire [63:0] ces_5_6_io_outs_left;
  wire  ces_5_6_io_lsbIns_1;
  wire  ces_5_6_io_lsbIns_2;
  wire  ces_5_6_io_lsbIns_3;
  wire  ces_5_6_io_lsbIns_4;
  wire  ces_5_6_io_lsbIns_5;
  wire  ces_5_6_io_lsbIns_6;
  wire  ces_5_6_io_lsbIns_7;
  wire  ces_5_6_io_lsbOuts_0;
  wire  ces_5_6_io_lsbOuts_1;
  wire  ces_5_6_io_lsbOuts_2;
  wire  ces_5_6_io_lsbOuts_3;
  wire  ces_5_6_io_lsbOuts_4;
  wire  ces_5_6_io_lsbOuts_5;
  wire  ces_5_6_io_lsbOuts_6;
  wire  ces_5_6_io_lsbOuts_7;
  wire  ces_5_7_clock;
  wire  ces_5_7_io_clockOutRight;
  wire [63:0] ces_5_7_io_ins_down;
  wire [63:0] ces_5_7_io_ins_right;
  wire [63:0] ces_5_7_io_ins_up;
  wire [63:0] ces_5_7_io_ins_left;
  wire [63:0] ces_5_7_io_outs_down;
  wire [63:0] ces_5_7_io_outs_right;
  wire [63:0] ces_5_7_io_outs_up;
  wire [63:0] ces_5_7_io_outs_left;
  wire  ces_5_7_io_lsbIns_1;
  wire  ces_5_7_io_lsbIns_2;
  wire  ces_5_7_io_lsbIns_3;
  wire  ces_5_7_io_lsbIns_4;
  wire  ces_5_7_io_lsbIns_5;
  wire  ces_5_7_io_lsbIns_6;
  wire  ces_5_7_io_lsbIns_7;
  wire  ces_5_7_io_lsbOuts_0;
  wire  ces_5_7_io_lsbOuts_1;
  wire  ces_5_7_io_lsbOuts_2;
  wire  ces_5_7_io_lsbOuts_3;
  wire  ces_5_7_io_lsbOuts_4;
  wire  ces_5_7_io_lsbOuts_5;
  wire  ces_5_7_io_lsbOuts_6;
  wire  ces_5_7_io_lsbOuts_7;
  wire  ces_6_0_clock;
  wire  ces_6_0_io_clockOutRight;
  wire [63:0] ces_6_0_io_ins_down;
  wire [63:0] ces_6_0_io_ins_right;
  wire [63:0] ces_6_0_io_ins_up;
  wire [63:0] ces_6_0_io_ins_left;
  wire [63:0] ces_6_0_io_outs_down;
  wire [63:0] ces_6_0_io_outs_right;
  wire [63:0] ces_6_0_io_outs_up;
  wire [63:0] ces_6_0_io_outs_left;
  wire  ces_6_0_io_lsbIns_1;
  wire  ces_6_0_io_lsbIns_2;
  wire  ces_6_0_io_lsbIns_3;
  wire  ces_6_0_io_lsbIns_4;
  wire  ces_6_0_io_lsbIns_5;
  wire  ces_6_0_io_lsbIns_6;
  wire  ces_6_0_io_lsbIns_7;
  wire  ces_6_0_io_lsbOuts_0;
  wire  ces_6_0_io_lsbOuts_1;
  wire  ces_6_0_io_lsbOuts_2;
  wire  ces_6_0_io_lsbOuts_3;
  wire  ces_6_0_io_lsbOuts_4;
  wire  ces_6_0_io_lsbOuts_5;
  wire  ces_6_0_io_lsbOuts_6;
  wire  ces_6_0_io_lsbOuts_7;
  wire  ces_6_1_clock;
  wire  ces_6_1_io_clockOutRight;
  wire [63:0] ces_6_1_io_ins_down;
  wire [63:0] ces_6_1_io_ins_right;
  wire [63:0] ces_6_1_io_ins_up;
  wire [63:0] ces_6_1_io_ins_left;
  wire [63:0] ces_6_1_io_outs_down;
  wire [63:0] ces_6_1_io_outs_right;
  wire [63:0] ces_6_1_io_outs_up;
  wire [63:0] ces_6_1_io_outs_left;
  wire  ces_6_1_io_lsbIns_1;
  wire  ces_6_1_io_lsbIns_2;
  wire  ces_6_1_io_lsbIns_3;
  wire  ces_6_1_io_lsbIns_4;
  wire  ces_6_1_io_lsbIns_5;
  wire  ces_6_1_io_lsbIns_6;
  wire  ces_6_1_io_lsbIns_7;
  wire  ces_6_1_io_lsbOuts_0;
  wire  ces_6_1_io_lsbOuts_1;
  wire  ces_6_1_io_lsbOuts_2;
  wire  ces_6_1_io_lsbOuts_3;
  wire  ces_6_1_io_lsbOuts_4;
  wire  ces_6_1_io_lsbOuts_5;
  wire  ces_6_1_io_lsbOuts_6;
  wire  ces_6_1_io_lsbOuts_7;
  wire  ces_6_2_clock;
  wire  ces_6_2_io_clockOutRight;
  wire [63:0] ces_6_2_io_ins_down;
  wire [63:0] ces_6_2_io_ins_right;
  wire [63:0] ces_6_2_io_ins_up;
  wire [63:0] ces_6_2_io_ins_left;
  wire [63:0] ces_6_2_io_outs_down;
  wire [63:0] ces_6_2_io_outs_right;
  wire [63:0] ces_6_2_io_outs_up;
  wire [63:0] ces_6_2_io_outs_left;
  wire  ces_6_2_io_lsbIns_1;
  wire  ces_6_2_io_lsbIns_2;
  wire  ces_6_2_io_lsbIns_3;
  wire  ces_6_2_io_lsbIns_4;
  wire  ces_6_2_io_lsbIns_5;
  wire  ces_6_2_io_lsbIns_6;
  wire  ces_6_2_io_lsbIns_7;
  wire  ces_6_2_io_lsbOuts_0;
  wire  ces_6_2_io_lsbOuts_1;
  wire  ces_6_2_io_lsbOuts_2;
  wire  ces_6_2_io_lsbOuts_3;
  wire  ces_6_2_io_lsbOuts_4;
  wire  ces_6_2_io_lsbOuts_5;
  wire  ces_6_2_io_lsbOuts_6;
  wire  ces_6_2_io_lsbOuts_7;
  wire  ces_6_3_clock;
  wire  ces_6_3_io_clockOutRight;
  wire [63:0] ces_6_3_io_ins_down;
  wire [63:0] ces_6_3_io_ins_right;
  wire [63:0] ces_6_3_io_ins_up;
  wire [63:0] ces_6_3_io_ins_left;
  wire [63:0] ces_6_3_io_outs_down;
  wire [63:0] ces_6_3_io_outs_right;
  wire [63:0] ces_6_3_io_outs_up;
  wire [63:0] ces_6_3_io_outs_left;
  wire  ces_6_3_io_lsbIns_1;
  wire  ces_6_3_io_lsbIns_2;
  wire  ces_6_3_io_lsbIns_3;
  wire  ces_6_3_io_lsbIns_4;
  wire  ces_6_3_io_lsbIns_5;
  wire  ces_6_3_io_lsbIns_6;
  wire  ces_6_3_io_lsbIns_7;
  wire  ces_6_3_io_lsbOuts_0;
  wire  ces_6_3_io_lsbOuts_1;
  wire  ces_6_3_io_lsbOuts_2;
  wire  ces_6_3_io_lsbOuts_3;
  wire  ces_6_3_io_lsbOuts_4;
  wire  ces_6_3_io_lsbOuts_5;
  wire  ces_6_3_io_lsbOuts_6;
  wire  ces_6_3_io_lsbOuts_7;
  wire  ces_6_4_clock;
  wire  ces_6_4_io_clockOutRight;
  wire [63:0] ces_6_4_io_ins_down;
  wire [63:0] ces_6_4_io_ins_right;
  wire [63:0] ces_6_4_io_ins_up;
  wire [63:0] ces_6_4_io_ins_left;
  wire [63:0] ces_6_4_io_outs_down;
  wire [63:0] ces_6_4_io_outs_right;
  wire [63:0] ces_6_4_io_outs_up;
  wire [63:0] ces_6_4_io_outs_left;
  wire  ces_6_4_io_lsbIns_1;
  wire  ces_6_4_io_lsbIns_2;
  wire  ces_6_4_io_lsbIns_3;
  wire  ces_6_4_io_lsbIns_4;
  wire  ces_6_4_io_lsbIns_5;
  wire  ces_6_4_io_lsbIns_6;
  wire  ces_6_4_io_lsbIns_7;
  wire  ces_6_4_io_lsbOuts_0;
  wire  ces_6_4_io_lsbOuts_1;
  wire  ces_6_4_io_lsbOuts_2;
  wire  ces_6_4_io_lsbOuts_3;
  wire  ces_6_4_io_lsbOuts_4;
  wire  ces_6_4_io_lsbOuts_5;
  wire  ces_6_4_io_lsbOuts_6;
  wire  ces_6_4_io_lsbOuts_7;
  wire  ces_6_5_clock;
  wire  ces_6_5_io_clockOutRight;
  wire [63:0] ces_6_5_io_ins_down;
  wire [63:0] ces_6_5_io_ins_right;
  wire [63:0] ces_6_5_io_ins_up;
  wire [63:0] ces_6_5_io_ins_left;
  wire [63:0] ces_6_5_io_outs_down;
  wire [63:0] ces_6_5_io_outs_right;
  wire [63:0] ces_6_5_io_outs_up;
  wire [63:0] ces_6_5_io_outs_left;
  wire  ces_6_5_io_lsbIns_1;
  wire  ces_6_5_io_lsbIns_2;
  wire  ces_6_5_io_lsbIns_3;
  wire  ces_6_5_io_lsbIns_4;
  wire  ces_6_5_io_lsbIns_5;
  wire  ces_6_5_io_lsbIns_6;
  wire  ces_6_5_io_lsbIns_7;
  wire  ces_6_5_io_lsbOuts_0;
  wire  ces_6_5_io_lsbOuts_1;
  wire  ces_6_5_io_lsbOuts_2;
  wire  ces_6_5_io_lsbOuts_3;
  wire  ces_6_5_io_lsbOuts_4;
  wire  ces_6_5_io_lsbOuts_5;
  wire  ces_6_5_io_lsbOuts_6;
  wire  ces_6_5_io_lsbOuts_7;
  wire  ces_6_6_clock;
  wire  ces_6_6_io_clockOutRight;
  wire [63:0] ces_6_6_io_ins_down;
  wire [63:0] ces_6_6_io_ins_right;
  wire [63:0] ces_6_6_io_ins_up;
  wire [63:0] ces_6_6_io_ins_left;
  wire [63:0] ces_6_6_io_outs_down;
  wire [63:0] ces_6_6_io_outs_right;
  wire [63:0] ces_6_6_io_outs_up;
  wire [63:0] ces_6_6_io_outs_left;
  wire  ces_6_6_io_lsbIns_1;
  wire  ces_6_6_io_lsbIns_2;
  wire  ces_6_6_io_lsbIns_3;
  wire  ces_6_6_io_lsbIns_4;
  wire  ces_6_6_io_lsbIns_5;
  wire  ces_6_6_io_lsbIns_6;
  wire  ces_6_6_io_lsbIns_7;
  wire  ces_6_6_io_lsbOuts_0;
  wire  ces_6_6_io_lsbOuts_1;
  wire  ces_6_6_io_lsbOuts_2;
  wire  ces_6_6_io_lsbOuts_3;
  wire  ces_6_6_io_lsbOuts_4;
  wire  ces_6_6_io_lsbOuts_5;
  wire  ces_6_6_io_lsbOuts_6;
  wire  ces_6_6_io_lsbOuts_7;
  wire  ces_6_7_clock;
  wire  ces_6_7_io_clockOutRight;
  wire [63:0] ces_6_7_io_ins_down;
  wire [63:0] ces_6_7_io_ins_right;
  wire [63:0] ces_6_7_io_ins_up;
  wire [63:0] ces_6_7_io_ins_left;
  wire [63:0] ces_6_7_io_outs_down;
  wire [63:0] ces_6_7_io_outs_right;
  wire [63:0] ces_6_7_io_outs_up;
  wire [63:0] ces_6_7_io_outs_left;
  wire  ces_6_7_io_lsbIns_1;
  wire  ces_6_7_io_lsbIns_2;
  wire  ces_6_7_io_lsbIns_3;
  wire  ces_6_7_io_lsbIns_4;
  wire  ces_6_7_io_lsbIns_5;
  wire  ces_6_7_io_lsbIns_6;
  wire  ces_6_7_io_lsbIns_7;
  wire  ces_6_7_io_lsbOuts_0;
  wire  ces_6_7_io_lsbOuts_1;
  wire  ces_6_7_io_lsbOuts_2;
  wire  ces_6_7_io_lsbOuts_3;
  wire  ces_6_7_io_lsbOuts_4;
  wire  ces_6_7_io_lsbOuts_5;
  wire  ces_6_7_io_lsbOuts_6;
  wire  ces_6_7_io_lsbOuts_7;
  wire  ces_7_0_clock;
  wire  ces_7_0_io_clockOutRight;
  wire [63:0] ces_7_0_io_ins_down;
  wire [63:0] ces_7_0_io_ins_right;
  wire [63:0] ces_7_0_io_ins_up;
  wire [63:0] ces_7_0_io_ins_left;
  wire [63:0] ces_7_0_io_outs_down;
  wire [63:0] ces_7_0_io_outs_right;
  wire [63:0] ces_7_0_io_outs_up;
  wire [63:0] ces_7_0_io_outs_left;
  wire  ces_7_0_io_lsbIns_1;
  wire  ces_7_0_io_lsbIns_2;
  wire  ces_7_0_io_lsbIns_3;
  wire  ces_7_0_io_lsbIns_4;
  wire  ces_7_0_io_lsbIns_5;
  wire  ces_7_0_io_lsbIns_6;
  wire  ces_7_0_io_lsbIns_7;
  wire  ces_7_0_io_lsbOuts_0;
  wire  ces_7_0_io_lsbOuts_1;
  wire  ces_7_0_io_lsbOuts_2;
  wire  ces_7_0_io_lsbOuts_3;
  wire  ces_7_0_io_lsbOuts_4;
  wire  ces_7_0_io_lsbOuts_5;
  wire  ces_7_0_io_lsbOuts_6;
  wire  ces_7_0_io_lsbOuts_7;
  wire  ces_7_1_clock;
  wire  ces_7_1_io_clockOutRight;
  wire [63:0] ces_7_1_io_ins_down;
  wire [63:0] ces_7_1_io_ins_right;
  wire [63:0] ces_7_1_io_ins_up;
  wire [63:0] ces_7_1_io_ins_left;
  wire [63:0] ces_7_1_io_outs_down;
  wire [63:0] ces_7_1_io_outs_right;
  wire [63:0] ces_7_1_io_outs_up;
  wire [63:0] ces_7_1_io_outs_left;
  wire  ces_7_1_io_lsbIns_1;
  wire  ces_7_1_io_lsbIns_2;
  wire  ces_7_1_io_lsbIns_3;
  wire  ces_7_1_io_lsbIns_4;
  wire  ces_7_1_io_lsbIns_5;
  wire  ces_7_1_io_lsbIns_6;
  wire  ces_7_1_io_lsbIns_7;
  wire  ces_7_1_io_lsbOuts_0;
  wire  ces_7_1_io_lsbOuts_1;
  wire  ces_7_1_io_lsbOuts_2;
  wire  ces_7_1_io_lsbOuts_3;
  wire  ces_7_1_io_lsbOuts_4;
  wire  ces_7_1_io_lsbOuts_5;
  wire  ces_7_1_io_lsbOuts_6;
  wire  ces_7_1_io_lsbOuts_7;
  wire  ces_7_2_clock;
  wire  ces_7_2_io_clockOutRight;
  wire [63:0] ces_7_2_io_ins_down;
  wire [63:0] ces_7_2_io_ins_right;
  wire [63:0] ces_7_2_io_ins_up;
  wire [63:0] ces_7_2_io_ins_left;
  wire [63:0] ces_7_2_io_outs_down;
  wire [63:0] ces_7_2_io_outs_right;
  wire [63:0] ces_7_2_io_outs_up;
  wire [63:0] ces_7_2_io_outs_left;
  wire  ces_7_2_io_lsbIns_1;
  wire  ces_7_2_io_lsbIns_2;
  wire  ces_7_2_io_lsbIns_3;
  wire  ces_7_2_io_lsbIns_4;
  wire  ces_7_2_io_lsbIns_5;
  wire  ces_7_2_io_lsbIns_6;
  wire  ces_7_2_io_lsbIns_7;
  wire  ces_7_2_io_lsbOuts_0;
  wire  ces_7_2_io_lsbOuts_1;
  wire  ces_7_2_io_lsbOuts_2;
  wire  ces_7_2_io_lsbOuts_3;
  wire  ces_7_2_io_lsbOuts_4;
  wire  ces_7_2_io_lsbOuts_5;
  wire  ces_7_2_io_lsbOuts_6;
  wire  ces_7_2_io_lsbOuts_7;
  wire  ces_7_3_clock;
  wire  ces_7_3_io_clockOutRight;
  wire [63:0] ces_7_3_io_ins_down;
  wire [63:0] ces_7_3_io_ins_right;
  wire [63:0] ces_7_3_io_ins_up;
  wire [63:0] ces_7_3_io_ins_left;
  wire [63:0] ces_7_3_io_outs_down;
  wire [63:0] ces_7_3_io_outs_right;
  wire [63:0] ces_7_3_io_outs_up;
  wire [63:0] ces_7_3_io_outs_left;
  wire  ces_7_3_io_lsbIns_1;
  wire  ces_7_3_io_lsbIns_2;
  wire  ces_7_3_io_lsbIns_3;
  wire  ces_7_3_io_lsbIns_4;
  wire  ces_7_3_io_lsbIns_5;
  wire  ces_7_3_io_lsbIns_6;
  wire  ces_7_3_io_lsbIns_7;
  wire  ces_7_3_io_lsbOuts_0;
  wire  ces_7_3_io_lsbOuts_1;
  wire  ces_7_3_io_lsbOuts_2;
  wire  ces_7_3_io_lsbOuts_3;
  wire  ces_7_3_io_lsbOuts_4;
  wire  ces_7_3_io_lsbOuts_5;
  wire  ces_7_3_io_lsbOuts_6;
  wire  ces_7_3_io_lsbOuts_7;
  wire  ces_7_4_clock;
  wire  ces_7_4_io_clockOutRight;
  wire [63:0] ces_7_4_io_ins_down;
  wire [63:0] ces_7_4_io_ins_right;
  wire [63:0] ces_7_4_io_ins_up;
  wire [63:0] ces_7_4_io_ins_left;
  wire [63:0] ces_7_4_io_outs_down;
  wire [63:0] ces_7_4_io_outs_right;
  wire [63:0] ces_7_4_io_outs_up;
  wire [63:0] ces_7_4_io_outs_left;
  wire  ces_7_4_io_lsbIns_1;
  wire  ces_7_4_io_lsbIns_2;
  wire  ces_7_4_io_lsbIns_3;
  wire  ces_7_4_io_lsbIns_4;
  wire  ces_7_4_io_lsbIns_5;
  wire  ces_7_4_io_lsbIns_6;
  wire  ces_7_4_io_lsbIns_7;
  wire  ces_7_4_io_lsbOuts_0;
  wire  ces_7_4_io_lsbOuts_1;
  wire  ces_7_4_io_lsbOuts_2;
  wire  ces_7_4_io_lsbOuts_3;
  wire  ces_7_4_io_lsbOuts_4;
  wire  ces_7_4_io_lsbOuts_5;
  wire  ces_7_4_io_lsbOuts_6;
  wire  ces_7_4_io_lsbOuts_7;
  wire  ces_7_5_clock;
  wire  ces_7_5_io_clockOutRight;
  wire [63:0] ces_7_5_io_ins_down;
  wire [63:0] ces_7_5_io_ins_right;
  wire [63:0] ces_7_5_io_ins_up;
  wire [63:0] ces_7_5_io_ins_left;
  wire [63:0] ces_7_5_io_outs_down;
  wire [63:0] ces_7_5_io_outs_right;
  wire [63:0] ces_7_5_io_outs_up;
  wire [63:0] ces_7_5_io_outs_left;
  wire  ces_7_5_io_lsbIns_1;
  wire  ces_7_5_io_lsbIns_2;
  wire  ces_7_5_io_lsbIns_3;
  wire  ces_7_5_io_lsbIns_4;
  wire  ces_7_5_io_lsbIns_5;
  wire  ces_7_5_io_lsbIns_6;
  wire  ces_7_5_io_lsbIns_7;
  wire  ces_7_5_io_lsbOuts_0;
  wire  ces_7_5_io_lsbOuts_1;
  wire  ces_7_5_io_lsbOuts_2;
  wire  ces_7_5_io_lsbOuts_3;
  wire  ces_7_5_io_lsbOuts_4;
  wire  ces_7_5_io_lsbOuts_5;
  wire  ces_7_5_io_lsbOuts_6;
  wire  ces_7_5_io_lsbOuts_7;
  wire  ces_7_6_clock;
  wire  ces_7_6_io_clockOutRight;
  wire [63:0] ces_7_6_io_ins_down;
  wire [63:0] ces_7_6_io_ins_right;
  wire [63:0] ces_7_6_io_ins_up;
  wire [63:0] ces_7_6_io_ins_left;
  wire [63:0] ces_7_6_io_outs_down;
  wire [63:0] ces_7_6_io_outs_right;
  wire [63:0] ces_7_6_io_outs_up;
  wire [63:0] ces_7_6_io_outs_left;
  wire  ces_7_6_io_lsbIns_1;
  wire  ces_7_6_io_lsbIns_2;
  wire  ces_7_6_io_lsbIns_3;
  wire  ces_7_6_io_lsbIns_4;
  wire  ces_7_6_io_lsbIns_5;
  wire  ces_7_6_io_lsbIns_6;
  wire  ces_7_6_io_lsbIns_7;
  wire  ces_7_6_io_lsbOuts_0;
  wire  ces_7_6_io_lsbOuts_1;
  wire  ces_7_6_io_lsbOuts_2;
  wire  ces_7_6_io_lsbOuts_3;
  wire  ces_7_6_io_lsbOuts_4;
  wire  ces_7_6_io_lsbOuts_5;
  wire  ces_7_6_io_lsbOuts_6;
  wire  ces_7_6_io_lsbOuts_7;
  wire  ces_7_7_clock;
  wire  ces_7_7_io_clockOutRight;
  wire [63:0] ces_7_7_io_ins_down;
  wire [63:0] ces_7_7_io_ins_right;
  wire [63:0] ces_7_7_io_ins_up;
  wire [63:0] ces_7_7_io_ins_left;
  wire [63:0] ces_7_7_io_outs_down;
  wire [63:0] ces_7_7_io_outs_right;
  wire [63:0] ces_7_7_io_outs_up;
  wire [63:0] ces_7_7_io_outs_left;
  wire  ces_7_7_io_lsbIns_1;
  wire  ces_7_7_io_lsbIns_2;
  wire  ces_7_7_io_lsbIns_3;
  wire  ces_7_7_io_lsbIns_4;
  wire  ces_7_7_io_lsbIns_5;
  wire  ces_7_7_io_lsbIns_6;
  wire  ces_7_7_io_lsbIns_7;
  wire  ces_7_7_io_lsbOuts_0;
  wire  ces_7_7_io_lsbOuts_1;
  wire  ces_7_7_io_lsbOuts_2;
  wire  ces_7_7_io_lsbOuts_3;
  wire  ces_7_7_io_lsbOuts_4;
  wire  ces_7_7_io_lsbOuts_5;
  wire  ces_7_7_io_lsbOuts_6;
  wire  ces_7_7_io_lsbOuts_7;
  reg  REG_0;
  reg  REG_1;
  reg  REG_2;
  reg  REG_3;
  reg  REG_4;
  reg  REG_5;
  reg  REG_6;
  reg  REG_7;
  reg  REG_8;
  reg  REG_9;
  reg  REG_10;
  reg  REG_11;
  reg  REG_12;
  reg  REG_13;
  reg  REG_14;
  reg  REG_15;
  reg  REG_16;
  reg  REG_17;
  reg  REG_18;
  reg  REG_19;
  reg  REG_20;
  reg  REG_21;
  reg  REG_22;
  reg  REG_23;
  reg  REG_24;
  reg  REG_25;
  reg  REG_26;
  reg  REG_27;
  reg  REG_28;
  reg  REG_29;
  reg  REG_30;
  reg  REG_31;
  reg  REG_32;
  reg  REG_33;
  reg  REG_34;
  reg  REG_35;
  reg  REG_36;
  reg  REG_37;
  reg  REG_38;
  reg  REG_39;
  reg  REG_40;
  reg  REG_41;
  reg  REG_42;
  reg  REG_43;
  reg  REG_44;
  reg  REG_45;
  reg  REG_46;
  reg  REG_47;
  reg  REG_48;
  reg  REG_49;
  reg  REG_50;
  reg  REG_51;
  reg  REG_52;
  reg  REG_53;
  reg  REG_54;
  reg  REG_55;
  reg  REG_56;
  reg  REG_57;
  reg  REG_58;
  reg  REG_59;
  reg  REG_60;
  reg  REG_61;
  reg  REG_62;
  reg  REG_63;
  Element ces_0_0 (
    .clock(ces_0_0_clock),
    .io_clockOutRight(ces_0_0_io_clockOutRight),
    .io_ins_down(ces_0_0_io_ins_down),
    .io_ins_right(ces_0_0_io_ins_right),
    .io_ins_up(ces_0_0_io_ins_up),
    .io_ins_left(ces_0_0_io_ins_left),
    .io_outs_down(ces_0_0_io_outs_down),
    .io_outs_right(ces_0_0_io_outs_right),
    .io_outs_up(ces_0_0_io_outs_up),
    .io_outs_left(ces_0_0_io_outs_left),
    .io_lsbIns_1(ces_0_0_io_lsbIns_1),
    .io_lsbIns_2(ces_0_0_io_lsbIns_2),
    .io_lsbIns_3(ces_0_0_io_lsbIns_3),
    .io_lsbIns_4(ces_0_0_io_lsbIns_4),
    .io_lsbIns_5(ces_0_0_io_lsbIns_5),
    .io_lsbIns_6(ces_0_0_io_lsbIns_6),
    .io_lsbIns_7(ces_0_0_io_lsbIns_7),
    .io_lsbOuts_0(ces_0_0_io_lsbOuts_0),
    .io_lsbOuts_1(ces_0_0_io_lsbOuts_1),
    .io_lsbOuts_2(ces_0_0_io_lsbOuts_2),
    .io_lsbOuts_3(ces_0_0_io_lsbOuts_3),
    .io_lsbOuts_4(ces_0_0_io_lsbOuts_4),
    .io_lsbOuts_5(ces_0_0_io_lsbOuts_5),
    .io_lsbOuts_6(ces_0_0_io_lsbOuts_6),
    .io_lsbOuts_7(ces_0_0_io_lsbOuts_7)
  );
  Element ces_0_1 (
    .clock(ces_0_1_clock),
    .io_clockOutRight(ces_0_1_io_clockOutRight),
    .io_ins_down(ces_0_1_io_ins_down),
    .io_ins_right(ces_0_1_io_ins_right),
    .io_ins_up(ces_0_1_io_ins_up),
    .io_ins_left(ces_0_1_io_ins_left),
    .io_outs_down(ces_0_1_io_outs_down),
    .io_outs_right(ces_0_1_io_outs_right),
    .io_outs_up(ces_0_1_io_outs_up),
    .io_outs_left(ces_0_1_io_outs_left),
    .io_lsbIns_1(ces_0_1_io_lsbIns_1),
    .io_lsbIns_2(ces_0_1_io_lsbIns_2),
    .io_lsbIns_3(ces_0_1_io_lsbIns_3),
    .io_lsbIns_4(ces_0_1_io_lsbIns_4),
    .io_lsbIns_5(ces_0_1_io_lsbIns_5),
    .io_lsbIns_6(ces_0_1_io_lsbIns_6),
    .io_lsbIns_7(ces_0_1_io_lsbIns_7),
    .io_lsbOuts_0(ces_0_1_io_lsbOuts_0),
    .io_lsbOuts_1(ces_0_1_io_lsbOuts_1),
    .io_lsbOuts_2(ces_0_1_io_lsbOuts_2),
    .io_lsbOuts_3(ces_0_1_io_lsbOuts_3),
    .io_lsbOuts_4(ces_0_1_io_lsbOuts_4),
    .io_lsbOuts_5(ces_0_1_io_lsbOuts_5),
    .io_lsbOuts_6(ces_0_1_io_lsbOuts_6),
    .io_lsbOuts_7(ces_0_1_io_lsbOuts_7)
  );
  Element ces_0_2 (
    .clock(ces_0_2_clock),
    .io_clockOutRight(ces_0_2_io_clockOutRight),
    .io_ins_down(ces_0_2_io_ins_down),
    .io_ins_right(ces_0_2_io_ins_right),
    .io_ins_up(ces_0_2_io_ins_up),
    .io_ins_left(ces_0_2_io_ins_left),
    .io_outs_down(ces_0_2_io_outs_down),
    .io_outs_right(ces_0_2_io_outs_right),
    .io_outs_up(ces_0_2_io_outs_up),
    .io_outs_left(ces_0_2_io_outs_left),
    .io_lsbIns_1(ces_0_2_io_lsbIns_1),
    .io_lsbIns_2(ces_0_2_io_lsbIns_2),
    .io_lsbIns_3(ces_0_2_io_lsbIns_3),
    .io_lsbIns_4(ces_0_2_io_lsbIns_4),
    .io_lsbIns_5(ces_0_2_io_lsbIns_5),
    .io_lsbIns_6(ces_0_2_io_lsbIns_6),
    .io_lsbIns_7(ces_0_2_io_lsbIns_7),
    .io_lsbOuts_0(ces_0_2_io_lsbOuts_0),
    .io_lsbOuts_1(ces_0_2_io_lsbOuts_1),
    .io_lsbOuts_2(ces_0_2_io_lsbOuts_2),
    .io_lsbOuts_3(ces_0_2_io_lsbOuts_3),
    .io_lsbOuts_4(ces_0_2_io_lsbOuts_4),
    .io_lsbOuts_5(ces_0_2_io_lsbOuts_5),
    .io_lsbOuts_6(ces_0_2_io_lsbOuts_6),
    .io_lsbOuts_7(ces_0_2_io_lsbOuts_7)
  );
  Element ces_0_3 (
    .clock(ces_0_3_clock),
    .io_clockOutRight(ces_0_3_io_clockOutRight),
    .io_ins_down(ces_0_3_io_ins_down),
    .io_ins_right(ces_0_3_io_ins_right),
    .io_ins_up(ces_0_3_io_ins_up),
    .io_ins_left(ces_0_3_io_ins_left),
    .io_outs_down(ces_0_3_io_outs_down),
    .io_outs_right(ces_0_3_io_outs_right),
    .io_outs_up(ces_0_3_io_outs_up),
    .io_outs_left(ces_0_3_io_outs_left),
    .io_lsbIns_1(ces_0_3_io_lsbIns_1),
    .io_lsbIns_2(ces_0_3_io_lsbIns_2),
    .io_lsbIns_3(ces_0_3_io_lsbIns_3),
    .io_lsbIns_4(ces_0_3_io_lsbIns_4),
    .io_lsbIns_5(ces_0_3_io_lsbIns_5),
    .io_lsbIns_6(ces_0_3_io_lsbIns_6),
    .io_lsbIns_7(ces_0_3_io_lsbIns_7),
    .io_lsbOuts_0(ces_0_3_io_lsbOuts_0),
    .io_lsbOuts_1(ces_0_3_io_lsbOuts_1),
    .io_lsbOuts_2(ces_0_3_io_lsbOuts_2),
    .io_lsbOuts_3(ces_0_3_io_lsbOuts_3),
    .io_lsbOuts_4(ces_0_3_io_lsbOuts_4),
    .io_lsbOuts_5(ces_0_3_io_lsbOuts_5),
    .io_lsbOuts_6(ces_0_3_io_lsbOuts_6),
    .io_lsbOuts_7(ces_0_3_io_lsbOuts_7)
  );
  Element ces_0_4 (
    .clock(ces_0_4_clock),
    .io_clockOutRight(ces_0_4_io_clockOutRight),
    .io_ins_down(ces_0_4_io_ins_down),
    .io_ins_right(ces_0_4_io_ins_right),
    .io_ins_up(ces_0_4_io_ins_up),
    .io_ins_left(ces_0_4_io_ins_left),
    .io_outs_down(ces_0_4_io_outs_down),
    .io_outs_right(ces_0_4_io_outs_right),
    .io_outs_up(ces_0_4_io_outs_up),
    .io_outs_left(ces_0_4_io_outs_left),
    .io_lsbIns_1(ces_0_4_io_lsbIns_1),
    .io_lsbIns_2(ces_0_4_io_lsbIns_2),
    .io_lsbIns_3(ces_0_4_io_lsbIns_3),
    .io_lsbIns_4(ces_0_4_io_lsbIns_4),
    .io_lsbIns_5(ces_0_4_io_lsbIns_5),
    .io_lsbIns_6(ces_0_4_io_lsbIns_6),
    .io_lsbIns_7(ces_0_4_io_lsbIns_7),
    .io_lsbOuts_0(ces_0_4_io_lsbOuts_0),
    .io_lsbOuts_1(ces_0_4_io_lsbOuts_1),
    .io_lsbOuts_2(ces_0_4_io_lsbOuts_2),
    .io_lsbOuts_3(ces_0_4_io_lsbOuts_3),
    .io_lsbOuts_4(ces_0_4_io_lsbOuts_4),
    .io_lsbOuts_5(ces_0_4_io_lsbOuts_5),
    .io_lsbOuts_6(ces_0_4_io_lsbOuts_6),
    .io_lsbOuts_7(ces_0_4_io_lsbOuts_7)
  );
  Element ces_0_5 (
    .clock(ces_0_5_clock),
    .io_clockOutRight(ces_0_5_io_clockOutRight),
    .io_ins_down(ces_0_5_io_ins_down),
    .io_ins_right(ces_0_5_io_ins_right),
    .io_ins_up(ces_0_5_io_ins_up),
    .io_ins_left(ces_0_5_io_ins_left),
    .io_outs_down(ces_0_5_io_outs_down),
    .io_outs_right(ces_0_5_io_outs_right),
    .io_outs_up(ces_0_5_io_outs_up),
    .io_outs_left(ces_0_5_io_outs_left),
    .io_lsbIns_1(ces_0_5_io_lsbIns_1),
    .io_lsbIns_2(ces_0_5_io_lsbIns_2),
    .io_lsbIns_3(ces_0_5_io_lsbIns_3),
    .io_lsbIns_4(ces_0_5_io_lsbIns_4),
    .io_lsbIns_5(ces_0_5_io_lsbIns_5),
    .io_lsbIns_6(ces_0_5_io_lsbIns_6),
    .io_lsbIns_7(ces_0_5_io_lsbIns_7),
    .io_lsbOuts_0(ces_0_5_io_lsbOuts_0),
    .io_lsbOuts_1(ces_0_5_io_lsbOuts_1),
    .io_lsbOuts_2(ces_0_5_io_lsbOuts_2),
    .io_lsbOuts_3(ces_0_5_io_lsbOuts_3),
    .io_lsbOuts_4(ces_0_5_io_lsbOuts_4),
    .io_lsbOuts_5(ces_0_5_io_lsbOuts_5),
    .io_lsbOuts_6(ces_0_5_io_lsbOuts_6),
    .io_lsbOuts_7(ces_0_5_io_lsbOuts_7)
  );
  Element ces_0_6 (
    .clock(ces_0_6_clock),
    .io_clockOutRight(ces_0_6_io_clockOutRight),
    .io_ins_down(ces_0_6_io_ins_down),
    .io_ins_right(ces_0_6_io_ins_right),
    .io_ins_up(ces_0_6_io_ins_up),
    .io_ins_left(ces_0_6_io_ins_left),
    .io_outs_down(ces_0_6_io_outs_down),
    .io_outs_right(ces_0_6_io_outs_right),
    .io_outs_up(ces_0_6_io_outs_up),
    .io_outs_left(ces_0_6_io_outs_left),
    .io_lsbIns_1(ces_0_6_io_lsbIns_1),
    .io_lsbIns_2(ces_0_6_io_lsbIns_2),
    .io_lsbIns_3(ces_0_6_io_lsbIns_3),
    .io_lsbIns_4(ces_0_6_io_lsbIns_4),
    .io_lsbIns_5(ces_0_6_io_lsbIns_5),
    .io_lsbIns_6(ces_0_6_io_lsbIns_6),
    .io_lsbIns_7(ces_0_6_io_lsbIns_7),
    .io_lsbOuts_0(ces_0_6_io_lsbOuts_0),
    .io_lsbOuts_1(ces_0_6_io_lsbOuts_1),
    .io_lsbOuts_2(ces_0_6_io_lsbOuts_2),
    .io_lsbOuts_3(ces_0_6_io_lsbOuts_3),
    .io_lsbOuts_4(ces_0_6_io_lsbOuts_4),
    .io_lsbOuts_5(ces_0_6_io_lsbOuts_5),
    .io_lsbOuts_6(ces_0_6_io_lsbOuts_6),
    .io_lsbOuts_7(ces_0_6_io_lsbOuts_7)
  );
  Element ces_0_7 (
    .clock(ces_0_7_clock),
    .io_clockOutRight(ces_0_7_io_clockOutRight),
    .io_ins_down(ces_0_7_io_ins_down),
    .io_ins_right(ces_0_7_io_ins_right),
    .io_ins_up(ces_0_7_io_ins_up),
    .io_ins_left(ces_0_7_io_ins_left),
    .io_outs_down(ces_0_7_io_outs_down),
    .io_outs_right(ces_0_7_io_outs_right),
    .io_outs_up(ces_0_7_io_outs_up),
    .io_outs_left(ces_0_7_io_outs_left),
    .io_lsbIns_1(ces_0_7_io_lsbIns_1),
    .io_lsbIns_2(ces_0_7_io_lsbIns_2),
    .io_lsbIns_3(ces_0_7_io_lsbIns_3),
    .io_lsbIns_4(ces_0_7_io_lsbIns_4),
    .io_lsbIns_5(ces_0_7_io_lsbIns_5),
    .io_lsbIns_6(ces_0_7_io_lsbIns_6),
    .io_lsbIns_7(ces_0_7_io_lsbIns_7),
    .io_lsbOuts_0(ces_0_7_io_lsbOuts_0),
    .io_lsbOuts_1(ces_0_7_io_lsbOuts_1),
    .io_lsbOuts_2(ces_0_7_io_lsbOuts_2),
    .io_lsbOuts_3(ces_0_7_io_lsbOuts_3),
    .io_lsbOuts_4(ces_0_7_io_lsbOuts_4),
    .io_lsbOuts_5(ces_0_7_io_lsbOuts_5),
    .io_lsbOuts_6(ces_0_7_io_lsbOuts_6),
    .io_lsbOuts_7(ces_0_7_io_lsbOuts_7)
  );
  Element ces_1_0 (
    .clock(ces_1_0_clock),
    .io_clockOutRight(ces_1_0_io_clockOutRight),
    .io_ins_down(ces_1_0_io_ins_down),
    .io_ins_right(ces_1_0_io_ins_right),
    .io_ins_up(ces_1_0_io_ins_up),
    .io_ins_left(ces_1_0_io_ins_left),
    .io_outs_down(ces_1_0_io_outs_down),
    .io_outs_right(ces_1_0_io_outs_right),
    .io_outs_up(ces_1_0_io_outs_up),
    .io_outs_left(ces_1_0_io_outs_left),
    .io_lsbIns_1(ces_1_0_io_lsbIns_1),
    .io_lsbIns_2(ces_1_0_io_lsbIns_2),
    .io_lsbIns_3(ces_1_0_io_lsbIns_3),
    .io_lsbIns_4(ces_1_0_io_lsbIns_4),
    .io_lsbIns_5(ces_1_0_io_lsbIns_5),
    .io_lsbIns_6(ces_1_0_io_lsbIns_6),
    .io_lsbIns_7(ces_1_0_io_lsbIns_7),
    .io_lsbOuts_0(ces_1_0_io_lsbOuts_0),
    .io_lsbOuts_1(ces_1_0_io_lsbOuts_1),
    .io_lsbOuts_2(ces_1_0_io_lsbOuts_2),
    .io_lsbOuts_3(ces_1_0_io_lsbOuts_3),
    .io_lsbOuts_4(ces_1_0_io_lsbOuts_4),
    .io_lsbOuts_5(ces_1_0_io_lsbOuts_5),
    .io_lsbOuts_6(ces_1_0_io_lsbOuts_6),
    .io_lsbOuts_7(ces_1_0_io_lsbOuts_7)
  );
  Element ces_1_1 (
    .clock(ces_1_1_clock),
    .io_clockOutRight(ces_1_1_io_clockOutRight),
    .io_ins_down(ces_1_1_io_ins_down),
    .io_ins_right(ces_1_1_io_ins_right),
    .io_ins_up(ces_1_1_io_ins_up),
    .io_ins_left(ces_1_1_io_ins_left),
    .io_outs_down(ces_1_1_io_outs_down),
    .io_outs_right(ces_1_1_io_outs_right),
    .io_outs_up(ces_1_1_io_outs_up),
    .io_outs_left(ces_1_1_io_outs_left),
    .io_lsbIns_1(ces_1_1_io_lsbIns_1),
    .io_lsbIns_2(ces_1_1_io_lsbIns_2),
    .io_lsbIns_3(ces_1_1_io_lsbIns_3),
    .io_lsbIns_4(ces_1_1_io_lsbIns_4),
    .io_lsbIns_5(ces_1_1_io_lsbIns_5),
    .io_lsbIns_6(ces_1_1_io_lsbIns_6),
    .io_lsbIns_7(ces_1_1_io_lsbIns_7),
    .io_lsbOuts_0(ces_1_1_io_lsbOuts_0),
    .io_lsbOuts_1(ces_1_1_io_lsbOuts_1),
    .io_lsbOuts_2(ces_1_1_io_lsbOuts_2),
    .io_lsbOuts_3(ces_1_1_io_lsbOuts_3),
    .io_lsbOuts_4(ces_1_1_io_lsbOuts_4),
    .io_lsbOuts_5(ces_1_1_io_lsbOuts_5),
    .io_lsbOuts_6(ces_1_1_io_lsbOuts_6),
    .io_lsbOuts_7(ces_1_1_io_lsbOuts_7)
  );
  Element ces_1_2 (
    .clock(ces_1_2_clock),
    .io_clockOutRight(ces_1_2_io_clockOutRight),
    .io_ins_down(ces_1_2_io_ins_down),
    .io_ins_right(ces_1_2_io_ins_right),
    .io_ins_up(ces_1_2_io_ins_up),
    .io_ins_left(ces_1_2_io_ins_left),
    .io_outs_down(ces_1_2_io_outs_down),
    .io_outs_right(ces_1_2_io_outs_right),
    .io_outs_up(ces_1_2_io_outs_up),
    .io_outs_left(ces_1_2_io_outs_left),
    .io_lsbIns_1(ces_1_2_io_lsbIns_1),
    .io_lsbIns_2(ces_1_2_io_lsbIns_2),
    .io_lsbIns_3(ces_1_2_io_lsbIns_3),
    .io_lsbIns_4(ces_1_2_io_lsbIns_4),
    .io_lsbIns_5(ces_1_2_io_lsbIns_5),
    .io_lsbIns_6(ces_1_2_io_lsbIns_6),
    .io_lsbIns_7(ces_1_2_io_lsbIns_7),
    .io_lsbOuts_0(ces_1_2_io_lsbOuts_0),
    .io_lsbOuts_1(ces_1_2_io_lsbOuts_1),
    .io_lsbOuts_2(ces_1_2_io_lsbOuts_2),
    .io_lsbOuts_3(ces_1_2_io_lsbOuts_3),
    .io_lsbOuts_4(ces_1_2_io_lsbOuts_4),
    .io_lsbOuts_5(ces_1_2_io_lsbOuts_5),
    .io_lsbOuts_6(ces_1_2_io_lsbOuts_6),
    .io_lsbOuts_7(ces_1_2_io_lsbOuts_7)
  );
  Element ces_1_3 (
    .clock(ces_1_3_clock),
    .io_clockOutRight(ces_1_3_io_clockOutRight),
    .io_ins_down(ces_1_3_io_ins_down),
    .io_ins_right(ces_1_3_io_ins_right),
    .io_ins_up(ces_1_3_io_ins_up),
    .io_ins_left(ces_1_3_io_ins_left),
    .io_outs_down(ces_1_3_io_outs_down),
    .io_outs_right(ces_1_3_io_outs_right),
    .io_outs_up(ces_1_3_io_outs_up),
    .io_outs_left(ces_1_3_io_outs_left),
    .io_lsbIns_1(ces_1_3_io_lsbIns_1),
    .io_lsbIns_2(ces_1_3_io_lsbIns_2),
    .io_lsbIns_3(ces_1_3_io_lsbIns_3),
    .io_lsbIns_4(ces_1_3_io_lsbIns_4),
    .io_lsbIns_5(ces_1_3_io_lsbIns_5),
    .io_lsbIns_6(ces_1_3_io_lsbIns_6),
    .io_lsbIns_7(ces_1_3_io_lsbIns_7),
    .io_lsbOuts_0(ces_1_3_io_lsbOuts_0),
    .io_lsbOuts_1(ces_1_3_io_lsbOuts_1),
    .io_lsbOuts_2(ces_1_3_io_lsbOuts_2),
    .io_lsbOuts_3(ces_1_3_io_lsbOuts_3),
    .io_lsbOuts_4(ces_1_3_io_lsbOuts_4),
    .io_lsbOuts_5(ces_1_3_io_lsbOuts_5),
    .io_lsbOuts_6(ces_1_3_io_lsbOuts_6),
    .io_lsbOuts_7(ces_1_3_io_lsbOuts_7)
  );
  Element ces_1_4 (
    .clock(ces_1_4_clock),
    .io_clockOutRight(ces_1_4_io_clockOutRight),
    .io_ins_down(ces_1_4_io_ins_down),
    .io_ins_right(ces_1_4_io_ins_right),
    .io_ins_up(ces_1_4_io_ins_up),
    .io_ins_left(ces_1_4_io_ins_left),
    .io_outs_down(ces_1_4_io_outs_down),
    .io_outs_right(ces_1_4_io_outs_right),
    .io_outs_up(ces_1_4_io_outs_up),
    .io_outs_left(ces_1_4_io_outs_left),
    .io_lsbIns_1(ces_1_4_io_lsbIns_1),
    .io_lsbIns_2(ces_1_4_io_lsbIns_2),
    .io_lsbIns_3(ces_1_4_io_lsbIns_3),
    .io_lsbIns_4(ces_1_4_io_lsbIns_4),
    .io_lsbIns_5(ces_1_4_io_lsbIns_5),
    .io_lsbIns_6(ces_1_4_io_lsbIns_6),
    .io_lsbIns_7(ces_1_4_io_lsbIns_7),
    .io_lsbOuts_0(ces_1_4_io_lsbOuts_0),
    .io_lsbOuts_1(ces_1_4_io_lsbOuts_1),
    .io_lsbOuts_2(ces_1_4_io_lsbOuts_2),
    .io_lsbOuts_3(ces_1_4_io_lsbOuts_3),
    .io_lsbOuts_4(ces_1_4_io_lsbOuts_4),
    .io_lsbOuts_5(ces_1_4_io_lsbOuts_5),
    .io_lsbOuts_6(ces_1_4_io_lsbOuts_6),
    .io_lsbOuts_7(ces_1_4_io_lsbOuts_7)
  );
  Element ces_1_5 (
    .clock(ces_1_5_clock),
    .io_clockOutRight(ces_1_5_io_clockOutRight),
    .io_ins_down(ces_1_5_io_ins_down),
    .io_ins_right(ces_1_5_io_ins_right),
    .io_ins_up(ces_1_5_io_ins_up),
    .io_ins_left(ces_1_5_io_ins_left),
    .io_outs_down(ces_1_5_io_outs_down),
    .io_outs_right(ces_1_5_io_outs_right),
    .io_outs_up(ces_1_5_io_outs_up),
    .io_outs_left(ces_1_5_io_outs_left),
    .io_lsbIns_1(ces_1_5_io_lsbIns_1),
    .io_lsbIns_2(ces_1_5_io_lsbIns_2),
    .io_lsbIns_3(ces_1_5_io_lsbIns_3),
    .io_lsbIns_4(ces_1_5_io_lsbIns_4),
    .io_lsbIns_5(ces_1_5_io_lsbIns_5),
    .io_lsbIns_6(ces_1_5_io_lsbIns_6),
    .io_lsbIns_7(ces_1_5_io_lsbIns_7),
    .io_lsbOuts_0(ces_1_5_io_lsbOuts_0),
    .io_lsbOuts_1(ces_1_5_io_lsbOuts_1),
    .io_lsbOuts_2(ces_1_5_io_lsbOuts_2),
    .io_lsbOuts_3(ces_1_5_io_lsbOuts_3),
    .io_lsbOuts_4(ces_1_5_io_lsbOuts_4),
    .io_lsbOuts_5(ces_1_5_io_lsbOuts_5),
    .io_lsbOuts_6(ces_1_5_io_lsbOuts_6),
    .io_lsbOuts_7(ces_1_5_io_lsbOuts_7)
  );
  Element ces_1_6 (
    .clock(ces_1_6_clock),
    .io_clockOutRight(ces_1_6_io_clockOutRight),
    .io_ins_down(ces_1_6_io_ins_down),
    .io_ins_right(ces_1_6_io_ins_right),
    .io_ins_up(ces_1_6_io_ins_up),
    .io_ins_left(ces_1_6_io_ins_left),
    .io_outs_down(ces_1_6_io_outs_down),
    .io_outs_right(ces_1_6_io_outs_right),
    .io_outs_up(ces_1_6_io_outs_up),
    .io_outs_left(ces_1_6_io_outs_left),
    .io_lsbIns_1(ces_1_6_io_lsbIns_1),
    .io_lsbIns_2(ces_1_6_io_lsbIns_2),
    .io_lsbIns_3(ces_1_6_io_lsbIns_3),
    .io_lsbIns_4(ces_1_6_io_lsbIns_4),
    .io_lsbIns_5(ces_1_6_io_lsbIns_5),
    .io_lsbIns_6(ces_1_6_io_lsbIns_6),
    .io_lsbIns_7(ces_1_6_io_lsbIns_7),
    .io_lsbOuts_0(ces_1_6_io_lsbOuts_0),
    .io_lsbOuts_1(ces_1_6_io_lsbOuts_1),
    .io_lsbOuts_2(ces_1_6_io_lsbOuts_2),
    .io_lsbOuts_3(ces_1_6_io_lsbOuts_3),
    .io_lsbOuts_4(ces_1_6_io_lsbOuts_4),
    .io_lsbOuts_5(ces_1_6_io_lsbOuts_5),
    .io_lsbOuts_6(ces_1_6_io_lsbOuts_6),
    .io_lsbOuts_7(ces_1_6_io_lsbOuts_7)
  );
  Element ces_1_7 (
    .clock(ces_1_7_clock),
    .io_clockOutRight(ces_1_7_io_clockOutRight),
    .io_ins_down(ces_1_7_io_ins_down),
    .io_ins_right(ces_1_7_io_ins_right),
    .io_ins_up(ces_1_7_io_ins_up),
    .io_ins_left(ces_1_7_io_ins_left),
    .io_outs_down(ces_1_7_io_outs_down),
    .io_outs_right(ces_1_7_io_outs_right),
    .io_outs_up(ces_1_7_io_outs_up),
    .io_outs_left(ces_1_7_io_outs_left),
    .io_lsbIns_1(ces_1_7_io_lsbIns_1),
    .io_lsbIns_2(ces_1_7_io_lsbIns_2),
    .io_lsbIns_3(ces_1_7_io_lsbIns_3),
    .io_lsbIns_4(ces_1_7_io_lsbIns_4),
    .io_lsbIns_5(ces_1_7_io_lsbIns_5),
    .io_lsbIns_6(ces_1_7_io_lsbIns_6),
    .io_lsbIns_7(ces_1_7_io_lsbIns_7),
    .io_lsbOuts_0(ces_1_7_io_lsbOuts_0),
    .io_lsbOuts_1(ces_1_7_io_lsbOuts_1),
    .io_lsbOuts_2(ces_1_7_io_lsbOuts_2),
    .io_lsbOuts_3(ces_1_7_io_lsbOuts_3),
    .io_lsbOuts_4(ces_1_7_io_lsbOuts_4),
    .io_lsbOuts_5(ces_1_7_io_lsbOuts_5),
    .io_lsbOuts_6(ces_1_7_io_lsbOuts_6),
    .io_lsbOuts_7(ces_1_7_io_lsbOuts_7)
  );
  Element ces_2_0 (
    .clock(ces_2_0_clock),
    .io_clockOutRight(ces_2_0_io_clockOutRight),
    .io_ins_down(ces_2_0_io_ins_down),
    .io_ins_right(ces_2_0_io_ins_right),
    .io_ins_up(ces_2_0_io_ins_up),
    .io_ins_left(ces_2_0_io_ins_left),
    .io_outs_down(ces_2_0_io_outs_down),
    .io_outs_right(ces_2_0_io_outs_right),
    .io_outs_up(ces_2_0_io_outs_up),
    .io_outs_left(ces_2_0_io_outs_left),
    .io_lsbIns_1(ces_2_0_io_lsbIns_1),
    .io_lsbIns_2(ces_2_0_io_lsbIns_2),
    .io_lsbIns_3(ces_2_0_io_lsbIns_3),
    .io_lsbIns_4(ces_2_0_io_lsbIns_4),
    .io_lsbIns_5(ces_2_0_io_lsbIns_5),
    .io_lsbIns_6(ces_2_0_io_lsbIns_6),
    .io_lsbIns_7(ces_2_0_io_lsbIns_7),
    .io_lsbOuts_0(ces_2_0_io_lsbOuts_0),
    .io_lsbOuts_1(ces_2_0_io_lsbOuts_1),
    .io_lsbOuts_2(ces_2_0_io_lsbOuts_2),
    .io_lsbOuts_3(ces_2_0_io_lsbOuts_3),
    .io_lsbOuts_4(ces_2_0_io_lsbOuts_4),
    .io_lsbOuts_5(ces_2_0_io_lsbOuts_5),
    .io_lsbOuts_6(ces_2_0_io_lsbOuts_6),
    .io_lsbOuts_7(ces_2_0_io_lsbOuts_7)
  );
  Element ces_2_1 (
    .clock(ces_2_1_clock),
    .io_clockOutRight(ces_2_1_io_clockOutRight),
    .io_ins_down(ces_2_1_io_ins_down),
    .io_ins_right(ces_2_1_io_ins_right),
    .io_ins_up(ces_2_1_io_ins_up),
    .io_ins_left(ces_2_1_io_ins_left),
    .io_outs_down(ces_2_1_io_outs_down),
    .io_outs_right(ces_2_1_io_outs_right),
    .io_outs_up(ces_2_1_io_outs_up),
    .io_outs_left(ces_2_1_io_outs_left),
    .io_lsbIns_1(ces_2_1_io_lsbIns_1),
    .io_lsbIns_2(ces_2_1_io_lsbIns_2),
    .io_lsbIns_3(ces_2_1_io_lsbIns_3),
    .io_lsbIns_4(ces_2_1_io_lsbIns_4),
    .io_lsbIns_5(ces_2_1_io_lsbIns_5),
    .io_lsbIns_6(ces_2_1_io_lsbIns_6),
    .io_lsbIns_7(ces_2_1_io_lsbIns_7),
    .io_lsbOuts_0(ces_2_1_io_lsbOuts_0),
    .io_lsbOuts_1(ces_2_1_io_lsbOuts_1),
    .io_lsbOuts_2(ces_2_1_io_lsbOuts_2),
    .io_lsbOuts_3(ces_2_1_io_lsbOuts_3),
    .io_lsbOuts_4(ces_2_1_io_lsbOuts_4),
    .io_lsbOuts_5(ces_2_1_io_lsbOuts_5),
    .io_lsbOuts_6(ces_2_1_io_lsbOuts_6),
    .io_lsbOuts_7(ces_2_1_io_lsbOuts_7)
  );
  Element ces_2_2 (
    .clock(ces_2_2_clock),
    .io_clockOutRight(ces_2_2_io_clockOutRight),
    .io_ins_down(ces_2_2_io_ins_down),
    .io_ins_right(ces_2_2_io_ins_right),
    .io_ins_up(ces_2_2_io_ins_up),
    .io_ins_left(ces_2_2_io_ins_left),
    .io_outs_down(ces_2_2_io_outs_down),
    .io_outs_right(ces_2_2_io_outs_right),
    .io_outs_up(ces_2_2_io_outs_up),
    .io_outs_left(ces_2_2_io_outs_left),
    .io_lsbIns_1(ces_2_2_io_lsbIns_1),
    .io_lsbIns_2(ces_2_2_io_lsbIns_2),
    .io_lsbIns_3(ces_2_2_io_lsbIns_3),
    .io_lsbIns_4(ces_2_2_io_lsbIns_4),
    .io_lsbIns_5(ces_2_2_io_lsbIns_5),
    .io_lsbIns_6(ces_2_2_io_lsbIns_6),
    .io_lsbIns_7(ces_2_2_io_lsbIns_7),
    .io_lsbOuts_0(ces_2_2_io_lsbOuts_0),
    .io_lsbOuts_1(ces_2_2_io_lsbOuts_1),
    .io_lsbOuts_2(ces_2_2_io_lsbOuts_2),
    .io_lsbOuts_3(ces_2_2_io_lsbOuts_3),
    .io_lsbOuts_4(ces_2_2_io_lsbOuts_4),
    .io_lsbOuts_5(ces_2_2_io_lsbOuts_5),
    .io_lsbOuts_6(ces_2_2_io_lsbOuts_6),
    .io_lsbOuts_7(ces_2_2_io_lsbOuts_7)
  );
  Element ces_2_3 (
    .clock(ces_2_3_clock),
    .io_clockOutRight(ces_2_3_io_clockOutRight),
    .io_ins_down(ces_2_3_io_ins_down),
    .io_ins_right(ces_2_3_io_ins_right),
    .io_ins_up(ces_2_3_io_ins_up),
    .io_ins_left(ces_2_3_io_ins_left),
    .io_outs_down(ces_2_3_io_outs_down),
    .io_outs_right(ces_2_3_io_outs_right),
    .io_outs_up(ces_2_3_io_outs_up),
    .io_outs_left(ces_2_3_io_outs_left),
    .io_lsbIns_1(ces_2_3_io_lsbIns_1),
    .io_lsbIns_2(ces_2_3_io_lsbIns_2),
    .io_lsbIns_3(ces_2_3_io_lsbIns_3),
    .io_lsbIns_4(ces_2_3_io_lsbIns_4),
    .io_lsbIns_5(ces_2_3_io_lsbIns_5),
    .io_lsbIns_6(ces_2_3_io_lsbIns_6),
    .io_lsbIns_7(ces_2_3_io_lsbIns_7),
    .io_lsbOuts_0(ces_2_3_io_lsbOuts_0),
    .io_lsbOuts_1(ces_2_3_io_lsbOuts_1),
    .io_lsbOuts_2(ces_2_3_io_lsbOuts_2),
    .io_lsbOuts_3(ces_2_3_io_lsbOuts_3),
    .io_lsbOuts_4(ces_2_3_io_lsbOuts_4),
    .io_lsbOuts_5(ces_2_3_io_lsbOuts_5),
    .io_lsbOuts_6(ces_2_3_io_lsbOuts_6),
    .io_lsbOuts_7(ces_2_3_io_lsbOuts_7)
  );
  Element ces_2_4 (
    .clock(ces_2_4_clock),
    .io_clockOutRight(ces_2_4_io_clockOutRight),
    .io_ins_down(ces_2_4_io_ins_down),
    .io_ins_right(ces_2_4_io_ins_right),
    .io_ins_up(ces_2_4_io_ins_up),
    .io_ins_left(ces_2_4_io_ins_left),
    .io_outs_down(ces_2_4_io_outs_down),
    .io_outs_right(ces_2_4_io_outs_right),
    .io_outs_up(ces_2_4_io_outs_up),
    .io_outs_left(ces_2_4_io_outs_left),
    .io_lsbIns_1(ces_2_4_io_lsbIns_1),
    .io_lsbIns_2(ces_2_4_io_lsbIns_2),
    .io_lsbIns_3(ces_2_4_io_lsbIns_3),
    .io_lsbIns_4(ces_2_4_io_lsbIns_4),
    .io_lsbIns_5(ces_2_4_io_lsbIns_5),
    .io_lsbIns_6(ces_2_4_io_lsbIns_6),
    .io_lsbIns_7(ces_2_4_io_lsbIns_7),
    .io_lsbOuts_0(ces_2_4_io_lsbOuts_0),
    .io_lsbOuts_1(ces_2_4_io_lsbOuts_1),
    .io_lsbOuts_2(ces_2_4_io_lsbOuts_2),
    .io_lsbOuts_3(ces_2_4_io_lsbOuts_3),
    .io_lsbOuts_4(ces_2_4_io_lsbOuts_4),
    .io_lsbOuts_5(ces_2_4_io_lsbOuts_5),
    .io_lsbOuts_6(ces_2_4_io_lsbOuts_6),
    .io_lsbOuts_7(ces_2_4_io_lsbOuts_7)
  );
  Element ces_2_5 (
    .clock(ces_2_5_clock),
    .io_clockOutRight(ces_2_5_io_clockOutRight),
    .io_ins_down(ces_2_5_io_ins_down),
    .io_ins_right(ces_2_5_io_ins_right),
    .io_ins_up(ces_2_5_io_ins_up),
    .io_ins_left(ces_2_5_io_ins_left),
    .io_outs_down(ces_2_5_io_outs_down),
    .io_outs_right(ces_2_5_io_outs_right),
    .io_outs_up(ces_2_5_io_outs_up),
    .io_outs_left(ces_2_5_io_outs_left),
    .io_lsbIns_1(ces_2_5_io_lsbIns_1),
    .io_lsbIns_2(ces_2_5_io_lsbIns_2),
    .io_lsbIns_3(ces_2_5_io_lsbIns_3),
    .io_lsbIns_4(ces_2_5_io_lsbIns_4),
    .io_lsbIns_5(ces_2_5_io_lsbIns_5),
    .io_lsbIns_6(ces_2_5_io_lsbIns_6),
    .io_lsbIns_7(ces_2_5_io_lsbIns_7),
    .io_lsbOuts_0(ces_2_5_io_lsbOuts_0),
    .io_lsbOuts_1(ces_2_5_io_lsbOuts_1),
    .io_lsbOuts_2(ces_2_5_io_lsbOuts_2),
    .io_lsbOuts_3(ces_2_5_io_lsbOuts_3),
    .io_lsbOuts_4(ces_2_5_io_lsbOuts_4),
    .io_lsbOuts_5(ces_2_5_io_lsbOuts_5),
    .io_lsbOuts_6(ces_2_5_io_lsbOuts_6),
    .io_lsbOuts_7(ces_2_5_io_lsbOuts_7)
  );
  Element ces_2_6 (
    .clock(ces_2_6_clock),
    .io_clockOutRight(ces_2_6_io_clockOutRight),
    .io_ins_down(ces_2_6_io_ins_down),
    .io_ins_right(ces_2_6_io_ins_right),
    .io_ins_up(ces_2_6_io_ins_up),
    .io_ins_left(ces_2_6_io_ins_left),
    .io_outs_down(ces_2_6_io_outs_down),
    .io_outs_right(ces_2_6_io_outs_right),
    .io_outs_up(ces_2_6_io_outs_up),
    .io_outs_left(ces_2_6_io_outs_left),
    .io_lsbIns_1(ces_2_6_io_lsbIns_1),
    .io_lsbIns_2(ces_2_6_io_lsbIns_2),
    .io_lsbIns_3(ces_2_6_io_lsbIns_3),
    .io_lsbIns_4(ces_2_6_io_lsbIns_4),
    .io_lsbIns_5(ces_2_6_io_lsbIns_5),
    .io_lsbIns_6(ces_2_6_io_lsbIns_6),
    .io_lsbIns_7(ces_2_6_io_lsbIns_7),
    .io_lsbOuts_0(ces_2_6_io_lsbOuts_0),
    .io_lsbOuts_1(ces_2_6_io_lsbOuts_1),
    .io_lsbOuts_2(ces_2_6_io_lsbOuts_2),
    .io_lsbOuts_3(ces_2_6_io_lsbOuts_3),
    .io_lsbOuts_4(ces_2_6_io_lsbOuts_4),
    .io_lsbOuts_5(ces_2_6_io_lsbOuts_5),
    .io_lsbOuts_6(ces_2_6_io_lsbOuts_6),
    .io_lsbOuts_7(ces_2_6_io_lsbOuts_7)
  );
  Element ces_2_7 (
    .clock(ces_2_7_clock),
    .io_clockOutRight(ces_2_7_io_clockOutRight),
    .io_ins_down(ces_2_7_io_ins_down),
    .io_ins_right(ces_2_7_io_ins_right),
    .io_ins_up(ces_2_7_io_ins_up),
    .io_ins_left(ces_2_7_io_ins_left),
    .io_outs_down(ces_2_7_io_outs_down),
    .io_outs_right(ces_2_7_io_outs_right),
    .io_outs_up(ces_2_7_io_outs_up),
    .io_outs_left(ces_2_7_io_outs_left),
    .io_lsbIns_1(ces_2_7_io_lsbIns_1),
    .io_lsbIns_2(ces_2_7_io_lsbIns_2),
    .io_lsbIns_3(ces_2_7_io_lsbIns_3),
    .io_lsbIns_4(ces_2_7_io_lsbIns_4),
    .io_lsbIns_5(ces_2_7_io_lsbIns_5),
    .io_lsbIns_6(ces_2_7_io_lsbIns_6),
    .io_lsbIns_7(ces_2_7_io_lsbIns_7),
    .io_lsbOuts_0(ces_2_7_io_lsbOuts_0),
    .io_lsbOuts_1(ces_2_7_io_lsbOuts_1),
    .io_lsbOuts_2(ces_2_7_io_lsbOuts_2),
    .io_lsbOuts_3(ces_2_7_io_lsbOuts_3),
    .io_lsbOuts_4(ces_2_7_io_lsbOuts_4),
    .io_lsbOuts_5(ces_2_7_io_lsbOuts_5),
    .io_lsbOuts_6(ces_2_7_io_lsbOuts_6),
    .io_lsbOuts_7(ces_2_7_io_lsbOuts_7)
  );
  Element ces_3_0 (
    .clock(ces_3_0_clock),
    .io_clockOutRight(ces_3_0_io_clockOutRight),
    .io_ins_down(ces_3_0_io_ins_down),
    .io_ins_right(ces_3_0_io_ins_right),
    .io_ins_up(ces_3_0_io_ins_up),
    .io_ins_left(ces_3_0_io_ins_left),
    .io_outs_down(ces_3_0_io_outs_down),
    .io_outs_right(ces_3_0_io_outs_right),
    .io_outs_up(ces_3_0_io_outs_up),
    .io_outs_left(ces_3_0_io_outs_left),
    .io_lsbIns_1(ces_3_0_io_lsbIns_1),
    .io_lsbIns_2(ces_3_0_io_lsbIns_2),
    .io_lsbIns_3(ces_3_0_io_lsbIns_3),
    .io_lsbIns_4(ces_3_0_io_lsbIns_4),
    .io_lsbIns_5(ces_3_0_io_lsbIns_5),
    .io_lsbIns_6(ces_3_0_io_lsbIns_6),
    .io_lsbIns_7(ces_3_0_io_lsbIns_7),
    .io_lsbOuts_0(ces_3_0_io_lsbOuts_0),
    .io_lsbOuts_1(ces_3_0_io_lsbOuts_1),
    .io_lsbOuts_2(ces_3_0_io_lsbOuts_2),
    .io_lsbOuts_3(ces_3_0_io_lsbOuts_3),
    .io_lsbOuts_4(ces_3_0_io_lsbOuts_4),
    .io_lsbOuts_5(ces_3_0_io_lsbOuts_5),
    .io_lsbOuts_6(ces_3_0_io_lsbOuts_6),
    .io_lsbOuts_7(ces_3_0_io_lsbOuts_7)
  );
  Element ces_3_1 (
    .clock(ces_3_1_clock),
    .io_clockOutRight(ces_3_1_io_clockOutRight),
    .io_ins_down(ces_3_1_io_ins_down),
    .io_ins_right(ces_3_1_io_ins_right),
    .io_ins_up(ces_3_1_io_ins_up),
    .io_ins_left(ces_3_1_io_ins_left),
    .io_outs_down(ces_3_1_io_outs_down),
    .io_outs_right(ces_3_1_io_outs_right),
    .io_outs_up(ces_3_1_io_outs_up),
    .io_outs_left(ces_3_1_io_outs_left),
    .io_lsbIns_1(ces_3_1_io_lsbIns_1),
    .io_lsbIns_2(ces_3_1_io_lsbIns_2),
    .io_lsbIns_3(ces_3_1_io_lsbIns_3),
    .io_lsbIns_4(ces_3_1_io_lsbIns_4),
    .io_lsbIns_5(ces_3_1_io_lsbIns_5),
    .io_lsbIns_6(ces_3_1_io_lsbIns_6),
    .io_lsbIns_7(ces_3_1_io_lsbIns_7),
    .io_lsbOuts_0(ces_3_1_io_lsbOuts_0),
    .io_lsbOuts_1(ces_3_1_io_lsbOuts_1),
    .io_lsbOuts_2(ces_3_1_io_lsbOuts_2),
    .io_lsbOuts_3(ces_3_1_io_lsbOuts_3),
    .io_lsbOuts_4(ces_3_1_io_lsbOuts_4),
    .io_lsbOuts_5(ces_3_1_io_lsbOuts_5),
    .io_lsbOuts_6(ces_3_1_io_lsbOuts_6),
    .io_lsbOuts_7(ces_3_1_io_lsbOuts_7)
  );
  Element ces_3_2 (
    .clock(ces_3_2_clock),
    .io_clockOutRight(ces_3_2_io_clockOutRight),
    .io_ins_down(ces_3_2_io_ins_down),
    .io_ins_right(ces_3_2_io_ins_right),
    .io_ins_up(ces_3_2_io_ins_up),
    .io_ins_left(ces_3_2_io_ins_left),
    .io_outs_down(ces_3_2_io_outs_down),
    .io_outs_right(ces_3_2_io_outs_right),
    .io_outs_up(ces_3_2_io_outs_up),
    .io_outs_left(ces_3_2_io_outs_left),
    .io_lsbIns_1(ces_3_2_io_lsbIns_1),
    .io_lsbIns_2(ces_3_2_io_lsbIns_2),
    .io_lsbIns_3(ces_3_2_io_lsbIns_3),
    .io_lsbIns_4(ces_3_2_io_lsbIns_4),
    .io_lsbIns_5(ces_3_2_io_lsbIns_5),
    .io_lsbIns_6(ces_3_2_io_lsbIns_6),
    .io_lsbIns_7(ces_3_2_io_lsbIns_7),
    .io_lsbOuts_0(ces_3_2_io_lsbOuts_0),
    .io_lsbOuts_1(ces_3_2_io_lsbOuts_1),
    .io_lsbOuts_2(ces_3_2_io_lsbOuts_2),
    .io_lsbOuts_3(ces_3_2_io_lsbOuts_3),
    .io_lsbOuts_4(ces_3_2_io_lsbOuts_4),
    .io_lsbOuts_5(ces_3_2_io_lsbOuts_5),
    .io_lsbOuts_6(ces_3_2_io_lsbOuts_6),
    .io_lsbOuts_7(ces_3_2_io_lsbOuts_7)
  );
  Element ces_3_3 (
    .clock(ces_3_3_clock),
    .io_clockOutRight(ces_3_3_io_clockOutRight),
    .io_ins_down(ces_3_3_io_ins_down),
    .io_ins_right(ces_3_3_io_ins_right),
    .io_ins_up(ces_3_3_io_ins_up),
    .io_ins_left(ces_3_3_io_ins_left),
    .io_outs_down(ces_3_3_io_outs_down),
    .io_outs_right(ces_3_3_io_outs_right),
    .io_outs_up(ces_3_3_io_outs_up),
    .io_outs_left(ces_3_3_io_outs_left),
    .io_lsbIns_1(ces_3_3_io_lsbIns_1),
    .io_lsbIns_2(ces_3_3_io_lsbIns_2),
    .io_lsbIns_3(ces_3_3_io_lsbIns_3),
    .io_lsbIns_4(ces_3_3_io_lsbIns_4),
    .io_lsbIns_5(ces_3_3_io_lsbIns_5),
    .io_lsbIns_6(ces_3_3_io_lsbIns_6),
    .io_lsbIns_7(ces_3_3_io_lsbIns_7),
    .io_lsbOuts_0(ces_3_3_io_lsbOuts_0),
    .io_lsbOuts_1(ces_3_3_io_lsbOuts_1),
    .io_lsbOuts_2(ces_3_3_io_lsbOuts_2),
    .io_lsbOuts_3(ces_3_3_io_lsbOuts_3),
    .io_lsbOuts_4(ces_3_3_io_lsbOuts_4),
    .io_lsbOuts_5(ces_3_3_io_lsbOuts_5),
    .io_lsbOuts_6(ces_3_3_io_lsbOuts_6),
    .io_lsbOuts_7(ces_3_3_io_lsbOuts_7)
  );
  Element ces_3_4 (
    .clock(ces_3_4_clock),
    .io_clockOutRight(ces_3_4_io_clockOutRight),
    .io_ins_down(ces_3_4_io_ins_down),
    .io_ins_right(ces_3_4_io_ins_right),
    .io_ins_up(ces_3_4_io_ins_up),
    .io_ins_left(ces_3_4_io_ins_left),
    .io_outs_down(ces_3_4_io_outs_down),
    .io_outs_right(ces_3_4_io_outs_right),
    .io_outs_up(ces_3_4_io_outs_up),
    .io_outs_left(ces_3_4_io_outs_left),
    .io_lsbIns_1(ces_3_4_io_lsbIns_1),
    .io_lsbIns_2(ces_3_4_io_lsbIns_2),
    .io_lsbIns_3(ces_3_4_io_lsbIns_3),
    .io_lsbIns_4(ces_3_4_io_lsbIns_4),
    .io_lsbIns_5(ces_3_4_io_lsbIns_5),
    .io_lsbIns_6(ces_3_4_io_lsbIns_6),
    .io_lsbIns_7(ces_3_4_io_lsbIns_7),
    .io_lsbOuts_0(ces_3_4_io_lsbOuts_0),
    .io_lsbOuts_1(ces_3_4_io_lsbOuts_1),
    .io_lsbOuts_2(ces_3_4_io_lsbOuts_2),
    .io_lsbOuts_3(ces_3_4_io_lsbOuts_3),
    .io_lsbOuts_4(ces_3_4_io_lsbOuts_4),
    .io_lsbOuts_5(ces_3_4_io_lsbOuts_5),
    .io_lsbOuts_6(ces_3_4_io_lsbOuts_6),
    .io_lsbOuts_7(ces_3_4_io_lsbOuts_7)
  );
  Element ces_3_5 (
    .clock(ces_3_5_clock),
    .io_clockOutRight(ces_3_5_io_clockOutRight),
    .io_ins_down(ces_3_5_io_ins_down),
    .io_ins_right(ces_3_5_io_ins_right),
    .io_ins_up(ces_3_5_io_ins_up),
    .io_ins_left(ces_3_5_io_ins_left),
    .io_outs_down(ces_3_5_io_outs_down),
    .io_outs_right(ces_3_5_io_outs_right),
    .io_outs_up(ces_3_5_io_outs_up),
    .io_outs_left(ces_3_5_io_outs_left),
    .io_lsbIns_1(ces_3_5_io_lsbIns_1),
    .io_lsbIns_2(ces_3_5_io_lsbIns_2),
    .io_lsbIns_3(ces_3_5_io_lsbIns_3),
    .io_lsbIns_4(ces_3_5_io_lsbIns_4),
    .io_lsbIns_5(ces_3_5_io_lsbIns_5),
    .io_lsbIns_6(ces_3_5_io_lsbIns_6),
    .io_lsbIns_7(ces_3_5_io_lsbIns_7),
    .io_lsbOuts_0(ces_3_5_io_lsbOuts_0),
    .io_lsbOuts_1(ces_3_5_io_lsbOuts_1),
    .io_lsbOuts_2(ces_3_5_io_lsbOuts_2),
    .io_lsbOuts_3(ces_3_5_io_lsbOuts_3),
    .io_lsbOuts_4(ces_3_5_io_lsbOuts_4),
    .io_lsbOuts_5(ces_3_5_io_lsbOuts_5),
    .io_lsbOuts_6(ces_3_5_io_lsbOuts_6),
    .io_lsbOuts_7(ces_3_5_io_lsbOuts_7)
  );
  Element ces_3_6 (
    .clock(ces_3_6_clock),
    .io_clockOutRight(ces_3_6_io_clockOutRight),
    .io_ins_down(ces_3_6_io_ins_down),
    .io_ins_right(ces_3_6_io_ins_right),
    .io_ins_up(ces_3_6_io_ins_up),
    .io_ins_left(ces_3_6_io_ins_left),
    .io_outs_down(ces_3_6_io_outs_down),
    .io_outs_right(ces_3_6_io_outs_right),
    .io_outs_up(ces_3_6_io_outs_up),
    .io_outs_left(ces_3_6_io_outs_left),
    .io_lsbIns_1(ces_3_6_io_lsbIns_1),
    .io_lsbIns_2(ces_3_6_io_lsbIns_2),
    .io_lsbIns_3(ces_3_6_io_lsbIns_3),
    .io_lsbIns_4(ces_3_6_io_lsbIns_4),
    .io_lsbIns_5(ces_3_6_io_lsbIns_5),
    .io_lsbIns_6(ces_3_6_io_lsbIns_6),
    .io_lsbIns_7(ces_3_6_io_lsbIns_7),
    .io_lsbOuts_0(ces_3_6_io_lsbOuts_0),
    .io_lsbOuts_1(ces_3_6_io_lsbOuts_1),
    .io_lsbOuts_2(ces_3_6_io_lsbOuts_2),
    .io_lsbOuts_3(ces_3_6_io_lsbOuts_3),
    .io_lsbOuts_4(ces_3_6_io_lsbOuts_4),
    .io_lsbOuts_5(ces_3_6_io_lsbOuts_5),
    .io_lsbOuts_6(ces_3_6_io_lsbOuts_6),
    .io_lsbOuts_7(ces_3_6_io_lsbOuts_7)
  );
  Element ces_3_7 (
    .clock(ces_3_7_clock),
    .io_clockOutRight(ces_3_7_io_clockOutRight),
    .io_ins_down(ces_3_7_io_ins_down),
    .io_ins_right(ces_3_7_io_ins_right),
    .io_ins_up(ces_3_7_io_ins_up),
    .io_ins_left(ces_3_7_io_ins_left),
    .io_outs_down(ces_3_7_io_outs_down),
    .io_outs_right(ces_3_7_io_outs_right),
    .io_outs_up(ces_3_7_io_outs_up),
    .io_outs_left(ces_3_7_io_outs_left),
    .io_lsbIns_1(ces_3_7_io_lsbIns_1),
    .io_lsbIns_2(ces_3_7_io_lsbIns_2),
    .io_lsbIns_3(ces_3_7_io_lsbIns_3),
    .io_lsbIns_4(ces_3_7_io_lsbIns_4),
    .io_lsbIns_5(ces_3_7_io_lsbIns_5),
    .io_lsbIns_6(ces_3_7_io_lsbIns_6),
    .io_lsbIns_7(ces_3_7_io_lsbIns_7),
    .io_lsbOuts_0(ces_3_7_io_lsbOuts_0),
    .io_lsbOuts_1(ces_3_7_io_lsbOuts_1),
    .io_lsbOuts_2(ces_3_7_io_lsbOuts_2),
    .io_lsbOuts_3(ces_3_7_io_lsbOuts_3),
    .io_lsbOuts_4(ces_3_7_io_lsbOuts_4),
    .io_lsbOuts_5(ces_3_7_io_lsbOuts_5),
    .io_lsbOuts_6(ces_3_7_io_lsbOuts_6),
    .io_lsbOuts_7(ces_3_7_io_lsbOuts_7)
  );
  Element ces_4_0 (
    .clock(ces_4_0_clock),
    .io_clockOutRight(ces_4_0_io_clockOutRight),
    .io_ins_down(ces_4_0_io_ins_down),
    .io_ins_right(ces_4_0_io_ins_right),
    .io_ins_up(ces_4_0_io_ins_up),
    .io_ins_left(ces_4_0_io_ins_left),
    .io_outs_down(ces_4_0_io_outs_down),
    .io_outs_right(ces_4_0_io_outs_right),
    .io_outs_up(ces_4_0_io_outs_up),
    .io_outs_left(ces_4_0_io_outs_left),
    .io_lsbIns_1(ces_4_0_io_lsbIns_1),
    .io_lsbIns_2(ces_4_0_io_lsbIns_2),
    .io_lsbIns_3(ces_4_0_io_lsbIns_3),
    .io_lsbIns_4(ces_4_0_io_lsbIns_4),
    .io_lsbIns_5(ces_4_0_io_lsbIns_5),
    .io_lsbIns_6(ces_4_0_io_lsbIns_6),
    .io_lsbIns_7(ces_4_0_io_lsbIns_7),
    .io_lsbOuts_0(ces_4_0_io_lsbOuts_0),
    .io_lsbOuts_1(ces_4_0_io_lsbOuts_1),
    .io_lsbOuts_2(ces_4_0_io_lsbOuts_2),
    .io_lsbOuts_3(ces_4_0_io_lsbOuts_3),
    .io_lsbOuts_4(ces_4_0_io_lsbOuts_4),
    .io_lsbOuts_5(ces_4_0_io_lsbOuts_5),
    .io_lsbOuts_6(ces_4_0_io_lsbOuts_6),
    .io_lsbOuts_7(ces_4_0_io_lsbOuts_7)
  );
  Element ces_4_1 (
    .clock(ces_4_1_clock),
    .io_clockOutRight(ces_4_1_io_clockOutRight),
    .io_ins_down(ces_4_1_io_ins_down),
    .io_ins_right(ces_4_1_io_ins_right),
    .io_ins_up(ces_4_1_io_ins_up),
    .io_ins_left(ces_4_1_io_ins_left),
    .io_outs_down(ces_4_1_io_outs_down),
    .io_outs_right(ces_4_1_io_outs_right),
    .io_outs_up(ces_4_1_io_outs_up),
    .io_outs_left(ces_4_1_io_outs_left),
    .io_lsbIns_1(ces_4_1_io_lsbIns_1),
    .io_lsbIns_2(ces_4_1_io_lsbIns_2),
    .io_lsbIns_3(ces_4_1_io_lsbIns_3),
    .io_lsbIns_4(ces_4_1_io_lsbIns_4),
    .io_lsbIns_5(ces_4_1_io_lsbIns_5),
    .io_lsbIns_6(ces_4_1_io_lsbIns_6),
    .io_lsbIns_7(ces_4_1_io_lsbIns_7),
    .io_lsbOuts_0(ces_4_1_io_lsbOuts_0),
    .io_lsbOuts_1(ces_4_1_io_lsbOuts_1),
    .io_lsbOuts_2(ces_4_1_io_lsbOuts_2),
    .io_lsbOuts_3(ces_4_1_io_lsbOuts_3),
    .io_lsbOuts_4(ces_4_1_io_lsbOuts_4),
    .io_lsbOuts_5(ces_4_1_io_lsbOuts_5),
    .io_lsbOuts_6(ces_4_1_io_lsbOuts_6),
    .io_lsbOuts_7(ces_4_1_io_lsbOuts_7)
  );
  Element ces_4_2 (
    .clock(ces_4_2_clock),
    .io_clockOutRight(ces_4_2_io_clockOutRight),
    .io_ins_down(ces_4_2_io_ins_down),
    .io_ins_right(ces_4_2_io_ins_right),
    .io_ins_up(ces_4_2_io_ins_up),
    .io_ins_left(ces_4_2_io_ins_left),
    .io_outs_down(ces_4_2_io_outs_down),
    .io_outs_right(ces_4_2_io_outs_right),
    .io_outs_up(ces_4_2_io_outs_up),
    .io_outs_left(ces_4_2_io_outs_left),
    .io_lsbIns_1(ces_4_2_io_lsbIns_1),
    .io_lsbIns_2(ces_4_2_io_lsbIns_2),
    .io_lsbIns_3(ces_4_2_io_lsbIns_3),
    .io_lsbIns_4(ces_4_2_io_lsbIns_4),
    .io_lsbIns_5(ces_4_2_io_lsbIns_5),
    .io_lsbIns_6(ces_4_2_io_lsbIns_6),
    .io_lsbIns_7(ces_4_2_io_lsbIns_7),
    .io_lsbOuts_0(ces_4_2_io_lsbOuts_0),
    .io_lsbOuts_1(ces_4_2_io_lsbOuts_1),
    .io_lsbOuts_2(ces_4_2_io_lsbOuts_2),
    .io_lsbOuts_3(ces_4_2_io_lsbOuts_3),
    .io_lsbOuts_4(ces_4_2_io_lsbOuts_4),
    .io_lsbOuts_5(ces_4_2_io_lsbOuts_5),
    .io_lsbOuts_6(ces_4_2_io_lsbOuts_6),
    .io_lsbOuts_7(ces_4_2_io_lsbOuts_7)
  );
  Element ces_4_3 (
    .clock(ces_4_3_clock),
    .io_clockOutRight(ces_4_3_io_clockOutRight),
    .io_ins_down(ces_4_3_io_ins_down),
    .io_ins_right(ces_4_3_io_ins_right),
    .io_ins_up(ces_4_3_io_ins_up),
    .io_ins_left(ces_4_3_io_ins_left),
    .io_outs_down(ces_4_3_io_outs_down),
    .io_outs_right(ces_4_3_io_outs_right),
    .io_outs_up(ces_4_3_io_outs_up),
    .io_outs_left(ces_4_3_io_outs_left),
    .io_lsbIns_1(ces_4_3_io_lsbIns_1),
    .io_lsbIns_2(ces_4_3_io_lsbIns_2),
    .io_lsbIns_3(ces_4_3_io_lsbIns_3),
    .io_lsbIns_4(ces_4_3_io_lsbIns_4),
    .io_lsbIns_5(ces_4_3_io_lsbIns_5),
    .io_lsbIns_6(ces_4_3_io_lsbIns_6),
    .io_lsbIns_7(ces_4_3_io_lsbIns_7),
    .io_lsbOuts_0(ces_4_3_io_lsbOuts_0),
    .io_lsbOuts_1(ces_4_3_io_lsbOuts_1),
    .io_lsbOuts_2(ces_4_3_io_lsbOuts_2),
    .io_lsbOuts_3(ces_4_3_io_lsbOuts_3),
    .io_lsbOuts_4(ces_4_3_io_lsbOuts_4),
    .io_lsbOuts_5(ces_4_3_io_lsbOuts_5),
    .io_lsbOuts_6(ces_4_3_io_lsbOuts_6),
    .io_lsbOuts_7(ces_4_3_io_lsbOuts_7)
  );
  Element ces_4_4 (
    .clock(ces_4_4_clock),
    .io_clockOutRight(ces_4_4_io_clockOutRight),
    .io_ins_down(ces_4_4_io_ins_down),
    .io_ins_right(ces_4_4_io_ins_right),
    .io_ins_up(ces_4_4_io_ins_up),
    .io_ins_left(ces_4_4_io_ins_left),
    .io_outs_down(ces_4_4_io_outs_down),
    .io_outs_right(ces_4_4_io_outs_right),
    .io_outs_up(ces_4_4_io_outs_up),
    .io_outs_left(ces_4_4_io_outs_left),
    .io_lsbIns_1(ces_4_4_io_lsbIns_1),
    .io_lsbIns_2(ces_4_4_io_lsbIns_2),
    .io_lsbIns_3(ces_4_4_io_lsbIns_3),
    .io_lsbIns_4(ces_4_4_io_lsbIns_4),
    .io_lsbIns_5(ces_4_4_io_lsbIns_5),
    .io_lsbIns_6(ces_4_4_io_lsbIns_6),
    .io_lsbIns_7(ces_4_4_io_lsbIns_7),
    .io_lsbOuts_0(ces_4_4_io_lsbOuts_0),
    .io_lsbOuts_1(ces_4_4_io_lsbOuts_1),
    .io_lsbOuts_2(ces_4_4_io_lsbOuts_2),
    .io_lsbOuts_3(ces_4_4_io_lsbOuts_3),
    .io_lsbOuts_4(ces_4_4_io_lsbOuts_4),
    .io_lsbOuts_5(ces_4_4_io_lsbOuts_5),
    .io_lsbOuts_6(ces_4_4_io_lsbOuts_6),
    .io_lsbOuts_7(ces_4_4_io_lsbOuts_7)
  );
  Element ces_4_5 (
    .clock(ces_4_5_clock),
    .io_clockOutRight(ces_4_5_io_clockOutRight),
    .io_ins_down(ces_4_5_io_ins_down),
    .io_ins_right(ces_4_5_io_ins_right),
    .io_ins_up(ces_4_5_io_ins_up),
    .io_ins_left(ces_4_5_io_ins_left),
    .io_outs_down(ces_4_5_io_outs_down),
    .io_outs_right(ces_4_5_io_outs_right),
    .io_outs_up(ces_4_5_io_outs_up),
    .io_outs_left(ces_4_5_io_outs_left),
    .io_lsbIns_1(ces_4_5_io_lsbIns_1),
    .io_lsbIns_2(ces_4_5_io_lsbIns_2),
    .io_lsbIns_3(ces_4_5_io_lsbIns_3),
    .io_lsbIns_4(ces_4_5_io_lsbIns_4),
    .io_lsbIns_5(ces_4_5_io_lsbIns_5),
    .io_lsbIns_6(ces_4_5_io_lsbIns_6),
    .io_lsbIns_7(ces_4_5_io_lsbIns_7),
    .io_lsbOuts_0(ces_4_5_io_lsbOuts_0),
    .io_lsbOuts_1(ces_4_5_io_lsbOuts_1),
    .io_lsbOuts_2(ces_4_5_io_lsbOuts_2),
    .io_lsbOuts_3(ces_4_5_io_lsbOuts_3),
    .io_lsbOuts_4(ces_4_5_io_lsbOuts_4),
    .io_lsbOuts_5(ces_4_5_io_lsbOuts_5),
    .io_lsbOuts_6(ces_4_5_io_lsbOuts_6),
    .io_lsbOuts_7(ces_4_5_io_lsbOuts_7)
  );
  Element ces_4_6 (
    .clock(ces_4_6_clock),
    .io_clockOutRight(ces_4_6_io_clockOutRight),
    .io_ins_down(ces_4_6_io_ins_down),
    .io_ins_right(ces_4_6_io_ins_right),
    .io_ins_up(ces_4_6_io_ins_up),
    .io_ins_left(ces_4_6_io_ins_left),
    .io_outs_down(ces_4_6_io_outs_down),
    .io_outs_right(ces_4_6_io_outs_right),
    .io_outs_up(ces_4_6_io_outs_up),
    .io_outs_left(ces_4_6_io_outs_left),
    .io_lsbIns_1(ces_4_6_io_lsbIns_1),
    .io_lsbIns_2(ces_4_6_io_lsbIns_2),
    .io_lsbIns_3(ces_4_6_io_lsbIns_3),
    .io_lsbIns_4(ces_4_6_io_lsbIns_4),
    .io_lsbIns_5(ces_4_6_io_lsbIns_5),
    .io_lsbIns_6(ces_4_6_io_lsbIns_6),
    .io_lsbIns_7(ces_4_6_io_lsbIns_7),
    .io_lsbOuts_0(ces_4_6_io_lsbOuts_0),
    .io_lsbOuts_1(ces_4_6_io_lsbOuts_1),
    .io_lsbOuts_2(ces_4_6_io_lsbOuts_2),
    .io_lsbOuts_3(ces_4_6_io_lsbOuts_3),
    .io_lsbOuts_4(ces_4_6_io_lsbOuts_4),
    .io_lsbOuts_5(ces_4_6_io_lsbOuts_5),
    .io_lsbOuts_6(ces_4_6_io_lsbOuts_6),
    .io_lsbOuts_7(ces_4_6_io_lsbOuts_7)
  );
  Element ces_4_7 (
    .clock(ces_4_7_clock),
    .io_clockOutRight(ces_4_7_io_clockOutRight),
    .io_ins_down(ces_4_7_io_ins_down),
    .io_ins_right(ces_4_7_io_ins_right),
    .io_ins_up(ces_4_7_io_ins_up),
    .io_ins_left(ces_4_7_io_ins_left),
    .io_outs_down(ces_4_7_io_outs_down),
    .io_outs_right(ces_4_7_io_outs_right),
    .io_outs_up(ces_4_7_io_outs_up),
    .io_outs_left(ces_4_7_io_outs_left),
    .io_lsbIns_1(ces_4_7_io_lsbIns_1),
    .io_lsbIns_2(ces_4_7_io_lsbIns_2),
    .io_lsbIns_3(ces_4_7_io_lsbIns_3),
    .io_lsbIns_4(ces_4_7_io_lsbIns_4),
    .io_lsbIns_5(ces_4_7_io_lsbIns_5),
    .io_lsbIns_6(ces_4_7_io_lsbIns_6),
    .io_lsbIns_7(ces_4_7_io_lsbIns_7),
    .io_lsbOuts_0(ces_4_7_io_lsbOuts_0),
    .io_lsbOuts_1(ces_4_7_io_lsbOuts_1),
    .io_lsbOuts_2(ces_4_7_io_lsbOuts_2),
    .io_lsbOuts_3(ces_4_7_io_lsbOuts_3),
    .io_lsbOuts_4(ces_4_7_io_lsbOuts_4),
    .io_lsbOuts_5(ces_4_7_io_lsbOuts_5),
    .io_lsbOuts_6(ces_4_7_io_lsbOuts_6),
    .io_lsbOuts_7(ces_4_7_io_lsbOuts_7)
  );
  Element ces_5_0 (
    .clock(ces_5_0_clock),
    .io_clockOutRight(ces_5_0_io_clockOutRight),
    .io_ins_down(ces_5_0_io_ins_down),
    .io_ins_right(ces_5_0_io_ins_right),
    .io_ins_up(ces_5_0_io_ins_up),
    .io_ins_left(ces_5_0_io_ins_left),
    .io_outs_down(ces_5_0_io_outs_down),
    .io_outs_right(ces_5_0_io_outs_right),
    .io_outs_up(ces_5_0_io_outs_up),
    .io_outs_left(ces_5_0_io_outs_left),
    .io_lsbIns_1(ces_5_0_io_lsbIns_1),
    .io_lsbIns_2(ces_5_0_io_lsbIns_2),
    .io_lsbIns_3(ces_5_0_io_lsbIns_3),
    .io_lsbIns_4(ces_5_0_io_lsbIns_4),
    .io_lsbIns_5(ces_5_0_io_lsbIns_5),
    .io_lsbIns_6(ces_5_0_io_lsbIns_6),
    .io_lsbIns_7(ces_5_0_io_lsbIns_7),
    .io_lsbOuts_0(ces_5_0_io_lsbOuts_0),
    .io_lsbOuts_1(ces_5_0_io_lsbOuts_1),
    .io_lsbOuts_2(ces_5_0_io_lsbOuts_2),
    .io_lsbOuts_3(ces_5_0_io_lsbOuts_3),
    .io_lsbOuts_4(ces_5_0_io_lsbOuts_4),
    .io_lsbOuts_5(ces_5_0_io_lsbOuts_5),
    .io_lsbOuts_6(ces_5_0_io_lsbOuts_6),
    .io_lsbOuts_7(ces_5_0_io_lsbOuts_7)
  );
  Element ces_5_1 (
    .clock(ces_5_1_clock),
    .io_clockOutRight(ces_5_1_io_clockOutRight),
    .io_ins_down(ces_5_1_io_ins_down),
    .io_ins_right(ces_5_1_io_ins_right),
    .io_ins_up(ces_5_1_io_ins_up),
    .io_ins_left(ces_5_1_io_ins_left),
    .io_outs_down(ces_5_1_io_outs_down),
    .io_outs_right(ces_5_1_io_outs_right),
    .io_outs_up(ces_5_1_io_outs_up),
    .io_outs_left(ces_5_1_io_outs_left),
    .io_lsbIns_1(ces_5_1_io_lsbIns_1),
    .io_lsbIns_2(ces_5_1_io_lsbIns_2),
    .io_lsbIns_3(ces_5_1_io_lsbIns_3),
    .io_lsbIns_4(ces_5_1_io_lsbIns_4),
    .io_lsbIns_5(ces_5_1_io_lsbIns_5),
    .io_lsbIns_6(ces_5_1_io_lsbIns_6),
    .io_lsbIns_7(ces_5_1_io_lsbIns_7),
    .io_lsbOuts_0(ces_5_1_io_lsbOuts_0),
    .io_lsbOuts_1(ces_5_1_io_lsbOuts_1),
    .io_lsbOuts_2(ces_5_1_io_lsbOuts_2),
    .io_lsbOuts_3(ces_5_1_io_lsbOuts_3),
    .io_lsbOuts_4(ces_5_1_io_lsbOuts_4),
    .io_lsbOuts_5(ces_5_1_io_lsbOuts_5),
    .io_lsbOuts_6(ces_5_1_io_lsbOuts_6),
    .io_lsbOuts_7(ces_5_1_io_lsbOuts_7)
  );
  Element ces_5_2 (
    .clock(ces_5_2_clock),
    .io_clockOutRight(ces_5_2_io_clockOutRight),
    .io_ins_down(ces_5_2_io_ins_down),
    .io_ins_right(ces_5_2_io_ins_right),
    .io_ins_up(ces_5_2_io_ins_up),
    .io_ins_left(ces_5_2_io_ins_left),
    .io_outs_down(ces_5_2_io_outs_down),
    .io_outs_right(ces_5_2_io_outs_right),
    .io_outs_up(ces_5_2_io_outs_up),
    .io_outs_left(ces_5_2_io_outs_left),
    .io_lsbIns_1(ces_5_2_io_lsbIns_1),
    .io_lsbIns_2(ces_5_2_io_lsbIns_2),
    .io_lsbIns_3(ces_5_2_io_lsbIns_3),
    .io_lsbIns_4(ces_5_2_io_lsbIns_4),
    .io_lsbIns_5(ces_5_2_io_lsbIns_5),
    .io_lsbIns_6(ces_5_2_io_lsbIns_6),
    .io_lsbIns_7(ces_5_2_io_lsbIns_7),
    .io_lsbOuts_0(ces_5_2_io_lsbOuts_0),
    .io_lsbOuts_1(ces_5_2_io_lsbOuts_1),
    .io_lsbOuts_2(ces_5_2_io_lsbOuts_2),
    .io_lsbOuts_3(ces_5_2_io_lsbOuts_3),
    .io_lsbOuts_4(ces_5_2_io_lsbOuts_4),
    .io_lsbOuts_5(ces_5_2_io_lsbOuts_5),
    .io_lsbOuts_6(ces_5_2_io_lsbOuts_6),
    .io_lsbOuts_7(ces_5_2_io_lsbOuts_7)
  );
  Element ces_5_3 (
    .clock(ces_5_3_clock),
    .io_clockOutRight(ces_5_3_io_clockOutRight),
    .io_ins_down(ces_5_3_io_ins_down),
    .io_ins_right(ces_5_3_io_ins_right),
    .io_ins_up(ces_5_3_io_ins_up),
    .io_ins_left(ces_5_3_io_ins_left),
    .io_outs_down(ces_5_3_io_outs_down),
    .io_outs_right(ces_5_3_io_outs_right),
    .io_outs_up(ces_5_3_io_outs_up),
    .io_outs_left(ces_5_3_io_outs_left),
    .io_lsbIns_1(ces_5_3_io_lsbIns_1),
    .io_lsbIns_2(ces_5_3_io_lsbIns_2),
    .io_lsbIns_3(ces_5_3_io_lsbIns_3),
    .io_lsbIns_4(ces_5_3_io_lsbIns_4),
    .io_lsbIns_5(ces_5_3_io_lsbIns_5),
    .io_lsbIns_6(ces_5_3_io_lsbIns_6),
    .io_lsbIns_7(ces_5_3_io_lsbIns_7),
    .io_lsbOuts_0(ces_5_3_io_lsbOuts_0),
    .io_lsbOuts_1(ces_5_3_io_lsbOuts_1),
    .io_lsbOuts_2(ces_5_3_io_lsbOuts_2),
    .io_lsbOuts_3(ces_5_3_io_lsbOuts_3),
    .io_lsbOuts_4(ces_5_3_io_lsbOuts_4),
    .io_lsbOuts_5(ces_5_3_io_lsbOuts_5),
    .io_lsbOuts_6(ces_5_3_io_lsbOuts_6),
    .io_lsbOuts_7(ces_5_3_io_lsbOuts_7)
  );
  Element ces_5_4 (
    .clock(ces_5_4_clock),
    .io_clockOutRight(ces_5_4_io_clockOutRight),
    .io_ins_down(ces_5_4_io_ins_down),
    .io_ins_right(ces_5_4_io_ins_right),
    .io_ins_up(ces_5_4_io_ins_up),
    .io_ins_left(ces_5_4_io_ins_left),
    .io_outs_down(ces_5_4_io_outs_down),
    .io_outs_right(ces_5_4_io_outs_right),
    .io_outs_up(ces_5_4_io_outs_up),
    .io_outs_left(ces_5_4_io_outs_left),
    .io_lsbIns_1(ces_5_4_io_lsbIns_1),
    .io_lsbIns_2(ces_5_4_io_lsbIns_2),
    .io_lsbIns_3(ces_5_4_io_lsbIns_3),
    .io_lsbIns_4(ces_5_4_io_lsbIns_4),
    .io_lsbIns_5(ces_5_4_io_lsbIns_5),
    .io_lsbIns_6(ces_5_4_io_lsbIns_6),
    .io_lsbIns_7(ces_5_4_io_lsbIns_7),
    .io_lsbOuts_0(ces_5_4_io_lsbOuts_0),
    .io_lsbOuts_1(ces_5_4_io_lsbOuts_1),
    .io_lsbOuts_2(ces_5_4_io_lsbOuts_2),
    .io_lsbOuts_3(ces_5_4_io_lsbOuts_3),
    .io_lsbOuts_4(ces_5_4_io_lsbOuts_4),
    .io_lsbOuts_5(ces_5_4_io_lsbOuts_5),
    .io_lsbOuts_6(ces_5_4_io_lsbOuts_6),
    .io_lsbOuts_7(ces_5_4_io_lsbOuts_7)
  );
  Element ces_5_5 (
    .clock(ces_5_5_clock),
    .io_clockOutRight(ces_5_5_io_clockOutRight),
    .io_ins_down(ces_5_5_io_ins_down),
    .io_ins_right(ces_5_5_io_ins_right),
    .io_ins_up(ces_5_5_io_ins_up),
    .io_ins_left(ces_5_5_io_ins_left),
    .io_outs_down(ces_5_5_io_outs_down),
    .io_outs_right(ces_5_5_io_outs_right),
    .io_outs_up(ces_5_5_io_outs_up),
    .io_outs_left(ces_5_5_io_outs_left),
    .io_lsbIns_1(ces_5_5_io_lsbIns_1),
    .io_lsbIns_2(ces_5_5_io_lsbIns_2),
    .io_lsbIns_3(ces_5_5_io_lsbIns_3),
    .io_lsbIns_4(ces_5_5_io_lsbIns_4),
    .io_lsbIns_5(ces_5_5_io_lsbIns_5),
    .io_lsbIns_6(ces_5_5_io_lsbIns_6),
    .io_lsbIns_7(ces_5_5_io_lsbIns_7),
    .io_lsbOuts_0(ces_5_5_io_lsbOuts_0),
    .io_lsbOuts_1(ces_5_5_io_lsbOuts_1),
    .io_lsbOuts_2(ces_5_5_io_lsbOuts_2),
    .io_lsbOuts_3(ces_5_5_io_lsbOuts_3),
    .io_lsbOuts_4(ces_5_5_io_lsbOuts_4),
    .io_lsbOuts_5(ces_5_5_io_lsbOuts_5),
    .io_lsbOuts_6(ces_5_5_io_lsbOuts_6),
    .io_lsbOuts_7(ces_5_5_io_lsbOuts_7)
  );
  Element ces_5_6 (
    .clock(ces_5_6_clock),
    .io_clockOutRight(ces_5_6_io_clockOutRight),
    .io_ins_down(ces_5_6_io_ins_down),
    .io_ins_right(ces_5_6_io_ins_right),
    .io_ins_up(ces_5_6_io_ins_up),
    .io_ins_left(ces_5_6_io_ins_left),
    .io_outs_down(ces_5_6_io_outs_down),
    .io_outs_right(ces_5_6_io_outs_right),
    .io_outs_up(ces_5_6_io_outs_up),
    .io_outs_left(ces_5_6_io_outs_left),
    .io_lsbIns_1(ces_5_6_io_lsbIns_1),
    .io_lsbIns_2(ces_5_6_io_lsbIns_2),
    .io_lsbIns_3(ces_5_6_io_lsbIns_3),
    .io_lsbIns_4(ces_5_6_io_lsbIns_4),
    .io_lsbIns_5(ces_5_6_io_lsbIns_5),
    .io_lsbIns_6(ces_5_6_io_lsbIns_6),
    .io_lsbIns_7(ces_5_6_io_lsbIns_7),
    .io_lsbOuts_0(ces_5_6_io_lsbOuts_0),
    .io_lsbOuts_1(ces_5_6_io_lsbOuts_1),
    .io_lsbOuts_2(ces_5_6_io_lsbOuts_2),
    .io_lsbOuts_3(ces_5_6_io_lsbOuts_3),
    .io_lsbOuts_4(ces_5_6_io_lsbOuts_4),
    .io_lsbOuts_5(ces_5_6_io_lsbOuts_5),
    .io_lsbOuts_6(ces_5_6_io_lsbOuts_6),
    .io_lsbOuts_7(ces_5_6_io_lsbOuts_7)
  );
  Element ces_5_7 (
    .clock(ces_5_7_clock),
    .io_clockOutRight(ces_5_7_io_clockOutRight),
    .io_ins_down(ces_5_7_io_ins_down),
    .io_ins_right(ces_5_7_io_ins_right),
    .io_ins_up(ces_5_7_io_ins_up),
    .io_ins_left(ces_5_7_io_ins_left),
    .io_outs_down(ces_5_7_io_outs_down),
    .io_outs_right(ces_5_7_io_outs_right),
    .io_outs_up(ces_5_7_io_outs_up),
    .io_outs_left(ces_5_7_io_outs_left),
    .io_lsbIns_1(ces_5_7_io_lsbIns_1),
    .io_lsbIns_2(ces_5_7_io_lsbIns_2),
    .io_lsbIns_3(ces_5_7_io_lsbIns_3),
    .io_lsbIns_4(ces_5_7_io_lsbIns_4),
    .io_lsbIns_5(ces_5_7_io_lsbIns_5),
    .io_lsbIns_6(ces_5_7_io_lsbIns_6),
    .io_lsbIns_7(ces_5_7_io_lsbIns_7),
    .io_lsbOuts_0(ces_5_7_io_lsbOuts_0),
    .io_lsbOuts_1(ces_5_7_io_lsbOuts_1),
    .io_lsbOuts_2(ces_5_7_io_lsbOuts_2),
    .io_lsbOuts_3(ces_5_7_io_lsbOuts_3),
    .io_lsbOuts_4(ces_5_7_io_lsbOuts_4),
    .io_lsbOuts_5(ces_5_7_io_lsbOuts_5),
    .io_lsbOuts_6(ces_5_7_io_lsbOuts_6),
    .io_lsbOuts_7(ces_5_7_io_lsbOuts_7)
  );
  Element ces_6_0 (
    .clock(ces_6_0_clock),
    .io_clockOutRight(ces_6_0_io_clockOutRight),
    .io_ins_down(ces_6_0_io_ins_down),
    .io_ins_right(ces_6_0_io_ins_right),
    .io_ins_up(ces_6_0_io_ins_up),
    .io_ins_left(ces_6_0_io_ins_left),
    .io_outs_down(ces_6_0_io_outs_down),
    .io_outs_right(ces_6_0_io_outs_right),
    .io_outs_up(ces_6_0_io_outs_up),
    .io_outs_left(ces_6_0_io_outs_left),
    .io_lsbIns_1(ces_6_0_io_lsbIns_1),
    .io_lsbIns_2(ces_6_0_io_lsbIns_2),
    .io_lsbIns_3(ces_6_0_io_lsbIns_3),
    .io_lsbIns_4(ces_6_0_io_lsbIns_4),
    .io_lsbIns_5(ces_6_0_io_lsbIns_5),
    .io_lsbIns_6(ces_6_0_io_lsbIns_6),
    .io_lsbIns_7(ces_6_0_io_lsbIns_7),
    .io_lsbOuts_0(ces_6_0_io_lsbOuts_0),
    .io_lsbOuts_1(ces_6_0_io_lsbOuts_1),
    .io_lsbOuts_2(ces_6_0_io_lsbOuts_2),
    .io_lsbOuts_3(ces_6_0_io_lsbOuts_3),
    .io_lsbOuts_4(ces_6_0_io_lsbOuts_4),
    .io_lsbOuts_5(ces_6_0_io_lsbOuts_5),
    .io_lsbOuts_6(ces_6_0_io_lsbOuts_6),
    .io_lsbOuts_7(ces_6_0_io_lsbOuts_7)
  );
  Element ces_6_1 (
    .clock(ces_6_1_clock),
    .io_clockOutRight(ces_6_1_io_clockOutRight),
    .io_ins_down(ces_6_1_io_ins_down),
    .io_ins_right(ces_6_1_io_ins_right),
    .io_ins_up(ces_6_1_io_ins_up),
    .io_ins_left(ces_6_1_io_ins_left),
    .io_outs_down(ces_6_1_io_outs_down),
    .io_outs_right(ces_6_1_io_outs_right),
    .io_outs_up(ces_6_1_io_outs_up),
    .io_outs_left(ces_6_1_io_outs_left),
    .io_lsbIns_1(ces_6_1_io_lsbIns_1),
    .io_lsbIns_2(ces_6_1_io_lsbIns_2),
    .io_lsbIns_3(ces_6_1_io_lsbIns_3),
    .io_lsbIns_4(ces_6_1_io_lsbIns_4),
    .io_lsbIns_5(ces_6_1_io_lsbIns_5),
    .io_lsbIns_6(ces_6_1_io_lsbIns_6),
    .io_lsbIns_7(ces_6_1_io_lsbIns_7),
    .io_lsbOuts_0(ces_6_1_io_lsbOuts_0),
    .io_lsbOuts_1(ces_6_1_io_lsbOuts_1),
    .io_lsbOuts_2(ces_6_1_io_lsbOuts_2),
    .io_lsbOuts_3(ces_6_1_io_lsbOuts_3),
    .io_lsbOuts_4(ces_6_1_io_lsbOuts_4),
    .io_lsbOuts_5(ces_6_1_io_lsbOuts_5),
    .io_lsbOuts_6(ces_6_1_io_lsbOuts_6),
    .io_lsbOuts_7(ces_6_1_io_lsbOuts_7)
  );
  Element ces_6_2 (
    .clock(ces_6_2_clock),
    .io_clockOutRight(ces_6_2_io_clockOutRight),
    .io_ins_down(ces_6_2_io_ins_down),
    .io_ins_right(ces_6_2_io_ins_right),
    .io_ins_up(ces_6_2_io_ins_up),
    .io_ins_left(ces_6_2_io_ins_left),
    .io_outs_down(ces_6_2_io_outs_down),
    .io_outs_right(ces_6_2_io_outs_right),
    .io_outs_up(ces_6_2_io_outs_up),
    .io_outs_left(ces_6_2_io_outs_left),
    .io_lsbIns_1(ces_6_2_io_lsbIns_1),
    .io_lsbIns_2(ces_6_2_io_lsbIns_2),
    .io_lsbIns_3(ces_6_2_io_lsbIns_3),
    .io_lsbIns_4(ces_6_2_io_lsbIns_4),
    .io_lsbIns_5(ces_6_2_io_lsbIns_5),
    .io_lsbIns_6(ces_6_2_io_lsbIns_6),
    .io_lsbIns_7(ces_6_2_io_lsbIns_7),
    .io_lsbOuts_0(ces_6_2_io_lsbOuts_0),
    .io_lsbOuts_1(ces_6_2_io_lsbOuts_1),
    .io_lsbOuts_2(ces_6_2_io_lsbOuts_2),
    .io_lsbOuts_3(ces_6_2_io_lsbOuts_3),
    .io_lsbOuts_4(ces_6_2_io_lsbOuts_4),
    .io_lsbOuts_5(ces_6_2_io_lsbOuts_5),
    .io_lsbOuts_6(ces_6_2_io_lsbOuts_6),
    .io_lsbOuts_7(ces_6_2_io_lsbOuts_7)
  );
  Element ces_6_3 (
    .clock(ces_6_3_clock),
    .io_clockOutRight(ces_6_3_io_clockOutRight),
    .io_ins_down(ces_6_3_io_ins_down),
    .io_ins_right(ces_6_3_io_ins_right),
    .io_ins_up(ces_6_3_io_ins_up),
    .io_ins_left(ces_6_3_io_ins_left),
    .io_outs_down(ces_6_3_io_outs_down),
    .io_outs_right(ces_6_3_io_outs_right),
    .io_outs_up(ces_6_3_io_outs_up),
    .io_outs_left(ces_6_3_io_outs_left),
    .io_lsbIns_1(ces_6_3_io_lsbIns_1),
    .io_lsbIns_2(ces_6_3_io_lsbIns_2),
    .io_lsbIns_3(ces_6_3_io_lsbIns_3),
    .io_lsbIns_4(ces_6_3_io_lsbIns_4),
    .io_lsbIns_5(ces_6_3_io_lsbIns_5),
    .io_lsbIns_6(ces_6_3_io_lsbIns_6),
    .io_lsbIns_7(ces_6_3_io_lsbIns_7),
    .io_lsbOuts_0(ces_6_3_io_lsbOuts_0),
    .io_lsbOuts_1(ces_6_3_io_lsbOuts_1),
    .io_lsbOuts_2(ces_6_3_io_lsbOuts_2),
    .io_lsbOuts_3(ces_6_3_io_lsbOuts_3),
    .io_lsbOuts_4(ces_6_3_io_lsbOuts_4),
    .io_lsbOuts_5(ces_6_3_io_lsbOuts_5),
    .io_lsbOuts_6(ces_6_3_io_lsbOuts_6),
    .io_lsbOuts_7(ces_6_3_io_lsbOuts_7)
  );
  Element ces_6_4 (
    .clock(ces_6_4_clock),
    .io_clockOutRight(ces_6_4_io_clockOutRight),
    .io_ins_down(ces_6_4_io_ins_down),
    .io_ins_right(ces_6_4_io_ins_right),
    .io_ins_up(ces_6_4_io_ins_up),
    .io_ins_left(ces_6_4_io_ins_left),
    .io_outs_down(ces_6_4_io_outs_down),
    .io_outs_right(ces_6_4_io_outs_right),
    .io_outs_up(ces_6_4_io_outs_up),
    .io_outs_left(ces_6_4_io_outs_left),
    .io_lsbIns_1(ces_6_4_io_lsbIns_1),
    .io_lsbIns_2(ces_6_4_io_lsbIns_2),
    .io_lsbIns_3(ces_6_4_io_lsbIns_3),
    .io_lsbIns_4(ces_6_4_io_lsbIns_4),
    .io_lsbIns_5(ces_6_4_io_lsbIns_5),
    .io_lsbIns_6(ces_6_4_io_lsbIns_6),
    .io_lsbIns_7(ces_6_4_io_lsbIns_7),
    .io_lsbOuts_0(ces_6_4_io_lsbOuts_0),
    .io_lsbOuts_1(ces_6_4_io_lsbOuts_1),
    .io_lsbOuts_2(ces_6_4_io_lsbOuts_2),
    .io_lsbOuts_3(ces_6_4_io_lsbOuts_3),
    .io_lsbOuts_4(ces_6_4_io_lsbOuts_4),
    .io_lsbOuts_5(ces_6_4_io_lsbOuts_5),
    .io_lsbOuts_6(ces_6_4_io_lsbOuts_6),
    .io_lsbOuts_7(ces_6_4_io_lsbOuts_7)
  );
  Element ces_6_5 (
    .clock(ces_6_5_clock),
    .io_clockOutRight(ces_6_5_io_clockOutRight),
    .io_ins_down(ces_6_5_io_ins_down),
    .io_ins_right(ces_6_5_io_ins_right),
    .io_ins_up(ces_6_5_io_ins_up),
    .io_ins_left(ces_6_5_io_ins_left),
    .io_outs_down(ces_6_5_io_outs_down),
    .io_outs_right(ces_6_5_io_outs_right),
    .io_outs_up(ces_6_5_io_outs_up),
    .io_outs_left(ces_6_5_io_outs_left),
    .io_lsbIns_1(ces_6_5_io_lsbIns_1),
    .io_lsbIns_2(ces_6_5_io_lsbIns_2),
    .io_lsbIns_3(ces_6_5_io_lsbIns_3),
    .io_lsbIns_4(ces_6_5_io_lsbIns_4),
    .io_lsbIns_5(ces_6_5_io_lsbIns_5),
    .io_lsbIns_6(ces_6_5_io_lsbIns_6),
    .io_lsbIns_7(ces_6_5_io_lsbIns_7),
    .io_lsbOuts_0(ces_6_5_io_lsbOuts_0),
    .io_lsbOuts_1(ces_6_5_io_lsbOuts_1),
    .io_lsbOuts_2(ces_6_5_io_lsbOuts_2),
    .io_lsbOuts_3(ces_6_5_io_lsbOuts_3),
    .io_lsbOuts_4(ces_6_5_io_lsbOuts_4),
    .io_lsbOuts_5(ces_6_5_io_lsbOuts_5),
    .io_lsbOuts_6(ces_6_5_io_lsbOuts_6),
    .io_lsbOuts_7(ces_6_5_io_lsbOuts_7)
  );
  Element ces_6_6 (
    .clock(ces_6_6_clock),
    .io_clockOutRight(ces_6_6_io_clockOutRight),
    .io_ins_down(ces_6_6_io_ins_down),
    .io_ins_right(ces_6_6_io_ins_right),
    .io_ins_up(ces_6_6_io_ins_up),
    .io_ins_left(ces_6_6_io_ins_left),
    .io_outs_down(ces_6_6_io_outs_down),
    .io_outs_right(ces_6_6_io_outs_right),
    .io_outs_up(ces_6_6_io_outs_up),
    .io_outs_left(ces_6_6_io_outs_left),
    .io_lsbIns_1(ces_6_6_io_lsbIns_1),
    .io_lsbIns_2(ces_6_6_io_lsbIns_2),
    .io_lsbIns_3(ces_6_6_io_lsbIns_3),
    .io_lsbIns_4(ces_6_6_io_lsbIns_4),
    .io_lsbIns_5(ces_6_6_io_lsbIns_5),
    .io_lsbIns_6(ces_6_6_io_lsbIns_6),
    .io_lsbIns_7(ces_6_6_io_lsbIns_7),
    .io_lsbOuts_0(ces_6_6_io_lsbOuts_0),
    .io_lsbOuts_1(ces_6_6_io_lsbOuts_1),
    .io_lsbOuts_2(ces_6_6_io_lsbOuts_2),
    .io_lsbOuts_3(ces_6_6_io_lsbOuts_3),
    .io_lsbOuts_4(ces_6_6_io_lsbOuts_4),
    .io_lsbOuts_5(ces_6_6_io_lsbOuts_5),
    .io_lsbOuts_6(ces_6_6_io_lsbOuts_6),
    .io_lsbOuts_7(ces_6_6_io_lsbOuts_7)
  );
  Element ces_6_7 (
    .clock(ces_6_7_clock),
    .io_clockOutRight(ces_6_7_io_clockOutRight),
    .io_ins_down(ces_6_7_io_ins_down),
    .io_ins_right(ces_6_7_io_ins_right),
    .io_ins_up(ces_6_7_io_ins_up),
    .io_ins_left(ces_6_7_io_ins_left),
    .io_outs_down(ces_6_7_io_outs_down),
    .io_outs_right(ces_6_7_io_outs_right),
    .io_outs_up(ces_6_7_io_outs_up),
    .io_outs_left(ces_6_7_io_outs_left),
    .io_lsbIns_1(ces_6_7_io_lsbIns_1),
    .io_lsbIns_2(ces_6_7_io_lsbIns_2),
    .io_lsbIns_3(ces_6_7_io_lsbIns_3),
    .io_lsbIns_4(ces_6_7_io_lsbIns_4),
    .io_lsbIns_5(ces_6_7_io_lsbIns_5),
    .io_lsbIns_6(ces_6_7_io_lsbIns_6),
    .io_lsbIns_7(ces_6_7_io_lsbIns_7),
    .io_lsbOuts_0(ces_6_7_io_lsbOuts_0),
    .io_lsbOuts_1(ces_6_7_io_lsbOuts_1),
    .io_lsbOuts_2(ces_6_7_io_lsbOuts_2),
    .io_lsbOuts_3(ces_6_7_io_lsbOuts_3),
    .io_lsbOuts_4(ces_6_7_io_lsbOuts_4),
    .io_lsbOuts_5(ces_6_7_io_lsbOuts_5),
    .io_lsbOuts_6(ces_6_7_io_lsbOuts_6),
    .io_lsbOuts_7(ces_6_7_io_lsbOuts_7)
  );
  Element ces_7_0 (
    .clock(ces_7_0_clock),
    .io_clockOutRight(ces_7_0_io_clockOutRight),
    .io_ins_down(ces_7_0_io_ins_down),
    .io_ins_right(ces_7_0_io_ins_right),
    .io_ins_up(ces_7_0_io_ins_up),
    .io_ins_left(ces_7_0_io_ins_left),
    .io_outs_down(ces_7_0_io_outs_down),
    .io_outs_right(ces_7_0_io_outs_right),
    .io_outs_up(ces_7_0_io_outs_up),
    .io_outs_left(ces_7_0_io_outs_left),
    .io_lsbIns_1(ces_7_0_io_lsbIns_1),
    .io_lsbIns_2(ces_7_0_io_lsbIns_2),
    .io_lsbIns_3(ces_7_0_io_lsbIns_3),
    .io_lsbIns_4(ces_7_0_io_lsbIns_4),
    .io_lsbIns_5(ces_7_0_io_lsbIns_5),
    .io_lsbIns_6(ces_7_0_io_lsbIns_6),
    .io_lsbIns_7(ces_7_0_io_lsbIns_7),
    .io_lsbOuts_0(ces_7_0_io_lsbOuts_0),
    .io_lsbOuts_1(ces_7_0_io_lsbOuts_1),
    .io_lsbOuts_2(ces_7_0_io_lsbOuts_2),
    .io_lsbOuts_3(ces_7_0_io_lsbOuts_3),
    .io_lsbOuts_4(ces_7_0_io_lsbOuts_4),
    .io_lsbOuts_5(ces_7_0_io_lsbOuts_5),
    .io_lsbOuts_6(ces_7_0_io_lsbOuts_6),
    .io_lsbOuts_7(ces_7_0_io_lsbOuts_7)
  );
  Element ces_7_1 (
    .clock(ces_7_1_clock),
    .io_clockOutRight(ces_7_1_io_clockOutRight),
    .io_ins_down(ces_7_1_io_ins_down),
    .io_ins_right(ces_7_1_io_ins_right),
    .io_ins_up(ces_7_1_io_ins_up),
    .io_ins_left(ces_7_1_io_ins_left),
    .io_outs_down(ces_7_1_io_outs_down),
    .io_outs_right(ces_7_1_io_outs_right),
    .io_outs_up(ces_7_1_io_outs_up),
    .io_outs_left(ces_7_1_io_outs_left),
    .io_lsbIns_1(ces_7_1_io_lsbIns_1),
    .io_lsbIns_2(ces_7_1_io_lsbIns_2),
    .io_lsbIns_3(ces_7_1_io_lsbIns_3),
    .io_lsbIns_4(ces_7_1_io_lsbIns_4),
    .io_lsbIns_5(ces_7_1_io_lsbIns_5),
    .io_lsbIns_6(ces_7_1_io_lsbIns_6),
    .io_lsbIns_7(ces_7_1_io_lsbIns_7),
    .io_lsbOuts_0(ces_7_1_io_lsbOuts_0),
    .io_lsbOuts_1(ces_7_1_io_lsbOuts_1),
    .io_lsbOuts_2(ces_7_1_io_lsbOuts_2),
    .io_lsbOuts_3(ces_7_1_io_lsbOuts_3),
    .io_lsbOuts_4(ces_7_1_io_lsbOuts_4),
    .io_lsbOuts_5(ces_7_1_io_lsbOuts_5),
    .io_lsbOuts_6(ces_7_1_io_lsbOuts_6),
    .io_lsbOuts_7(ces_7_1_io_lsbOuts_7)
  );
  Element ces_7_2 (
    .clock(ces_7_2_clock),
    .io_clockOutRight(ces_7_2_io_clockOutRight),
    .io_ins_down(ces_7_2_io_ins_down),
    .io_ins_right(ces_7_2_io_ins_right),
    .io_ins_up(ces_7_2_io_ins_up),
    .io_ins_left(ces_7_2_io_ins_left),
    .io_outs_down(ces_7_2_io_outs_down),
    .io_outs_right(ces_7_2_io_outs_right),
    .io_outs_up(ces_7_2_io_outs_up),
    .io_outs_left(ces_7_2_io_outs_left),
    .io_lsbIns_1(ces_7_2_io_lsbIns_1),
    .io_lsbIns_2(ces_7_2_io_lsbIns_2),
    .io_lsbIns_3(ces_7_2_io_lsbIns_3),
    .io_lsbIns_4(ces_7_2_io_lsbIns_4),
    .io_lsbIns_5(ces_7_2_io_lsbIns_5),
    .io_lsbIns_6(ces_7_2_io_lsbIns_6),
    .io_lsbIns_7(ces_7_2_io_lsbIns_7),
    .io_lsbOuts_0(ces_7_2_io_lsbOuts_0),
    .io_lsbOuts_1(ces_7_2_io_lsbOuts_1),
    .io_lsbOuts_2(ces_7_2_io_lsbOuts_2),
    .io_lsbOuts_3(ces_7_2_io_lsbOuts_3),
    .io_lsbOuts_4(ces_7_2_io_lsbOuts_4),
    .io_lsbOuts_5(ces_7_2_io_lsbOuts_5),
    .io_lsbOuts_6(ces_7_2_io_lsbOuts_6),
    .io_lsbOuts_7(ces_7_2_io_lsbOuts_7)
  );
  Element ces_7_3 (
    .clock(ces_7_3_clock),
    .io_clockOutRight(ces_7_3_io_clockOutRight),
    .io_ins_down(ces_7_3_io_ins_down),
    .io_ins_right(ces_7_3_io_ins_right),
    .io_ins_up(ces_7_3_io_ins_up),
    .io_ins_left(ces_7_3_io_ins_left),
    .io_outs_down(ces_7_3_io_outs_down),
    .io_outs_right(ces_7_3_io_outs_right),
    .io_outs_up(ces_7_3_io_outs_up),
    .io_outs_left(ces_7_3_io_outs_left),
    .io_lsbIns_1(ces_7_3_io_lsbIns_1),
    .io_lsbIns_2(ces_7_3_io_lsbIns_2),
    .io_lsbIns_3(ces_7_3_io_lsbIns_3),
    .io_lsbIns_4(ces_7_3_io_lsbIns_4),
    .io_lsbIns_5(ces_7_3_io_lsbIns_5),
    .io_lsbIns_6(ces_7_3_io_lsbIns_6),
    .io_lsbIns_7(ces_7_3_io_lsbIns_7),
    .io_lsbOuts_0(ces_7_3_io_lsbOuts_0),
    .io_lsbOuts_1(ces_7_3_io_lsbOuts_1),
    .io_lsbOuts_2(ces_7_3_io_lsbOuts_2),
    .io_lsbOuts_3(ces_7_3_io_lsbOuts_3),
    .io_lsbOuts_4(ces_7_3_io_lsbOuts_4),
    .io_lsbOuts_5(ces_7_3_io_lsbOuts_5),
    .io_lsbOuts_6(ces_7_3_io_lsbOuts_6),
    .io_lsbOuts_7(ces_7_3_io_lsbOuts_7)
  );
  Element ces_7_4 (
    .clock(ces_7_4_clock),
    .io_clockOutRight(ces_7_4_io_clockOutRight),
    .io_ins_down(ces_7_4_io_ins_down),
    .io_ins_right(ces_7_4_io_ins_right),
    .io_ins_up(ces_7_4_io_ins_up),
    .io_ins_left(ces_7_4_io_ins_left),
    .io_outs_down(ces_7_4_io_outs_down),
    .io_outs_right(ces_7_4_io_outs_right),
    .io_outs_up(ces_7_4_io_outs_up),
    .io_outs_left(ces_7_4_io_outs_left),
    .io_lsbIns_1(ces_7_4_io_lsbIns_1),
    .io_lsbIns_2(ces_7_4_io_lsbIns_2),
    .io_lsbIns_3(ces_7_4_io_lsbIns_3),
    .io_lsbIns_4(ces_7_4_io_lsbIns_4),
    .io_lsbIns_5(ces_7_4_io_lsbIns_5),
    .io_lsbIns_6(ces_7_4_io_lsbIns_6),
    .io_lsbIns_7(ces_7_4_io_lsbIns_7),
    .io_lsbOuts_0(ces_7_4_io_lsbOuts_0),
    .io_lsbOuts_1(ces_7_4_io_lsbOuts_1),
    .io_lsbOuts_2(ces_7_4_io_lsbOuts_2),
    .io_lsbOuts_3(ces_7_4_io_lsbOuts_3),
    .io_lsbOuts_4(ces_7_4_io_lsbOuts_4),
    .io_lsbOuts_5(ces_7_4_io_lsbOuts_5),
    .io_lsbOuts_6(ces_7_4_io_lsbOuts_6),
    .io_lsbOuts_7(ces_7_4_io_lsbOuts_7)
  );
  Element ces_7_5 (
    .clock(ces_7_5_clock),
    .io_clockOutRight(ces_7_5_io_clockOutRight),
    .io_ins_down(ces_7_5_io_ins_down),
    .io_ins_right(ces_7_5_io_ins_right),
    .io_ins_up(ces_7_5_io_ins_up),
    .io_ins_left(ces_7_5_io_ins_left),
    .io_outs_down(ces_7_5_io_outs_down),
    .io_outs_right(ces_7_5_io_outs_right),
    .io_outs_up(ces_7_5_io_outs_up),
    .io_outs_left(ces_7_5_io_outs_left),
    .io_lsbIns_1(ces_7_5_io_lsbIns_1),
    .io_lsbIns_2(ces_7_5_io_lsbIns_2),
    .io_lsbIns_3(ces_7_5_io_lsbIns_3),
    .io_lsbIns_4(ces_7_5_io_lsbIns_4),
    .io_lsbIns_5(ces_7_5_io_lsbIns_5),
    .io_lsbIns_6(ces_7_5_io_lsbIns_6),
    .io_lsbIns_7(ces_7_5_io_lsbIns_7),
    .io_lsbOuts_0(ces_7_5_io_lsbOuts_0),
    .io_lsbOuts_1(ces_7_5_io_lsbOuts_1),
    .io_lsbOuts_2(ces_7_5_io_lsbOuts_2),
    .io_lsbOuts_3(ces_7_5_io_lsbOuts_3),
    .io_lsbOuts_4(ces_7_5_io_lsbOuts_4),
    .io_lsbOuts_5(ces_7_5_io_lsbOuts_5),
    .io_lsbOuts_6(ces_7_5_io_lsbOuts_6),
    .io_lsbOuts_7(ces_7_5_io_lsbOuts_7)
  );
  Element ces_7_6 (
    .clock(ces_7_6_clock),
    .io_clockOutRight(ces_7_6_io_clockOutRight),
    .io_ins_down(ces_7_6_io_ins_down),
    .io_ins_right(ces_7_6_io_ins_right),
    .io_ins_up(ces_7_6_io_ins_up),
    .io_ins_left(ces_7_6_io_ins_left),
    .io_outs_down(ces_7_6_io_outs_down),
    .io_outs_right(ces_7_6_io_outs_right),
    .io_outs_up(ces_7_6_io_outs_up),
    .io_outs_left(ces_7_6_io_outs_left),
    .io_lsbIns_1(ces_7_6_io_lsbIns_1),
    .io_lsbIns_2(ces_7_6_io_lsbIns_2),
    .io_lsbIns_3(ces_7_6_io_lsbIns_3),
    .io_lsbIns_4(ces_7_6_io_lsbIns_4),
    .io_lsbIns_5(ces_7_6_io_lsbIns_5),
    .io_lsbIns_6(ces_7_6_io_lsbIns_6),
    .io_lsbIns_7(ces_7_6_io_lsbIns_7),
    .io_lsbOuts_0(ces_7_6_io_lsbOuts_0),
    .io_lsbOuts_1(ces_7_6_io_lsbOuts_1),
    .io_lsbOuts_2(ces_7_6_io_lsbOuts_2),
    .io_lsbOuts_3(ces_7_6_io_lsbOuts_3),
    .io_lsbOuts_4(ces_7_6_io_lsbOuts_4),
    .io_lsbOuts_5(ces_7_6_io_lsbOuts_5),
    .io_lsbOuts_6(ces_7_6_io_lsbOuts_6),
    .io_lsbOuts_7(ces_7_6_io_lsbOuts_7)
  );
  Element ces_7_7 (
    .clock(ces_7_7_clock),
    .io_clockOutRight(ces_7_7_io_clockOutRight),
    .io_ins_down(ces_7_7_io_ins_down),
    .io_ins_right(ces_7_7_io_ins_right),
    .io_ins_up(ces_7_7_io_ins_up),
    .io_ins_left(ces_7_7_io_ins_left),
    .io_outs_down(ces_7_7_io_outs_down),
    .io_outs_right(ces_7_7_io_outs_right),
    .io_outs_up(ces_7_7_io_outs_up),
    .io_outs_left(ces_7_7_io_outs_left),
    .io_lsbIns_1(ces_7_7_io_lsbIns_1),
    .io_lsbIns_2(ces_7_7_io_lsbIns_2),
    .io_lsbIns_3(ces_7_7_io_lsbIns_3),
    .io_lsbIns_4(ces_7_7_io_lsbIns_4),
    .io_lsbIns_5(ces_7_7_io_lsbIns_5),
    .io_lsbIns_6(ces_7_7_io_lsbIns_6),
    .io_lsbIns_7(ces_7_7_io_lsbIns_7),
    .io_lsbOuts_0(ces_7_7_io_lsbOuts_0),
    .io_lsbOuts_1(ces_7_7_io_lsbOuts_1),
    .io_lsbOuts_2(ces_7_7_io_lsbOuts_2),
    .io_lsbOuts_3(ces_7_7_io_lsbOuts_3),
    .io_lsbOuts_4(ces_7_7_io_lsbOuts_4),
    .io_lsbOuts_5(ces_7_7_io_lsbOuts_5),
    .io_lsbOuts_6(ces_7_7_io_lsbOuts_6),
    .io_lsbOuts_7(ces_7_7_io_lsbOuts_7)
  );
  assign io_outs_down_0 = ces_0_0_io_outs_down;
  assign io_outs_down_1 = ces_0_1_io_outs_down;
  assign io_outs_down_2 = ces_0_2_io_outs_down;
  assign io_outs_down_3 = ces_0_3_io_outs_down;
  assign io_outs_down_4 = ces_0_4_io_outs_down;
  assign io_outs_down_5 = ces_0_5_io_outs_down;
  assign io_outs_down_6 = ces_0_6_io_outs_down;
  assign io_outs_down_7 = ces_0_7_io_outs_down;
  assign io_outs_up_0 = ces_7_0_io_outs_up;
  assign io_outs_up_1 = ces_7_1_io_outs_up;
  assign io_outs_up_2 = ces_7_2_io_outs_up;
  assign io_outs_up_3 = ces_7_3_io_outs_up;
  assign io_outs_up_4 = ces_7_4_io_outs_up;
  assign io_outs_up_5 = ces_7_5_io_outs_up;
  assign io_outs_up_6 = ces_7_6_io_outs_up;
  assign io_outs_up_7 = ces_7_7_io_outs_up;
  assign io_outs_right_0 = ces_0_7_io_outs_right;
  assign io_outs_right_1 = ces_1_7_io_outs_right;
  assign io_outs_right_2 = ces_2_7_io_outs_right;
  assign io_outs_right_3 = ces_3_7_io_outs_right;
  assign io_outs_right_4 = ces_4_7_io_outs_right;
  assign io_outs_right_5 = ces_5_7_io_outs_right;
  assign io_outs_right_6 = ces_6_7_io_outs_right;
  assign io_outs_right_7 = ces_7_7_io_outs_right;
  assign io_outs_left_0 = ces_0_0_io_outs_left;
  assign io_outs_left_1 = ces_1_0_io_outs_left;
  assign io_outs_left_2 = ces_2_0_io_outs_left;
  assign io_outs_left_3 = ces_3_0_io_outs_left;
  assign io_outs_left_4 = ces_4_0_io_outs_left;
  assign io_outs_left_5 = ces_5_0_io_outs_left;
  assign io_outs_left_6 = ces_6_0_io_outs_left;
  assign io_outs_left_7 = ces_7_0_io_outs_left;
  assign io_lsbs_0 = REG_0;
  assign io_lsbs_1 = REG_1;
  assign io_lsbs_2 = REG_2;
  assign io_lsbs_3 = REG_3;
  assign io_lsbs_4 = REG_4;
  assign io_lsbs_5 = REG_5;
  assign io_lsbs_6 = REG_6;
  assign io_lsbs_7 = REG_7;
  assign io_lsbs_8 = REG_8;
  assign io_lsbs_9 = REG_9;
  assign io_lsbs_10 = REG_10;
  assign io_lsbs_11 = REG_11;
  assign io_lsbs_12 = REG_12;
  assign io_lsbs_13 = REG_13;
  assign io_lsbs_14 = REG_14;
  assign io_lsbs_15 = REG_15;
  assign io_lsbs_16 = REG_16;
  assign io_lsbs_17 = REG_17;
  assign io_lsbs_18 = REG_18;
  assign io_lsbs_19 = REG_19;
  assign io_lsbs_20 = REG_20;
  assign io_lsbs_21 = REG_21;
  assign io_lsbs_22 = REG_22;
  assign io_lsbs_23 = REG_23;
  assign io_lsbs_24 = REG_24;
  assign io_lsbs_25 = REG_25;
  assign io_lsbs_26 = REG_26;
  assign io_lsbs_27 = REG_27;
  assign io_lsbs_28 = REG_28;
  assign io_lsbs_29 = REG_29;
  assign io_lsbs_30 = REG_30;
  assign io_lsbs_31 = REG_31;
  assign io_lsbs_32 = REG_32;
  assign io_lsbs_33 = REG_33;
  assign io_lsbs_34 = REG_34;
  assign io_lsbs_35 = REG_35;
  assign io_lsbs_36 = REG_36;
  assign io_lsbs_37 = REG_37;
  assign io_lsbs_38 = REG_38;
  assign io_lsbs_39 = REG_39;
  assign io_lsbs_40 = REG_40;
  assign io_lsbs_41 = REG_41;
  assign io_lsbs_42 = REG_42;
  assign io_lsbs_43 = REG_43;
  assign io_lsbs_44 = REG_44;
  assign io_lsbs_45 = REG_45;
  assign io_lsbs_46 = REG_46;
  assign io_lsbs_47 = REG_47;
  assign io_lsbs_48 = REG_48;
  assign io_lsbs_49 = REG_49;
  assign io_lsbs_50 = REG_50;
  assign io_lsbs_51 = REG_51;
  assign io_lsbs_52 = REG_52;
  assign io_lsbs_53 = REG_53;
  assign io_lsbs_54 = REG_54;
  assign io_lsbs_55 = REG_55;
  assign io_lsbs_56 = REG_56;
  assign io_lsbs_57 = REG_57;
  assign io_lsbs_58 = REG_58;
  assign io_lsbs_59 = REG_59;
  assign io_lsbs_60 = REG_60;
  assign io_lsbs_61 = REG_61;
  assign io_lsbs_62 = REG_62;
  assign io_lsbs_63 = REG_63;
  assign ces_0_0_clock = clock;
  assign ces_0_0_io_ins_down = ces_1_0_io_outs_down;
  assign ces_0_0_io_ins_right = io_ins_right_0;
  assign ces_0_0_io_ins_up = io_ins_up_0;
  assign ces_0_0_io_ins_left = ces_0_1_io_outs_left;
  assign ces_0_0_io_lsbIns_1 = 1'h0;
  assign ces_0_0_io_lsbIns_2 = 1'h0;
  assign ces_0_0_io_lsbIns_3 = 1'h0;
  assign ces_0_0_io_lsbIns_4 = 1'h0;
  assign ces_0_0_io_lsbIns_5 = 1'h0;
  assign ces_0_0_io_lsbIns_6 = 1'h0;
  assign ces_0_0_io_lsbIns_7 = 1'h0;
  assign ces_0_1_clock = ces_0_0_io_clockOutRight;
  assign ces_0_1_io_ins_down = ces_1_1_io_outs_down;
  assign ces_0_1_io_ins_right = ces_0_0_io_outs_right;
  assign ces_0_1_io_ins_up = io_ins_up_1;
  assign ces_0_1_io_ins_left = ces_0_2_io_outs_left;
  assign ces_0_1_io_lsbIns_1 = ces_0_0_io_lsbOuts_1;
  assign ces_0_1_io_lsbIns_2 = ces_0_0_io_lsbOuts_2;
  assign ces_0_1_io_lsbIns_3 = ces_0_0_io_lsbOuts_3;
  assign ces_0_1_io_lsbIns_4 = ces_0_0_io_lsbOuts_4;
  assign ces_0_1_io_lsbIns_5 = ces_0_0_io_lsbOuts_5;
  assign ces_0_1_io_lsbIns_6 = ces_0_0_io_lsbOuts_6;
  assign ces_0_1_io_lsbIns_7 = ces_0_0_io_lsbOuts_7;
  assign ces_0_2_clock = ces_0_1_io_clockOutRight;
  assign ces_0_2_io_ins_down = ces_1_2_io_outs_down;
  assign ces_0_2_io_ins_right = ces_0_1_io_outs_right;
  assign ces_0_2_io_ins_up = io_ins_up_2;
  assign ces_0_2_io_ins_left = ces_0_3_io_outs_left;
  assign ces_0_2_io_lsbIns_1 = ces_0_1_io_lsbOuts_1;
  assign ces_0_2_io_lsbIns_2 = ces_0_1_io_lsbOuts_2;
  assign ces_0_2_io_lsbIns_3 = ces_0_1_io_lsbOuts_3;
  assign ces_0_2_io_lsbIns_4 = ces_0_1_io_lsbOuts_4;
  assign ces_0_2_io_lsbIns_5 = ces_0_1_io_lsbOuts_5;
  assign ces_0_2_io_lsbIns_6 = ces_0_1_io_lsbOuts_6;
  assign ces_0_2_io_lsbIns_7 = ces_0_1_io_lsbOuts_7;
  assign ces_0_3_clock = ces_0_2_io_clockOutRight;
  assign ces_0_3_io_ins_down = ces_1_3_io_outs_down;
  assign ces_0_3_io_ins_right = ces_0_2_io_outs_right;
  assign ces_0_3_io_ins_up = io_ins_up_3;
  assign ces_0_3_io_ins_left = ces_0_4_io_outs_left;
  assign ces_0_3_io_lsbIns_1 = ces_0_2_io_lsbOuts_1;
  assign ces_0_3_io_lsbIns_2 = ces_0_2_io_lsbOuts_2;
  assign ces_0_3_io_lsbIns_3 = ces_0_2_io_lsbOuts_3;
  assign ces_0_3_io_lsbIns_4 = ces_0_2_io_lsbOuts_4;
  assign ces_0_3_io_lsbIns_5 = ces_0_2_io_lsbOuts_5;
  assign ces_0_3_io_lsbIns_6 = ces_0_2_io_lsbOuts_6;
  assign ces_0_3_io_lsbIns_7 = ces_0_2_io_lsbOuts_7;
  assign ces_0_4_clock = ces_0_3_io_clockOutRight;
  assign ces_0_4_io_ins_down = ces_1_4_io_outs_down;
  assign ces_0_4_io_ins_right = ces_0_3_io_outs_right;
  assign ces_0_4_io_ins_up = io_ins_up_4;
  assign ces_0_4_io_ins_left = ces_0_5_io_outs_left;
  assign ces_0_4_io_lsbIns_1 = ces_0_3_io_lsbOuts_1;
  assign ces_0_4_io_lsbIns_2 = ces_0_3_io_lsbOuts_2;
  assign ces_0_4_io_lsbIns_3 = ces_0_3_io_lsbOuts_3;
  assign ces_0_4_io_lsbIns_4 = ces_0_3_io_lsbOuts_4;
  assign ces_0_4_io_lsbIns_5 = ces_0_3_io_lsbOuts_5;
  assign ces_0_4_io_lsbIns_6 = ces_0_3_io_lsbOuts_6;
  assign ces_0_4_io_lsbIns_7 = ces_0_3_io_lsbOuts_7;
  assign ces_0_5_clock = ces_0_4_io_clockOutRight;
  assign ces_0_5_io_ins_down = ces_1_5_io_outs_down;
  assign ces_0_5_io_ins_right = ces_0_4_io_outs_right;
  assign ces_0_5_io_ins_up = io_ins_up_5;
  assign ces_0_5_io_ins_left = ces_0_6_io_outs_left;
  assign ces_0_5_io_lsbIns_1 = ces_0_4_io_lsbOuts_1;
  assign ces_0_5_io_lsbIns_2 = ces_0_4_io_lsbOuts_2;
  assign ces_0_5_io_lsbIns_3 = ces_0_4_io_lsbOuts_3;
  assign ces_0_5_io_lsbIns_4 = ces_0_4_io_lsbOuts_4;
  assign ces_0_5_io_lsbIns_5 = ces_0_4_io_lsbOuts_5;
  assign ces_0_5_io_lsbIns_6 = ces_0_4_io_lsbOuts_6;
  assign ces_0_5_io_lsbIns_7 = ces_0_4_io_lsbOuts_7;
  assign ces_0_6_clock = ces_0_5_io_clockOutRight;
  assign ces_0_6_io_ins_down = ces_1_6_io_outs_down;
  assign ces_0_6_io_ins_right = ces_0_5_io_outs_right;
  assign ces_0_6_io_ins_up = io_ins_up_6;
  assign ces_0_6_io_ins_left = ces_0_7_io_outs_left;
  assign ces_0_6_io_lsbIns_1 = ces_0_5_io_lsbOuts_1;
  assign ces_0_6_io_lsbIns_2 = ces_0_5_io_lsbOuts_2;
  assign ces_0_6_io_lsbIns_3 = ces_0_5_io_lsbOuts_3;
  assign ces_0_6_io_lsbIns_4 = ces_0_5_io_lsbOuts_4;
  assign ces_0_6_io_lsbIns_5 = ces_0_5_io_lsbOuts_5;
  assign ces_0_6_io_lsbIns_6 = ces_0_5_io_lsbOuts_6;
  assign ces_0_6_io_lsbIns_7 = ces_0_5_io_lsbOuts_7;
  assign ces_0_7_clock = ces_0_6_io_clockOutRight;
  assign ces_0_7_io_ins_down = ces_1_7_io_outs_down;
  assign ces_0_7_io_ins_right = ces_0_6_io_outs_right;
  assign ces_0_7_io_ins_up = io_ins_up_7;
  assign ces_0_7_io_ins_left = io_ins_left_0;
  assign ces_0_7_io_lsbIns_1 = ces_0_6_io_lsbOuts_1;
  assign ces_0_7_io_lsbIns_2 = ces_0_6_io_lsbOuts_2;
  assign ces_0_7_io_lsbIns_3 = ces_0_6_io_lsbOuts_3;
  assign ces_0_7_io_lsbIns_4 = ces_0_6_io_lsbOuts_4;
  assign ces_0_7_io_lsbIns_5 = ces_0_6_io_lsbOuts_5;
  assign ces_0_7_io_lsbIns_6 = ces_0_6_io_lsbOuts_6;
  assign ces_0_7_io_lsbIns_7 = ces_0_6_io_lsbOuts_7;
  assign ces_1_0_clock = clock;
  assign ces_1_0_io_ins_down = ces_2_0_io_outs_down;
  assign ces_1_0_io_ins_right = io_ins_right_1;
  assign ces_1_0_io_ins_up = ces_0_0_io_outs_up;
  assign ces_1_0_io_ins_left = ces_1_1_io_outs_left;
  assign ces_1_0_io_lsbIns_1 = 1'h0;
  assign ces_1_0_io_lsbIns_2 = 1'h0;
  assign ces_1_0_io_lsbIns_3 = 1'h0;
  assign ces_1_0_io_lsbIns_4 = 1'h0;
  assign ces_1_0_io_lsbIns_5 = 1'h0;
  assign ces_1_0_io_lsbIns_6 = 1'h0;
  assign ces_1_0_io_lsbIns_7 = 1'h0;
  assign ces_1_1_clock = ces_1_0_io_clockOutRight;
  assign ces_1_1_io_ins_down = ces_2_1_io_outs_down;
  assign ces_1_1_io_ins_right = ces_1_0_io_outs_right;
  assign ces_1_1_io_ins_up = ces_0_1_io_outs_up;
  assign ces_1_1_io_ins_left = ces_1_2_io_outs_left;
  assign ces_1_1_io_lsbIns_1 = ces_1_0_io_lsbOuts_1;
  assign ces_1_1_io_lsbIns_2 = ces_1_0_io_lsbOuts_2;
  assign ces_1_1_io_lsbIns_3 = ces_1_0_io_lsbOuts_3;
  assign ces_1_1_io_lsbIns_4 = ces_1_0_io_lsbOuts_4;
  assign ces_1_1_io_lsbIns_5 = ces_1_0_io_lsbOuts_5;
  assign ces_1_1_io_lsbIns_6 = ces_1_0_io_lsbOuts_6;
  assign ces_1_1_io_lsbIns_7 = ces_1_0_io_lsbOuts_7;
  assign ces_1_2_clock = ces_1_1_io_clockOutRight;
  assign ces_1_2_io_ins_down = ces_2_2_io_outs_down;
  assign ces_1_2_io_ins_right = ces_1_1_io_outs_right;
  assign ces_1_2_io_ins_up = ces_0_2_io_outs_up;
  assign ces_1_2_io_ins_left = ces_1_3_io_outs_left;
  assign ces_1_2_io_lsbIns_1 = ces_1_1_io_lsbOuts_1;
  assign ces_1_2_io_lsbIns_2 = ces_1_1_io_lsbOuts_2;
  assign ces_1_2_io_lsbIns_3 = ces_1_1_io_lsbOuts_3;
  assign ces_1_2_io_lsbIns_4 = ces_1_1_io_lsbOuts_4;
  assign ces_1_2_io_lsbIns_5 = ces_1_1_io_lsbOuts_5;
  assign ces_1_2_io_lsbIns_6 = ces_1_1_io_lsbOuts_6;
  assign ces_1_2_io_lsbIns_7 = ces_1_1_io_lsbOuts_7;
  assign ces_1_3_clock = ces_1_2_io_clockOutRight;
  assign ces_1_3_io_ins_down = ces_2_3_io_outs_down;
  assign ces_1_3_io_ins_right = ces_1_2_io_outs_right;
  assign ces_1_3_io_ins_up = ces_0_3_io_outs_up;
  assign ces_1_3_io_ins_left = ces_1_4_io_outs_left;
  assign ces_1_3_io_lsbIns_1 = ces_1_2_io_lsbOuts_1;
  assign ces_1_3_io_lsbIns_2 = ces_1_2_io_lsbOuts_2;
  assign ces_1_3_io_lsbIns_3 = ces_1_2_io_lsbOuts_3;
  assign ces_1_3_io_lsbIns_4 = ces_1_2_io_lsbOuts_4;
  assign ces_1_3_io_lsbIns_5 = ces_1_2_io_lsbOuts_5;
  assign ces_1_3_io_lsbIns_6 = ces_1_2_io_lsbOuts_6;
  assign ces_1_3_io_lsbIns_7 = ces_1_2_io_lsbOuts_7;
  assign ces_1_4_clock = ces_1_3_io_clockOutRight;
  assign ces_1_4_io_ins_down = ces_2_4_io_outs_down;
  assign ces_1_4_io_ins_right = ces_1_3_io_outs_right;
  assign ces_1_4_io_ins_up = ces_0_4_io_outs_up;
  assign ces_1_4_io_ins_left = ces_1_5_io_outs_left;
  assign ces_1_4_io_lsbIns_1 = ces_1_3_io_lsbOuts_1;
  assign ces_1_4_io_lsbIns_2 = ces_1_3_io_lsbOuts_2;
  assign ces_1_4_io_lsbIns_3 = ces_1_3_io_lsbOuts_3;
  assign ces_1_4_io_lsbIns_4 = ces_1_3_io_lsbOuts_4;
  assign ces_1_4_io_lsbIns_5 = ces_1_3_io_lsbOuts_5;
  assign ces_1_4_io_lsbIns_6 = ces_1_3_io_lsbOuts_6;
  assign ces_1_4_io_lsbIns_7 = ces_1_3_io_lsbOuts_7;
  assign ces_1_5_clock = ces_1_4_io_clockOutRight;
  assign ces_1_5_io_ins_down = ces_2_5_io_outs_down;
  assign ces_1_5_io_ins_right = ces_1_4_io_outs_right;
  assign ces_1_5_io_ins_up = ces_0_5_io_outs_up;
  assign ces_1_5_io_ins_left = ces_1_6_io_outs_left;
  assign ces_1_5_io_lsbIns_1 = ces_1_4_io_lsbOuts_1;
  assign ces_1_5_io_lsbIns_2 = ces_1_4_io_lsbOuts_2;
  assign ces_1_5_io_lsbIns_3 = ces_1_4_io_lsbOuts_3;
  assign ces_1_5_io_lsbIns_4 = ces_1_4_io_lsbOuts_4;
  assign ces_1_5_io_lsbIns_5 = ces_1_4_io_lsbOuts_5;
  assign ces_1_5_io_lsbIns_6 = ces_1_4_io_lsbOuts_6;
  assign ces_1_5_io_lsbIns_7 = ces_1_4_io_lsbOuts_7;
  assign ces_1_6_clock = ces_1_5_io_clockOutRight;
  assign ces_1_6_io_ins_down = ces_2_6_io_outs_down;
  assign ces_1_6_io_ins_right = ces_1_5_io_outs_right;
  assign ces_1_6_io_ins_up = ces_0_6_io_outs_up;
  assign ces_1_6_io_ins_left = ces_1_7_io_outs_left;
  assign ces_1_6_io_lsbIns_1 = ces_1_5_io_lsbOuts_1;
  assign ces_1_6_io_lsbIns_2 = ces_1_5_io_lsbOuts_2;
  assign ces_1_6_io_lsbIns_3 = ces_1_5_io_lsbOuts_3;
  assign ces_1_6_io_lsbIns_4 = ces_1_5_io_lsbOuts_4;
  assign ces_1_6_io_lsbIns_5 = ces_1_5_io_lsbOuts_5;
  assign ces_1_6_io_lsbIns_6 = ces_1_5_io_lsbOuts_6;
  assign ces_1_6_io_lsbIns_7 = ces_1_5_io_lsbOuts_7;
  assign ces_1_7_clock = ces_1_6_io_clockOutRight;
  assign ces_1_7_io_ins_down = ces_2_7_io_outs_down;
  assign ces_1_7_io_ins_right = ces_1_6_io_outs_right;
  assign ces_1_7_io_ins_up = ces_0_7_io_outs_up;
  assign ces_1_7_io_ins_left = io_ins_left_1;
  assign ces_1_7_io_lsbIns_1 = ces_1_6_io_lsbOuts_1;
  assign ces_1_7_io_lsbIns_2 = ces_1_6_io_lsbOuts_2;
  assign ces_1_7_io_lsbIns_3 = ces_1_6_io_lsbOuts_3;
  assign ces_1_7_io_lsbIns_4 = ces_1_6_io_lsbOuts_4;
  assign ces_1_7_io_lsbIns_5 = ces_1_6_io_lsbOuts_5;
  assign ces_1_7_io_lsbIns_6 = ces_1_6_io_lsbOuts_6;
  assign ces_1_7_io_lsbIns_7 = ces_1_6_io_lsbOuts_7;
  assign ces_2_0_clock = clock;
  assign ces_2_0_io_ins_down = ces_3_0_io_outs_down;
  assign ces_2_0_io_ins_right = io_ins_right_2;
  assign ces_2_0_io_ins_up = ces_1_0_io_outs_up;
  assign ces_2_0_io_ins_left = ces_2_1_io_outs_left;
  assign ces_2_0_io_lsbIns_1 = 1'h0;
  assign ces_2_0_io_lsbIns_2 = 1'h0;
  assign ces_2_0_io_lsbIns_3 = 1'h0;
  assign ces_2_0_io_lsbIns_4 = 1'h0;
  assign ces_2_0_io_lsbIns_5 = 1'h0;
  assign ces_2_0_io_lsbIns_6 = 1'h0;
  assign ces_2_0_io_lsbIns_7 = 1'h0;
  assign ces_2_1_clock = ces_2_0_io_clockOutRight;
  assign ces_2_1_io_ins_down = ces_3_1_io_outs_down;
  assign ces_2_1_io_ins_right = ces_2_0_io_outs_right;
  assign ces_2_1_io_ins_up = ces_1_1_io_outs_up;
  assign ces_2_1_io_ins_left = ces_2_2_io_outs_left;
  assign ces_2_1_io_lsbIns_1 = ces_2_0_io_lsbOuts_1;
  assign ces_2_1_io_lsbIns_2 = ces_2_0_io_lsbOuts_2;
  assign ces_2_1_io_lsbIns_3 = ces_2_0_io_lsbOuts_3;
  assign ces_2_1_io_lsbIns_4 = ces_2_0_io_lsbOuts_4;
  assign ces_2_1_io_lsbIns_5 = ces_2_0_io_lsbOuts_5;
  assign ces_2_1_io_lsbIns_6 = ces_2_0_io_lsbOuts_6;
  assign ces_2_1_io_lsbIns_7 = ces_2_0_io_lsbOuts_7;
  assign ces_2_2_clock = ces_2_1_io_clockOutRight;
  assign ces_2_2_io_ins_down = ces_3_2_io_outs_down;
  assign ces_2_2_io_ins_right = ces_2_1_io_outs_right;
  assign ces_2_2_io_ins_up = ces_1_2_io_outs_up;
  assign ces_2_2_io_ins_left = ces_2_3_io_outs_left;
  assign ces_2_2_io_lsbIns_1 = ces_2_1_io_lsbOuts_1;
  assign ces_2_2_io_lsbIns_2 = ces_2_1_io_lsbOuts_2;
  assign ces_2_2_io_lsbIns_3 = ces_2_1_io_lsbOuts_3;
  assign ces_2_2_io_lsbIns_4 = ces_2_1_io_lsbOuts_4;
  assign ces_2_2_io_lsbIns_5 = ces_2_1_io_lsbOuts_5;
  assign ces_2_2_io_lsbIns_6 = ces_2_1_io_lsbOuts_6;
  assign ces_2_2_io_lsbIns_7 = ces_2_1_io_lsbOuts_7;
  assign ces_2_3_clock = ces_2_2_io_clockOutRight;
  assign ces_2_3_io_ins_down = ces_3_3_io_outs_down;
  assign ces_2_3_io_ins_right = ces_2_2_io_outs_right;
  assign ces_2_3_io_ins_up = ces_1_3_io_outs_up;
  assign ces_2_3_io_ins_left = ces_2_4_io_outs_left;
  assign ces_2_3_io_lsbIns_1 = ces_2_2_io_lsbOuts_1;
  assign ces_2_3_io_lsbIns_2 = ces_2_2_io_lsbOuts_2;
  assign ces_2_3_io_lsbIns_3 = ces_2_2_io_lsbOuts_3;
  assign ces_2_3_io_lsbIns_4 = ces_2_2_io_lsbOuts_4;
  assign ces_2_3_io_lsbIns_5 = ces_2_2_io_lsbOuts_5;
  assign ces_2_3_io_lsbIns_6 = ces_2_2_io_lsbOuts_6;
  assign ces_2_3_io_lsbIns_7 = ces_2_2_io_lsbOuts_7;
  assign ces_2_4_clock = ces_2_3_io_clockOutRight;
  assign ces_2_4_io_ins_down = ces_3_4_io_outs_down;
  assign ces_2_4_io_ins_right = ces_2_3_io_outs_right;
  assign ces_2_4_io_ins_up = ces_1_4_io_outs_up;
  assign ces_2_4_io_ins_left = ces_2_5_io_outs_left;
  assign ces_2_4_io_lsbIns_1 = ces_2_3_io_lsbOuts_1;
  assign ces_2_4_io_lsbIns_2 = ces_2_3_io_lsbOuts_2;
  assign ces_2_4_io_lsbIns_3 = ces_2_3_io_lsbOuts_3;
  assign ces_2_4_io_lsbIns_4 = ces_2_3_io_lsbOuts_4;
  assign ces_2_4_io_lsbIns_5 = ces_2_3_io_lsbOuts_5;
  assign ces_2_4_io_lsbIns_6 = ces_2_3_io_lsbOuts_6;
  assign ces_2_4_io_lsbIns_7 = ces_2_3_io_lsbOuts_7;
  assign ces_2_5_clock = ces_2_4_io_clockOutRight;
  assign ces_2_5_io_ins_down = ces_3_5_io_outs_down;
  assign ces_2_5_io_ins_right = ces_2_4_io_outs_right;
  assign ces_2_5_io_ins_up = ces_1_5_io_outs_up;
  assign ces_2_5_io_ins_left = ces_2_6_io_outs_left;
  assign ces_2_5_io_lsbIns_1 = ces_2_4_io_lsbOuts_1;
  assign ces_2_5_io_lsbIns_2 = ces_2_4_io_lsbOuts_2;
  assign ces_2_5_io_lsbIns_3 = ces_2_4_io_lsbOuts_3;
  assign ces_2_5_io_lsbIns_4 = ces_2_4_io_lsbOuts_4;
  assign ces_2_5_io_lsbIns_5 = ces_2_4_io_lsbOuts_5;
  assign ces_2_5_io_lsbIns_6 = ces_2_4_io_lsbOuts_6;
  assign ces_2_5_io_lsbIns_7 = ces_2_4_io_lsbOuts_7;
  assign ces_2_6_clock = ces_2_5_io_clockOutRight;
  assign ces_2_6_io_ins_down = ces_3_6_io_outs_down;
  assign ces_2_6_io_ins_right = ces_2_5_io_outs_right;
  assign ces_2_6_io_ins_up = ces_1_6_io_outs_up;
  assign ces_2_6_io_ins_left = ces_2_7_io_outs_left;
  assign ces_2_6_io_lsbIns_1 = ces_2_5_io_lsbOuts_1;
  assign ces_2_6_io_lsbIns_2 = ces_2_5_io_lsbOuts_2;
  assign ces_2_6_io_lsbIns_3 = ces_2_5_io_lsbOuts_3;
  assign ces_2_6_io_lsbIns_4 = ces_2_5_io_lsbOuts_4;
  assign ces_2_6_io_lsbIns_5 = ces_2_5_io_lsbOuts_5;
  assign ces_2_6_io_lsbIns_6 = ces_2_5_io_lsbOuts_6;
  assign ces_2_6_io_lsbIns_7 = ces_2_5_io_lsbOuts_7;
  assign ces_2_7_clock = ces_2_6_io_clockOutRight;
  assign ces_2_7_io_ins_down = ces_3_7_io_outs_down;
  assign ces_2_7_io_ins_right = ces_2_6_io_outs_right;
  assign ces_2_7_io_ins_up = ces_1_7_io_outs_up;
  assign ces_2_7_io_ins_left = io_ins_left_2;
  assign ces_2_7_io_lsbIns_1 = ces_2_6_io_lsbOuts_1;
  assign ces_2_7_io_lsbIns_2 = ces_2_6_io_lsbOuts_2;
  assign ces_2_7_io_lsbIns_3 = ces_2_6_io_lsbOuts_3;
  assign ces_2_7_io_lsbIns_4 = ces_2_6_io_lsbOuts_4;
  assign ces_2_7_io_lsbIns_5 = ces_2_6_io_lsbOuts_5;
  assign ces_2_7_io_lsbIns_6 = ces_2_6_io_lsbOuts_6;
  assign ces_2_7_io_lsbIns_7 = ces_2_6_io_lsbOuts_7;
  assign ces_3_0_clock = clock;
  assign ces_3_0_io_ins_down = ces_4_0_io_outs_down;
  assign ces_3_0_io_ins_right = io_ins_right_3;
  assign ces_3_0_io_ins_up = ces_2_0_io_outs_up;
  assign ces_3_0_io_ins_left = ces_3_1_io_outs_left;
  assign ces_3_0_io_lsbIns_1 = 1'h0;
  assign ces_3_0_io_lsbIns_2 = 1'h0;
  assign ces_3_0_io_lsbIns_3 = 1'h0;
  assign ces_3_0_io_lsbIns_4 = 1'h0;
  assign ces_3_0_io_lsbIns_5 = 1'h0;
  assign ces_3_0_io_lsbIns_6 = 1'h0;
  assign ces_3_0_io_lsbIns_7 = 1'h0;
  assign ces_3_1_clock = ces_3_0_io_clockOutRight;
  assign ces_3_1_io_ins_down = ces_4_1_io_outs_down;
  assign ces_3_1_io_ins_right = ces_3_0_io_outs_right;
  assign ces_3_1_io_ins_up = ces_2_1_io_outs_up;
  assign ces_3_1_io_ins_left = ces_3_2_io_outs_left;
  assign ces_3_1_io_lsbIns_1 = ces_3_0_io_lsbOuts_1;
  assign ces_3_1_io_lsbIns_2 = ces_3_0_io_lsbOuts_2;
  assign ces_3_1_io_lsbIns_3 = ces_3_0_io_lsbOuts_3;
  assign ces_3_1_io_lsbIns_4 = ces_3_0_io_lsbOuts_4;
  assign ces_3_1_io_lsbIns_5 = ces_3_0_io_lsbOuts_5;
  assign ces_3_1_io_lsbIns_6 = ces_3_0_io_lsbOuts_6;
  assign ces_3_1_io_lsbIns_7 = ces_3_0_io_lsbOuts_7;
  assign ces_3_2_clock = ces_3_1_io_clockOutRight;
  assign ces_3_2_io_ins_down = ces_4_2_io_outs_down;
  assign ces_3_2_io_ins_right = ces_3_1_io_outs_right;
  assign ces_3_2_io_ins_up = ces_2_2_io_outs_up;
  assign ces_3_2_io_ins_left = ces_3_3_io_outs_left;
  assign ces_3_2_io_lsbIns_1 = ces_3_1_io_lsbOuts_1;
  assign ces_3_2_io_lsbIns_2 = ces_3_1_io_lsbOuts_2;
  assign ces_3_2_io_lsbIns_3 = ces_3_1_io_lsbOuts_3;
  assign ces_3_2_io_lsbIns_4 = ces_3_1_io_lsbOuts_4;
  assign ces_3_2_io_lsbIns_5 = ces_3_1_io_lsbOuts_5;
  assign ces_3_2_io_lsbIns_6 = ces_3_1_io_lsbOuts_6;
  assign ces_3_2_io_lsbIns_7 = ces_3_1_io_lsbOuts_7;
  assign ces_3_3_clock = ces_3_2_io_clockOutRight;
  assign ces_3_3_io_ins_down = ces_4_3_io_outs_down;
  assign ces_3_3_io_ins_right = ces_3_2_io_outs_right;
  assign ces_3_3_io_ins_up = ces_2_3_io_outs_up;
  assign ces_3_3_io_ins_left = ces_3_4_io_outs_left;
  assign ces_3_3_io_lsbIns_1 = ces_3_2_io_lsbOuts_1;
  assign ces_3_3_io_lsbIns_2 = ces_3_2_io_lsbOuts_2;
  assign ces_3_3_io_lsbIns_3 = ces_3_2_io_lsbOuts_3;
  assign ces_3_3_io_lsbIns_4 = ces_3_2_io_lsbOuts_4;
  assign ces_3_3_io_lsbIns_5 = ces_3_2_io_lsbOuts_5;
  assign ces_3_3_io_lsbIns_6 = ces_3_2_io_lsbOuts_6;
  assign ces_3_3_io_lsbIns_7 = ces_3_2_io_lsbOuts_7;
  assign ces_3_4_clock = ces_3_3_io_clockOutRight;
  assign ces_3_4_io_ins_down = ces_4_4_io_outs_down;
  assign ces_3_4_io_ins_right = ces_3_3_io_outs_right;
  assign ces_3_4_io_ins_up = ces_2_4_io_outs_up;
  assign ces_3_4_io_ins_left = ces_3_5_io_outs_left;
  assign ces_3_4_io_lsbIns_1 = ces_3_3_io_lsbOuts_1;
  assign ces_3_4_io_lsbIns_2 = ces_3_3_io_lsbOuts_2;
  assign ces_3_4_io_lsbIns_3 = ces_3_3_io_lsbOuts_3;
  assign ces_3_4_io_lsbIns_4 = ces_3_3_io_lsbOuts_4;
  assign ces_3_4_io_lsbIns_5 = ces_3_3_io_lsbOuts_5;
  assign ces_3_4_io_lsbIns_6 = ces_3_3_io_lsbOuts_6;
  assign ces_3_4_io_lsbIns_7 = ces_3_3_io_lsbOuts_7;
  assign ces_3_5_clock = ces_3_4_io_clockOutRight;
  assign ces_3_5_io_ins_down = ces_4_5_io_outs_down;
  assign ces_3_5_io_ins_right = ces_3_4_io_outs_right;
  assign ces_3_5_io_ins_up = ces_2_5_io_outs_up;
  assign ces_3_5_io_ins_left = ces_3_6_io_outs_left;
  assign ces_3_5_io_lsbIns_1 = ces_3_4_io_lsbOuts_1;
  assign ces_3_5_io_lsbIns_2 = ces_3_4_io_lsbOuts_2;
  assign ces_3_5_io_lsbIns_3 = ces_3_4_io_lsbOuts_3;
  assign ces_3_5_io_lsbIns_4 = ces_3_4_io_lsbOuts_4;
  assign ces_3_5_io_lsbIns_5 = ces_3_4_io_lsbOuts_5;
  assign ces_3_5_io_lsbIns_6 = ces_3_4_io_lsbOuts_6;
  assign ces_3_5_io_lsbIns_7 = ces_3_4_io_lsbOuts_7;
  assign ces_3_6_clock = ces_3_5_io_clockOutRight;
  assign ces_3_6_io_ins_down = ces_4_6_io_outs_down;
  assign ces_3_6_io_ins_right = ces_3_5_io_outs_right;
  assign ces_3_6_io_ins_up = ces_2_6_io_outs_up;
  assign ces_3_6_io_ins_left = ces_3_7_io_outs_left;
  assign ces_3_6_io_lsbIns_1 = ces_3_5_io_lsbOuts_1;
  assign ces_3_6_io_lsbIns_2 = ces_3_5_io_lsbOuts_2;
  assign ces_3_6_io_lsbIns_3 = ces_3_5_io_lsbOuts_3;
  assign ces_3_6_io_lsbIns_4 = ces_3_5_io_lsbOuts_4;
  assign ces_3_6_io_lsbIns_5 = ces_3_5_io_lsbOuts_5;
  assign ces_3_6_io_lsbIns_6 = ces_3_5_io_lsbOuts_6;
  assign ces_3_6_io_lsbIns_7 = ces_3_5_io_lsbOuts_7;
  assign ces_3_7_clock = ces_3_6_io_clockOutRight;
  assign ces_3_7_io_ins_down = ces_4_7_io_outs_down;
  assign ces_3_7_io_ins_right = ces_3_6_io_outs_right;
  assign ces_3_7_io_ins_up = ces_2_7_io_outs_up;
  assign ces_3_7_io_ins_left = io_ins_left_3;
  assign ces_3_7_io_lsbIns_1 = ces_3_6_io_lsbOuts_1;
  assign ces_3_7_io_lsbIns_2 = ces_3_6_io_lsbOuts_2;
  assign ces_3_7_io_lsbIns_3 = ces_3_6_io_lsbOuts_3;
  assign ces_3_7_io_lsbIns_4 = ces_3_6_io_lsbOuts_4;
  assign ces_3_7_io_lsbIns_5 = ces_3_6_io_lsbOuts_5;
  assign ces_3_7_io_lsbIns_6 = ces_3_6_io_lsbOuts_6;
  assign ces_3_7_io_lsbIns_7 = ces_3_6_io_lsbOuts_7;
  assign ces_4_0_clock = clock;
  assign ces_4_0_io_ins_down = ces_5_0_io_outs_down;
  assign ces_4_0_io_ins_right = io_ins_right_4;
  assign ces_4_0_io_ins_up = ces_3_0_io_outs_up;
  assign ces_4_0_io_ins_left = ces_4_1_io_outs_left;
  assign ces_4_0_io_lsbIns_1 = 1'h0;
  assign ces_4_0_io_lsbIns_2 = 1'h0;
  assign ces_4_0_io_lsbIns_3 = 1'h0;
  assign ces_4_0_io_lsbIns_4 = 1'h0;
  assign ces_4_0_io_lsbIns_5 = 1'h0;
  assign ces_4_0_io_lsbIns_6 = 1'h0;
  assign ces_4_0_io_lsbIns_7 = 1'h0;
  assign ces_4_1_clock = ces_4_0_io_clockOutRight;
  assign ces_4_1_io_ins_down = ces_5_1_io_outs_down;
  assign ces_4_1_io_ins_right = ces_4_0_io_outs_right;
  assign ces_4_1_io_ins_up = ces_3_1_io_outs_up;
  assign ces_4_1_io_ins_left = ces_4_2_io_outs_left;
  assign ces_4_1_io_lsbIns_1 = ces_4_0_io_lsbOuts_1;
  assign ces_4_1_io_lsbIns_2 = ces_4_0_io_lsbOuts_2;
  assign ces_4_1_io_lsbIns_3 = ces_4_0_io_lsbOuts_3;
  assign ces_4_1_io_lsbIns_4 = ces_4_0_io_lsbOuts_4;
  assign ces_4_1_io_lsbIns_5 = ces_4_0_io_lsbOuts_5;
  assign ces_4_1_io_lsbIns_6 = ces_4_0_io_lsbOuts_6;
  assign ces_4_1_io_lsbIns_7 = ces_4_0_io_lsbOuts_7;
  assign ces_4_2_clock = ces_4_1_io_clockOutRight;
  assign ces_4_2_io_ins_down = ces_5_2_io_outs_down;
  assign ces_4_2_io_ins_right = ces_4_1_io_outs_right;
  assign ces_4_2_io_ins_up = ces_3_2_io_outs_up;
  assign ces_4_2_io_ins_left = ces_4_3_io_outs_left;
  assign ces_4_2_io_lsbIns_1 = ces_4_1_io_lsbOuts_1;
  assign ces_4_2_io_lsbIns_2 = ces_4_1_io_lsbOuts_2;
  assign ces_4_2_io_lsbIns_3 = ces_4_1_io_lsbOuts_3;
  assign ces_4_2_io_lsbIns_4 = ces_4_1_io_lsbOuts_4;
  assign ces_4_2_io_lsbIns_5 = ces_4_1_io_lsbOuts_5;
  assign ces_4_2_io_lsbIns_6 = ces_4_1_io_lsbOuts_6;
  assign ces_4_2_io_lsbIns_7 = ces_4_1_io_lsbOuts_7;
  assign ces_4_3_clock = ces_4_2_io_clockOutRight;
  assign ces_4_3_io_ins_down = ces_5_3_io_outs_down;
  assign ces_4_3_io_ins_right = ces_4_2_io_outs_right;
  assign ces_4_3_io_ins_up = ces_3_3_io_outs_up;
  assign ces_4_3_io_ins_left = ces_4_4_io_outs_left;
  assign ces_4_3_io_lsbIns_1 = ces_4_2_io_lsbOuts_1;
  assign ces_4_3_io_lsbIns_2 = ces_4_2_io_lsbOuts_2;
  assign ces_4_3_io_lsbIns_3 = ces_4_2_io_lsbOuts_3;
  assign ces_4_3_io_lsbIns_4 = ces_4_2_io_lsbOuts_4;
  assign ces_4_3_io_lsbIns_5 = ces_4_2_io_lsbOuts_5;
  assign ces_4_3_io_lsbIns_6 = ces_4_2_io_lsbOuts_6;
  assign ces_4_3_io_lsbIns_7 = ces_4_2_io_lsbOuts_7;
  assign ces_4_4_clock = ces_4_3_io_clockOutRight;
  assign ces_4_4_io_ins_down = ces_5_4_io_outs_down;
  assign ces_4_4_io_ins_right = ces_4_3_io_outs_right;
  assign ces_4_4_io_ins_up = ces_3_4_io_outs_up;
  assign ces_4_4_io_ins_left = ces_4_5_io_outs_left;
  assign ces_4_4_io_lsbIns_1 = ces_4_3_io_lsbOuts_1;
  assign ces_4_4_io_lsbIns_2 = ces_4_3_io_lsbOuts_2;
  assign ces_4_4_io_lsbIns_3 = ces_4_3_io_lsbOuts_3;
  assign ces_4_4_io_lsbIns_4 = ces_4_3_io_lsbOuts_4;
  assign ces_4_4_io_lsbIns_5 = ces_4_3_io_lsbOuts_5;
  assign ces_4_4_io_lsbIns_6 = ces_4_3_io_lsbOuts_6;
  assign ces_4_4_io_lsbIns_7 = ces_4_3_io_lsbOuts_7;
  assign ces_4_5_clock = ces_4_4_io_clockOutRight;
  assign ces_4_5_io_ins_down = ces_5_5_io_outs_down;
  assign ces_4_5_io_ins_right = ces_4_4_io_outs_right;
  assign ces_4_5_io_ins_up = ces_3_5_io_outs_up;
  assign ces_4_5_io_ins_left = ces_4_6_io_outs_left;
  assign ces_4_5_io_lsbIns_1 = ces_4_4_io_lsbOuts_1;
  assign ces_4_5_io_lsbIns_2 = ces_4_4_io_lsbOuts_2;
  assign ces_4_5_io_lsbIns_3 = ces_4_4_io_lsbOuts_3;
  assign ces_4_5_io_lsbIns_4 = ces_4_4_io_lsbOuts_4;
  assign ces_4_5_io_lsbIns_5 = ces_4_4_io_lsbOuts_5;
  assign ces_4_5_io_lsbIns_6 = ces_4_4_io_lsbOuts_6;
  assign ces_4_5_io_lsbIns_7 = ces_4_4_io_lsbOuts_7;
  assign ces_4_6_clock = ces_4_5_io_clockOutRight;
  assign ces_4_6_io_ins_down = ces_5_6_io_outs_down;
  assign ces_4_6_io_ins_right = ces_4_5_io_outs_right;
  assign ces_4_6_io_ins_up = ces_3_6_io_outs_up;
  assign ces_4_6_io_ins_left = ces_4_7_io_outs_left;
  assign ces_4_6_io_lsbIns_1 = ces_4_5_io_lsbOuts_1;
  assign ces_4_6_io_lsbIns_2 = ces_4_5_io_lsbOuts_2;
  assign ces_4_6_io_lsbIns_3 = ces_4_5_io_lsbOuts_3;
  assign ces_4_6_io_lsbIns_4 = ces_4_5_io_lsbOuts_4;
  assign ces_4_6_io_lsbIns_5 = ces_4_5_io_lsbOuts_5;
  assign ces_4_6_io_lsbIns_6 = ces_4_5_io_lsbOuts_6;
  assign ces_4_6_io_lsbIns_7 = ces_4_5_io_lsbOuts_7;
  assign ces_4_7_clock = ces_4_6_io_clockOutRight;
  assign ces_4_7_io_ins_down = ces_5_7_io_outs_down;
  assign ces_4_7_io_ins_right = ces_4_6_io_outs_right;
  assign ces_4_7_io_ins_up = ces_3_7_io_outs_up;
  assign ces_4_7_io_ins_left = io_ins_left_4;
  assign ces_4_7_io_lsbIns_1 = ces_4_6_io_lsbOuts_1;
  assign ces_4_7_io_lsbIns_2 = ces_4_6_io_lsbOuts_2;
  assign ces_4_7_io_lsbIns_3 = ces_4_6_io_lsbOuts_3;
  assign ces_4_7_io_lsbIns_4 = ces_4_6_io_lsbOuts_4;
  assign ces_4_7_io_lsbIns_5 = ces_4_6_io_lsbOuts_5;
  assign ces_4_7_io_lsbIns_6 = ces_4_6_io_lsbOuts_6;
  assign ces_4_7_io_lsbIns_7 = ces_4_6_io_lsbOuts_7;
  assign ces_5_0_clock = clock;
  assign ces_5_0_io_ins_down = ces_6_0_io_outs_down;
  assign ces_5_0_io_ins_right = io_ins_right_5;
  assign ces_5_0_io_ins_up = ces_4_0_io_outs_up;
  assign ces_5_0_io_ins_left = ces_5_1_io_outs_left;
  assign ces_5_0_io_lsbIns_1 = 1'h0;
  assign ces_5_0_io_lsbIns_2 = 1'h0;
  assign ces_5_0_io_lsbIns_3 = 1'h0;
  assign ces_5_0_io_lsbIns_4 = 1'h0;
  assign ces_5_0_io_lsbIns_5 = 1'h0;
  assign ces_5_0_io_lsbIns_6 = 1'h0;
  assign ces_5_0_io_lsbIns_7 = 1'h0;
  assign ces_5_1_clock = ces_5_0_io_clockOutRight;
  assign ces_5_1_io_ins_down = ces_6_1_io_outs_down;
  assign ces_5_1_io_ins_right = ces_5_0_io_outs_right;
  assign ces_5_1_io_ins_up = ces_4_1_io_outs_up;
  assign ces_5_1_io_ins_left = ces_5_2_io_outs_left;
  assign ces_5_1_io_lsbIns_1 = ces_5_0_io_lsbOuts_1;
  assign ces_5_1_io_lsbIns_2 = ces_5_0_io_lsbOuts_2;
  assign ces_5_1_io_lsbIns_3 = ces_5_0_io_lsbOuts_3;
  assign ces_5_1_io_lsbIns_4 = ces_5_0_io_lsbOuts_4;
  assign ces_5_1_io_lsbIns_5 = ces_5_0_io_lsbOuts_5;
  assign ces_5_1_io_lsbIns_6 = ces_5_0_io_lsbOuts_6;
  assign ces_5_1_io_lsbIns_7 = ces_5_0_io_lsbOuts_7;
  assign ces_5_2_clock = ces_5_1_io_clockOutRight;
  assign ces_5_2_io_ins_down = ces_6_2_io_outs_down;
  assign ces_5_2_io_ins_right = ces_5_1_io_outs_right;
  assign ces_5_2_io_ins_up = ces_4_2_io_outs_up;
  assign ces_5_2_io_ins_left = ces_5_3_io_outs_left;
  assign ces_5_2_io_lsbIns_1 = ces_5_1_io_lsbOuts_1;
  assign ces_5_2_io_lsbIns_2 = ces_5_1_io_lsbOuts_2;
  assign ces_5_2_io_lsbIns_3 = ces_5_1_io_lsbOuts_3;
  assign ces_5_2_io_lsbIns_4 = ces_5_1_io_lsbOuts_4;
  assign ces_5_2_io_lsbIns_5 = ces_5_1_io_lsbOuts_5;
  assign ces_5_2_io_lsbIns_6 = ces_5_1_io_lsbOuts_6;
  assign ces_5_2_io_lsbIns_7 = ces_5_1_io_lsbOuts_7;
  assign ces_5_3_clock = ces_5_2_io_clockOutRight;
  assign ces_5_3_io_ins_down = ces_6_3_io_outs_down;
  assign ces_5_3_io_ins_right = ces_5_2_io_outs_right;
  assign ces_5_3_io_ins_up = ces_4_3_io_outs_up;
  assign ces_5_3_io_ins_left = ces_5_4_io_outs_left;
  assign ces_5_3_io_lsbIns_1 = ces_5_2_io_lsbOuts_1;
  assign ces_5_3_io_lsbIns_2 = ces_5_2_io_lsbOuts_2;
  assign ces_5_3_io_lsbIns_3 = ces_5_2_io_lsbOuts_3;
  assign ces_5_3_io_lsbIns_4 = ces_5_2_io_lsbOuts_4;
  assign ces_5_3_io_lsbIns_5 = ces_5_2_io_lsbOuts_5;
  assign ces_5_3_io_lsbIns_6 = ces_5_2_io_lsbOuts_6;
  assign ces_5_3_io_lsbIns_7 = ces_5_2_io_lsbOuts_7;
  assign ces_5_4_clock = ces_5_3_io_clockOutRight;
  assign ces_5_4_io_ins_down = ces_6_4_io_outs_down;
  assign ces_5_4_io_ins_right = ces_5_3_io_outs_right;
  assign ces_5_4_io_ins_up = ces_4_4_io_outs_up;
  assign ces_5_4_io_ins_left = ces_5_5_io_outs_left;
  assign ces_5_4_io_lsbIns_1 = ces_5_3_io_lsbOuts_1;
  assign ces_5_4_io_lsbIns_2 = ces_5_3_io_lsbOuts_2;
  assign ces_5_4_io_lsbIns_3 = ces_5_3_io_lsbOuts_3;
  assign ces_5_4_io_lsbIns_4 = ces_5_3_io_lsbOuts_4;
  assign ces_5_4_io_lsbIns_5 = ces_5_3_io_lsbOuts_5;
  assign ces_5_4_io_lsbIns_6 = ces_5_3_io_lsbOuts_6;
  assign ces_5_4_io_lsbIns_7 = ces_5_3_io_lsbOuts_7;
  assign ces_5_5_clock = ces_5_4_io_clockOutRight;
  assign ces_5_5_io_ins_down = ces_6_5_io_outs_down;
  assign ces_5_5_io_ins_right = ces_5_4_io_outs_right;
  assign ces_5_5_io_ins_up = ces_4_5_io_outs_up;
  assign ces_5_5_io_ins_left = ces_5_6_io_outs_left;
  assign ces_5_5_io_lsbIns_1 = ces_5_4_io_lsbOuts_1;
  assign ces_5_5_io_lsbIns_2 = ces_5_4_io_lsbOuts_2;
  assign ces_5_5_io_lsbIns_3 = ces_5_4_io_lsbOuts_3;
  assign ces_5_5_io_lsbIns_4 = ces_5_4_io_lsbOuts_4;
  assign ces_5_5_io_lsbIns_5 = ces_5_4_io_lsbOuts_5;
  assign ces_5_5_io_lsbIns_6 = ces_5_4_io_lsbOuts_6;
  assign ces_5_5_io_lsbIns_7 = ces_5_4_io_lsbOuts_7;
  assign ces_5_6_clock = ces_5_5_io_clockOutRight;
  assign ces_5_6_io_ins_down = ces_6_6_io_outs_down;
  assign ces_5_6_io_ins_right = ces_5_5_io_outs_right;
  assign ces_5_6_io_ins_up = ces_4_6_io_outs_up;
  assign ces_5_6_io_ins_left = ces_5_7_io_outs_left;
  assign ces_5_6_io_lsbIns_1 = ces_5_5_io_lsbOuts_1;
  assign ces_5_6_io_lsbIns_2 = ces_5_5_io_lsbOuts_2;
  assign ces_5_6_io_lsbIns_3 = ces_5_5_io_lsbOuts_3;
  assign ces_5_6_io_lsbIns_4 = ces_5_5_io_lsbOuts_4;
  assign ces_5_6_io_lsbIns_5 = ces_5_5_io_lsbOuts_5;
  assign ces_5_6_io_lsbIns_6 = ces_5_5_io_lsbOuts_6;
  assign ces_5_6_io_lsbIns_7 = ces_5_5_io_lsbOuts_7;
  assign ces_5_7_clock = ces_5_6_io_clockOutRight;
  assign ces_5_7_io_ins_down = ces_6_7_io_outs_down;
  assign ces_5_7_io_ins_right = ces_5_6_io_outs_right;
  assign ces_5_7_io_ins_up = ces_4_7_io_outs_up;
  assign ces_5_7_io_ins_left = io_ins_left_5;
  assign ces_5_7_io_lsbIns_1 = ces_5_6_io_lsbOuts_1;
  assign ces_5_7_io_lsbIns_2 = ces_5_6_io_lsbOuts_2;
  assign ces_5_7_io_lsbIns_3 = ces_5_6_io_lsbOuts_3;
  assign ces_5_7_io_lsbIns_4 = ces_5_6_io_lsbOuts_4;
  assign ces_5_7_io_lsbIns_5 = ces_5_6_io_lsbOuts_5;
  assign ces_5_7_io_lsbIns_6 = ces_5_6_io_lsbOuts_6;
  assign ces_5_7_io_lsbIns_7 = ces_5_6_io_lsbOuts_7;
  assign ces_6_0_clock = clock;
  assign ces_6_0_io_ins_down = ces_7_0_io_outs_down;
  assign ces_6_0_io_ins_right = io_ins_right_6;
  assign ces_6_0_io_ins_up = ces_5_0_io_outs_up;
  assign ces_6_0_io_ins_left = ces_6_1_io_outs_left;
  assign ces_6_0_io_lsbIns_1 = 1'h0;
  assign ces_6_0_io_lsbIns_2 = 1'h0;
  assign ces_6_0_io_lsbIns_3 = 1'h0;
  assign ces_6_0_io_lsbIns_4 = 1'h0;
  assign ces_6_0_io_lsbIns_5 = 1'h0;
  assign ces_6_0_io_lsbIns_6 = 1'h0;
  assign ces_6_0_io_lsbIns_7 = 1'h0;
  assign ces_6_1_clock = ces_6_0_io_clockOutRight;
  assign ces_6_1_io_ins_down = ces_7_1_io_outs_down;
  assign ces_6_1_io_ins_right = ces_6_0_io_outs_right;
  assign ces_6_1_io_ins_up = ces_5_1_io_outs_up;
  assign ces_6_1_io_ins_left = ces_6_2_io_outs_left;
  assign ces_6_1_io_lsbIns_1 = ces_6_0_io_lsbOuts_1;
  assign ces_6_1_io_lsbIns_2 = ces_6_0_io_lsbOuts_2;
  assign ces_6_1_io_lsbIns_3 = ces_6_0_io_lsbOuts_3;
  assign ces_6_1_io_lsbIns_4 = ces_6_0_io_lsbOuts_4;
  assign ces_6_1_io_lsbIns_5 = ces_6_0_io_lsbOuts_5;
  assign ces_6_1_io_lsbIns_6 = ces_6_0_io_lsbOuts_6;
  assign ces_6_1_io_lsbIns_7 = ces_6_0_io_lsbOuts_7;
  assign ces_6_2_clock = ces_6_1_io_clockOutRight;
  assign ces_6_2_io_ins_down = ces_7_2_io_outs_down;
  assign ces_6_2_io_ins_right = ces_6_1_io_outs_right;
  assign ces_6_2_io_ins_up = ces_5_2_io_outs_up;
  assign ces_6_2_io_ins_left = ces_6_3_io_outs_left;
  assign ces_6_2_io_lsbIns_1 = ces_6_1_io_lsbOuts_1;
  assign ces_6_2_io_lsbIns_2 = ces_6_1_io_lsbOuts_2;
  assign ces_6_2_io_lsbIns_3 = ces_6_1_io_lsbOuts_3;
  assign ces_6_2_io_lsbIns_4 = ces_6_1_io_lsbOuts_4;
  assign ces_6_2_io_lsbIns_5 = ces_6_1_io_lsbOuts_5;
  assign ces_6_2_io_lsbIns_6 = ces_6_1_io_lsbOuts_6;
  assign ces_6_2_io_lsbIns_7 = ces_6_1_io_lsbOuts_7;
  assign ces_6_3_clock = ces_6_2_io_clockOutRight;
  assign ces_6_3_io_ins_down = ces_7_3_io_outs_down;
  assign ces_6_3_io_ins_right = ces_6_2_io_outs_right;
  assign ces_6_3_io_ins_up = ces_5_3_io_outs_up;
  assign ces_6_3_io_ins_left = ces_6_4_io_outs_left;
  assign ces_6_3_io_lsbIns_1 = ces_6_2_io_lsbOuts_1;
  assign ces_6_3_io_lsbIns_2 = ces_6_2_io_lsbOuts_2;
  assign ces_6_3_io_lsbIns_3 = ces_6_2_io_lsbOuts_3;
  assign ces_6_3_io_lsbIns_4 = ces_6_2_io_lsbOuts_4;
  assign ces_6_3_io_lsbIns_5 = ces_6_2_io_lsbOuts_5;
  assign ces_6_3_io_lsbIns_6 = ces_6_2_io_lsbOuts_6;
  assign ces_6_3_io_lsbIns_7 = ces_6_2_io_lsbOuts_7;
  assign ces_6_4_clock = ces_6_3_io_clockOutRight;
  assign ces_6_4_io_ins_down = ces_7_4_io_outs_down;
  assign ces_6_4_io_ins_right = ces_6_3_io_outs_right;
  assign ces_6_4_io_ins_up = ces_5_4_io_outs_up;
  assign ces_6_4_io_ins_left = ces_6_5_io_outs_left;
  assign ces_6_4_io_lsbIns_1 = ces_6_3_io_lsbOuts_1;
  assign ces_6_4_io_lsbIns_2 = ces_6_3_io_lsbOuts_2;
  assign ces_6_4_io_lsbIns_3 = ces_6_3_io_lsbOuts_3;
  assign ces_6_4_io_lsbIns_4 = ces_6_3_io_lsbOuts_4;
  assign ces_6_4_io_lsbIns_5 = ces_6_3_io_lsbOuts_5;
  assign ces_6_4_io_lsbIns_6 = ces_6_3_io_lsbOuts_6;
  assign ces_6_4_io_lsbIns_7 = ces_6_3_io_lsbOuts_7;
  assign ces_6_5_clock = ces_6_4_io_clockOutRight;
  assign ces_6_5_io_ins_down = ces_7_5_io_outs_down;
  assign ces_6_5_io_ins_right = ces_6_4_io_outs_right;
  assign ces_6_5_io_ins_up = ces_5_5_io_outs_up;
  assign ces_6_5_io_ins_left = ces_6_6_io_outs_left;
  assign ces_6_5_io_lsbIns_1 = ces_6_4_io_lsbOuts_1;
  assign ces_6_5_io_lsbIns_2 = ces_6_4_io_lsbOuts_2;
  assign ces_6_5_io_lsbIns_3 = ces_6_4_io_lsbOuts_3;
  assign ces_6_5_io_lsbIns_4 = ces_6_4_io_lsbOuts_4;
  assign ces_6_5_io_lsbIns_5 = ces_6_4_io_lsbOuts_5;
  assign ces_6_5_io_lsbIns_6 = ces_6_4_io_lsbOuts_6;
  assign ces_6_5_io_lsbIns_7 = ces_6_4_io_lsbOuts_7;
  assign ces_6_6_clock = ces_6_5_io_clockOutRight;
  assign ces_6_6_io_ins_down = ces_7_6_io_outs_down;
  assign ces_6_6_io_ins_right = ces_6_5_io_outs_right;
  assign ces_6_6_io_ins_up = ces_5_6_io_outs_up;
  assign ces_6_6_io_ins_left = ces_6_7_io_outs_left;
  assign ces_6_6_io_lsbIns_1 = ces_6_5_io_lsbOuts_1;
  assign ces_6_6_io_lsbIns_2 = ces_6_5_io_lsbOuts_2;
  assign ces_6_6_io_lsbIns_3 = ces_6_5_io_lsbOuts_3;
  assign ces_6_6_io_lsbIns_4 = ces_6_5_io_lsbOuts_4;
  assign ces_6_6_io_lsbIns_5 = ces_6_5_io_lsbOuts_5;
  assign ces_6_6_io_lsbIns_6 = ces_6_5_io_lsbOuts_6;
  assign ces_6_6_io_lsbIns_7 = ces_6_5_io_lsbOuts_7;
  assign ces_6_7_clock = ces_6_6_io_clockOutRight;
  assign ces_6_7_io_ins_down = ces_7_7_io_outs_down;
  assign ces_6_7_io_ins_right = ces_6_6_io_outs_right;
  assign ces_6_7_io_ins_up = ces_5_7_io_outs_up;
  assign ces_6_7_io_ins_left = io_ins_left_6;
  assign ces_6_7_io_lsbIns_1 = ces_6_6_io_lsbOuts_1;
  assign ces_6_7_io_lsbIns_2 = ces_6_6_io_lsbOuts_2;
  assign ces_6_7_io_lsbIns_3 = ces_6_6_io_lsbOuts_3;
  assign ces_6_7_io_lsbIns_4 = ces_6_6_io_lsbOuts_4;
  assign ces_6_7_io_lsbIns_5 = ces_6_6_io_lsbOuts_5;
  assign ces_6_7_io_lsbIns_6 = ces_6_6_io_lsbOuts_6;
  assign ces_6_7_io_lsbIns_7 = ces_6_6_io_lsbOuts_7;
  assign ces_7_0_clock = clock;
  assign ces_7_0_io_ins_down = io_ins_down_0;
  assign ces_7_0_io_ins_right = io_ins_right_7;
  assign ces_7_0_io_ins_up = ces_6_0_io_outs_up;
  assign ces_7_0_io_ins_left = ces_7_1_io_outs_left;
  assign ces_7_0_io_lsbIns_1 = 1'h0;
  assign ces_7_0_io_lsbIns_2 = 1'h0;
  assign ces_7_0_io_lsbIns_3 = 1'h0;
  assign ces_7_0_io_lsbIns_4 = 1'h0;
  assign ces_7_0_io_lsbIns_5 = 1'h0;
  assign ces_7_0_io_lsbIns_6 = 1'h0;
  assign ces_7_0_io_lsbIns_7 = 1'h0;
  assign ces_7_1_clock = ces_7_0_io_clockOutRight;
  assign ces_7_1_io_ins_down = io_ins_down_1;
  assign ces_7_1_io_ins_right = ces_7_0_io_outs_right;
  assign ces_7_1_io_ins_up = ces_6_1_io_outs_up;
  assign ces_7_1_io_ins_left = ces_7_2_io_outs_left;
  assign ces_7_1_io_lsbIns_1 = ces_7_0_io_lsbOuts_1;
  assign ces_7_1_io_lsbIns_2 = ces_7_0_io_lsbOuts_2;
  assign ces_7_1_io_lsbIns_3 = ces_7_0_io_lsbOuts_3;
  assign ces_7_1_io_lsbIns_4 = ces_7_0_io_lsbOuts_4;
  assign ces_7_1_io_lsbIns_5 = ces_7_0_io_lsbOuts_5;
  assign ces_7_1_io_lsbIns_6 = ces_7_0_io_lsbOuts_6;
  assign ces_7_1_io_lsbIns_7 = ces_7_0_io_lsbOuts_7;
  assign ces_7_2_clock = ces_7_1_io_clockOutRight;
  assign ces_7_2_io_ins_down = io_ins_down_2;
  assign ces_7_2_io_ins_right = ces_7_1_io_outs_right;
  assign ces_7_2_io_ins_up = ces_6_2_io_outs_up;
  assign ces_7_2_io_ins_left = ces_7_3_io_outs_left;
  assign ces_7_2_io_lsbIns_1 = ces_7_1_io_lsbOuts_1;
  assign ces_7_2_io_lsbIns_2 = ces_7_1_io_lsbOuts_2;
  assign ces_7_2_io_lsbIns_3 = ces_7_1_io_lsbOuts_3;
  assign ces_7_2_io_lsbIns_4 = ces_7_1_io_lsbOuts_4;
  assign ces_7_2_io_lsbIns_5 = ces_7_1_io_lsbOuts_5;
  assign ces_7_2_io_lsbIns_6 = ces_7_1_io_lsbOuts_6;
  assign ces_7_2_io_lsbIns_7 = ces_7_1_io_lsbOuts_7;
  assign ces_7_3_clock = ces_7_2_io_clockOutRight;
  assign ces_7_3_io_ins_down = io_ins_down_3;
  assign ces_7_3_io_ins_right = ces_7_2_io_outs_right;
  assign ces_7_3_io_ins_up = ces_6_3_io_outs_up;
  assign ces_7_3_io_ins_left = ces_7_4_io_outs_left;
  assign ces_7_3_io_lsbIns_1 = ces_7_2_io_lsbOuts_1;
  assign ces_7_3_io_lsbIns_2 = ces_7_2_io_lsbOuts_2;
  assign ces_7_3_io_lsbIns_3 = ces_7_2_io_lsbOuts_3;
  assign ces_7_3_io_lsbIns_4 = ces_7_2_io_lsbOuts_4;
  assign ces_7_3_io_lsbIns_5 = ces_7_2_io_lsbOuts_5;
  assign ces_7_3_io_lsbIns_6 = ces_7_2_io_lsbOuts_6;
  assign ces_7_3_io_lsbIns_7 = ces_7_2_io_lsbOuts_7;
  assign ces_7_4_clock = ces_7_3_io_clockOutRight;
  assign ces_7_4_io_ins_down = io_ins_down_4;
  assign ces_7_4_io_ins_right = ces_7_3_io_outs_right;
  assign ces_7_4_io_ins_up = ces_6_4_io_outs_up;
  assign ces_7_4_io_ins_left = ces_7_5_io_outs_left;
  assign ces_7_4_io_lsbIns_1 = ces_7_3_io_lsbOuts_1;
  assign ces_7_4_io_lsbIns_2 = ces_7_3_io_lsbOuts_2;
  assign ces_7_4_io_lsbIns_3 = ces_7_3_io_lsbOuts_3;
  assign ces_7_4_io_lsbIns_4 = ces_7_3_io_lsbOuts_4;
  assign ces_7_4_io_lsbIns_5 = ces_7_3_io_lsbOuts_5;
  assign ces_7_4_io_lsbIns_6 = ces_7_3_io_lsbOuts_6;
  assign ces_7_4_io_lsbIns_7 = ces_7_3_io_lsbOuts_7;
  assign ces_7_5_clock = ces_7_4_io_clockOutRight;
  assign ces_7_5_io_ins_down = io_ins_down_5;
  assign ces_7_5_io_ins_right = ces_7_4_io_outs_right;
  assign ces_7_5_io_ins_up = ces_6_5_io_outs_up;
  assign ces_7_5_io_ins_left = ces_7_6_io_outs_left;
  assign ces_7_5_io_lsbIns_1 = ces_7_4_io_lsbOuts_1;
  assign ces_7_5_io_lsbIns_2 = ces_7_4_io_lsbOuts_2;
  assign ces_7_5_io_lsbIns_3 = ces_7_4_io_lsbOuts_3;
  assign ces_7_5_io_lsbIns_4 = ces_7_4_io_lsbOuts_4;
  assign ces_7_5_io_lsbIns_5 = ces_7_4_io_lsbOuts_5;
  assign ces_7_5_io_lsbIns_6 = ces_7_4_io_lsbOuts_6;
  assign ces_7_5_io_lsbIns_7 = ces_7_4_io_lsbOuts_7;
  assign ces_7_6_clock = ces_7_5_io_clockOutRight;
  assign ces_7_6_io_ins_down = io_ins_down_6;
  assign ces_7_6_io_ins_right = ces_7_5_io_outs_right;
  assign ces_7_6_io_ins_up = ces_6_6_io_outs_up;
  assign ces_7_6_io_ins_left = ces_7_7_io_outs_left;
  assign ces_7_6_io_lsbIns_1 = ces_7_5_io_lsbOuts_1;
  assign ces_7_6_io_lsbIns_2 = ces_7_5_io_lsbOuts_2;
  assign ces_7_6_io_lsbIns_3 = ces_7_5_io_lsbOuts_3;
  assign ces_7_6_io_lsbIns_4 = ces_7_5_io_lsbOuts_4;
  assign ces_7_6_io_lsbIns_5 = ces_7_5_io_lsbOuts_5;
  assign ces_7_6_io_lsbIns_6 = ces_7_5_io_lsbOuts_6;
  assign ces_7_6_io_lsbIns_7 = ces_7_5_io_lsbOuts_7;
  assign ces_7_7_clock = ces_7_6_io_clockOutRight;
  assign ces_7_7_io_ins_down = io_ins_down_7;
  assign ces_7_7_io_ins_right = ces_7_6_io_outs_right;
  assign ces_7_7_io_ins_up = ces_6_7_io_outs_up;
  assign ces_7_7_io_ins_left = io_ins_left_7;
  assign ces_7_7_io_lsbIns_1 = ces_7_6_io_lsbOuts_1;
  assign ces_7_7_io_lsbIns_2 = ces_7_6_io_lsbOuts_2;
  assign ces_7_7_io_lsbIns_3 = ces_7_6_io_lsbOuts_3;
  assign ces_7_7_io_lsbIns_4 = ces_7_6_io_lsbOuts_4;
  assign ces_7_7_io_lsbIns_5 = ces_7_6_io_lsbOuts_5;
  assign ces_7_7_io_lsbIns_6 = ces_7_6_io_lsbOuts_6;
  assign ces_7_7_io_lsbIns_7 = ces_7_6_io_lsbOuts_7;
  always @(posedge ces_0_7_io_clockOutRight) begin
    REG_0 <= ces_0_7_io_lsbOuts_0;
    REG_1 <= ces_0_7_io_lsbOuts_1;
    REG_2 <= ces_0_7_io_lsbOuts_2;
    REG_3 <= ces_0_7_io_lsbOuts_3;
    REG_4 <= ces_0_7_io_lsbOuts_4;
    REG_5 <= ces_0_7_io_lsbOuts_5;
    REG_6 <= ces_0_7_io_lsbOuts_6;
    REG_7 <= ces_0_7_io_lsbOuts_7;
    REG_8 <= ces_1_7_io_lsbOuts_0;
    REG_9 <= ces_1_7_io_lsbOuts_1;
    REG_10 <= ces_1_7_io_lsbOuts_2;
    REG_11 <= ces_1_7_io_lsbOuts_3;
    REG_12 <= ces_1_7_io_lsbOuts_4;
    REG_13 <= ces_1_7_io_lsbOuts_5;
    REG_14 <= ces_1_7_io_lsbOuts_6;
    REG_15 <= ces_1_7_io_lsbOuts_7;
    REG_16 <= ces_2_7_io_lsbOuts_0;
    REG_17 <= ces_2_7_io_lsbOuts_1;
    REG_18 <= ces_2_7_io_lsbOuts_2;
    REG_19 <= ces_2_7_io_lsbOuts_3;
    REG_20 <= ces_2_7_io_lsbOuts_4;
    REG_21 <= ces_2_7_io_lsbOuts_5;
    REG_22 <= ces_2_7_io_lsbOuts_6;
    REG_23 <= ces_2_7_io_lsbOuts_7;
    REG_24 <= ces_3_7_io_lsbOuts_0;
    REG_25 <= ces_3_7_io_lsbOuts_1;
    REG_26 <= ces_3_7_io_lsbOuts_2;
    REG_27 <= ces_3_7_io_lsbOuts_3;
    REG_28 <= ces_3_7_io_lsbOuts_4;
    REG_29 <= ces_3_7_io_lsbOuts_5;
    REG_30 <= ces_3_7_io_lsbOuts_6;
    REG_31 <= ces_3_7_io_lsbOuts_7;
    REG_32 <= ces_4_7_io_lsbOuts_0;
    REG_33 <= ces_4_7_io_lsbOuts_1;
    REG_34 <= ces_4_7_io_lsbOuts_2;
    REG_35 <= ces_4_7_io_lsbOuts_3;
    REG_36 <= ces_4_7_io_lsbOuts_4;
    REG_37 <= ces_4_7_io_lsbOuts_5;
    REG_38 <= ces_4_7_io_lsbOuts_6;
    REG_39 <= ces_4_7_io_lsbOuts_7;
    REG_40 <= ces_5_7_io_lsbOuts_0;
    REG_41 <= ces_5_7_io_lsbOuts_1;
    REG_42 <= ces_5_7_io_lsbOuts_2;
    REG_43 <= ces_5_7_io_lsbOuts_3;
    REG_44 <= ces_5_7_io_lsbOuts_4;
    REG_45 <= ces_5_7_io_lsbOuts_5;
    REG_46 <= ces_5_7_io_lsbOuts_6;
    REG_47 <= ces_5_7_io_lsbOuts_7;
    REG_48 <= ces_6_7_io_lsbOuts_0;
    REG_49 <= ces_6_7_io_lsbOuts_1;
    REG_50 <= ces_6_7_io_lsbOuts_2;
    REG_51 <= ces_6_7_io_lsbOuts_3;
    REG_52 <= ces_6_7_io_lsbOuts_4;
    REG_53 <= ces_6_7_io_lsbOuts_5;
    REG_54 <= ces_6_7_io_lsbOuts_6;
    REG_55 <= ces_6_7_io_lsbOuts_7;
    REG_56 <= ces_7_7_io_lsbOuts_0;
    REG_57 <= ces_7_7_io_lsbOuts_1;
    REG_58 <= ces_7_7_io_lsbOuts_2;
    REG_59 <= ces_7_7_io_lsbOuts_3;
    REG_60 <= ces_7_7_io_lsbOuts_4;
    REG_61 <= ces_7_7_io_lsbOuts_5;
    REG_62 <= ces_7_7_io_lsbOuts_6;
    REG_63 <= ces_7_7_io_lsbOuts_7;
  end
endmodule
