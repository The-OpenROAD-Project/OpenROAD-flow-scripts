module MockArray(
  input        clock,
  input        reset,
  input  [7:0] io_insHorizontal_0_0,
  input  [7:0] io_insHorizontal_0_1,
  input  [7:0] io_insHorizontal_0_2,
  input  [7:0] io_insHorizontal_0_3,
  input  [7:0] io_insHorizontal_0_4,
  input  [7:0] io_insHorizontal_0_5,
  input  [7:0] io_insHorizontal_0_6,
  input  [7:0] io_insHorizontal_0_7,
  input  [7:0] io_insHorizontal_0_8,
  input  [7:0] io_insHorizontal_0_9,
  input  [7:0] io_insHorizontal_0_10,
  input  [7:0] io_insHorizontal_0_11,
  input  [7:0] io_insHorizontal_0_12,
  input  [7:0] io_insHorizontal_0_13,
  input  [7:0] io_insHorizontal_0_14,
  input  [7:0] io_insHorizontal_0_15,
  input  [7:0] io_insHorizontal_0_16,
  input  [7:0] io_insHorizontal_0_17,
  input  [7:0] io_insHorizontal_0_18,
  input  [7:0] io_insHorizontal_0_19,
  input  [7:0] io_insHorizontal_0_20,
  input  [7:0] io_insHorizontal_0_21,
  input  [7:0] io_insHorizontal_0_22,
  input  [7:0] io_insHorizontal_0_23,
  input  [7:0] io_insHorizontal_0_24,
  input  [7:0] io_insHorizontal_0_25,
  input  [7:0] io_insHorizontal_0_26,
  input  [7:0] io_insHorizontal_0_27,
  input  [7:0] io_insHorizontal_0_28,
  input  [7:0] io_insHorizontal_0_29,
  input  [7:0] io_insHorizontal_0_30,
  input  [7:0] io_insHorizontal_0_31,
  input  [7:0] io_insHorizontal_1_0,
  input  [7:0] io_insHorizontal_1_1,
  input  [7:0] io_insHorizontal_1_2,
  input  [7:0] io_insHorizontal_1_3,
  input  [7:0] io_insHorizontal_1_4,
  input  [7:0] io_insHorizontal_1_5,
  input  [7:0] io_insHorizontal_1_6,
  input  [7:0] io_insHorizontal_1_7,
  input  [7:0] io_insHorizontal_1_8,
  input  [7:0] io_insHorizontal_1_9,
  input  [7:0] io_insHorizontal_1_10,
  input  [7:0] io_insHorizontal_1_11,
  input  [7:0] io_insHorizontal_1_12,
  input  [7:0] io_insHorizontal_1_13,
  input  [7:0] io_insHorizontal_1_14,
  input  [7:0] io_insHorizontal_1_15,
  input  [7:0] io_insHorizontal_1_16,
  input  [7:0] io_insHorizontal_1_17,
  input  [7:0] io_insHorizontal_1_18,
  input  [7:0] io_insHorizontal_1_19,
  input  [7:0] io_insHorizontal_1_20,
  input  [7:0] io_insHorizontal_1_21,
  input  [7:0] io_insHorizontal_1_22,
  input  [7:0] io_insHorizontal_1_23,
  input  [7:0] io_insHorizontal_1_24,
  input  [7:0] io_insHorizontal_1_25,
  input  [7:0] io_insHorizontal_1_26,
  input  [7:0] io_insHorizontal_1_27,
  input  [7:0] io_insHorizontal_1_28,
  input  [7:0] io_insHorizontal_1_29,
  input  [7:0] io_insHorizontal_1_30,
  input  [7:0] io_insHorizontal_1_31,
  output [7:0] io_outsHorizontal_0_0,
  output [7:0] io_outsHorizontal_0_1,
  output [7:0] io_outsHorizontal_0_2,
  output [7:0] io_outsHorizontal_0_3,
  output [7:0] io_outsHorizontal_0_4,
  output [7:0] io_outsHorizontal_0_5,
  output [7:0] io_outsHorizontal_0_6,
  output [7:0] io_outsHorizontal_0_7,
  output [7:0] io_outsHorizontal_0_8,
  output [7:0] io_outsHorizontal_0_9,
  output [7:0] io_outsHorizontal_0_10,
  output [7:0] io_outsHorizontal_0_11,
  output [7:0] io_outsHorizontal_0_12,
  output [7:0] io_outsHorizontal_0_13,
  output [7:0] io_outsHorizontal_0_14,
  output [7:0] io_outsHorizontal_0_15,
  output [7:0] io_outsHorizontal_0_16,
  output [7:0] io_outsHorizontal_0_17,
  output [7:0] io_outsHorizontal_0_18,
  output [7:0] io_outsHorizontal_0_19,
  output [7:0] io_outsHorizontal_0_20,
  output [7:0] io_outsHorizontal_0_21,
  output [7:0] io_outsHorizontal_0_22,
  output [7:0] io_outsHorizontal_0_23,
  output [7:0] io_outsHorizontal_0_24,
  output [7:0] io_outsHorizontal_0_25,
  output [7:0] io_outsHorizontal_0_26,
  output [7:0] io_outsHorizontal_0_27,
  output [7:0] io_outsHorizontal_0_28,
  output [7:0] io_outsHorizontal_0_29,
  output [7:0] io_outsHorizontal_0_30,
  output [7:0] io_outsHorizontal_0_31,
  output [7:0] io_outsHorizontal_1_0,
  output [7:0] io_outsHorizontal_1_1,
  output [7:0] io_outsHorizontal_1_2,
  output [7:0] io_outsHorizontal_1_3,
  output [7:0] io_outsHorizontal_1_4,
  output [7:0] io_outsHorizontal_1_5,
  output [7:0] io_outsHorizontal_1_6,
  output [7:0] io_outsHorizontal_1_7,
  output [7:0] io_outsHorizontal_1_8,
  output [7:0] io_outsHorizontal_1_9,
  output [7:0] io_outsHorizontal_1_10,
  output [7:0] io_outsHorizontal_1_11,
  output [7:0] io_outsHorizontal_1_12,
  output [7:0] io_outsHorizontal_1_13,
  output [7:0] io_outsHorizontal_1_14,
  output [7:0] io_outsHorizontal_1_15,
  output [7:0] io_outsHorizontal_1_16,
  output [7:0] io_outsHorizontal_1_17,
  output [7:0] io_outsHorizontal_1_18,
  output [7:0] io_outsHorizontal_1_19,
  output [7:0] io_outsHorizontal_1_20,
  output [7:0] io_outsHorizontal_1_21,
  output [7:0] io_outsHorizontal_1_22,
  output [7:0] io_outsHorizontal_1_23,
  output [7:0] io_outsHorizontal_1_24,
  output [7:0] io_outsHorizontal_1_25,
  output [7:0] io_outsHorizontal_1_26,
  output [7:0] io_outsHorizontal_1_27,
  output [7:0] io_outsHorizontal_1_28,
  output [7:0] io_outsHorizontal_1_29,
  output [7:0] io_outsHorizontal_1_30,
  output [7:0] io_outsHorizontal_1_31,
  input  [7:0] io_insVertical_0_0,
  input  [7:0] io_insVertical_1_0,
  output [7:0] io_outsVertical_0_0,
  output [7:0] io_outsVertical_1_0,
  output       io_lsbs_0,
  output       io_lsbs_1,
  output       io_lsbs_2,
  output       io_lsbs_3,
  output       io_lsbs_4,
  output       io_lsbs_5,
  output       io_lsbs_6,
  output       io_lsbs_7,
  output       io_lsbs_8,
  output       io_lsbs_9,
  output       io_lsbs_10,
  output       io_lsbs_11,
  output       io_lsbs_12,
  output       io_lsbs_13,
  output       io_lsbs_14,
  output       io_lsbs_15,
  output       io_lsbs_16,
  output       io_lsbs_17,
  output       io_lsbs_18,
  output       io_lsbs_19,
  output       io_lsbs_20,
  output       io_lsbs_21,
  output       io_lsbs_22,
  output       io_lsbs_23,
  output       io_lsbs_24,
  output       io_lsbs_25,
  output       io_lsbs_26,
  output       io_lsbs_27,
  output       io_lsbs_28,
  output       io_lsbs_29,
  output       io_lsbs_30,
  output       io_lsbs_31
);
  wire  ces_0_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_1_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_2_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_3_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_4_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_5_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_6_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_7_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_8_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_9_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_10_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_11_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_12_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_13_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_14_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_15_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_16_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_17_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_18_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_19_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_20_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_21_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_22_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_23_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_24_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_25_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_26_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_27_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_28_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_29_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_30_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_31_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_31_io_outs_3; // @[MockArray.scala 36:52]
  Element ces_0_0 ( // @[MockArray.scala 36:52]
    .clock(ces_0_0_clock),
    .io_ins_0(ces_0_0_io_ins_0),
    .io_ins_1(ces_0_0_io_ins_1),
    .io_ins_2(ces_0_0_io_ins_2),
    .io_ins_3(ces_0_0_io_ins_3),
    .io_outs_0(ces_0_0_io_outs_0),
    .io_outs_1(ces_0_0_io_outs_1),
    .io_outs_2(ces_0_0_io_outs_2),
    .io_outs_3(ces_0_0_io_outs_3)
  );
  Element ces_0_1 ( // @[MockArray.scala 36:52]
    .clock(ces_0_1_clock),
    .io_ins_0(ces_0_1_io_ins_0),
    .io_ins_1(ces_0_1_io_ins_1),
    .io_ins_2(ces_0_1_io_ins_2),
    .io_ins_3(ces_0_1_io_ins_3),
    .io_outs_0(ces_0_1_io_outs_0),
    .io_outs_1(ces_0_1_io_outs_1),
    .io_outs_2(ces_0_1_io_outs_2),
    .io_outs_3(ces_0_1_io_outs_3)
  );
  Element ces_0_2 ( // @[MockArray.scala 36:52]
    .clock(ces_0_2_clock),
    .io_ins_0(ces_0_2_io_ins_0),
    .io_ins_1(ces_0_2_io_ins_1),
    .io_ins_2(ces_0_2_io_ins_2),
    .io_ins_3(ces_0_2_io_ins_3),
    .io_outs_0(ces_0_2_io_outs_0),
    .io_outs_1(ces_0_2_io_outs_1),
    .io_outs_2(ces_0_2_io_outs_2),
    .io_outs_3(ces_0_2_io_outs_3)
  );
  Element ces_0_3 ( // @[MockArray.scala 36:52]
    .clock(ces_0_3_clock),
    .io_ins_0(ces_0_3_io_ins_0),
    .io_ins_1(ces_0_3_io_ins_1),
    .io_ins_2(ces_0_3_io_ins_2),
    .io_ins_3(ces_0_3_io_ins_3),
    .io_outs_0(ces_0_3_io_outs_0),
    .io_outs_1(ces_0_3_io_outs_1),
    .io_outs_2(ces_0_3_io_outs_2),
    .io_outs_3(ces_0_3_io_outs_3)
  );
  Element ces_0_4 ( // @[MockArray.scala 36:52]
    .clock(ces_0_4_clock),
    .io_ins_0(ces_0_4_io_ins_0),
    .io_ins_1(ces_0_4_io_ins_1),
    .io_ins_2(ces_0_4_io_ins_2),
    .io_ins_3(ces_0_4_io_ins_3),
    .io_outs_0(ces_0_4_io_outs_0),
    .io_outs_1(ces_0_4_io_outs_1),
    .io_outs_2(ces_0_4_io_outs_2),
    .io_outs_3(ces_0_4_io_outs_3)
  );
  Element ces_0_5 ( // @[MockArray.scala 36:52]
    .clock(ces_0_5_clock),
    .io_ins_0(ces_0_5_io_ins_0),
    .io_ins_1(ces_0_5_io_ins_1),
    .io_ins_2(ces_0_5_io_ins_2),
    .io_ins_3(ces_0_5_io_ins_3),
    .io_outs_0(ces_0_5_io_outs_0),
    .io_outs_1(ces_0_5_io_outs_1),
    .io_outs_2(ces_0_5_io_outs_2),
    .io_outs_3(ces_0_5_io_outs_3)
  );
  Element ces_0_6 ( // @[MockArray.scala 36:52]
    .clock(ces_0_6_clock),
    .io_ins_0(ces_0_6_io_ins_0),
    .io_ins_1(ces_0_6_io_ins_1),
    .io_ins_2(ces_0_6_io_ins_2),
    .io_ins_3(ces_0_6_io_ins_3),
    .io_outs_0(ces_0_6_io_outs_0),
    .io_outs_1(ces_0_6_io_outs_1),
    .io_outs_2(ces_0_6_io_outs_2),
    .io_outs_3(ces_0_6_io_outs_3)
  );
  Element ces_0_7 ( // @[MockArray.scala 36:52]
    .clock(ces_0_7_clock),
    .io_ins_0(ces_0_7_io_ins_0),
    .io_ins_1(ces_0_7_io_ins_1),
    .io_ins_2(ces_0_7_io_ins_2),
    .io_ins_3(ces_0_7_io_ins_3),
    .io_outs_0(ces_0_7_io_outs_0),
    .io_outs_1(ces_0_7_io_outs_1),
    .io_outs_2(ces_0_7_io_outs_2),
    .io_outs_3(ces_0_7_io_outs_3)
  );
  Element ces_0_8 ( // @[MockArray.scala 36:52]
    .clock(ces_0_8_clock),
    .io_ins_0(ces_0_8_io_ins_0),
    .io_ins_1(ces_0_8_io_ins_1),
    .io_ins_2(ces_0_8_io_ins_2),
    .io_ins_3(ces_0_8_io_ins_3),
    .io_outs_0(ces_0_8_io_outs_0),
    .io_outs_1(ces_0_8_io_outs_1),
    .io_outs_2(ces_0_8_io_outs_2),
    .io_outs_3(ces_0_8_io_outs_3)
  );
  Element ces_0_9 ( // @[MockArray.scala 36:52]
    .clock(ces_0_9_clock),
    .io_ins_0(ces_0_9_io_ins_0),
    .io_ins_1(ces_0_9_io_ins_1),
    .io_ins_2(ces_0_9_io_ins_2),
    .io_ins_3(ces_0_9_io_ins_3),
    .io_outs_0(ces_0_9_io_outs_0),
    .io_outs_1(ces_0_9_io_outs_1),
    .io_outs_2(ces_0_9_io_outs_2),
    .io_outs_3(ces_0_9_io_outs_3)
  );
  Element ces_0_10 ( // @[MockArray.scala 36:52]
    .clock(ces_0_10_clock),
    .io_ins_0(ces_0_10_io_ins_0),
    .io_ins_1(ces_0_10_io_ins_1),
    .io_ins_2(ces_0_10_io_ins_2),
    .io_ins_3(ces_0_10_io_ins_3),
    .io_outs_0(ces_0_10_io_outs_0),
    .io_outs_1(ces_0_10_io_outs_1),
    .io_outs_2(ces_0_10_io_outs_2),
    .io_outs_3(ces_0_10_io_outs_3)
  );
  Element ces_0_11 ( // @[MockArray.scala 36:52]
    .clock(ces_0_11_clock),
    .io_ins_0(ces_0_11_io_ins_0),
    .io_ins_1(ces_0_11_io_ins_1),
    .io_ins_2(ces_0_11_io_ins_2),
    .io_ins_3(ces_0_11_io_ins_3),
    .io_outs_0(ces_0_11_io_outs_0),
    .io_outs_1(ces_0_11_io_outs_1),
    .io_outs_2(ces_0_11_io_outs_2),
    .io_outs_3(ces_0_11_io_outs_3)
  );
  Element ces_0_12 ( // @[MockArray.scala 36:52]
    .clock(ces_0_12_clock),
    .io_ins_0(ces_0_12_io_ins_0),
    .io_ins_1(ces_0_12_io_ins_1),
    .io_ins_2(ces_0_12_io_ins_2),
    .io_ins_3(ces_0_12_io_ins_3),
    .io_outs_0(ces_0_12_io_outs_0),
    .io_outs_1(ces_0_12_io_outs_1),
    .io_outs_2(ces_0_12_io_outs_2),
    .io_outs_3(ces_0_12_io_outs_3)
  );
  Element ces_0_13 ( // @[MockArray.scala 36:52]
    .clock(ces_0_13_clock),
    .io_ins_0(ces_0_13_io_ins_0),
    .io_ins_1(ces_0_13_io_ins_1),
    .io_ins_2(ces_0_13_io_ins_2),
    .io_ins_3(ces_0_13_io_ins_3),
    .io_outs_0(ces_0_13_io_outs_0),
    .io_outs_1(ces_0_13_io_outs_1),
    .io_outs_2(ces_0_13_io_outs_2),
    .io_outs_3(ces_0_13_io_outs_3)
  );
  Element ces_0_14 ( // @[MockArray.scala 36:52]
    .clock(ces_0_14_clock),
    .io_ins_0(ces_0_14_io_ins_0),
    .io_ins_1(ces_0_14_io_ins_1),
    .io_ins_2(ces_0_14_io_ins_2),
    .io_ins_3(ces_0_14_io_ins_3),
    .io_outs_0(ces_0_14_io_outs_0),
    .io_outs_1(ces_0_14_io_outs_1),
    .io_outs_2(ces_0_14_io_outs_2),
    .io_outs_3(ces_0_14_io_outs_3)
  );
  Element ces_0_15 ( // @[MockArray.scala 36:52]
    .clock(ces_0_15_clock),
    .io_ins_0(ces_0_15_io_ins_0),
    .io_ins_1(ces_0_15_io_ins_1),
    .io_ins_2(ces_0_15_io_ins_2),
    .io_ins_3(ces_0_15_io_ins_3),
    .io_outs_0(ces_0_15_io_outs_0),
    .io_outs_1(ces_0_15_io_outs_1),
    .io_outs_2(ces_0_15_io_outs_2),
    .io_outs_3(ces_0_15_io_outs_3)
  );
  Element ces_0_16 ( // @[MockArray.scala 36:52]
    .clock(ces_0_16_clock),
    .io_ins_0(ces_0_16_io_ins_0),
    .io_ins_1(ces_0_16_io_ins_1),
    .io_ins_2(ces_0_16_io_ins_2),
    .io_ins_3(ces_0_16_io_ins_3),
    .io_outs_0(ces_0_16_io_outs_0),
    .io_outs_1(ces_0_16_io_outs_1),
    .io_outs_2(ces_0_16_io_outs_2),
    .io_outs_3(ces_0_16_io_outs_3)
  );
  Element ces_0_17 ( // @[MockArray.scala 36:52]
    .clock(ces_0_17_clock),
    .io_ins_0(ces_0_17_io_ins_0),
    .io_ins_1(ces_0_17_io_ins_1),
    .io_ins_2(ces_0_17_io_ins_2),
    .io_ins_3(ces_0_17_io_ins_3),
    .io_outs_0(ces_0_17_io_outs_0),
    .io_outs_1(ces_0_17_io_outs_1),
    .io_outs_2(ces_0_17_io_outs_2),
    .io_outs_3(ces_0_17_io_outs_3)
  );
  Element ces_0_18 ( // @[MockArray.scala 36:52]
    .clock(ces_0_18_clock),
    .io_ins_0(ces_0_18_io_ins_0),
    .io_ins_1(ces_0_18_io_ins_1),
    .io_ins_2(ces_0_18_io_ins_2),
    .io_ins_3(ces_0_18_io_ins_3),
    .io_outs_0(ces_0_18_io_outs_0),
    .io_outs_1(ces_0_18_io_outs_1),
    .io_outs_2(ces_0_18_io_outs_2),
    .io_outs_3(ces_0_18_io_outs_3)
  );
  Element ces_0_19 ( // @[MockArray.scala 36:52]
    .clock(ces_0_19_clock),
    .io_ins_0(ces_0_19_io_ins_0),
    .io_ins_1(ces_0_19_io_ins_1),
    .io_ins_2(ces_0_19_io_ins_2),
    .io_ins_3(ces_0_19_io_ins_3),
    .io_outs_0(ces_0_19_io_outs_0),
    .io_outs_1(ces_0_19_io_outs_1),
    .io_outs_2(ces_0_19_io_outs_2),
    .io_outs_3(ces_0_19_io_outs_3)
  );
  Element ces_0_20 ( // @[MockArray.scala 36:52]
    .clock(ces_0_20_clock),
    .io_ins_0(ces_0_20_io_ins_0),
    .io_ins_1(ces_0_20_io_ins_1),
    .io_ins_2(ces_0_20_io_ins_2),
    .io_ins_3(ces_0_20_io_ins_3),
    .io_outs_0(ces_0_20_io_outs_0),
    .io_outs_1(ces_0_20_io_outs_1),
    .io_outs_2(ces_0_20_io_outs_2),
    .io_outs_3(ces_0_20_io_outs_3)
  );
  Element ces_0_21 ( // @[MockArray.scala 36:52]
    .clock(ces_0_21_clock),
    .io_ins_0(ces_0_21_io_ins_0),
    .io_ins_1(ces_0_21_io_ins_1),
    .io_ins_2(ces_0_21_io_ins_2),
    .io_ins_3(ces_0_21_io_ins_3),
    .io_outs_0(ces_0_21_io_outs_0),
    .io_outs_1(ces_0_21_io_outs_1),
    .io_outs_2(ces_0_21_io_outs_2),
    .io_outs_3(ces_0_21_io_outs_3)
  );
  Element ces_0_22 ( // @[MockArray.scala 36:52]
    .clock(ces_0_22_clock),
    .io_ins_0(ces_0_22_io_ins_0),
    .io_ins_1(ces_0_22_io_ins_1),
    .io_ins_2(ces_0_22_io_ins_2),
    .io_ins_3(ces_0_22_io_ins_3),
    .io_outs_0(ces_0_22_io_outs_0),
    .io_outs_1(ces_0_22_io_outs_1),
    .io_outs_2(ces_0_22_io_outs_2),
    .io_outs_3(ces_0_22_io_outs_3)
  );
  Element ces_0_23 ( // @[MockArray.scala 36:52]
    .clock(ces_0_23_clock),
    .io_ins_0(ces_0_23_io_ins_0),
    .io_ins_1(ces_0_23_io_ins_1),
    .io_ins_2(ces_0_23_io_ins_2),
    .io_ins_3(ces_0_23_io_ins_3),
    .io_outs_0(ces_0_23_io_outs_0),
    .io_outs_1(ces_0_23_io_outs_1),
    .io_outs_2(ces_0_23_io_outs_2),
    .io_outs_3(ces_0_23_io_outs_3)
  );
  Element ces_0_24 ( // @[MockArray.scala 36:52]
    .clock(ces_0_24_clock),
    .io_ins_0(ces_0_24_io_ins_0),
    .io_ins_1(ces_0_24_io_ins_1),
    .io_ins_2(ces_0_24_io_ins_2),
    .io_ins_3(ces_0_24_io_ins_3),
    .io_outs_0(ces_0_24_io_outs_0),
    .io_outs_1(ces_0_24_io_outs_1),
    .io_outs_2(ces_0_24_io_outs_2),
    .io_outs_3(ces_0_24_io_outs_3)
  );
  Element ces_0_25 ( // @[MockArray.scala 36:52]
    .clock(ces_0_25_clock),
    .io_ins_0(ces_0_25_io_ins_0),
    .io_ins_1(ces_0_25_io_ins_1),
    .io_ins_2(ces_0_25_io_ins_2),
    .io_ins_3(ces_0_25_io_ins_3),
    .io_outs_0(ces_0_25_io_outs_0),
    .io_outs_1(ces_0_25_io_outs_1),
    .io_outs_2(ces_0_25_io_outs_2),
    .io_outs_3(ces_0_25_io_outs_3)
  );
  Element ces_0_26 ( // @[MockArray.scala 36:52]
    .clock(ces_0_26_clock),
    .io_ins_0(ces_0_26_io_ins_0),
    .io_ins_1(ces_0_26_io_ins_1),
    .io_ins_2(ces_0_26_io_ins_2),
    .io_ins_3(ces_0_26_io_ins_3),
    .io_outs_0(ces_0_26_io_outs_0),
    .io_outs_1(ces_0_26_io_outs_1),
    .io_outs_2(ces_0_26_io_outs_2),
    .io_outs_3(ces_0_26_io_outs_3)
  );
  Element ces_0_27 ( // @[MockArray.scala 36:52]
    .clock(ces_0_27_clock),
    .io_ins_0(ces_0_27_io_ins_0),
    .io_ins_1(ces_0_27_io_ins_1),
    .io_ins_2(ces_0_27_io_ins_2),
    .io_ins_3(ces_0_27_io_ins_3),
    .io_outs_0(ces_0_27_io_outs_0),
    .io_outs_1(ces_0_27_io_outs_1),
    .io_outs_2(ces_0_27_io_outs_2),
    .io_outs_3(ces_0_27_io_outs_3)
  );
  Element ces_0_28 ( // @[MockArray.scala 36:52]
    .clock(ces_0_28_clock),
    .io_ins_0(ces_0_28_io_ins_0),
    .io_ins_1(ces_0_28_io_ins_1),
    .io_ins_2(ces_0_28_io_ins_2),
    .io_ins_3(ces_0_28_io_ins_3),
    .io_outs_0(ces_0_28_io_outs_0),
    .io_outs_1(ces_0_28_io_outs_1),
    .io_outs_2(ces_0_28_io_outs_2),
    .io_outs_3(ces_0_28_io_outs_3)
  );
  Element ces_0_29 ( // @[MockArray.scala 36:52]
    .clock(ces_0_29_clock),
    .io_ins_0(ces_0_29_io_ins_0),
    .io_ins_1(ces_0_29_io_ins_1),
    .io_ins_2(ces_0_29_io_ins_2),
    .io_ins_3(ces_0_29_io_ins_3),
    .io_outs_0(ces_0_29_io_outs_0),
    .io_outs_1(ces_0_29_io_outs_1),
    .io_outs_2(ces_0_29_io_outs_2),
    .io_outs_3(ces_0_29_io_outs_3)
  );
  Element ces_0_30 ( // @[MockArray.scala 36:52]
    .clock(ces_0_30_clock),
    .io_ins_0(ces_0_30_io_ins_0),
    .io_ins_1(ces_0_30_io_ins_1),
    .io_ins_2(ces_0_30_io_ins_2),
    .io_ins_3(ces_0_30_io_ins_3),
    .io_outs_0(ces_0_30_io_outs_0),
    .io_outs_1(ces_0_30_io_outs_1),
    .io_outs_2(ces_0_30_io_outs_2),
    .io_outs_3(ces_0_30_io_outs_3)
  );
  Element ces_0_31 ( // @[MockArray.scala 36:52]
    .clock(ces_0_31_clock),
    .io_ins_0(ces_0_31_io_ins_0),
    .io_ins_1(ces_0_31_io_ins_1),
    .io_ins_2(ces_0_31_io_ins_2),
    .io_ins_3(ces_0_31_io_ins_3),
    .io_outs_0(ces_0_31_io_outs_0),
    .io_outs_1(ces_0_31_io_outs_1),
    .io_outs_2(ces_0_31_io_outs_2),
    .io_outs_3(ces_0_31_io_outs_3)
  );
  assign io_outsHorizontal_0_0 = ces_0_0_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_1 = ces_0_1_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_2 = ces_0_2_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_3 = ces_0_3_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_4 = ces_0_4_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_5 = ces_0_5_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_6 = ces_0_6_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_7 = ces_0_7_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_8 = ces_0_8_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_9 = ces_0_9_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_10 = ces_0_10_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_11 = ces_0_11_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_12 = ces_0_12_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_13 = ces_0_13_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_14 = ces_0_14_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_15 = ces_0_15_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_16 = ces_0_16_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_17 = ces_0_17_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_18 = ces_0_18_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_19 = ces_0_19_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_20 = ces_0_20_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_21 = ces_0_21_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_22 = ces_0_22_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_23 = ces_0_23_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_24 = ces_0_24_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_25 = ces_0_25_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_26 = ces_0_26_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_27 = ces_0_27_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_28 = ces_0_28_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_29 = ces_0_29_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_30 = ces_0_30_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_31 = ces_0_31_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_1_0 = ces_0_0_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_1 = ces_0_1_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_2 = ces_0_2_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_3 = ces_0_3_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_4 = ces_0_4_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_5 = ces_0_5_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_6 = ces_0_6_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_7 = ces_0_7_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_8 = ces_0_8_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_9 = ces_0_9_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_10 = ces_0_10_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_11 = ces_0_11_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_12 = ces_0_12_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_13 = ces_0_13_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_14 = ces_0_14_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_15 = ces_0_15_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_16 = ces_0_16_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_17 = ces_0_17_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_18 = ces_0_18_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_19 = ces_0_19_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_20 = ces_0_20_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_21 = ces_0_21_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_22 = ces_0_22_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_23 = ces_0_23_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_24 = ces_0_24_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_25 = ces_0_25_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_26 = ces_0_26_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_27 = ces_0_27_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_28 = ces_0_28_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_29 = ces_0_29_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_30 = ces_0_30_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_31 = ces_0_31_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_0 = ces_0_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_1_0 = ces_0_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_lsbs_0 = ces_0_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1 = ces_0_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_2 = ces_0_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_3 = ces_0_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_4 = ces_0_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_5 = ces_0_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_6 = ces_0_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_7 = ces_0_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_8 = ces_0_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_9 = ces_0_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_10 = ces_0_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_11 = ces_0_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_12 = ces_0_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_13 = ces_0_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_14 = ces_0_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_15 = ces_0_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_16 = ces_0_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_17 = ces_0_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_18 = ces_0_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_19 = ces_0_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_20 = ces_0_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_21 = ces_0_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_22 = ces_0_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_23 = ces_0_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_24 = ces_0_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_25 = ces_0_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_26 = ces_0_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_27 = ces_0_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_28 = ces_0_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_29 = ces_0_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_30 = ces_0_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_31 = ces_0_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign ces_0_0_clock = clock;
  assign ces_0_0_io_ins_0 = io_insHorizontal_0_0; // @[MockArray.scala 44:87]
  assign ces_0_0_io_ins_1 = ces_0_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_0_io_ins_2 = io_insHorizontal_1_0; // @[MockArray.scala 46:87]
  assign ces_0_0_io_ins_3 = io_insVertical_1_0; // @[MockArray.scala 47:87]
  assign ces_0_1_clock = clock;
  assign ces_0_1_io_ins_0 = io_insHorizontal_0_1; // @[MockArray.scala 44:87]
  assign ces_0_1_io_ins_1 = ces_0_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_1_io_ins_2 = io_insHorizontal_1_1; // @[MockArray.scala 46:87]
  assign ces_0_1_io_ins_3 = ces_0_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_2_clock = clock;
  assign ces_0_2_io_ins_0 = io_insHorizontal_0_2; // @[MockArray.scala 44:87]
  assign ces_0_2_io_ins_1 = ces_0_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_2_io_ins_2 = io_insHorizontal_1_2; // @[MockArray.scala 46:87]
  assign ces_0_2_io_ins_3 = ces_0_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_3_clock = clock;
  assign ces_0_3_io_ins_0 = io_insHorizontal_0_3; // @[MockArray.scala 44:87]
  assign ces_0_3_io_ins_1 = ces_0_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_3_io_ins_2 = io_insHorizontal_1_3; // @[MockArray.scala 46:87]
  assign ces_0_3_io_ins_3 = ces_0_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_4_clock = clock;
  assign ces_0_4_io_ins_0 = io_insHorizontal_0_4; // @[MockArray.scala 44:87]
  assign ces_0_4_io_ins_1 = ces_0_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_4_io_ins_2 = io_insHorizontal_1_4; // @[MockArray.scala 46:87]
  assign ces_0_4_io_ins_3 = ces_0_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_5_clock = clock;
  assign ces_0_5_io_ins_0 = io_insHorizontal_0_5; // @[MockArray.scala 44:87]
  assign ces_0_5_io_ins_1 = ces_0_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_5_io_ins_2 = io_insHorizontal_1_5; // @[MockArray.scala 46:87]
  assign ces_0_5_io_ins_3 = ces_0_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_6_clock = clock;
  assign ces_0_6_io_ins_0 = io_insHorizontal_0_6; // @[MockArray.scala 44:87]
  assign ces_0_6_io_ins_1 = ces_0_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_6_io_ins_2 = io_insHorizontal_1_6; // @[MockArray.scala 46:87]
  assign ces_0_6_io_ins_3 = ces_0_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_7_clock = clock;
  assign ces_0_7_io_ins_0 = io_insHorizontal_0_7; // @[MockArray.scala 44:87]
  assign ces_0_7_io_ins_1 = ces_0_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_7_io_ins_2 = io_insHorizontal_1_7; // @[MockArray.scala 46:87]
  assign ces_0_7_io_ins_3 = ces_0_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_8_clock = clock;
  assign ces_0_8_io_ins_0 = io_insHorizontal_0_8; // @[MockArray.scala 44:87]
  assign ces_0_8_io_ins_1 = ces_0_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_8_io_ins_2 = io_insHorizontal_1_8; // @[MockArray.scala 46:87]
  assign ces_0_8_io_ins_3 = ces_0_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_9_clock = clock;
  assign ces_0_9_io_ins_0 = io_insHorizontal_0_9; // @[MockArray.scala 44:87]
  assign ces_0_9_io_ins_1 = ces_0_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_9_io_ins_2 = io_insHorizontal_1_9; // @[MockArray.scala 46:87]
  assign ces_0_9_io_ins_3 = ces_0_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_10_clock = clock;
  assign ces_0_10_io_ins_0 = io_insHorizontal_0_10; // @[MockArray.scala 44:87]
  assign ces_0_10_io_ins_1 = ces_0_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_10_io_ins_2 = io_insHorizontal_1_10; // @[MockArray.scala 46:87]
  assign ces_0_10_io_ins_3 = ces_0_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_11_clock = clock;
  assign ces_0_11_io_ins_0 = io_insHorizontal_0_11; // @[MockArray.scala 44:87]
  assign ces_0_11_io_ins_1 = ces_0_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_11_io_ins_2 = io_insHorizontal_1_11; // @[MockArray.scala 46:87]
  assign ces_0_11_io_ins_3 = ces_0_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_12_clock = clock;
  assign ces_0_12_io_ins_0 = io_insHorizontal_0_12; // @[MockArray.scala 44:87]
  assign ces_0_12_io_ins_1 = ces_0_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_12_io_ins_2 = io_insHorizontal_1_12; // @[MockArray.scala 46:87]
  assign ces_0_12_io_ins_3 = ces_0_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_13_clock = clock;
  assign ces_0_13_io_ins_0 = io_insHorizontal_0_13; // @[MockArray.scala 44:87]
  assign ces_0_13_io_ins_1 = ces_0_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_13_io_ins_2 = io_insHorizontal_1_13; // @[MockArray.scala 46:87]
  assign ces_0_13_io_ins_3 = ces_0_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_14_clock = clock;
  assign ces_0_14_io_ins_0 = io_insHorizontal_0_14; // @[MockArray.scala 44:87]
  assign ces_0_14_io_ins_1 = ces_0_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_14_io_ins_2 = io_insHorizontal_1_14; // @[MockArray.scala 46:87]
  assign ces_0_14_io_ins_3 = ces_0_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_15_clock = clock;
  assign ces_0_15_io_ins_0 = io_insHorizontal_0_15; // @[MockArray.scala 44:87]
  assign ces_0_15_io_ins_1 = ces_0_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_15_io_ins_2 = io_insHorizontal_1_15; // @[MockArray.scala 46:87]
  assign ces_0_15_io_ins_3 = ces_0_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_16_clock = clock;
  assign ces_0_16_io_ins_0 = io_insHorizontal_0_16; // @[MockArray.scala 44:87]
  assign ces_0_16_io_ins_1 = ces_0_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_16_io_ins_2 = io_insHorizontal_1_16; // @[MockArray.scala 46:87]
  assign ces_0_16_io_ins_3 = ces_0_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_17_clock = clock;
  assign ces_0_17_io_ins_0 = io_insHorizontal_0_17; // @[MockArray.scala 44:87]
  assign ces_0_17_io_ins_1 = ces_0_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_17_io_ins_2 = io_insHorizontal_1_17; // @[MockArray.scala 46:87]
  assign ces_0_17_io_ins_3 = ces_0_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_18_clock = clock;
  assign ces_0_18_io_ins_0 = io_insHorizontal_0_18; // @[MockArray.scala 44:87]
  assign ces_0_18_io_ins_1 = ces_0_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_18_io_ins_2 = io_insHorizontal_1_18; // @[MockArray.scala 46:87]
  assign ces_0_18_io_ins_3 = ces_0_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_19_clock = clock;
  assign ces_0_19_io_ins_0 = io_insHorizontal_0_19; // @[MockArray.scala 44:87]
  assign ces_0_19_io_ins_1 = ces_0_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_19_io_ins_2 = io_insHorizontal_1_19; // @[MockArray.scala 46:87]
  assign ces_0_19_io_ins_3 = ces_0_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_20_clock = clock;
  assign ces_0_20_io_ins_0 = io_insHorizontal_0_20; // @[MockArray.scala 44:87]
  assign ces_0_20_io_ins_1 = ces_0_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_20_io_ins_2 = io_insHorizontal_1_20; // @[MockArray.scala 46:87]
  assign ces_0_20_io_ins_3 = ces_0_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_21_clock = clock;
  assign ces_0_21_io_ins_0 = io_insHorizontal_0_21; // @[MockArray.scala 44:87]
  assign ces_0_21_io_ins_1 = ces_0_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_21_io_ins_2 = io_insHorizontal_1_21; // @[MockArray.scala 46:87]
  assign ces_0_21_io_ins_3 = ces_0_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_22_clock = clock;
  assign ces_0_22_io_ins_0 = io_insHorizontal_0_22; // @[MockArray.scala 44:87]
  assign ces_0_22_io_ins_1 = ces_0_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_22_io_ins_2 = io_insHorizontal_1_22; // @[MockArray.scala 46:87]
  assign ces_0_22_io_ins_3 = ces_0_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_23_clock = clock;
  assign ces_0_23_io_ins_0 = io_insHorizontal_0_23; // @[MockArray.scala 44:87]
  assign ces_0_23_io_ins_1 = ces_0_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_23_io_ins_2 = io_insHorizontal_1_23; // @[MockArray.scala 46:87]
  assign ces_0_23_io_ins_3 = ces_0_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_24_clock = clock;
  assign ces_0_24_io_ins_0 = io_insHorizontal_0_24; // @[MockArray.scala 44:87]
  assign ces_0_24_io_ins_1 = ces_0_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_24_io_ins_2 = io_insHorizontal_1_24; // @[MockArray.scala 46:87]
  assign ces_0_24_io_ins_3 = ces_0_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_25_clock = clock;
  assign ces_0_25_io_ins_0 = io_insHorizontal_0_25; // @[MockArray.scala 44:87]
  assign ces_0_25_io_ins_1 = ces_0_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_25_io_ins_2 = io_insHorizontal_1_25; // @[MockArray.scala 46:87]
  assign ces_0_25_io_ins_3 = ces_0_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_26_clock = clock;
  assign ces_0_26_io_ins_0 = io_insHorizontal_0_26; // @[MockArray.scala 44:87]
  assign ces_0_26_io_ins_1 = ces_0_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_26_io_ins_2 = io_insHorizontal_1_26; // @[MockArray.scala 46:87]
  assign ces_0_26_io_ins_3 = ces_0_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_27_clock = clock;
  assign ces_0_27_io_ins_0 = io_insHorizontal_0_27; // @[MockArray.scala 44:87]
  assign ces_0_27_io_ins_1 = ces_0_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_27_io_ins_2 = io_insHorizontal_1_27; // @[MockArray.scala 46:87]
  assign ces_0_27_io_ins_3 = ces_0_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_28_clock = clock;
  assign ces_0_28_io_ins_0 = io_insHorizontal_0_28; // @[MockArray.scala 44:87]
  assign ces_0_28_io_ins_1 = ces_0_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_28_io_ins_2 = io_insHorizontal_1_28; // @[MockArray.scala 46:87]
  assign ces_0_28_io_ins_3 = ces_0_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_29_clock = clock;
  assign ces_0_29_io_ins_0 = io_insHorizontal_0_29; // @[MockArray.scala 44:87]
  assign ces_0_29_io_ins_1 = ces_0_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_29_io_ins_2 = io_insHorizontal_1_29; // @[MockArray.scala 46:87]
  assign ces_0_29_io_ins_3 = ces_0_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_30_clock = clock;
  assign ces_0_30_io_ins_0 = io_insHorizontal_0_30; // @[MockArray.scala 44:87]
  assign ces_0_30_io_ins_1 = ces_0_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_30_io_ins_2 = io_insHorizontal_1_30; // @[MockArray.scala 46:87]
  assign ces_0_30_io_ins_3 = ces_0_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_31_clock = clock;
  assign ces_0_31_io_ins_0 = io_insHorizontal_0_31; // @[MockArray.scala 44:87]
  assign ces_0_31_io_ins_1 = io_insVertical_0_0; // @[MockArray.scala 45:87]
  assign ces_0_31_io_ins_2 = io_insHorizontal_1_31; // @[MockArray.scala 46:87]
  assign ces_0_31_io_ins_3 = ces_0_30_io_outs_1; // @[MockArray.scala 63:19]
endmodule
