(* blackbox *) module AND2x2_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module AND2x4_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module AND2x6_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module AND3x1_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module AND3x2_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module AND3x4_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module AND4x1_ASAP7_75t_R (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module AND4x2_ASAP7_75t_R (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module AND5x1_ASAP7_75t_R (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module AND5x2_ASAP7_75t_R (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module FAx1_ASAP7_75t_R (CON, SN, A, B, CI);
	output CON, SN;
	input A, B, CI;
endmodule
(* blackbox *) module HAxp5_ASAP7_75t_R (CON, SN, A, B);
	output CON, SN;
	input A, B;
endmodule
(* blackbox *) module MAJIxp5_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module MAJx2_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module MAJx3_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NAND2x1_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2x1p5_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2x2_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2xp33_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2xp5_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND2xp67_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NAND3x1_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NAND3x2_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NAND3xp33_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NAND4xp25_ASAP7_75t_R (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module NAND4xp75_ASAP7_75t_R (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module NAND5xp2_ASAP7_75t_R (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module NOR2x1_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR2x1p5_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR2x2_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR2xp33_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR2xp67_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module NOR3x1_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NOR3x2_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NOR3xp33_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module NOR4xp25_ASAP7_75t_R (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module NOR4xp75_ASAP7_75t_R (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module NOR5xp2_ASAP7_75t_R (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module OR2x2_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module OR2x4_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module OR2x6_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module OR3x1_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module OR3x2_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module OR3x4_ASAP7_75t_R (Y, A, B, C);
	output Y;
	input A, B, C;
endmodule
(* blackbox *) module OR4x1_ASAP7_75t_R (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module OR4x2_ASAP7_75t_R (Y, A, B, C, D);
	output Y;
	input A, B, C, D;
endmodule
(* blackbox *) module OR5x1_ASAP7_75t_R (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module OR5x2_ASAP7_75t_R (Y, A, B, C, D, E);
	output Y;
	input A, B, C, D, E;
endmodule
(* blackbox *) module TIEHIx1_ASAP7_75t_R (H);
	output H;
endmodule
(* blackbox *) module TIELOx1_ASAP7_75t_R (L);
	output L;
endmodule
(* blackbox *) module XNOR2x1_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XNOR2x2_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XNOR2xp5_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XOR2x1_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XOR2x2_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
(* blackbox *) module XOR2xp5_ASAP7_75t_R (Y, A, B);
	output Y;
	input A, B;
endmodule
