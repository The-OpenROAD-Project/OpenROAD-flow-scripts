

module ibex_fetch_fifo
(
  clk_i,
  rst_ni,
  clear_i,
  in_addr_i,
  in_rdata_i,
  in_valid_i,
  in_ready_o,
  out_valid_o,
  out_ready_i,
  out_rdata_o,
  out_addr_o,
  out_valid_stored_o
);

  input [31:0] in_addr_i;
  input [31:0] in_rdata_i;
  output [31:0] out_rdata_o;
  output [31:0] out_addr_o;
  input clk_i;
  input rst_ni;
  input clear_i;
  input in_valid_i;
  input out_ready_i;
  output in_ready_o;
  output out_valid_o;
  output out_valid_stored_o;
  wire [31:0] out_rdata_o,out_addr_o,rdata;
  wire in_ready_o,out_valid_o,out_valid_stored_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,
  N12,N13,N14,N15,N16,N17,N18,N19,valid,N20,valid_unaligned,N21,N22,N23,
  addr_int_0__31_,addr_int_0__30_,addr_int_0__29_,addr_int_0__28_,addr_int_0__27_,
  addr_int_0__26_,addr_int_0__25_,addr_int_0__24_,addr_int_0__23_,addr_int_0__22_,
  addr_int_0__21_,addr_int_0__20_,addr_int_0__19_,addr_int_0__18_,addr_int_0__17_,
  addr_int_0__16_,addr_int_0__15_,addr_int_0__14_,addr_int_0__13_,addr_int_0__12_,
  addr_int_0__11_,addr_int_0__10_,addr_int_0__9_,addr_int_0__8_,addr_int_0__7_,
  addr_int_0__6_,addr_int_0__5_,addr_int_0__4_,addr_int_0__3_,addr_int_0__2_,addr_int_0__1_,
  addr_int_0__0_,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,
  N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,
  N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,
  N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,
  N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,
  N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,
  N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,
  N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,
  N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,
  N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
  N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,
  N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,
  N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,
  N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,
  N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,
  N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,
  N356,N357,N358,N359,N360,addr_n_0__31_,addr_n_0__30_,addr_n_0__29_,addr_n_0__28_,
  addr_n_0__27_,addr_n_0__26_,addr_n_0__25_,addr_n_0__24_,addr_n_0__23_,
  addr_n_0__22_,addr_n_0__21_,addr_n_0__20_,addr_n_0__19_,addr_n_0__18_,addr_n_0__17_,
  addr_n_0__16_,addr_n_0__15_,addr_n_0__14_,addr_n_0__13_,addr_n_0__12_,addr_n_0__11_,
  addr_n_0__10_,addr_n_0__9_,addr_n_0__8_,addr_n_0__7_,addr_n_0__6_,addr_n_0__5_,
  addr_n_0__4_,addr_n_0__3_,addr_n_0__2_,addr_n_0__1_,addr_n_0__0_,N361,N362,N363,N364,
  N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,
  N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,
  N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,
  N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,
  N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,
  N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,
  N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,
  N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,
  N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508;
  wire [31:16] rdata_unaligned;
  wire [95:0] rdata_int,rdata_n;
  wire [2:0] valid_int,valid_n;
  wire [31:2] addr_next;
  reg [2:0] valid_q;
  reg addr_q_0__31_,addr_q_0__30_,addr_q_0__29_,addr_q_0__28_,addr_q_0__27_,
  addr_q_0__26_,addr_q_0__25_,addr_q_0__24_,addr_q_0__23_,addr_q_0__22_,addr_q_0__21_,
  addr_q_0__20_,addr_q_0__19_,addr_q_0__18_,addr_q_0__17_,addr_q_0__16_,addr_q_0__15_,
  addr_q_0__14_,addr_q_0__13_,addr_q_0__12_,addr_q_0__11_,addr_q_0__10_,
  addr_q_0__9_,addr_q_0__8_,addr_q_0__7_,addr_q_0__6_,addr_q_0__5_,addr_q_0__4_,addr_q_0__3_,
  addr_q_0__2_,addr_q_0__1_,addr_q_0__0_;
  reg [95:0] rdata_q;

  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      valid_q[2] <= 1'b0;
    end else if(1'b1) begin
      valid_q[2] <= N501;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      valid_q[1] <= 1'b0;
    end else if(1'b1) begin
      valid_q[1] <= N500;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      valid_q[0] <= 1'b0;
    end else if(1'b1) begin
      valid_q[0] <= N499;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__31_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__31_ <= addr_n_0__31_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__30_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__30_ <= addr_n_0__30_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__29_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__29_ <= addr_n_0__29_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__28_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__28_ <= addr_n_0__28_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__27_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__27_ <= addr_n_0__27_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__26_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__26_ <= addr_n_0__26_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__25_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__25_ <= addr_n_0__25_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__24_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__24_ <= addr_n_0__24_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__23_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__23_ <= addr_n_0__23_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__22_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__22_ <= addr_n_0__22_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__21_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__21_ <= addr_n_0__21_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__20_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__20_ <= addr_n_0__20_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__19_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__19_ <= addr_n_0__19_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__18_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__18_ <= addr_n_0__18_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__17_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__17_ <= addr_n_0__17_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__16_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__16_ <= addr_n_0__16_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__15_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__15_ <= addr_n_0__15_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__14_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__14_ <= addr_n_0__14_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__13_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__13_ <= addr_n_0__13_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__12_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__12_ <= addr_n_0__12_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__11_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__11_ <= addr_n_0__11_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__10_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__10_ <= addr_n_0__10_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__9_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__9_ <= addr_n_0__9_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__8_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__8_ <= addr_n_0__8_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__7_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__7_ <= addr_n_0__7_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__6_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__6_ <= addr_n_0__6_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__5_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__5_ <= addr_n_0__5_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__4_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__4_ <= addr_n_0__4_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__3_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__3_ <= addr_n_0__3_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__2_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__2_ <= addr_n_0__2_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__1_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__1_ <= addr_n_0__1_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      addr_q_0__0_ <= 1'b0;
    end else if(N498) begin
      addr_q_0__0_ <= addr_n_0__0_;
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[95] <= 1'b0;
    end else if(N498) begin
      rdata_q[95] <= rdata_n[95];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[94] <= 1'b0;
    end else if(N498) begin
      rdata_q[94] <= rdata_n[94];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[93] <= 1'b0;
    end else if(N498) begin
      rdata_q[93] <= rdata_n[93];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[92] <= 1'b0;
    end else if(N498) begin
      rdata_q[92] <= rdata_n[92];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[91] <= 1'b0;
    end else if(N498) begin
      rdata_q[91] <= rdata_n[91];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[90] <= 1'b0;
    end else if(N498) begin
      rdata_q[90] <= rdata_n[90];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[89] <= 1'b0;
    end else if(N498) begin
      rdata_q[89] <= rdata_n[89];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[88] <= 1'b0;
    end else if(N498) begin
      rdata_q[88] <= rdata_n[88];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[87] <= 1'b0;
    end else if(N498) begin
      rdata_q[87] <= rdata_n[87];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[86] <= 1'b0;
    end else if(N498) begin
      rdata_q[86] <= rdata_n[86];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[85] <= 1'b0;
    end else if(N498) begin
      rdata_q[85] <= rdata_n[85];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[84] <= 1'b0;
    end else if(N498) begin
      rdata_q[84] <= rdata_n[84];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[83] <= 1'b0;
    end else if(N498) begin
      rdata_q[83] <= rdata_n[83];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[82] <= 1'b0;
    end else if(N498) begin
      rdata_q[82] <= rdata_n[82];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[81] <= 1'b0;
    end else if(N498) begin
      rdata_q[81] <= rdata_n[81];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[80] <= 1'b0;
    end else if(N498) begin
      rdata_q[80] <= rdata_n[80];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[79] <= 1'b0;
    end else if(N498) begin
      rdata_q[79] <= rdata_n[79];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[78] <= 1'b0;
    end else if(N498) begin
      rdata_q[78] <= rdata_n[78];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[77] <= 1'b0;
    end else if(N498) begin
      rdata_q[77] <= rdata_n[77];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[76] <= 1'b0;
    end else if(N498) begin
      rdata_q[76] <= rdata_n[76];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[75] <= 1'b0;
    end else if(N498) begin
      rdata_q[75] <= rdata_n[75];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[74] <= 1'b0;
    end else if(N498) begin
      rdata_q[74] <= rdata_n[74];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[73] <= 1'b0;
    end else if(N498) begin
      rdata_q[73] <= rdata_n[73];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[72] <= 1'b0;
    end else if(N498) begin
      rdata_q[72] <= rdata_n[72];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[71] <= 1'b0;
    end else if(N498) begin
      rdata_q[71] <= rdata_n[71];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[70] <= 1'b0;
    end else if(N498) begin
      rdata_q[70] <= rdata_n[70];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[69] <= 1'b0;
    end else if(N498) begin
      rdata_q[69] <= rdata_n[69];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[68] <= 1'b0;
    end else if(N498) begin
      rdata_q[68] <= rdata_n[68];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[67] <= 1'b0;
    end else if(N498) begin
      rdata_q[67] <= rdata_n[67];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[66] <= 1'b0;
    end else if(N498) begin
      rdata_q[66] <= rdata_n[66];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[65] <= 1'b0;
    end else if(N498) begin
      rdata_q[65] <= rdata_n[65];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[64] <= 1'b0;
    end else if(N498) begin
      rdata_q[64] <= rdata_n[64];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[63] <= 1'b0;
    end else if(N498) begin
      rdata_q[63] <= rdata_n[63];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[62] <= 1'b0;
    end else if(N498) begin
      rdata_q[62] <= rdata_n[62];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[61] <= 1'b0;
    end else if(N498) begin
      rdata_q[61] <= rdata_n[61];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[60] <= 1'b0;
    end else if(N498) begin
      rdata_q[60] <= rdata_n[60];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[59] <= 1'b0;
    end else if(N498) begin
      rdata_q[59] <= rdata_n[59];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[58] <= 1'b0;
    end else if(N498) begin
      rdata_q[58] <= rdata_n[58];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[57] <= 1'b0;
    end else if(N498) begin
      rdata_q[57] <= rdata_n[57];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[56] <= 1'b0;
    end else if(N498) begin
      rdata_q[56] <= rdata_n[56];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[55] <= 1'b0;
    end else if(N498) begin
      rdata_q[55] <= rdata_n[55];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[54] <= 1'b0;
    end else if(N498) begin
      rdata_q[54] <= rdata_n[54];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[53] <= 1'b0;
    end else if(N498) begin
      rdata_q[53] <= rdata_n[53];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[52] <= 1'b0;
    end else if(N498) begin
      rdata_q[52] <= rdata_n[52];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[51] <= 1'b0;
    end else if(N498) begin
      rdata_q[51] <= rdata_n[51];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[50] <= 1'b0;
    end else if(N498) begin
      rdata_q[50] <= rdata_n[50];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[49] <= 1'b0;
    end else if(N498) begin
      rdata_q[49] <= rdata_n[49];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[48] <= 1'b0;
    end else if(N498) begin
      rdata_q[48] <= rdata_n[48];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[47] <= 1'b0;
    end else if(N498) begin
      rdata_q[47] <= rdata_n[47];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[46] <= 1'b0;
    end else if(N498) begin
      rdata_q[46] <= rdata_n[46];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[45] <= 1'b0;
    end else if(N498) begin
      rdata_q[45] <= rdata_n[45];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[44] <= 1'b0;
    end else if(N498) begin
      rdata_q[44] <= rdata_n[44];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[43] <= 1'b0;
    end else if(N498) begin
      rdata_q[43] <= rdata_n[43];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[42] <= 1'b0;
    end else if(N498) begin
      rdata_q[42] <= rdata_n[42];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[41] <= 1'b0;
    end else if(N498) begin
      rdata_q[41] <= rdata_n[41];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[40] <= 1'b0;
    end else if(N498) begin
      rdata_q[40] <= rdata_n[40];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[39] <= 1'b0;
    end else if(N498) begin
      rdata_q[39] <= rdata_n[39];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[38] <= 1'b0;
    end else if(N498) begin
      rdata_q[38] <= rdata_n[38];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[37] <= 1'b0;
    end else if(N498) begin
      rdata_q[37] <= rdata_n[37];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[36] <= 1'b0;
    end else if(N498) begin
      rdata_q[36] <= rdata_n[36];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[35] <= 1'b0;
    end else if(N498) begin
      rdata_q[35] <= rdata_n[35];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[34] <= 1'b0;
    end else if(N498) begin
      rdata_q[34] <= rdata_n[34];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[33] <= 1'b0;
    end else if(N498) begin
      rdata_q[33] <= rdata_n[33];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[32] <= 1'b0;
    end else if(N498) begin
      rdata_q[32] <= rdata_n[32];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[31] <= 1'b0;
    end else if(N498) begin
      rdata_q[31] <= rdata_n[31];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[30] <= 1'b0;
    end else if(N498) begin
      rdata_q[30] <= rdata_n[30];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[29] <= 1'b0;
    end else if(N498) begin
      rdata_q[29] <= rdata_n[29];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[28] <= 1'b0;
    end else if(N498) begin
      rdata_q[28] <= rdata_n[28];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[27] <= 1'b0;
    end else if(N498) begin
      rdata_q[27] <= rdata_n[27];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[26] <= 1'b0;
    end else if(N498) begin
      rdata_q[26] <= rdata_n[26];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[25] <= 1'b0;
    end else if(N498) begin
      rdata_q[25] <= rdata_n[25];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[24] <= 1'b0;
    end else if(N498) begin
      rdata_q[24] <= rdata_n[24];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[23] <= 1'b0;
    end else if(N498) begin
      rdata_q[23] <= rdata_n[23];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[22] <= 1'b0;
    end else if(N498) begin
      rdata_q[22] <= rdata_n[22];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[21] <= 1'b0;
    end else if(N498) begin
      rdata_q[21] <= rdata_n[21];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[20] <= 1'b0;
    end else if(N498) begin
      rdata_q[20] <= rdata_n[20];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[19] <= 1'b0;
    end else if(N498) begin
      rdata_q[19] <= rdata_n[19];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[18] <= 1'b0;
    end else if(N498) begin
      rdata_q[18] <= rdata_n[18];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[17] <= 1'b0;
    end else if(N498) begin
      rdata_q[17] <= rdata_n[17];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[16] <= 1'b0;
    end else if(N498) begin
      rdata_q[16] <= rdata_n[16];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[15] <= 1'b0;
    end else if(N498) begin
      rdata_q[15] <= rdata_n[15];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[14] <= 1'b0;
    end else if(N498) begin
      rdata_q[14] <= rdata_n[14];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[13] <= 1'b0;
    end else if(N498) begin
      rdata_q[13] <= rdata_n[13];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[12] <= 1'b0;
    end else if(N498) begin
      rdata_q[12] <= rdata_n[12];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[11] <= 1'b0;
    end else if(N498) begin
      rdata_q[11] <= rdata_n[11];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[10] <= 1'b0;
    end else if(N498) begin
      rdata_q[10] <= rdata_n[10];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[9] <= 1'b0;
    end else if(N498) begin
      rdata_q[9] <= rdata_n[9];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[8] <= 1'b0;
    end else if(N498) begin
      rdata_q[8] <= rdata_n[8];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[7] <= 1'b0;
    end else if(N498) begin
      rdata_q[7] <= rdata_n[7];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[6] <= 1'b0;
    end else if(N498) begin
      rdata_q[6] <= rdata_n[6];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[5] <= 1'b0;
    end else if(N498) begin
      rdata_q[5] <= rdata_n[5];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[4] <= 1'b0;
    end else if(N498) begin
      rdata_q[4] <= rdata_n[4];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[3] <= 1'b0;
    end else if(N498) begin
      rdata_q[3] <= rdata_n[3];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[2] <= 1'b0;
    end else if(N498) begin
      rdata_q[2] <= rdata_n[2];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[1] <= 1'b0;
    end else if(N498) begin
      rdata_q[1] <= rdata_n[1];
    end 
  end


  always @(posedge clk_i or posedge N497) begin
    if(N497) begin
      rdata_q[0] <= 1'b0;
    end else if(N498) begin
      rdata_q[0] <= rdata_n[0];
    end 
  end

  assign N502 = rdata_q[16] & rdata_q[17];
  assign N503 = ~N502;
  assign N504 = rdata[0] & rdata[1];
  assign N505 = ~N504;
  assign N506 = rdata[16] & rdata[17];
  assign N507 = ~N506;
  assign addr_next = { addr_int_0__31_, addr_int_0__30_, addr_int_0__29_, addr_int_0__28_, addr_int_0__27_, addr_int_0__26_, addr_int_0__25_, addr_int_0__24_, addr_int_0__23_, addr_int_0__22_, addr_int_0__21_, addr_int_0__20_, addr_int_0__19_, addr_int_0__18_, addr_int_0__17_, addr_int_0__16_, addr_int_0__15_, addr_int_0__14_, addr_int_0__13_, addr_int_0__12_, addr_int_0__11_, addr_int_0__10_, addr_int_0__9_, addr_int_0__8_, addr_int_0__7_, addr_int_0__6_, addr_int_0__5_, addr_int_0__4_, addr_int_0__3_, addr_int_0__2_ } + 1'b1;
  assign rdata = (N0)? rdata_q[31:0] : 
                 (N19)? in_rdata_i : 1'b0;
  assign N0 = valid_q[0];
  assign rdata_unaligned = (N1)? rdata_q[47:32] : 
                           (N20)? in_rdata_i[15:0] : 1'b0;
  assign N1 = valid_q[1];
  assign N22 = (N2)? valid : 
               (N3)? valid_unaligned : 1'b0;
  assign N2 = N507;
  assign N3 = N506;
  assign out_rdata_o = (N4)? { rdata_unaligned, rdata[31:16] } : 
                       (N21)? rdata : 1'b0;
  assign N4 = out_addr_o[1];
  assign out_valid_o = (N4)? N22 : 
                       (N21)? valid : 1'b0;
  assign out_addr_o = (N0)? { addr_q_0__31_, addr_q_0__30_, addr_q_0__29_, addr_q_0__28_, addr_q_0__27_, addr_q_0__26_, addr_q_0__25_, addr_q_0__24_, addr_q_0__23_, addr_q_0__22_, addr_q_0__21_, addr_q_0__20_, addr_q_0__19_, addr_q_0__18_, addr_q_0__17_, addr_q_0__16_, addr_q_0__15_, addr_q_0__14_, addr_q_0__13_, addr_q_0__12_, addr_q_0__11_, addr_q_0__10_, addr_q_0__9_, addr_q_0__8_, addr_q_0__7_, addr_q_0__6_, addr_q_0__5_, addr_q_0__4_, addr_q_0__3_, addr_q_0__2_, addr_q_0__1_, addr_q_0__0_ } : 
                      (N19)? in_addr_i : 1'b0;
  assign N23 = (N5)? 1'b1 : 
               (N6)? valid_q[1] : 1'b0;
  assign N5 = N503;
  assign N6 = N502;
  assign out_valid_stored_o = (N4)? N23 : 
                              (N21)? valid_q[0] : 1'b0;
  assign { N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26 } = (N7)? in_addr_i : 
                                                                                                                                                                              (N0)? { addr_q_0__31_, addr_q_0__30_, addr_q_0__29_, addr_q_0__28_, addr_q_0__27_, addr_q_0__26_, addr_q_0__25_, addr_q_0__24_, addr_q_0__23_, addr_q_0__22_, addr_q_0__21_, addr_q_0__20_, addr_q_0__19_, addr_q_0__18_, addr_q_0__17_, addr_q_0__16_, addr_q_0__15_, addr_q_0__14_, addr_q_0__13_, addr_q_0__12_, addr_q_0__11_, addr_q_0__10_, addr_q_0__9_, addr_q_0__8_, addr_q_0__7_, addr_q_0__6_, addr_q_0__5_, addr_q_0__4_, addr_q_0__3_, addr_q_0__2_, addr_q_0__1_, addr_q_0__0_ } : 1'b0;
  assign N7 = N25;
  assign { N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58 } = (N7)? in_rdata_i : 
                                                                                                                                                                              (N0)? rdata_q[31:0] : 1'b0;
  assign N90 = (N7)? 1'b1 : 
               (N0)? valid_q[0] : 1'b0;
  assign { N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92 } = (N8)? in_rdata_i : 
                                                                                                                                                                                                      (N1)? rdata_q[63:32] : 1'b0;
  assign N8 = N91;
  assign N124 = (N8)? 1'b1 : 
                (N1)? valid_q[1] : 1'b0;
  assign N125 = (N8)? 1'b0 : 
                (N1)? valid_q[0] : 1'b0;
  assign { N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128 } = (N9)? in_rdata_i : 
                                                                                                                                                                                                              (N10)? rdata_q[95:64] : 1'b0;
  assign N9 = N127;
  assign N10 = valid_q[2];
  assign N160 = (N9)? 1'b1 : 
                (N10)? valid_q[2] : 1'b0;
  assign { N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162 } = (N11)? { N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128 } : 
                                                                                                                                                                                                              (N161)? rdata_q[95:64] : 1'b0;
  assign N11 = N125;
  assign N194 = (N11)? N160 : 
                (N161)? valid_q[2] : 1'b0;
  assign { N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195 } = (N11)? { N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162 } : 
                                                                                                                                                                                                              (N12)? rdata_q[95:64] : 1'b0;
  assign N12 = N126;
  assign N227 = (N11)? N194 : 
                (N12)? valid_q[2] : 1'b0;
  assign { N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229 } = (N0)? { N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N228)? rdata_q[95:32] : 1'b0;
  assign { N294, N293 } = (N0)? { N227, N124 } : 
                          (N228)? valid_q[2:1] : 1'b0;
  assign { N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295 } = (N0)? { N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N7)? rdata_q[95:32] : 1'b0;
  assign { N360, N359 } = (N0)? { N294, N293 } : 
                          (N7)? valid_q[2:1] : 1'b0;
  assign valid_int = (N13)? { N360, N359, N90 } : 
                     (N14)? valid_q : 1'b0;
  assign N13 = in_valid_i;
  assign N14 = N24;
  assign { addr_int_0__31_, addr_int_0__30_, addr_int_0__29_, addr_int_0__28_, addr_int_0__27_, addr_int_0__26_, addr_int_0__25_, addr_int_0__24_, addr_int_0__23_, addr_int_0__22_, addr_int_0__21_, addr_int_0__20_, addr_int_0__19_, addr_int_0__18_, addr_int_0__17_, addr_int_0__16_, addr_int_0__15_, addr_int_0__14_, addr_int_0__13_, addr_int_0__12_, addr_int_0__11_, addr_int_0__10_, addr_int_0__9_, addr_int_0__8_, addr_int_0__7_, addr_int_0__6_, addr_int_0__5_, addr_int_0__4_, addr_int_0__3_, addr_int_0__2_, addr_int_0__1_, addr_int_0__0_ } = (N13)? { N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N14)? { addr_q_0__31_, addr_q_0__30_, addr_q_0__29_, addr_q_0__28_, addr_q_0__27_, addr_q_0__26_, addr_q_0__25_, addr_q_0__24_, addr_q_0__23_, addr_q_0__22_, addr_q_0__21_, addr_q_0__20_, addr_q_0__19_, addr_q_0__18_, addr_q_0__17_, addr_q_0__16_, addr_q_0__15_, addr_q_0__14_, addr_q_0__13_, addr_q_0__12_, addr_q_0__11_, addr_q_0__10_, addr_q_0__9_, addr_q_0__8_, addr_q_0__7_, addr_q_0__6_, addr_q_0__5_, addr_q_0__4_, addr_q_0__3_, addr_q_0__2_, addr_q_0__1_, addr_q_0__0_ } : 1'b0;
  assign rdata_int = (N13)? { N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58 } : 
                     (N14)? rdata_q : 1'b0;
  assign { N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365 } = (N15)? { addr_next, N506 } : 
                                                                                                                                                                                                        (N496)? { addr_int_0__31_, addr_int_0__30_, addr_int_0__29_, addr_int_0__28_, addr_int_0__27_, addr_int_0__26_, addr_int_0__25_, addr_int_0__24_, addr_int_0__23_, addr_int_0__22_, addr_int_0__21_, addr_int_0__20_, addr_int_0__19_, addr_int_0__18_, addr_int_0__17_, addr_int_0__16_, addr_int_0__15_, addr_int_0__14_, addr_int_0__13_, addr_int_0__12_, addr_int_0__11_, addr_int_0__10_, addr_int_0__9_, addr_int_0__8_, addr_int_0__7_, addr_int_0__6_, addr_int_0__5_, addr_int_0__4_, addr_int_0__3_, addr_int_0__2_, 1'b1 } : 
                                                                                                                                                                                                        (N364)? { addr_next, 1'b0 } : 1'b0;
  assign N15 = addr_int_0__1_;
  assign { N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396 } = (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rdata_int[95:32] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N496)? rdata_int : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N364)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, rdata_int[95:32] } : 1'b0;
  assign { N494, N493, N492 } = (N15)? { 1'b0, valid_int[2:1] } : 
                                (N496)? valid_int : 
                                (N364)? { 1'b0, valid_int[2:1] } : 1'b0;
  assign valid_n = (N16)? { N494, N493, N492 } : 
                   (N362)? valid_int : 1'b0;
  assign N16 = N361;
  assign { addr_n_0__31_, addr_n_0__30_, addr_n_0__29_, addr_n_0__28_, addr_n_0__27_, addr_n_0__26_, addr_n_0__25_, addr_n_0__24_, addr_n_0__23_, addr_n_0__22_, addr_n_0__21_, addr_n_0__20_, addr_n_0__19_, addr_n_0__18_, addr_n_0__17_, addr_n_0__16_, addr_n_0__15_, addr_n_0__14_, addr_n_0__13_, addr_n_0__12_, addr_n_0__11_, addr_n_0__10_, addr_n_0__9_, addr_n_0__8_, addr_n_0__7_, addr_n_0__6_, addr_n_0__5_, addr_n_0__4_, addr_n_0__3_, addr_n_0__2_, addr_n_0__1_, addr_n_0__0_ } = (N16)? { N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N362)? { addr_int_0__31_, addr_int_0__30_, addr_int_0__29_, addr_int_0__28_, addr_int_0__27_, addr_int_0__26_, addr_int_0__25_, addr_int_0__24_, addr_int_0__23_, addr_int_0__22_, addr_int_0__21_, addr_int_0__20_, addr_int_0__19_, addr_int_0__18_, addr_int_0__17_, addr_int_0__16_, addr_int_0__15_, addr_int_0__14_, addr_int_0__13_, addr_int_0__12_, addr_int_0__11_, addr_int_0__10_, addr_int_0__9_, addr_int_0__8_, addr_int_0__7_, addr_int_0__6_, addr_int_0__5_, addr_int_0__4_, addr_int_0__3_, addr_int_0__2_, addr_int_0__1_, addr_int_0__0_ } : 1'b0;
  assign rdata_n = (N16)? { N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396 } : 
                   (N362)? rdata_int : 1'b0;
  assign { N501, N500, N499 } = (N17)? { 1'b0, 1'b0, 1'b0 } : 
                                (N18)? valid_n : 1'b0;
  assign N17 = clear_i;
  assign N18 = N498;
  assign N19 = ~valid_q[0];
  assign valid = valid_q[0] | in_valid_i;
  assign N20 = ~valid_q[1];
  assign valid_unaligned = valid_q[1] | N508;
  assign N508 = valid_q[0] & in_valid_i;
  assign N21 = ~out_addr_o[1];
  assign in_ready_o = ~valid_q[1];
  assign N24 = ~in_valid_i;
  assign N25 = ~valid_q[0];
  assign N91 = ~valid_q[1];
  assign N126 = ~N125;
  assign N127 = ~valid_q[2];
  assign N161 = ~N125;
  assign N228 = ~valid_q[0];
  assign N361 = out_ready_i & out_valid_o;
  assign N362 = ~N361;
  assign N363 = N505 | addr_int_0__1_;
  assign N364 = ~N363;
  assign N495 = ~addr_int_0__1_;
  assign N496 = N505 & N495;
  assign N497 = ~rst_ni;
  assign N498 = ~clear_i;

endmodule



module ibex_prefetch_buffer
(
  clk_i,
  rst_ni,
  req_i,
  branch_i,
  addr_i,
  ready_i,
  valid_o,
  rdata_o,
  addr_o,
  instr_req_o,
  instr_gnt_i,
  instr_addr_o,
  instr_rdata_i,
  instr_rvalid_i,
  busy_o
);

  input [31:0] addr_i;
  output [31:0] rdata_o;
  output [31:0] addr_o;
  output [31:0] instr_addr_o;
  input [31:0] instr_rdata_i;
  input clk_i;
  input rst_ni;
  input req_i;
  input branch_i;
  input ready_i;
  input instr_gnt_i;
  input instr_rvalid_i;
  output valid_o;
  output instr_req_o;
  output busy_o;
  wire [31:0] rdata_o,addr_o,instr_addr_o,fetch_addr;
  wire valid_o,instr_req_o,busy_o,N0,N1,N2,N3,N4,N5,N6,N7,fifo_valid,fifo_ready,N8,
  addr_valid,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,
  N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,
  N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,
  N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,
  N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,
  N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,
  N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,
  N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,
  N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,
  N170,N171,N172,N173;
  wire [1:0] pf_fsm_ns,instr_addr;
  reg [31:0] instr_addr_q;
  reg [1:0] pf_fsm_cs;
  assign instr_addr_o[0] = 1'b0;
  assign instr_addr_o[1] = 1'b0;

  ibex_fetch_fifo
  fifo_i
  (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .clear_i(branch_i),
    .in_addr_i(instr_addr_q),
    .in_rdata_i(instr_rdata_i),
    .in_valid_i(fifo_valid),
    .in_ready_o(fifo_ready),
    .out_valid_o(valid_o),
    .out_ready_i(ready_i),
    .out_rdata_o(rdata_o),
    .out_addr_o(addr_o)
  );

  assign N11 = N9 & N10;
  assign N12 = pf_fsm_cs[1] | N10;
  assign N14 = N9 | pf_fsm_cs[0];
  assign N16 = pf_fsm_cs[1] & pf_fsm_cs[0];

  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[31] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[31] <= instr_addr_o[31];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[30] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[30] <= instr_addr_o[30];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[29] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[29] <= instr_addr_o[29];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[28] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[28] <= instr_addr_o[28];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[27] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[27] <= instr_addr_o[27];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[26] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[26] <= instr_addr_o[26];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[25] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[25] <= instr_addr_o[25];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[24] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[24] <= instr_addr_o[24];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[23] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[23] <= instr_addr_o[23];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[22] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[22] <= instr_addr_o[22];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[21] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[21] <= instr_addr_o[21];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[20] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[20] <= instr_addr_o[20];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[19] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[19] <= instr_addr_o[19];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[18] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[18] <= instr_addr_o[18];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[17] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[17] <= instr_addr_o[17];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[16] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[16] <= instr_addr_o[16];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[15] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[15] <= instr_addr_o[15];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[14] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[14] <= instr_addr_o[14];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[13] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[13] <= instr_addr_o[13];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[12] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[12] <= instr_addr_o[12];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[11] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[11] <= instr_addr_o[11];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[10] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[10] <= instr_addr_o[10];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[9] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[9] <= instr_addr_o[9];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[8] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[8] <= instr_addr_o[8];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[7] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[7] <= instr_addr_o[7];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[6] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[6] <= instr_addr_o[6];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[5] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[5] <= instr_addr_o[5];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[4] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[4] <= instr_addr_o[4];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[3] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[3] <= instr_addr_o[3];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[2] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[2] <= instr_addr_o[2];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[1] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[1] <= instr_addr[1];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      instr_addr_q[0] <= 1'b0;
    end else if(addr_valid) begin
      instr_addr_q[0] <= instr_addr[0];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      pf_fsm_cs[1] <= 1'b0;
    end else if(N171) begin
      pf_fsm_cs[1] <= pf_fsm_ns[1];
    end 
  end


  always @(posedge clk_i or posedge N169) begin
    if(N169) begin
      pf_fsm_cs[0] <= 1'b0;
    end else if(N171) begin
      pf_fsm_cs[0] <= pf_fsm_ns[0];
    end 
  end

  assign N172 = pf_fsm_cs[0] | pf_fsm_cs[1];
  assign fetch_addr = { instr_addr_q[31:2], 1'b0, 1'b0 } + { 1'b1, 1'b0, 1'b0 };
  assign { N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18 } = (N0)? addr_i : 
                                                                                                                                                                              (N1)? fetch_addr : 1'b0;
  assign N0 = N165;
  assign N1 = N17;
  assign { N52, N51 } = (N2)? { instr_gnt_i, N86 } : 
                        (N50)? pf_fsm_cs : 1'b0;
  assign N2 = N8;
  assign { N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53 } = (N3)? addr_i : 
                                                                                                                                                                              (N1)? instr_addr_q : 1'b0;
  assign N3 = N85;
  assign { N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87 } = (N0)? addr_i : 
                                                                                                                                                                                                 (N1)? fetch_addr : 1'b0;
  assign N124 = (N4)? 1'b1 : 
                (N123)? 1'b0 : 
                (N5)? 1'b0 : 1'b0;
  assign N4 = instr_rvalid_i;
  assign N5 = 1'b0;
  assign N125 = (N4)? 1'b1 : 
                (N168)? 1'b1 : 
                (N122)? 1'b0 : 1'b0;
  assign { N127, N126 } = (N4)? { instr_gnt_i, N86 } : 
                          (N168)? { 1'b1, 1'b1 } : 
                          (N122)? pf_fsm_cs : 1'b0;
  assign { N129, N128 } = (N2)? { N127, N126 } : 
                          (N167)? { 1'b0, 1'b0 } : 
                          (N120)? pf_fsm_cs : 1'b0;
  assign N130 = (N2)? N124 : 
                (N50)? 1'b0 : 
                (N5)? 1'b0 : 1'b0;
  assign N131 = (N2)? N124 : 
                (N167)? 1'b1 : 
                (N120)? 1'b0 : 1'b0;
  assign N132 = (N2)? N125 : 
                (N50)? 1'b0 : 
                (N5)? 1'b0 : 1'b0;
  assign { N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133 } = (N0)? addr_i : 
                                                                                                                                                                                                              (N1)? instr_addr_q : 1'b0;
  assign { instr_addr_o[31:2], instr_addr } = (N6)? { N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18 } : 
                                              (N13)? { N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53 } : 
                                              (N15)? { N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87 } : 
                                              (N7)? { N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133 } : 1'b0;
  assign N6 = N11;
  assign N7 = N16;
  assign instr_req_o = (N6)? N8 : 
                       (N13)? 1'b1 : 
                       (N15)? N130 : 
                       (N7)? instr_rvalid_i : 1'b0;
  assign pf_fsm_ns = (N6)? { N52, N51 } : 
                     (N13)? { instr_gnt_i, N86 } : 
                     (N15)? { N129, N128 } : 
                     (N7)? { instr_gnt_i, N86 } : 1'b0;
  assign addr_valid = (N6)? N8 : 
                      (N13)? N85 : 
                      (N15)? N132 : 
                      (N7)? N165 : 1'b0;
  assign fifo_valid = (N6)? 1'b0 : 
                      (N13)? 1'b0 : 
                      (N15)? N131 : 
                      (N7)? 1'b0 : 1'b0;
  assign busy_o = N172 | instr_req_o;
  assign N8 = req_i & N173;
  assign N173 = fifo_ready | branch_i;
  assign N9 = ~pf_fsm_cs[1];
  assign N10 = ~pf_fsm_cs[0];
  assign N13 = ~N12;
  assign N15 = ~N14;
  assign N17 = ~branch_i;
  assign N165 = branch_i;
  assign N50 = ~N8;
  assign N85 = branch_i;
  assign N86 = ~instr_gnt_i;
  assign N119 = instr_rvalid_i | N8;
  assign N120 = ~N119;
  assign N121 = N165 | instr_rvalid_i;
  assign N122 = ~N121;
  assign N123 = ~instr_rvalid_i;
  assign N166 = ~instr_rvalid_i;
  assign N167 = instr_rvalid_i & N50;
  assign N168 = N165 & N123;
  assign N169 = ~rst_ni;
  assign N170 = N166 & N16;
  assign N171 = ~N170;

endmodule



module ibex_compressed_decoder
(
  instr_i,
  instr_o,
  is_compressed_o,
  illegal_instr_o
);

  input [31:0] instr_i;
  output [31:0] instr_o;
  output is_compressed_o;
  output illegal_instr_o;
  wire [31:0] instr_o;
  wire is_compressed_o,illegal_instr_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,
  N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,
  N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,
  N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,
  N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,
  N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,
  N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,
  N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,
  N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,
  N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,
  N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,
  N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,
  N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,
  N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,
  N239,N240,N241,N242,N243,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,
  N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,
  N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282;
  assign N26 = N24 & N25;
  assign N27 = instr_i[1] | N25;
  assign N29 = N24 | instr_i[0];
  assign N31 = instr_i[1] & instr_i[0];
  assign N34 = N83 & N33;
  assign N35 = instr_i[15] | N33;
  assign N37 = instr_i[15] & instr_i[14];
  assign N38 = N83 | instr_i[14];
  assign N65 = N62 & N63;
  assign N66 = N65 & N64;
  assign N67 = instr_i[15] | instr_i[14];
  assign N68 = N67 | N64;
  assign N69 = N62 | instr_i[14];
  assign N70 = N69 | N64;
  assign N72 = instr_i[15] | N63;
  assign N73 = N72 | instr_i[13];
  assign N75 = N72 | N64;
  assign N77 = N69 | instr_i[13];
  assign N79 = N62 | N63;
  assign N80 = N79 | instr_i[13];
  assign N81 = N37 & instr_i[13];
  assign N106 = N103 & N104;
  assign N107 = N106 & N105;
  assign N108 = instr_i[12] | instr_i[6];
  assign N109 = N108 | N105;
  assign N111 = instr_i[12] | N104;
  assign N112 = N111 | instr_i[5];
  assign N114 = N111 | N105;
  assign N116 = N103 | instr_i[6];
  assign N117 = N116 | instr_i[5];
  assign N118 = N116 | N105;
  assign N119 = N103 | N104;
  assign N120 = N119 | instr_i[5];
  assign N121 = instr_i[12] & instr_i[6];
  assign N122 = N121 & instr_i[5];
  assign N243 = instr_i[0] & instr_i[1];
  assign is_compressed_o = ~N243;
  assign N245 = ~instr_i[8];
  assign N246 = instr_i[10] | instr_i[11];
  assign N247 = instr_i[9] | N246;
  assign N248 = N245 | N247;
  assign N249 = instr_i[7] | N248;
  assign N250 = ~N249;
  assign N251 = instr_i[6] | instr_i[12];
  assign N252 = instr_i[5] | N251;
  assign N253 = instr_i[4] | N252;
  assign N254 = instr_i[3] | N253;
  assign N255 = instr_i[2] | N254;
  assign N256 = ~N255;
  assign N257 = instr_i[8] | N247;
  assign N258 = instr_i[7] | N257;
  assign N259 = ~N258;
  assign N260 = instr_i[11] | instr_i[12];
  assign N261 = instr_i[10] | N260;
  assign N262 = instr_i[9] | N261;
  assign N263 = instr_i[8] | N262;
  assign N264 = instr_i[7] | N263;
  assign N265 = instr_i[6] | N264;
  assign N266 = instr_i[5] | N265;
  assign N267 = ~N266;
  assign N268 = instr_i[5] | instr_i[6];
  assign N269 = instr_i[4] | N268;
  assign N270 = instr_i[3] | N269;
  assign N271 = instr_i[2] | N270;
  assign N272 = ~instr_i[12];
  assign N100 = ~instr_i[11];
  assign N101 = instr_i[11] & N0;
  assign N0 = ~instr_i[10];
  assign N102 = instr_i[11] & N1;
  assign N1 = ~N101;
  assign { N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40 } = (N2)? { instr_i[10:7], instr_i[11:11], instr_i[5:5], instr_i[6:6], 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, instr_i[4:2], 1'b0, 1'b1 } : 
                                                                                                                  (N3)? { 1'b0, 1'b0, 1'b0, instr_i[5:5], instr_i[11:10], instr_i[6:6], 1'b0, 1'b0, instr_i[9:7], 1'b1, 1'b0, 1'b1, instr_i[4:2], 1'b0, 1'b0 } : 
                                                                                                                  (N4)? { 1'b0, 1'b0, 1'b0, instr_i[5:5], 1'b0, 1'b1, instr_i[4:2], instr_i[9:7], 1'b1, instr_i[11:10], instr_i[6:6], 1'b0, 1'b0, 1'b1, 1'b0 } : 1'b0;
  assign N2 = N34;
  assign N3 = N36;
  assign N4 = N37;
  assign N60 = (N2)? N267 : 
               (N3)? 1'b0 : 
               (N4)? 1'b0 : 
               (N5)? 1'b1 : 1'b0;
  assign N5 = N39;
  assign N61 = (N6)? N60 : 
               (N7)? 1'b1 : 1'b0;
  assign N6 = N32;
  assign N7 = instr_i[13];
  assign { N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84 } = (N8)? { instr_i[4:3], instr_i[5:5], instr_i[2:2], instr_i[6:6], 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                                                                              (N9)? { instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[6:2], instr_i[11:7] } : 1'b0;
  assign N8 = N250;
  assign N9 = N249;
  assign { N127, N126, N125, N124 } = (N10)? { 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                      (N110)? { 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                      (N113)? { 1'b0, 1'b1, 1'b1, 1'b0 } : 
                                      (N115)? { 1'b0, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N10 = N107;
  assign N128 = (N10)? 1'b0 : 
                (N110)? 1'b0 : 
                (N113)? 1'b0 : 
                (N115)? 1'b0 : 
                (N123)? 1'b1 : 1'b0;
  assign { N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129 } = (N11)? { 1'b0, instr_i[10:10], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, instr_i[6:5], 1'b1, 1'b0, 1'b1, 1'b0 } : 
                                                                                            (N12)? { instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[6:5], 1'b1, 1'b1, 1'b1, 1'b0 } : 
                                                                                            (N13)? { 1'b0, N127, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, N126, N125, N124, 1'b1 } : 1'b0;
  assign N11 = N100;
  assign N12 = N101;
  assign N13 = N102;
  assign N142 = (N11)? instr_i[12] : 
                (N12)? 1'b0 : 
                (N13)? N128 : 1'b0;
  assign { N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143 } = (N14)? { instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[6:2], instr_i[11:7], 1'b0, 1'b0, 1'b0, instr_i[11:7], 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                                                                                                                                                                                  (N71)? { instr_i[12:12], instr_i[8:8], instr_i[10:9], instr_i[6:6], instr_i[7:7], instr_i[2:2], instr_i[11:11], instr_i[5:3], instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[12:12], 1'b0, 1'b0, 1'b0, 1'b0, N83, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                                                                                                                                                                                                  (N74)? { instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[6:2], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, instr_i[11:7], 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                                                                                                                                                                                  (N76)? { instr_i[12:12], instr_i[12:12], instr_i[12:12], N99, N98, N97, N96, N95, N94, N94, N94, N94, N94, N94, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, 1'b0, N249, 1'b1, 1'b0, N249 } : 
                                                                                                                                                                                                  (N78)? { N141, N140, N139, N138, N137, N136, N135, N134, N133, instr_i[4:2], 1'b0, 1'b1, instr_i[9:7], N132, N131, N130, 1'b0, 1'b1, instr_i[9:7], 1'b0, N129, 1'b1, 1'b0, 1'b0 } : 
                                                                                                                                                                                                  (N82)? { instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[12:12], instr_i[6:5], instr_i[2:2], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, instr_i[9:7], 1'b0, 1'b0, instr_i[13:13], instr_i[11:10], instr_i[4:3], instr_i[12:12], 1'b1, 1'b1, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N14 = N66;
  assign N173 = (N14)? 1'b0 : 
                (N71)? 1'b0 : 
                (N74)? 1'b0 : 
                (N76)? N256 : 
                (N78)? N142 : 
                (N82)? 1'b0 : 1'b0;
  assign N179 = ~N271;
  assign { N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180 } = (N15)? { instr_i[6:2], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, instr_i[11:7] } : 
                                                                                                        (N178)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, instr_i[11:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N15 = N271;
  assign N195 = (N15)? 1'b0 : 
                (N178)? N259 : 1'b0;
  assign N196 = (N16)? N195 : 
                (N17)? 1'b0 : 
                (N18)? 1'b0 : 
                (N18)? 1'b0 : 1'b0;
  assign N16 = N272;
  assign N17 = instr_i[12];
  assign N18 = 1'b0;
  assign { N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197 } = (N16)? { N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N271, N179 } : 
                                                                                                                          (N240)? { instr_i[6:2], instr_i[11:7], instr_i[11:7], 1'b0, 1'b1, 1'b0 } : 
                                                                                                                          (N242)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                                                                                                                          (N177)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, instr_i[11:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1 } : 1'b0;
  assign { N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215 } = (N14)? { 1'b0, 1'b0, 1'b0, instr_i[6:2], instr_i[11:7], 1'b0, 1'b1, instr_i[11:7], 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                                                                                                                                              (N74)? { instr_i[3:2], instr_i[12:12], instr_i[6:4], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, instr_i[11:7], 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                              (N78)? { 1'b0, 1'b0, 1'b0, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, 1'b0, 1'b0, N204, N203, N202, N201, N200, N199, 1'b1, N198, N197 } : 
                                                                                                                                                              (N19)? { instr_i[8:7], instr_i[12:12], instr_i[6:2], 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, instr_i[11:9], 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 1'b0;
  assign N19 = N275;
  assign N239 = (N14)? instr_i[12] : 
                (N74)? N259 : 
                (N78)? N196 : 
                (N19)? 1'b0 : 
                (N174)? 1'b1 : 1'b0;
  assign illegal_instr_o = (N20)? N61 : 
                           (N21)? N173 : 
                           (N22)? N239 : 
                           (N23)? 1'b0 : 1'b0;
  assign N20 = N26;
  assign N21 = N28;
  assign N22 = N30;
  assign N23 = N31;
  assign instr_o = (N20)? { 1'b0, 1'b0, N59, N58, N57, N56, instr_i[12:12], N55, N54, N53, N52, N51, 1'b0, N47, N50, N49, N48, 1'b0, N47, 1'b0, N46, N45, N44, N43, N42, 1'b0, N41, N40, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                   (N21)? { N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, 1'b1, 1'b1 } : 
                   (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, 1'b0, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, 1'b0, N215, 1'b1, 1'b1 } : 
                   (N23)? instr_i : 1'b0;
  assign N24 = ~instr_i[1];
  assign N25 = ~instr_i[0];
  assign N28 = ~N27;
  assign N30 = ~N29;
  assign N32 = ~instr_i[13];
  assign N33 = ~instr_i[14];
  assign N36 = ~N35;
  assign N39 = ~N38;
  assign N62 = ~instr_i[15];
  assign N63 = ~instr_i[14];
  assign N64 = ~instr_i[13];
  assign N71 = N273 | N274;
  assign N273 = ~N68;
  assign N274 = ~N70;
  assign N74 = ~N73;
  assign N76 = ~N75;
  assign N78 = ~N77;
  assign N82 = N275 | N81;
  assign N275 = ~N80;
  assign N83 = ~instr_i[15];
  assign N103 = ~instr_i[12];
  assign N104 = ~instr_i[6];
  assign N105 = ~instr_i[5];
  assign N110 = ~N109;
  assign N113 = ~N112;
  assign N115 = ~N114;
  assign N123 = N280 | N122;
  assign N280 = N278 | N279;
  assign N278 = N276 | N277;
  assign N276 = ~N117;
  assign N277 = ~N118;
  assign N279 = ~N120;
  assign N174 = N282 | N81;
  assign N282 = N281 | N274;
  assign N281 = N273 | N76;
  assign N175 = N271 | N272;
  assign N176 = N259 | N175;
  assign N177 = ~N176;
  assign N178 = ~N271;
  assign N240 = N271 & instr_i[12];
  assign N241 = instr_i[12] & N178;
  assign N242 = N259 & N241;

endmodule



module ibex_if_stage_1a110800_1a110808
(
  clk_i,
  rst_ni,
  boot_addr_i,
  req_i,
  instr_req_o,
  instr_addr_o,
  instr_gnt_i,
  instr_rvalid_i,
  instr_rdata_i,
  instr_valid_id_o,
  instr_new_id_o,
  instr_rdata_id_o,
  instr_rdata_c_id_o,
  instr_is_compressed_id_o,
  illegal_c_insn_id_o,
  pc_if_o,
  pc_id_o,
  instr_valid_clear_i,
  pc_set_i,
  csr_mepc_i,
  csr_depc_i,
  pc_mux_i,
  exc_pc_mux_i,
  exc_cause,
  jump_target_ex_i,
  csr_mtvec_o,
  id_in_ready_i,
  if_busy_o,
  perf_imiss_o
);

  input [31:0] boot_addr_i;
  output [31:0] instr_addr_o;
  input [31:0] instr_rdata_i;
  output [31:0] instr_rdata_id_o;
  output [15:0] instr_rdata_c_id_o;
  output [31:0] pc_if_o;
  output [31:0] pc_id_o;
  input [31:0] csr_mepc_i;
  input [31:0] csr_depc_i;
  input [2:0] pc_mux_i;
  input [1:0] exc_pc_mux_i;
  input [5:0] exc_cause;
  input [31:0] jump_target_ex_i;
  output [31:0] csr_mtvec_o;
  input clk_i;
  input rst_ni;
  input req_i;
  input instr_gnt_i;
  input instr_rvalid_i;
  input instr_valid_clear_i;
  input pc_set_i;
  input id_in_ready_i;
  output instr_req_o;
  output instr_valid_id_o;
  output instr_new_id_o;
  output instr_is_compressed_id_o;
  output illegal_c_insn_id_o;
  output if_busy_o;
  output perf_imiss_o;
  wire [31:0] instr_addr_o,pc_if_o,csr_mtvec_o,fetch_rdata,instr_decompressed;
  wire instr_req_o,if_busy_o,perf_imiss_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,
  N13,N14,N15,N16,N17,N18,exc_pc_6,exc_pc_5,exc_pc_4,exc_pc_3,exc_pc_2,N19,N20,N21,
  N22,N23,N24,N25,branch_req,fetch_ready,fetch_valid,N26,offset_in_init_d,
  have_instr,N27,N28,N29,N30,if_id_pipe_reg_we,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  instr_is_compressed_int,illegal_c_insn,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51;
  wire [31:8] exc_pc;
  wire [31:1] fetch_addr_n;
  reg offset_in_init_q,illegal_c_insn_id_o,instr_new_id_o,instr_valid_id_o,
  instr_is_compressed_id_o;
  reg [31:0] pc_id_o,instr_rdata_id_o;
  reg [15:0] instr_rdata_c_id_o;
  assign csr_mtvec_o[0] = 1'b1;
  assign csr_mtvec_o[1] = 1'b0;
  assign csr_mtvec_o[2] = 1'b0;
  assign csr_mtvec_o[3] = 1'b0;
  assign csr_mtvec_o[4] = 1'b0;
  assign csr_mtvec_o[5] = 1'b0;
  assign csr_mtvec_o[6] = 1'b0;
  assign csr_mtvec_o[7] = 1'b0;
  assign csr_mtvec_o[31] = boot_addr_i[31];
  assign csr_mtvec_o[30] = boot_addr_i[30];
  assign csr_mtvec_o[29] = boot_addr_i[29];
  assign csr_mtvec_o[28] = boot_addr_i[28];
  assign csr_mtvec_o[27] = boot_addr_i[27];
  assign csr_mtvec_o[26] = boot_addr_i[26];
  assign csr_mtvec_o[25] = boot_addr_i[25];
  assign csr_mtvec_o[24] = boot_addr_i[24];
  assign csr_mtvec_o[23] = boot_addr_i[23];
  assign csr_mtvec_o[22] = boot_addr_i[22];
  assign csr_mtvec_o[21] = boot_addr_i[21];
  assign csr_mtvec_o[20] = boot_addr_i[20];
  assign csr_mtvec_o[19] = boot_addr_i[19];
  assign csr_mtvec_o[18] = boot_addr_i[18];
  assign csr_mtvec_o[17] = boot_addr_i[17];
  assign csr_mtvec_o[16] = boot_addr_i[16];
  assign csr_mtvec_o[15] = boot_addr_i[15];
  assign csr_mtvec_o[14] = boot_addr_i[14];
  assign csr_mtvec_o[13] = boot_addr_i[13];
  assign csr_mtvec_o[12] = boot_addr_i[12];
  assign csr_mtvec_o[11] = boot_addr_i[11];
  assign csr_mtvec_o[10] = boot_addr_i[10];
  assign csr_mtvec_o[9] = boot_addr_i[9];
  assign csr_mtvec_o[8] = boot_addr_i[8];
  assign N13 = N11 & N12;
  assign N14 = exc_pc_mux_i[1] | N12;
  assign N16 = N11 | exc_pc_mux_i[0];
  assign N18 = exc_pc_mux_i[1] & exc_pc_mux_i[0];
  assign N21 = ~pc_mux_i[2];

  ibex_prefetch_buffer
  prefetch_buffer_i
  (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .req_i(req_i),
    .branch_i(branch_req),
    .addr_i({ fetch_addr_n, 1'b0 }),
    .ready_i(fetch_ready),
    .valid_o(fetch_valid),
    .rdata_o(fetch_rdata),
    .addr_o(pc_if_o),
    .instr_req_o(instr_req_o),
    .instr_gnt_i(instr_gnt_i),
    .instr_addr_o(instr_addr_o),
    .instr_rdata_i(instr_rdata_i),
    .instr_rvalid_i(instr_rvalid_i),
    .busy_o(if_busy_o)
  );


  always @(posedge clk_i or posedge N26) begin
    if(N26) begin
      offset_in_init_q <= 1'b1;
    end else if(N49) begin
      offset_in_init_q <= offset_in_init_d;
    end 
  end


  ibex_compressed_decoder
  compressed_decoder_i
  (
    .instr_i(fetch_rdata),
    .instr_o(instr_decompressed),
    .is_compressed_o(instr_is_compressed_int),
    .illegal_instr_o(illegal_c_insn)
  );


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      illegal_c_insn_id_o <= 1'b0;
    end else if(N44) begin
      illegal_c_insn_id_o <= illegal_c_insn;
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[31] <= 1'b0;
    end else if(N44) begin
      pc_id_o[31] <= pc_if_o[31];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[30] <= 1'b0;
    end else if(N44) begin
      pc_id_o[30] <= pc_if_o[30];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[29] <= 1'b0;
    end else if(N44) begin
      pc_id_o[29] <= pc_if_o[29];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[28] <= 1'b0;
    end else if(N44) begin
      pc_id_o[28] <= pc_if_o[28];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[27] <= 1'b0;
    end else if(N44) begin
      pc_id_o[27] <= pc_if_o[27];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[26] <= 1'b0;
    end else if(N44) begin
      pc_id_o[26] <= pc_if_o[26];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[25] <= 1'b0;
    end else if(N44) begin
      pc_id_o[25] <= pc_if_o[25];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[24] <= 1'b0;
    end else if(N44) begin
      pc_id_o[24] <= pc_if_o[24];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[23] <= 1'b0;
    end else if(N44) begin
      pc_id_o[23] <= pc_if_o[23];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[22] <= 1'b0;
    end else if(N44) begin
      pc_id_o[22] <= pc_if_o[22];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[21] <= 1'b0;
    end else if(N44) begin
      pc_id_o[21] <= pc_if_o[21];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[20] <= 1'b0;
    end else if(N44) begin
      pc_id_o[20] <= pc_if_o[20];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[19] <= 1'b0;
    end else if(N44) begin
      pc_id_o[19] <= pc_if_o[19];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[18] <= 1'b0;
    end else if(N44) begin
      pc_id_o[18] <= pc_if_o[18];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[17] <= 1'b0;
    end else if(N44) begin
      pc_id_o[17] <= pc_if_o[17];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[16] <= 1'b0;
    end else if(N44) begin
      pc_id_o[16] <= pc_if_o[16];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[15] <= 1'b0;
    end else if(N44) begin
      pc_id_o[15] <= pc_if_o[15];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[14] <= 1'b0;
    end else if(N44) begin
      pc_id_o[14] <= pc_if_o[14];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[13] <= 1'b0;
    end else if(N44) begin
      pc_id_o[13] <= pc_if_o[13];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[12] <= 1'b0;
    end else if(N44) begin
      pc_id_o[12] <= pc_if_o[12];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[11] <= 1'b0;
    end else if(N44) begin
      pc_id_o[11] <= pc_if_o[11];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[10] <= 1'b0;
    end else if(N44) begin
      pc_id_o[10] <= pc_if_o[10];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[9] <= 1'b0;
    end else if(N44) begin
      pc_id_o[9] <= pc_if_o[9];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[8] <= 1'b0;
    end else if(N44) begin
      pc_id_o[8] <= pc_if_o[8];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[7] <= 1'b0;
    end else if(N44) begin
      pc_id_o[7] <= pc_if_o[7];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[6] <= 1'b0;
    end else if(N44) begin
      pc_id_o[6] <= pc_if_o[6];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[5] <= 1'b0;
    end else if(N44) begin
      pc_id_o[5] <= pc_if_o[5];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[4] <= 1'b0;
    end else if(N44) begin
      pc_id_o[4] <= pc_if_o[4];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[3] <= 1'b0;
    end else if(N44) begin
      pc_id_o[3] <= pc_if_o[3];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[2] <= 1'b0;
    end else if(N44) begin
      pc_id_o[2] <= pc_if_o[2];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[1] <= 1'b0;
    end else if(N44) begin
      pc_id_o[1] <= pc_if_o[1];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      pc_id_o[0] <= 1'b0;
    end else if(N44) begin
      pc_id_o[0] <= pc_if_o[0];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_new_id_o <= 1'b0;
    end else if(1'b1) begin
      instr_new_id_o <= if_id_pipe_reg_we;
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_valid_id_o <= 1'b0;
    end else if(N43) begin
      instr_valid_id_o <= if_id_pipe_reg_we;
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[31] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[31] <= instr_decompressed[31];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[30] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[30] <= instr_decompressed[30];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[29] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[29] <= instr_decompressed[29];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[28] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[28] <= instr_decompressed[28];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[27] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[27] <= instr_decompressed[27];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[26] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[26] <= instr_decompressed[26];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[25] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[25] <= instr_decompressed[25];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[24] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[24] <= instr_decompressed[24];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[23] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[23] <= instr_decompressed[23];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[22] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[22] <= instr_decompressed[22];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[21] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[21] <= instr_decompressed[21];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[20] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[20] <= instr_decompressed[20];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[19] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[19] <= instr_decompressed[19];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[18] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[18] <= instr_decompressed[18];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[17] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[17] <= instr_decompressed[17];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[16] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[16] <= instr_decompressed[16];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[15] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[15] <= instr_decompressed[15];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[14] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[14] <= instr_decompressed[14];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[13] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[13] <= instr_decompressed[13];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[12] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[12] <= instr_decompressed[12];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[11] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[11] <= instr_decompressed[11];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[10] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[10] <= instr_decompressed[10];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[9] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[9] <= instr_decompressed[9];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[8] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[8] <= instr_decompressed[8];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[7] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[7] <= instr_decompressed[7];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[6] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[6] <= instr_decompressed[6];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[5] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[5] <= instr_decompressed[5];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[4] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[4] <= instr_decompressed[4];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[3] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[3] <= instr_decompressed[3];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[2] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[2] <= instr_decompressed[2];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[1] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[1] <= instr_decompressed[1];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_id_o[0] <= 1'b0;
    end else if(N44) begin
      instr_rdata_id_o[0] <= instr_decompressed[0];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_c_id_o[15] <= 1'b0;
    end else if(N44) begin
      instr_rdata_c_id_o[15] <= fetch_rdata[15];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_c_id_o[14] <= 1'b0;
    end else if(N44) begin
      instr_rdata_c_id_o[14] <= fetch_rdata[14];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_c_id_o[13] <= 1'b0;
    end else if(N44) begin
      instr_rdata_c_id_o[13] <= fetch_rdata[13];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_c_id_o[12] <= 1'b0;
    end else if(N44) begin
      instr_rdata_c_id_o[12] <= fetch_rdata[12];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_c_id_o[11] <= 1'b0;
    end else if(N44) begin
      instr_rdata_c_id_o[11] <= fetch_rdata[11];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_c_id_o[10] <= 1'b0;
    end else if(N44) begin
      instr_rdata_c_id_o[10] <= fetch_rdata[10];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_c_id_o[9] <= 1'b0;
    end else if(N44) begin
      instr_rdata_c_id_o[9] <= fetch_rdata[9];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_c_id_o[8] <= 1'b0;
    end else if(N44) begin
      instr_rdata_c_id_o[8] <= fetch_rdata[8];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_c_id_o[7] <= 1'b0;
    end else if(N44) begin
      instr_rdata_c_id_o[7] <= fetch_rdata[7];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_c_id_o[6] <= 1'b0;
    end else if(N44) begin
      instr_rdata_c_id_o[6] <= fetch_rdata[6];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_c_id_o[5] <= 1'b0;
    end else if(N44) begin
      instr_rdata_c_id_o[5] <= fetch_rdata[5];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_c_id_o[4] <= 1'b0;
    end else if(N44) begin
      instr_rdata_c_id_o[4] <= fetch_rdata[4];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_c_id_o[3] <= 1'b0;
    end else if(N44) begin
      instr_rdata_c_id_o[3] <= fetch_rdata[3];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_c_id_o[2] <= 1'b0;
    end else if(N44) begin
      instr_rdata_c_id_o[2] <= fetch_rdata[2];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_c_id_o[1] <= 1'b0;
    end else if(N44) begin
      instr_rdata_c_id_o[1] <= fetch_rdata[1];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_rdata_c_id_o[0] <= 1'b0;
    end else if(N44) begin
      instr_rdata_c_id_o[0] <= fetch_rdata[0];
    end 
  end


  always @(posedge clk_i or posedge N40) begin
    if(N40) begin
      instr_is_compressed_id_o <= 1'b0;
    end else if(N44) begin
      instr_is_compressed_id_o <= instr_is_compressed_int;
    end 
  end

  assign { exc_pc, exc_pc_6, exc_pc_5, exc_pc_4, exc_pc_3, exc_pc_2 } = (N0)? { boot_addr_i[31:8], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                        (N1)? { boot_addr_i[31:8], exc_cause[4:0] } : 
                                                                        (N2)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                        (N3)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 1'b0;
  assign N0 = N13;
  assign N1 = N15;
  assign N2 = N17;
  assign N3 = N18;
  assign fetch_addr_n = (N22)? { boot_addr_i[31:8], 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                        (N23)? jump_target_ex_i[31:1] : 
                        (N24)? { exc_pc, 1'b0, exc_pc_6, exc_pc_5, exc_pc_4, exc_pc_3, exc_pc_2, 1'b0 } : 
                        (N25)? csr_mepc_i[31:1] : 
                        (N4)? csr_depc_i[31:1] : 1'b0;
  assign N4 = pc_mux_i[2];
  assign N33 = (N5)? 1'b0 : 
               (N32)? offset_in_init_q : 1'b0;
  assign N5 = N31;
  assign N34 = (N6)? 1'b0 : 
               (N39)? N33 : 
               (N28)? offset_in_init_q : 1'b0;
  assign N6 = offset_in_init_q;
  assign N36 = (N6)? N30 : 
               (N35)? 1'b0 : 
               (N7)? 1'b0 : 1'b0;
  assign N7 = 1'b0;
  assign N37 = (N6)? 1'b0 : 
               (N39)? 1'b1 : 
               (N28)? 1'b0 : 1'b0;
  assign fetch_ready = (N6)? 1'b0 : 
                       (N39)? N31 : 
                       (N28)? 1'b0 : 1'b0;
  assign have_instr = (N8)? 1'b0 : 
                      (N9)? N37 : 1'b0;
  assign N8 = pc_set_i;
  assign N9 = N38;
  assign branch_req = (N8)? 1'b1 : 
                      (N9)? N36 : 1'b0;
  assign offset_in_init_d = (N8)? 1'b0 : 
                            (N9)? N34 : 1'b0;
  assign N43 = (N10)? 1'b1 : 
               (N46)? 1'b1 : 
               (N42)? 1'b0 : 1'b0;
  assign N10 = if_id_pipe_reg_we;
  assign N44 = (N10)? 1'b1 : 
               (N46)? 1'b0 : 
               (N42)? 1'b0 : 1'b0;
  assign N11 = ~exc_pc_mux_i[1];
  assign N12 = ~exc_pc_mux_i[0];
  assign N15 = ~N14;
  assign N17 = ~N16;
  assign N19 = ~pc_mux_i[1];
  assign N20 = ~pc_mux_i[0];
  assign N22 = N50 & N20;
  assign N50 = N21 & N19;
  assign N23 = N19 & pc_mux_i[0];
  assign N24 = pc_mux_i[1] & N20;
  assign N25 = pc_mux_i[1] & pc_mux_i[0];
  assign N26 = ~rst_ni;
  assign N27 = fetch_valid | offset_in_init_q;
  assign N28 = ~N27;
  assign N29 = ~req_i;
  assign N30 = req_i;
  assign N31 = req_i & if_id_pipe_reg_we;
  assign N32 = ~N31;
  assign N35 = ~offset_in_init_q;
  assign N38 = ~pc_set_i;
  assign N39 = fetch_valid & N35;
  assign perf_imiss_o = N51 | branch_req;
  assign N51 = ~fetch_valid;
  assign if_id_pipe_reg_we = have_instr & id_in_ready_i;
  assign N40 = ~rst_ni;
  assign N41 = instr_valid_clear_i | if_id_pipe_reg_we;
  assign N42 = ~N41;
  assign N45 = ~if_id_pipe_reg_we;
  assign N46 = instr_valid_clear_i & N45;
  assign N47 = offset_in_init_q & N38;
  assign N48 = N29 & N47;
  assign N49 = ~N48;

endmodule



module ibex_register_file_0
(
  clk_i,
  rst_ni,
  test_en_i,
  raddr_a_i,
  rdata_a_o,
  raddr_b_i,
  rdata_b_o,
  waddr_a_i,
  wdata_a_i,
  we_a_i
);

  input [4:0] raddr_a_i;
  output [31:0] rdata_a_o;
  input [4:0] raddr_b_i;
  output [31:0] rdata_b_o;
  input [4:0] waddr_a_i;
  input [31:0] wdata_a_i;
  input clk_i;
  input rst_ni;
  input test_en_i;
  input we_a_i;
  wire [31:0] rdata_a_o,rdata_b_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289;
  wire [31:1] we_a_dec;
  reg [991:0] rf_reg_tmp;

  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[991] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[991] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[990] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[990] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[989] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[989] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[988] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[988] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[987] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[987] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[986] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[986] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[985] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[985] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[984] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[984] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[983] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[983] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[982] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[982] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[981] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[981] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[980] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[980] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[979] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[979] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[978] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[978] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[977] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[977] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[976] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[976] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[975] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[975] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[974] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[974] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[973] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[973] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[972] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[972] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[971] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[971] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[970] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[970] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[969] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[969] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[968] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[968] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[967] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[967] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[966] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[966] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[965] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[965] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[964] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[964] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[963] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[963] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[962] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[962] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[961] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[961] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[960] <= 1'b0;
    end else if(we_a_dec[31]) begin
      rf_reg_tmp[960] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[959] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[959] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[958] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[958] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[957] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[957] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[956] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[956] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[955] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[955] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[954] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[954] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[953] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[953] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[952] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[952] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[951] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[951] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[950] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[950] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[949] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[949] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[948] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[948] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[947] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[947] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[946] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[946] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[945] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[945] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[944] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[944] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[943] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[943] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[942] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[942] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[941] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[941] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[940] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[940] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[939] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[939] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[938] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[938] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[937] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[937] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[936] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[936] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[935] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[935] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[934] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[934] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[933] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[933] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[932] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[932] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[931] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[931] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[930] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[930] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[929] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[929] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[928] <= 1'b0;
    end else if(we_a_dec[30]) begin
      rf_reg_tmp[928] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[927] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[927] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[926] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[926] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[925] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[925] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[924] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[924] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[923] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[923] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[922] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[922] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[921] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[921] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[920] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[920] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[919] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[919] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[918] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[918] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[917] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[917] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[916] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[916] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[915] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[915] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[914] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[914] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[913] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[913] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[912] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[912] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[911] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[911] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[910] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[910] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[909] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[909] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[908] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[908] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[907] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[907] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[906] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[906] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[905] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[905] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[904] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[904] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[903] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[903] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[902] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[902] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[901] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[901] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[900] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[900] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[899] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[899] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[898] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[898] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[897] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[897] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[896] <= 1'b0;
    end else if(we_a_dec[29]) begin
      rf_reg_tmp[896] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[895] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[895] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[894] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[894] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[893] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[893] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[892] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[892] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[891] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[891] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[890] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[890] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[889] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[889] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[888] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[888] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[887] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[887] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[886] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[886] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[885] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[885] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[884] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[884] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[883] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[883] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[882] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[882] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[881] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[881] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[880] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[880] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[879] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[879] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[878] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[878] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[877] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[877] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[876] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[876] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[875] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[875] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[874] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[874] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[873] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[873] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[872] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[872] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[871] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[871] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[870] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[870] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[869] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[869] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[868] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[868] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[867] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[867] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[866] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[866] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[865] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[865] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[864] <= 1'b0;
    end else if(we_a_dec[28]) begin
      rf_reg_tmp[864] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[863] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[863] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[862] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[862] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[861] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[861] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[860] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[860] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[859] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[859] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[858] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[858] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[857] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[857] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[856] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[856] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[855] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[855] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[854] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[854] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[853] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[853] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[852] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[852] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[851] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[851] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[850] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[850] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[849] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[849] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[848] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[848] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[847] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[847] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[846] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[846] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[845] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[845] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[844] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[844] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[843] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[843] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[842] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[842] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[841] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[841] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[840] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[840] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[839] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[839] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[838] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[838] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[837] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[837] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[836] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[836] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[835] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[835] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[834] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[834] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[833] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[833] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[832] <= 1'b0;
    end else if(we_a_dec[27]) begin
      rf_reg_tmp[832] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[831] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[831] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[830] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[830] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[829] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[829] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[828] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[828] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[827] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[827] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[826] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[826] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[825] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[825] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[824] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[824] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[823] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[823] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[822] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[822] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[821] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[821] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[820] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[820] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[819] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[819] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[818] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[818] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[817] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[817] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[816] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[816] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[815] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[815] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[814] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[814] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[813] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[813] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[812] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[812] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[811] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[811] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[810] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[810] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[809] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[809] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[808] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[808] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[807] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[807] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[806] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[806] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[805] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[805] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[804] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[804] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[803] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[803] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[802] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[802] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[801] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[801] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[800] <= 1'b0;
    end else if(we_a_dec[26]) begin
      rf_reg_tmp[800] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[799] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[799] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[798] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[798] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[797] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[797] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[796] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[796] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[795] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[795] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[794] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[794] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[793] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[793] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[792] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[792] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[791] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[791] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[790] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[790] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[789] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[789] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[788] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[788] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[787] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[787] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[786] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[786] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[785] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[785] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[784] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[784] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[783] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[783] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[782] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[782] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[781] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[781] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[780] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[780] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[779] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[779] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[778] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[778] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[777] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[777] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[776] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[776] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[775] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[775] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[774] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[774] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[773] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[773] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[772] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[772] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[771] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[771] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[770] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[770] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[769] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[769] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[768] <= 1'b0;
    end else if(we_a_dec[25]) begin
      rf_reg_tmp[768] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[767] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[767] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[766] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[766] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[765] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[765] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[764] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[764] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[763] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[763] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[762] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[762] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[761] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[761] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[760] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[760] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[759] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[759] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[758] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[758] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[757] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[757] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[756] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[756] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[755] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[755] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[754] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[754] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[753] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[753] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[752] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[752] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[751] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[751] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[750] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[750] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[749] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[749] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[748] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[748] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[747] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[747] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[746] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[746] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[745] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[745] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[744] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[744] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[743] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[743] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[742] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[742] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[741] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[741] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[740] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[740] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[739] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[739] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[738] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[738] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[737] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[737] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[736] <= 1'b0;
    end else if(we_a_dec[24]) begin
      rf_reg_tmp[736] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[735] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[735] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[734] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[734] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[733] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[733] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[732] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[732] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[731] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[731] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[730] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[730] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[729] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[729] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[728] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[728] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[727] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[727] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[726] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[726] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[725] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[725] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[724] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[724] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[723] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[723] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[722] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[722] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[721] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[721] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[720] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[720] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[719] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[719] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[718] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[718] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[717] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[717] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[716] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[716] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[715] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[715] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[714] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[714] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[713] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[713] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[712] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[712] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[711] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[711] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[710] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[710] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[709] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[709] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[708] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[708] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[707] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[707] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[706] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[706] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[705] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[705] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[704] <= 1'b0;
    end else if(we_a_dec[23]) begin
      rf_reg_tmp[704] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[703] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[703] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[702] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[702] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[701] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[701] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[700] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[700] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[699] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[699] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[698] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[698] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[697] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[697] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[696] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[696] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[695] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[695] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[694] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[694] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[693] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[693] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[692] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[692] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[691] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[691] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[690] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[690] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[689] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[689] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[688] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[688] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[687] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[687] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[686] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[686] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[685] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[685] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[684] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[684] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[683] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[683] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[682] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[682] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[681] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[681] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[680] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[680] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[679] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[679] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[678] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[678] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[677] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[677] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[676] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[676] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[675] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[675] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[674] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[674] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[673] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[673] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[672] <= 1'b0;
    end else if(we_a_dec[22]) begin
      rf_reg_tmp[672] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[671] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[671] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[670] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[670] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[669] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[669] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[668] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[668] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[667] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[667] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[666] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[666] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[665] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[665] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[664] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[664] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[663] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[663] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[662] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[662] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[661] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[661] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[660] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[660] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[659] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[659] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[658] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[658] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[657] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[657] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[656] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[656] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[655] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[655] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[654] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[654] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[653] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[653] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[652] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[652] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[651] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[651] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[650] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[650] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[649] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[649] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[648] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[648] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[647] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[647] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[646] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[646] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[645] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[645] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[644] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[644] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[643] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[643] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[642] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[642] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[641] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[641] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[640] <= 1'b0;
    end else if(we_a_dec[21]) begin
      rf_reg_tmp[640] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[639] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[639] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[638] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[638] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[637] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[637] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[636] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[636] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[635] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[635] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[634] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[634] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[633] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[633] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[632] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[632] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[631] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[631] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[630] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[630] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[629] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[629] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[628] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[628] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[627] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[627] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[626] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[626] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[625] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[625] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[624] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[624] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[623] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[623] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[622] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[622] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[621] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[621] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[620] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[620] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[619] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[619] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[618] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[618] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[617] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[617] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[616] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[616] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[615] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[615] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[614] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[614] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[613] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[613] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[612] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[612] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[611] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[611] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[610] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[610] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[609] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[609] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[608] <= 1'b0;
    end else if(we_a_dec[20]) begin
      rf_reg_tmp[608] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[607] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[607] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[606] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[606] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[605] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[605] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[604] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[604] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[603] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[603] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[602] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[602] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[601] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[601] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[600] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[600] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[599] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[599] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[598] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[598] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[597] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[597] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[596] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[596] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[595] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[595] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[594] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[594] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[593] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[593] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[592] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[592] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[591] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[591] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[590] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[590] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[589] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[589] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[588] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[588] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[587] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[587] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[586] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[586] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[585] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[585] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[584] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[584] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[583] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[583] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[582] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[582] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[581] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[581] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[580] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[580] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[579] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[579] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[578] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[578] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[577] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[577] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[576] <= 1'b0;
    end else if(we_a_dec[19]) begin
      rf_reg_tmp[576] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[575] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[575] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[574] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[574] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[573] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[573] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[572] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[572] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[571] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[571] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[570] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[570] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[569] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[569] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[568] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[568] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[567] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[567] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[566] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[566] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[565] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[565] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[564] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[564] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[563] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[563] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[562] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[562] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[561] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[561] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[560] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[560] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[559] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[559] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[558] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[558] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[557] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[557] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[556] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[556] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[555] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[555] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[554] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[554] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[553] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[553] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[552] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[552] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[551] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[551] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[550] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[550] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[549] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[549] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[548] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[548] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[547] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[547] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[546] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[546] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[545] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[545] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[544] <= 1'b0;
    end else if(we_a_dec[18]) begin
      rf_reg_tmp[544] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[543] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[543] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[542] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[542] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[541] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[541] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[540] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[540] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[539] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[539] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[538] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[538] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[537] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[537] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[536] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[536] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[535] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[535] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[534] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[534] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[533] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[533] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[532] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[532] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[531] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[531] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[530] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[530] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[529] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[529] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[528] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[528] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[527] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[527] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[526] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[526] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[525] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[525] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[524] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[524] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[523] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[523] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[522] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[522] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[521] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[521] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[520] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[520] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[519] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[519] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[518] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[518] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[517] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[517] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[516] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[516] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[515] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[515] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[514] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[514] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[513] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[513] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[512] <= 1'b0;
    end else if(we_a_dec[17]) begin
      rf_reg_tmp[512] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[511] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[511] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[510] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[510] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[509] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[509] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[508] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[508] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[507] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[507] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[506] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[506] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[505] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[505] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[504] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[504] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[503] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[503] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[502] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[502] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[501] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[501] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[500] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[500] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[499] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[499] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[498] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[498] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[497] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[497] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[496] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[496] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[495] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[495] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[494] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[494] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[493] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[493] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[492] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[492] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[491] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[491] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[490] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[490] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[489] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[489] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[488] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[488] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[487] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[487] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[486] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[486] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[485] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[485] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[484] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[484] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[483] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[483] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[482] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[482] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[481] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[481] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[480] <= 1'b0;
    end else if(we_a_dec[16]) begin
      rf_reg_tmp[480] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[479] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[479] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[478] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[478] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[477] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[477] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[476] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[476] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[475] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[475] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[474] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[474] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[473] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[473] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[472] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[472] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[471] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[471] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[470] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[470] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[469] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[469] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[468] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[468] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[467] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[467] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[466] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[466] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[465] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[465] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[464] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[464] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[463] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[463] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[462] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[462] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[461] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[461] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[460] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[460] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[459] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[459] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[458] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[458] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[457] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[457] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[456] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[456] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[455] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[455] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[454] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[454] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[453] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[453] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[452] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[452] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[451] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[451] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[450] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[450] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[449] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[449] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[448] <= 1'b0;
    end else if(we_a_dec[15]) begin
      rf_reg_tmp[448] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[447] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[447] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[446] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[446] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[445] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[445] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[444] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[444] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[443] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[443] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[442] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[442] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[441] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[441] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[440] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[440] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[439] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[439] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[438] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[438] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[437] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[437] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[436] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[436] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[435] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[435] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[434] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[434] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[433] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[433] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[432] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[432] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[431] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[431] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[430] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[430] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[429] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[429] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[428] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[428] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[427] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[427] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[426] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[426] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[425] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[425] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[424] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[424] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[423] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[423] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[422] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[422] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[421] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[421] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[420] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[420] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[419] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[419] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[418] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[418] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[417] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[417] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[416] <= 1'b0;
    end else if(we_a_dec[14]) begin
      rf_reg_tmp[416] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[415] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[415] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[414] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[414] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[413] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[413] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[412] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[412] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[411] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[411] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[410] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[410] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[409] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[409] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[408] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[408] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[407] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[407] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[406] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[406] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[405] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[405] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[404] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[404] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[403] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[403] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[402] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[402] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[401] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[401] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[400] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[400] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[399] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[399] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[398] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[398] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[397] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[397] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[396] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[396] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[395] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[395] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[394] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[394] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[393] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[393] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[392] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[392] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[391] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[391] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[390] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[390] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[389] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[389] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[388] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[388] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[387] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[387] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[386] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[386] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[385] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[385] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[384] <= 1'b0;
    end else if(we_a_dec[13]) begin
      rf_reg_tmp[384] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[383] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[383] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[382] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[382] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[381] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[381] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[380] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[380] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[379] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[379] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[378] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[378] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[377] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[377] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[376] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[376] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[375] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[375] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[374] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[374] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[373] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[373] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[372] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[372] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[371] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[371] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[370] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[370] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[369] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[369] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[368] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[368] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[367] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[367] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[366] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[366] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[365] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[365] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[364] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[364] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[363] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[363] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[362] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[362] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[361] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[361] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[360] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[360] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[359] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[359] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[358] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[358] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[357] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[357] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[356] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[356] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[355] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[355] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[354] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[354] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[353] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[353] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[352] <= 1'b0;
    end else if(we_a_dec[12]) begin
      rf_reg_tmp[352] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[351] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[351] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[350] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[350] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[349] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[349] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[348] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[348] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[347] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[347] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[346] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[346] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[345] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[345] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[344] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[344] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[343] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[343] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[342] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[342] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[341] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[341] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[340] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[340] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[339] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[339] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[338] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[338] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[337] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[337] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[336] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[336] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[335] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[335] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[334] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[334] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[333] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[333] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[332] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[332] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[331] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[331] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[330] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[330] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[329] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[329] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[328] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[328] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[327] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[327] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[326] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[326] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[325] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[325] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[324] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[324] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[323] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[323] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[322] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[322] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[321] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[321] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[320] <= 1'b0;
    end else if(we_a_dec[11]) begin
      rf_reg_tmp[320] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[319] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[319] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[318] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[318] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[317] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[317] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[316] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[316] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[315] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[315] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[314] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[314] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[313] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[313] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[312] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[312] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[311] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[311] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[310] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[310] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[309] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[309] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[308] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[308] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[307] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[307] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[306] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[306] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[305] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[305] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[304] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[304] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[303] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[303] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[302] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[302] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[301] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[301] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[300] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[300] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[299] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[299] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[298] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[298] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[297] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[297] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[296] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[296] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[295] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[295] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[294] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[294] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[293] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[293] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[292] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[292] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[291] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[291] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[290] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[290] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[289] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[289] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[288] <= 1'b0;
    end else if(we_a_dec[10]) begin
      rf_reg_tmp[288] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[287] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[287] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[286] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[286] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[285] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[285] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[284] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[284] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[283] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[283] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[282] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[282] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[281] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[281] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[280] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[280] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[279] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[279] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[278] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[278] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[277] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[277] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[276] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[276] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[275] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[275] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[274] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[274] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[273] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[273] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[272] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[272] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[271] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[271] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[270] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[270] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[269] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[269] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[268] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[268] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[267] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[267] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[266] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[266] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[265] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[265] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[264] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[264] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[263] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[263] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[262] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[262] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[261] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[261] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[260] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[260] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[259] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[259] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[258] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[258] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[257] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[257] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[256] <= 1'b0;
    end else if(we_a_dec[9]) begin
      rf_reg_tmp[256] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[255] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[255] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[254] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[254] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[253] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[253] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[252] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[252] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[251] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[251] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[250] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[250] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[249] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[249] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[248] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[248] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[247] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[247] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[246] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[246] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[245] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[245] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[244] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[244] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[243] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[243] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[242] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[242] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[241] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[241] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[240] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[240] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[239] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[239] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[238] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[238] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[237] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[237] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[236] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[236] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[235] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[235] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[234] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[234] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[233] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[233] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[232] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[232] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[231] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[231] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[230] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[230] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[229] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[229] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[228] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[228] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[227] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[227] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[226] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[226] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[225] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[225] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[224] <= 1'b0;
    end else if(we_a_dec[8]) begin
      rf_reg_tmp[224] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[223] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[223] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[222] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[222] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[221] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[221] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[220] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[220] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[219] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[219] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[218] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[218] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[217] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[217] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[216] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[216] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[215] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[215] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[214] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[214] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[213] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[213] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[212] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[212] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[211] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[211] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[210] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[210] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[209] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[209] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[208] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[208] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[207] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[207] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[206] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[206] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[205] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[205] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[204] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[204] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[203] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[203] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[202] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[202] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[201] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[201] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[200] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[200] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[199] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[199] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[198] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[198] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[197] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[197] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[196] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[196] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[195] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[195] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[194] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[194] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[193] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[193] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[192] <= 1'b0;
    end else if(we_a_dec[7]) begin
      rf_reg_tmp[192] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[191] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[191] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[190] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[190] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[189] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[189] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[188] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[188] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[187] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[187] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[186] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[186] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[185] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[185] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[184] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[184] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[183] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[183] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[182] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[182] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[181] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[181] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[180] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[180] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[179] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[179] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[178] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[178] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[177] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[177] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[176] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[176] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[175] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[175] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[174] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[174] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[173] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[173] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[172] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[172] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[171] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[171] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[170] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[170] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[169] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[169] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[168] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[168] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[167] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[167] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[166] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[166] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[165] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[165] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[164] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[164] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[163] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[163] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[162] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[162] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[161] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[161] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[160] <= 1'b0;
    end else if(we_a_dec[6]) begin
      rf_reg_tmp[160] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[159] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[159] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[158] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[158] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[157] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[157] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[156] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[156] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[155] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[155] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[154] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[154] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[153] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[153] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[152] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[152] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[151] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[151] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[150] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[150] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[149] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[149] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[148] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[148] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[147] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[147] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[146] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[146] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[145] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[145] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[144] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[144] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[143] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[143] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[142] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[142] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[141] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[141] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[140] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[140] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[139] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[139] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[138] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[138] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[137] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[137] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[136] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[136] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[135] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[135] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[134] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[134] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[133] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[133] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[132] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[132] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[131] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[131] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[130] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[130] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[129] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[129] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[128] <= 1'b0;
    end else if(we_a_dec[5]) begin
      rf_reg_tmp[128] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[127] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[127] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[126] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[126] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[125] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[125] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[124] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[124] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[123] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[123] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[122] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[122] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[121] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[121] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[120] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[120] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[119] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[119] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[118] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[118] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[117] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[117] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[116] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[116] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[115] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[115] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[114] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[114] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[113] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[113] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[112] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[112] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[111] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[111] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[110] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[110] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[109] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[109] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[108] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[108] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[107] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[107] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[106] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[106] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[105] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[105] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[104] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[104] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[103] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[103] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[102] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[102] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[101] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[101] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[100] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[100] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[99] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[99] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[98] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[98] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[97] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[97] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[96] <= 1'b0;
    end else if(we_a_dec[4]) begin
      rf_reg_tmp[96] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[95] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[95] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[94] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[94] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[93] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[93] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[92] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[92] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[91] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[91] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[90] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[90] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[89] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[89] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[88] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[88] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[87] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[87] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[86] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[86] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[85] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[85] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[84] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[84] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[83] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[83] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[82] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[82] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[81] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[81] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[80] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[80] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[79] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[79] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[78] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[78] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[77] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[77] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[76] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[76] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[75] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[75] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[74] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[74] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[73] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[73] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[72] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[72] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[71] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[71] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[70] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[70] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[69] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[69] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[68] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[68] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[67] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[67] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[66] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[66] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[65] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[65] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[64] <= 1'b0;
    end else if(we_a_dec[3]) begin
      rf_reg_tmp[64] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[63] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[63] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[62] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[62] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[61] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[61] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[60] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[60] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[59] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[59] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[58] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[58] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[57] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[57] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[56] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[56] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[55] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[55] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[54] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[54] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[53] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[53] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[52] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[52] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[51] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[51] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[50] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[50] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[49] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[49] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[48] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[48] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[47] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[47] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[46] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[46] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[45] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[45] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[44] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[44] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[43] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[43] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[42] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[42] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[41] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[41] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[40] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[40] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[39] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[39] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[38] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[38] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[37] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[37] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[36] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[36] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[35] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[35] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[34] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[34] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[33] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[33] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[32] <= 1'b0;
    end else if(we_a_dec[2]) begin
      rf_reg_tmp[32] <= wdata_a_i[0];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[31] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[31] <= wdata_a_i[31];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[30] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[30] <= wdata_a_i[30];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[29] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[29] <= wdata_a_i[29];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[28] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[28] <= wdata_a_i[28];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[27] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[27] <= wdata_a_i[27];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[26] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[26] <= wdata_a_i[26];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[25] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[25] <= wdata_a_i[25];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[24] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[24] <= wdata_a_i[24];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[23] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[23] <= wdata_a_i[23];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[22] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[22] <= wdata_a_i[22];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[21] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[21] <= wdata_a_i[21];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[20] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[20] <= wdata_a_i[20];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[19] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[19] <= wdata_a_i[19];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[18] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[18] <= wdata_a_i[18];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[17] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[17] <= wdata_a_i[17];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[16] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[16] <= wdata_a_i[16];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[15] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[15] <= wdata_a_i[15];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[14] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[14] <= wdata_a_i[14];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[13] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[13] <= wdata_a_i[13];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[12] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[12] <= wdata_a_i[12];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[11] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[11] <= wdata_a_i[11];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[10] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[10] <= wdata_a_i[10];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[9] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[9] <= wdata_a_i[9];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[8] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[8] <= wdata_a_i[8];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[7] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[7] <= wdata_a_i[7];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[6] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[6] <= wdata_a_i[6];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[5] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[5] <= wdata_a_i[5];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[4] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[4] <= wdata_a_i[4];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[3] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[3] <= wdata_a_i[3];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[2] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[2] <= wdata_a_i[2];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[1] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[1] <= wdata_a_i[1];
    end 
  end


  always @(posedge clk_i or posedge N62) begin
    if(N62) begin
      rf_reg_tmp[0] <= 1'b0;
    end else if(we_a_dec[1]) begin
      rf_reg_tmp[0] <= wdata_a_i[0];
    end 
  end

  assign rdata_a_o[31] = (N96)? 1'b0 : 
                         (N98)? rf_reg_tmp[31] : 
                         (N100)? rf_reg_tmp[63] : 
                         (N102)? rf_reg_tmp[95] : 
                         (N104)? rf_reg_tmp[127] : 
                         (N106)? rf_reg_tmp[159] : 
                         (N108)? rf_reg_tmp[191] : 
                         (N110)? rf_reg_tmp[223] : 
                         (N112)? rf_reg_tmp[255] : 
                         (N114)? rf_reg_tmp[287] : 
                         (N116)? rf_reg_tmp[319] : 
                         (N118)? rf_reg_tmp[351] : 
                         (N120)? rf_reg_tmp[383] : 
                         (N122)? rf_reg_tmp[415] : 
                         (N124)? rf_reg_tmp[447] : 
                         (N126)? rf_reg_tmp[479] : 
                         (N97)? rf_reg_tmp[511] : 
                         (N99)? rf_reg_tmp[543] : 
                         (N101)? rf_reg_tmp[575] : 
                         (N103)? rf_reg_tmp[607] : 
                         (N105)? rf_reg_tmp[639] : 
                         (N107)? rf_reg_tmp[671] : 
                         (N109)? rf_reg_tmp[703] : 
                         (N111)? rf_reg_tmp[735] : 
                         (N113)? rf_reg_tmp[767] : 
                         (N115)? rf_reg_tmp[799] : 
                         (N117)? rf_reg_tmp[831] : 
                         (N119)? rf_reg_tmp[863] : 
                         (N121)? rf_reg_tmp[895] : 
                         (N123)? rf_reg_tmp[927] : 
                         (N125)? rf_reg_tmp[959] : 
                         (N127)? rf_reg_tmp[991] : 1'b0;
  assign rdata_a_o[30] = (N96)? 1'b0 : 
                         (N98)? rf_reg_tmp[30] : 
                         (N100)? rf_reg_tmp[62] : 
                         (N102)? rf_reg_tmp[94] : 
                         (N104)? rf_reg_tmp[126] : 
                         (N106)? rf_reg_tmp[158] : 
                         (N108)? rf_reg_tmp[190] : 
                         (N110)? rf_reg_tmp[222] : 
                         (N112)? rf_reg_tmp[254] : 
                         (N114)? rf_reg_tmp[286] : 
                         (N116)? rf_reg_tmp[318] : 
                         (N118)? rf_reg_tmp[350] : 
                         (N120)? rf_reg_tmp[382] : 
                         (N122)? rf_reg_tmp[414] : 
                         (N124)? rf_reg_tmp[446] : 
                         (N126)? rf_reg_tmp[478] : 
                         (N97)? rf_reg_tmp[510] : 
                         (N99)? rf_reg_tmp[542] : 
                         (N101)? rf_reg_tmp[574] : 
                         (N103)? rf_reg_tmp[606] : 
                         (N105)? rf_reg_tmp[638] : 
                         (N107)? rf_reg_tmp[670] : 
                         (N109)? rf_reg_tmp[702] : 
                         (N111)? rf_reg_tmp[734] : 
                         (N113)? rf_reg_tmp[766] : 
                         (N115)? rf_reg_tmp[798] : 
                         (N117)? rf_reg_tmp[830] : 
                         (N119)? rf_reg_tmp[862] : 
                         (N121)? rf_reg_tmp[894] : 
                         (N123)? rf_reg_tmp[926] : 
                         (N125)? rf_reg_tmp[958] : 
                         (N127)? rf_reg_tmp[990] : 1'b0;
  assign rdata_a_o[29] = (N96)? 1'b0 : 
                         (N98)? rf_reg_tmp[29] : 
                         (N100)? rf_reg_tmp[61] : 
                         (N102)? rf_reg_tmp[93] : 
                         (N104)? rf_reg_tmp[125] : 
                         (N106)? rf_reg_tmp[157] : 
                         (N108)? rf_reg_tmp[189] : 
                         (N110)? rf_reg_tmp[221] : 
                         (N112)? rf_reg_tmp[253] : 
                         (N114)? rf_reg_tmp[285] : 
                         (N116)? rf_reg_tmp[317] : 
                         (N118)? rf_reg_tmp[349] : 
                         (N120)? rf_reg_tmp[381] : 
                         (N122)? rf_reg_tmp[413] : 
                         (N124)? rf_reg_tmp[445] : 
                         (N126)? rf_reg_tmp[477] : 
                         (N97)? rf_reg_tmp[509] : 
                         (N99)? rf_reg_tmp[541] : 
                         (N101)? rf_reg_tmp[573] : 
                         (N103)? rf_reg_tmp[605] : 
                         (N105)? rf_reg_tmp[637] : 
                         (N107)? rf_reg_tmp[669] : 
                         (N109)? rf_reg_tmp[701] : 
                         (N111)? rf_reg_tmp[733] : 
                         (N113)? rf_reg_tmp[765] : 
                         (N115)? rf_reg_tmp[797] : 
                         (N117)? rf_reg_tmp[829] : 
                         (N119)? rf_reg_tmp[861] : 
                         (N121)? rf_reg_tmp[893] : 
                         (N123)? rf_reg_tmp[925] : 
                         (N125)? rf_reg_tmp[957] : 
                         (N127)? rf_reg_tmp[989] : 1'b0;
  assign rdata_a_o[28] = (N96)? 1'b0 : 
                         (N98)? rf_reg_tmp[28] : 
                         (N100)? rf_reg_tmp[60] : 
                         (N102)? rf_reg_tmp[92] : 
                         (N104)? rf_reg_tmp[124] : 
                         (N106)? rf_reg_tmp[156] : 
                         (N108)? rf_reg_tmp[188] : 
                         (N110)? rf_reg_tmp[220] : 
                         (N112)? rf_reg_tmp[252] : 
                         (N114)? rf_reg_tmp[284] : 
                         (N116)? rf_reg_tmp[316] : 
                         (N118)? rf_reg_tmp[348] : 
                         (N120)? rf_reg_tmp[380] : 
                         (N122)? rf_reg_tmp[412] : 
                         (N124)? rf_reg_tmp[444] : 
                         (N126)? rf_reg_tmp[476] : 
                         (N97)? rf_reg_tmp[508] : 
                         (N99)? rf_reg_tmp[540] : 
                         (N101)? rf_reg_tmp[572] : 
                         (N103)? rf_reg_tmp[604] : 
                         (N105)? rf_reg_tmp[636] : 
                         (N107)? rf_reg_tmp[668] : 
                         (N109)? rf_reg_tmp[700] : 
                         (N111)? rf_reg_tmp[732] : 
                         (N113)? rf_reg_tmp[764] : 
                         (N115)? rf_reg_tmp[796] : 
                         (N117)? rf_reg_tmp[828] : 
                         (N119)? rf_reg_tmp[860] : 
                         (N121)? rf_reg_tmp[892] : 
                         (N123)? rf_reg_tmp[924] : 
                         (N125)? rf_reg_tmp[956] : 
                         (N127)? rf_reg_tmp[988] : 1'b0;
  assign rdata_a_o[27] = (N96)? 1'b0 : 
                         (N98)? rf_reg_tmp[27] : 
                         (N100)? rf_reg_tmp[59] : 
                         (N102)? rf_reg_tmp[91] : 
                         (N104)? rf_reg_tmp[123] : 
                         (N106)? rf_reg_tmp[155] : 
                         (N108)? rf_reg_tmp[187] : 
                         (N110)? rf_reg_tmp[219] : 
                         (N112)? rf_reg_tmp[251] : 
                         (N114)? rf_reg_tmp[283] : 
                         (N116)? rf_reg_tmp[315] : 
                         (N118)? rf_reg_tmp[347] : 
                         (N120)? rf_reg_tmp[379] : 
                         (N122)? rf_reg_tmp[411] : 
                         (N124)? rf_reg_tmp[443] : 
                         (N126)? rf_reg_tmp[475] : 
                         (N97)? rf_reg_tmp[507] : 
                         (N99)? rf_reg_tmp[539] : 
                         (N101)? rf_reg_tmp[571] : 
                         (N103)? rf_reg_tmp[603] : 
                         (N105)? rf_reg_tmp[635] : 
                         (N107)? rf_reg_tmp[667] : 
                         (N109)? rf_reg_tmp[699] : 
                         (N111)? rf_reg_tmp[731] : 
                         (N113)? rf_reg_tmp[763] : 
                         (N115)? rf_reg_tmp[795] : 
                         (N117)? rf_reg_tmp[827] : 
                         (N119)? rf_reg_tmp[859] : 
                         (N121)? rf_reg_tmp[891] : 
                         (N123)? rf_reg_tmp[923] : 
                         (N125)? rf_reg_tmp[955] : 
                         (N127)? rf_reg_tmp[987] : 1'b0;
  assign rdata_a_o[26] = (N96)? 1'b0 : 
                         (N98)? rf_reg_tmp[26] : 
                         (N100)? rf_reg_tmp[58] : 
                         (N102)? rf_reg_tmp[90] : 
                         (N104)? rf_reg_tmp[122] : 
                         (N106)? rf_reg_tmp[154] : 
                         (N108)? rf_reg_tmp[186] : 
                         (N110)? rf_reg_tmp[218] : 
                         (N112)? rf_reg_tmp[250] : 
                         (N114)? rf_reg_tmp[282] : 
                         (N116)? rf_reg_tmp[314] : 
                         (N118)? rf_reg_tmp[346] : 
                         (N120)? rf_reg_tmp[378] : 
                         (N122)? rf_reg_tmp[410] : 
                         (N124)? rf_reg_tmp[442] : 
                         (N126)? rf_reg_tmp[474] : 
                         (N97)? rf_reg_tmp[506] : 
                         (N99)? rf_reg_tmp[538] : 
                         (N101)? rf_reg_tmp[570] : 
                         (N103)? rf_reg_tmp[602] : 
                         (N105)? rf_reg_tmp[634] : 
                         (N107)? rf_reg_tmp[666] : 
                         (N109)? rf_reg_tmp[698] : 
                         (N111)? rf_reg_tmp[730] : 
                         (N113)? rf_reg_tmp[762] : 
                         (N115)? rf_reg_tmp[794] : 
                         (N117)? rf_reg_tmp[826] : 
                         (N119)? rf_reg_tmp[858] : 
                         (N121)? rf_reg_tmp[890] : 
                         (N123)? rf_reg_tmp[922] : 
                         (N125)? rf_reg_tmp[954] : 
                         (N127)? rf_reg_tmp[986] : 1'b0;
  assign rdata_a_o[25] = (N96)? 1'b0 : 
                         (N98)? rf_reg_tmp[25] : 
                         (N100)? rf_reg_tmp[57] : 
                         (N102)? rf_reg_tmp[89] : 
                         (N104)? rf_reg_tmp[121] : 
                         (N106)? rf_reg_tmp[153] : 
                         (N108)? rf_reg_tmp[185] : 
                         (N110)? rf_reg_tmp[217] : 
                         (N112)? rf_reg_tmp[249] : 
                         (N114)? rf_reg_tmp[281] : 
                         (N116)? rf_reg_tmp[313] : 
                         (N118)? rf_reg_tmp[345] : 
                         (N120)? rf_reg_tmp[377] : 
                         (N122)? rf_reg_tmp[409] : 
                         (N124)? rf_reg_tmp[441] : 
                         (N126)? rf_reg_tmp[473] : 
                         (N97)? rf_reg_tmp[505] : 
                         (N99)? rf_reg_tmp[537] : 
                         (N101)? rf_reg_tmp[569] : 
                         (N103)? rf_reg_tmp[601] : 
                         (N105)? rf_reg_tmp[633] : 
                         (N107)? rf_reg_tmp[665] : 
                         (N109)? rf_reg_tmp[697] : 
                         (N111)? rf_reg_tmp[729] : 
                         (N113)? rf_reg_tmp[761] : 
                         (N115)? rf_reg_tmp[793] : 
                         (N117)? rf_reg_tmp[825] : 
                         (N119)? rf_reg_tmp[857] : 
                         (N121)? rf_reg_tmp[889] : 
                         (N123)? rf_reg_tmp[921] : 
                         (N125)? rf_reg_tmp[953] : 
                         (N127)? rf_reg_tmp[985] : 1'b0;
  assign rdata_a_o[24] = (N96)? 1'b0 : 
                         (N98)? rf_reg_tmp[24] : 
                         (N100)? rf_reg_tmp[56] : 
                         (N102)? rf_reg_tmp[88] : 
                         (N104)? rf_reg_tmp[120] : 
                         (N106)? rf_reg_tmp[152] : 
                         (N108)? rf_reg_tmp[184] : 
                         (N110)? rf_reg_tmp[216] : 
                         (N112)? rf_reg_tmp[248] : 
                         (N114)? rf_reg_tmp[280] : 
                         (N116)? rf_reg_tmp[312] : 
                         (N118)? rf_reg_tmp[344] : 
                         (N120)? rf_reg_tmp[376] : 
                         (N122)? rf_reg_tmp[408] : 
                         (N124)? rf_reg_tmp[440] : 
                         (N126)? rf_reg_tmp[472] : 
                         (N97)? rf_reg_tmp[504] : 
                         (N99)? rf_reg_tmp[536] : 
                         (N101)? rf_reg_tmp[568] : 
                         (N103)? rf_reg_tmp[600] : 
                         (N105)? rf_reg_tmp[632] : 
                         (N107)? rf_reg_tmp[664] : 
                         (N109)? rf_reg_tmp[696] : 
                         (N111)? rf_reg_tmp[728] : 
                         (N113)? rf_reg_tmp[760] : 
                         (N115)? rf_reg_tmp[792] : 
                         (N117)? rf_reg_tmp[824] : 
                         (N119)? rf_reg_tmp[856] : 
                         (N121)? rf_reg_tmp[888] : 
                         (N123)? rf_reg_tmp[920] : 
                         (N125)? rf_reg_tmp[952] : 
                         (N127)? rf_reg_tmp[984] : 1'b0;
  assign rdata_a_o[23] = (N96)? 1'b0 : 
                         (N98)? rf_reg_tmp[23] : 
                         (N100)? rf_reg_tmp[55] : 
                         (N102)? rf_reg_tmp[87] : 
                         (N104)? rf_reg_tmp[119] : 
                         (N106)? rf_reg_tmp[151] : 
                         (N108)? rf_reg_tmp[183] : 
                         (N110)? rf_reg_tmp[215] : 
                         (N112)? rf_reg_tmp[247] : 
                         (N114)? rf_reg_tmp[279] : 
                         (N116)? rf_reg_tmp[311] : 
                         (N118)? rf_reg_tmp[343] : 
                         (N120)? rf_reg_tmp[375] : 
                         (N122)? rf_reg_tmp[407] : 
                         (N124)? rf_reg_tmp[439] : 
                         (N126)? rf_reg_tmp[471] : 
                         (N97)? rf_reg_tmp[503] : 
                         (N99)? rf_reg_tmp[535] : 
                         (N101)? rf_reg_tmp[567] : 
                         (N103)? rf_reg_tmp[599] : 
                         (N105)? rf_reg_tmp[631] : 
                         (N107)? rf_reg_tmp[663] : 
                         (N109)? rf_reg_tmp[695] : 
                         (N111)? rf_reg_tmp[727] : 
                         (N113)? rf_reg_tmp[759] : 
                         (N115)? rf_reg_tmp[791] : 
                         (N117)? rf_reg_tmp[823] : 
                         (N119)? rf_reg_tmp[855] : 
                         (N121)? rf_reg_tmp[887] : 
                         (N123)? rf_reg_tmp[919] : 
                         (N125)? rf_reg_tmp[951] : 
                         (N127)? rf_reg_tmp[983] : 1'b0;
  assign rdata_a_o[22] = (N96)? 1'b0 : 
                         (N98)? rf_reg_tmp[22] : 
                         (N100)? rf_reg_tmp[54] : 
                         (N102)? rf_reg_tmp[86] : 
                         (N104)? rf_reg_tmp[118] : 
                         (N106)? rf_reg_tmp[150] : 
                         (N108)? rf_reg_tmp[182] : 
                         (N110)? rf_reg_tmp[214] : 
                         (N112)? rf_reg_tmp[246] : 
                         (N114)? rf_reg_tmp[278] : 
                         (N116)? rf_reg_tmp[310] : 
                         (N118)? rf_reg_tmp[342] : 
                         (N120)? rf_reg_tmp[374] : 
                         (N122)? rf_reg_tmp[406] : 
                         (N124)? rf_reg_tmp[438] : 
                         (N126)? rf_reg_tmp[470] : 
                         (N97)? rf_reg_tmp[502] : 
                         (N99)? rf_reg_tmp[534] : 
                         (N101)? rf_reg_tmp[566] : 
                         (N103)? rf_reg_tmp[598] : 
                         (N105)? rf_reg_tmp[630] : 
                         (N107)? rf_reg_tmp[662] : 
                         (N109)? rf_reg_tmp[694] : 
                         (N111)? rf_reg_tmp[726] : 
                         (N113)? rf_reg_tmp[758] : 
                         (N115)? rf_reg_tmp[790] : 
                         (N117)? rf_reg_tmp[822] : 
                         (N119)? rf_reg_tmp[854] : 
                         (N121)? rf_reg_tmp[886] : 
                         (N123)? rf_reg_tmp[918] : 
                         (N125)? rf_reg_tmp[950] : 
                         (N127)? rf_reg_tmp[982] : 1'b0;
  assign rdata_a_o[21] = (N96)? 1'b0 : 
                         (N98)? rf_reg_tmp[21] : 
                         (N100)? rf_reg_tmp[53] : 
                         (N102)? rf_reg_tmp[85] : 
                         (N104)? rf_reg_tmp[117] : 
                         (N106)? rf_reg_tmp[149] : 
                         (N108)? rf_reg_tmp[181] : 
                         (N110)? rf_reg_tmp[213] : 
                         (N112)? rf_reg_tmp[245] : 
                         (N114)? rf_reg_tmp[277] : 
                         (N116)? rf_reg_tmp[309] : 
                         (N118)? rf_reg_tmp[341] : 
                         (N120)? rf_reg_tmp[373] : 
                         (N122)? rf_reg_tmp[405] : 
                         (N124)? rf_reg_tmp[437] : 
                         (N126)? rf_reg_tmp[469] : 
                         (N97)? rf_reg_tmp[501] : 
                         (N99)? rf_reg_tmp[533] : 
                         (N101)? rf_reg_tmp[565] : 
                         (N103)? rf_reg_tmp[597] : 
                         (N105)? rf_reg_tmp[629] : 
                         (N107)? rf_reg_tmp[661] : 
                         (N109)? rf_reg_tmp[693] : 
                         (N111)? rf_reg_tmp[725] : 
                         (N113)? rf_reg_tmp[757] : 
                         (N115)? rf_reg_tmp[789] : 
                         (N117)? rf_reg_tmp[821] : 
                         (N119)? rf_reg_tmp[853] : 
                         (N121)? rf_reg_tmp[885] : 
                         (N123)? rf_reg_tmp[917] : 
                         (N125)? rf_reg_tmp[949] : 
                         (N127)? rf_reg_tmp[981] : 1'b0;
  assign rdata_a_o[20] = (N96)? 1'b0 : 
                         (N98)? rf_reg_tmp[20] : 
                         (N100)? rf_reg_tmp[52] : 
                         (N102)? rf_reg_tmp[84] : 
                         (N104)? rf_reg_tmp[116] : 
                         (N106)? rf_reg_tmp[148] : 
                         (N108)? rf_reg_tmp[180] : 
                         (N110)? rf_reg_tmp[212] : 
                         (N112)? rf_reg_tmp[244] : 
                         (N114)? rf_reg_tmp[276] : 
                         (N116)? rf_reg_tmp[308] : 
                         (N118)? rf_reg_tmp[340] : 
                         (N120)? rf_reg_tmp[372] : 
                         (N122)? rf_reg_tmp[404] : 
                         (N124)? rf_reg_tmp[436] : 
                         (N126)? rf_reg_tmp[468] : 
                         (N97)? rf_reg_tmp[500] : 
                         (N99)? rf_reg_tmp[532] : 
                         (N101)? rf_reg_tmp[564] : 
                         (N103)? rf_reg_tmp[596] : 
                         (N105)? rf_reg_tmp[628] : 
                         (N107)? rf_reg_tmp[660] : 
                         (N109)? rf_reg_tmp[692] : 
                         (N111)? rf_reg_tmp[724] : 
                         (N113)? rf_reg_tmp[756] : 
                         (N115)? rf_reg_tmp[788] : 
                         (N117)? rf_reg_tmp[820] : 
                         (N119)? rf_reg_tmp[852] : 
                         (N121)? rf_reg_tmp[884] : 
                         (N123)? rf_reg_tmp[916] : 
                         (N125)? rf_reg_tmp[948] : 
                         (N127)? rf_reg_tmp[980] : 1'b0;
  assign rdata_a_o[19] = (N96)? 1'b0 : 
                         (N98)? rf_reg_tmp[19] : 
                         (N100)? rf_reg_tmp[51] : 
                         (N102)? rf_reg_tmp[83] : 
                         (N104)? rf_reg_tmp[115] : 
                         (N106)? rf_reg_tmp[147] : 
                         (N108)? rf_reg_tmp[179] : 
                         (N110)? rf_reg_tmp[211] : 
                         (N112)? rf_reg_tmp[243] : 
                         (N114)? rf_reg_tmp[275] : 
                         (N116)? rf_reg_tmp[307] : 
                         (N118)? rf_reg_tmp[339] : 
                         (N120)? rf_reg_tmp[371] : 
                         (N122)? rf_reg_tmp[403] : 
                         (N124)? rf_reg_tmp[435] : 
                         (N126)? rf_reg_tmp[467] : 
                         (N97)? rf_reg_tmp[499] : 
                         (N99)? rf_reg_tmp[531] : 
                         (N101)? rf_reg_tmp[563] : 
                         (N103)? rf_reg_tmp[595] : 
                         (N105)? rf_reg_tmp[627] : 
                         (N107)? rf_reg_tmp[659] : 
                         (N109)? rf_reg_tmp[691] : 
                         (N111)? rf_reg_tmp[723] : 
                         (N113)? rf_reg_tmp[755] : 
                         (N115)? rf_reg_tmp[787] : 
                         (N117)? rf_reg_tmp[819] : 
                         (N119)? rf_reg_tmp[851] : 
                         (N121)? rf_reg_tmp[883] : 
                         (N123)? rf_reg_tmp[915] : 
                         (N125)? rf_reg_tmp[947] : 
                         (N127)? rf_reg_tmp[979] : 1'b0;
  assign rdata_a_o[18] = (N96)? 1'b0 : 
                         (N98)? rf_reg_tmp[18] : 
                         (N100)? rf_reg_tmp[50] : 
                         (N102)? rf_reg_tmp[82] : 
                         (N104)? rf_reg_tmp[114] : 
                         (N106)? rf_reg_tmp[146] : 
                         (N108)? rf_reg_tmp[178] : 
                         (N110)? rf_reg_tmp[210] : 
                         (N112)? rf_reg_tmp[242] : 
                         (N114)? rf_reg_tmp[274] : 
                         (N116)? rf_reg_tmp[306] : 
                         (N118)? rf_reg_tmp[338] : 
                         (N120)? rf_reg_tmp[370] : 
                         (N122)? rf_reg_tmp[402] : 
                         (N124)? rf_reg_tmp[434] : 
                         (N126)? rf_reg_tmp[466] : 
                         (N97)? rf_reg_tmp[498] : 
                         (N99)? rf_reg_tmp[530] : 
                         (N101)? rf_reg_tmp[562] : 
                         (N103)? rf_reg_tmp[594] : 
                         (N105)? rf_reg_tmp[626] : 
                         (N107)? rf_reg_tmp[658] : 
                         (N109)? rf_reg_tmp[690] : 
                         (N111)? rf_reg_tmp[722] : 
                         (N113)? rf_reg_tmp[754] : 
                         (N115)? rf_reg_tmp[786] : 
                         (N117)? rf_reg_tmp[818] : 
                         (N119)? rf_reg_tmp[850] : 
                         (N121)? rf_reg_tmp[882] : 
                         (N123)? rf_reg_tmp[914] : 
                         (N125)? rf_reg_tmp[946] : 
                         (N127)? rf_reg_tmp[978] : 1'b0;
  assign rdata_a_o[17] = (N96)? 1'b0 : 
                         (N98)? rf_reg_tmp[17] : 
                         (N100)? rf_reg_tmp[49] : 
                         (N102)? rf_reg_tmp[81] : 
                         (N104)? rf_reg_tmp[113] : 
                         (N106)? rf_reg_tmp[145] : 
                         (N108)? rf_reg_tmp[177] : 
                         (N110)? rf_reg_tmp[209] : 
                         (N112)? rf_reg_tmp[241] : 
                         (N114)? rf_reg_tmp[273] : 
                         (N116)? rf_reg_tmp[305] : 
                         (N118)? rf_reg_tmp[337] : 
                         (N120)? rf_reg_tmp[369] : 
                         (N122)? rf_reg_tmp[401] : 
                         (N124)? rf_reg_tmp[433] : 
                         (N126)? rf_reg_tmp[465] : 
                         (N97)? rf_reg_tmp[497] : 
                         (N99)? rf_reg_tmp[529] : 
                         (N101)? rf_reg_tmp[561] : 
                         (N103)? rf_reg_tmp[593] : 
                         (N105)? rf_reg_tmp[625] : 
                         (N107)? rf_reg_tmp[657] : 
                         (N109)? rf_reg_tmp[689] : 
                         (N111)? rf_reg_tmp[721] : 
                         (N113)? rf_reg_tmp[753] : 
                         (N115)? rf_reg_tmp[785] : 
                         (N117)? rf_reg_tmp[817] : 
                         (N119)? rf_reg_tmp[849] : 
                         (N121)? rf_reg_tmp[881] : 
                         (N123)? rf_reg_tmp[913] : 
                         (N125)? rf_reg_tmp[945] : 
                         (N127)? rf_reg_tmp[977] : 1'b0;
  assign rdata_a_o[16] = (N96)? 1'b0 : 
                         (N98)? rf_reg_tmp[16] : 
                         (N100)? rf_reg_tmp[48] : 
                         (N102)? rf_reg_tmp[80] : 
                         (N104)? rf_reg_tmp[112] : 
                         (N106)? rf_reg_tmp[144] : 
                         (N108)? rf_reg_tmp[176] : 
                         (N110)? rf_reg_tmp[208] : 
                         (N112)? rf_reg_tmp[240] : 
                         (N114)? rf_reg_tmp[272] : 
                         (N116)? rf_reg_tmp[304] : 
                         (N118)? rf_reg_tmp[336] : 
                         (N120)? rf_reg_tmp[368] : 
                         (N122)? rf_reg_tmp[400] : 
                         (N124)? rf_reg_tmp[432] : 
                         (N126)? rf_reg_tmp[464] : 
                         (N97)? rf_reg_tmp[496] : 
                         (N99)? rf_reg_tmp[528] : 
                         (N101)? rf_reg_tmp[560] : 
                         (N103)? rf_reg_tmp[592] : 
                         (N105)? rf_reg_tmp[624] : 
                         (N107)? rf_reg_tmp[656] : 
                         (N109)? rf_reg_tmp[688] : 
                         (N111)? rf_reg_tmp[720] : 
                         (N113)? rf_reg_tmp[752] : 
                         (N115)? rf_reg_tmp[784] : 
                         (N117)? rf_reg_tmp[816] : 
                         (N119)? rf_reg_tmp[848] : 
                         (N121)? rf_reg_tmp[880] : 
                         (N123)? rf_reg_tmp[912] : 
                         (N125)? rf_reg_tmp[944] : 
                         (N127)? rf_reg_tmp[976] : 1'b0;
  assign rdata_a_o[15] = (N96)? 1'b0 : 
                         (N98)? rf_reg_tmp[15] : 
                         (N100)? rf_reg_tmp[47] : 
                         (N102)? rf_reg_tmp[79] : 
                         (N104)? rf_reg_tmp[111] : 
                         (N106)? rf_reg_tmp[143] : 
                         (N108)? rf_reg_tmp[175] : 
                         (N110)? rf_reg_tmp[207] : 
                         (N112)? rf_reg_tmp[239] : 
                         (N114)? rf_reg_tmp[271] : 
                         (N116)? rf_reg_tmp[303] : 
                         (N118)? rf_reg_tmp[335] : 
                         (N120)? rf_reg_tmp[367] : 
                         (N122)? rf_reg_tmp[399] : 
                         (N124)? rf_reg_tmp[431] : 
                         (N126)? rf_reg_tmp[463] : 
                         (N97)? rf_reg_tmp[495] : 
                         (N99)? rf_reg_tmp[527] : 
                         (N101)? rf_reg_tmp[559] : 
                         (N103)? rf_reg_tmp[591] : 
                         (N105)? rf_reg_tmp[623] : 
                         (N107)? rf_reg_tmp[655] : 
                         (N109)? rf_reg_tmp[687] : 
                         (N111)? rf_reg_tmp[719] : 
                         (N113)? rf_reg_tmp[751] : 
                         (N115)? rf_reg_tmp[783] : 
                         (N117)? rf_reg_tmp[815] : 
                         (N119)? rf_reg_tmp[847] : 
                         (N121)? rf_reg_tmp[879] : 
                         (N123)? rf_reg_tmp[911] : 
                         (N125)? rf_reg_tmp[943] : 
                         (N127)? rf_reg_tmp[975] : 1'b0;
  assign rdata_a_o[14] = (N96)? 1'b0 : 
                         (N98)? rf_reg_tmp[14] : 
                         (N100)? rf_reg_tmp[46] : 
                         (N102)? rf_reg_tmp[78] : 
                         (N104)? rf_reg_tmp[110] : 
                         (N106)? rf_reg_tmp[142] : 
                         (N108)? rf_reg_tmp[174] : 
                         (N110)? rf_reg_tmp[206] : 
                         (N112)? rf_reg_tmp[238] : 
                         (N114)? rf_reg_tmp[270] : 
                         (N116)? rf_reg_tmp[302] : 
                         (N118)? rf_reg_tmp[334] : 
                         (N120)? rf_reg_tmp[366] : 
                         (N122)? rf_reg_tmp[398] : 
                         (N124)? rf_reg_tmp[430] : 
                         (N126)? rf_reg_tmp[462] : 
                         (N97)? rf_reg_tmp[494] : 
                         (N99)? rf_reg_tmp[526] : 
                         (N101)? rf_reg_tmp[558] : 
                         (N103)? rf_reg_tmp[590] : 
                         (N105)? rf_reg_tmp[622] : 
                         (N107)? rf_reg_tmp[654] : 
                         (N109)? rf_reg_tmp[686] : 
                         (N111)? rf_reg_tmp[718] : 
                         (N113)? rf_reg_tmp[750] : 
                         (N115)? rf_reg_tmp[782] : 
                         (N117)? rf_reg_tmp[814] : 
                         (N119)? rf_reg_tmp[846] : 
                         (N121)? rf_reg_tmp[878] : 
                         (N123)? rf_reg_tmp[910] : 
                         (N125)? rf_reg_tmp[942] : 
                         (N127)? rf_reg_tmp[974] : 1'b0;
  assign rdata_a_o[13] = (N96)? 1'b0 : 
                         (N98)? rf_reg_tmp[13] : 
                         (N100)? rf_reg_tmp[45] : 
                         (N102)? rf_reg_tmp[77] : 
                         (N104)? rf_reg_tmp[109] : 
                         (N106)? rf_reg_tmp[141] : 
                         (N108)? rf_reg_tmp[173] : 
                         (N110)? rf_reg_tmp[205] : 
                         (N112)? rf_reg_tmp[237] : 
                         (N114)? rf_reg_tmp[269] : 
                         (N116)? rf_reg_tmp[301] : 
                         (N118)? rf_reg_tmp[333] : 
                         (N120)? rf_reg_tmp[365] : 
                         (N122)? rf_reg_tmp[397] : 
                         (N124)? rf_reg_tmp[429] : 
                         (N126)? rf_reg_tmp[461] : 
                         (N97)? rf_reg_tmp[493] : 
                         (N99)? rf_reg_tmp[525] : 
                         (N101)? rf_reg_tmp[557] : 
                         (N103)? rf_reg_tmp[589] : 
                         (N105)? rf_reg_tmp[621] : 
                         (N107)? rf_reg_tmp[653] : 
                         (N109)? rf_reg_tmp[685] : 
                         (N111)? rf_reg_tmp[717] : 
                         (N113)? rf_reg_tmp[749] : 
                         (N115)? rf_reg_tmp[781] : 
                         (N117)? rf_reg_tmp[813] : 
                         (N119)? rf_reg_tmp[845] : 
                         (N121)? rf_reg_tmp[877] : 
                         (N123)? rf_reg_tmp[909] : 
                         (N125)? rf_reg_tmp[941] : 
                         (N127)? rf_reg_tmp[973] : 1'b0;
  assign rdata_a_o[12] = (N96)? 1'b0 : 
                         (N98)? rf_reg_tmp[12] : 
                         (N100)? rf_reg_tmp[44] : 
                         (N102)? rf_reg_tmp[76] : 
                         (N104)? rf_reg_tmp[108] : 
                         (N106)? rf_reg_tmp[140] : 
                         (N108)? rf_reg_tmp[172] : 
                         (N110)? rf_reg_tmp[204] : 
                         (N112)? rf_reg_tmp[236] : 
                         (N114)? rf_reg_tmp[268] : 
                         (N116)? rf_reg_tmp[300] : 
                         (N118)? rf_reg_tmp[332] : 
                         (N120)? rf_reg_tmp[364] : 
                         (N122)? rf_reg_tmp[396] : 
                         (N124)? rf_reg_tmp[428] : 
                         (N126)? rf_reg_tmp[460] : 
                         (N97)? rf_reg_tmp[492] : 
                         (N99)? rf_reg_tmp[524] : 
                         (N101)? rf_reg_tmp[556] : 
                         (N103)? rf_reg_tmp[588] : 
                         (N105)? rf_reg_tmp[620] : 
                         (N107)? rf_reg_tmp[652] : 
                         (N109)? rf_reg_tmp[684] : 
                         (N111)? rf_reg_tmp[716] : 
                         (N113)? rf_reg_tmp[748] : 
                         (N115)? rf_reg_tmp[780] : 
                         (N117)? rf_reg_tmp[812] : 
                         (N119)? rf_reg_tmp[844] : 
                         (N121)? rf_reg_tmp[876] : 
                         (N123)? rf_reg_tmp[908] : 
                         (N125)? rf_reg_tmp[940] : 
                         (N127)? rf_reg_tmp[972] : 1'b0;
  assign rdata_a_o[11] = (N96)? 1'b0 : 
                         (N98)? rf_reg_tmp[11] : 
                         (N100)? rf_reg_tmp[43] : 
                         (N102)? rf_reg_tmp[75] : 
                         (N104)? rf_reg_tmp[107] : 
                         (N106)? rf_reg_tmp[139] : 
                         (N108)? rf_reg_tmp[171] : 
                         (N110)? rf_reg_tmp[203] : 
                         (N112)? rf_reg_tmp[235] : 
                         (N114)? rf_reg_tmp[267] : 
                         (N116)? rf_reg_tmp[299] : 
                         (N118)? rf_reg_tmp[331] : 
                         (N120)? rf_reg_tmp[363] : 
                         (N122)? rf_reg_tmp[395] : 
                         (N124)? rf_reg_tmp[427] : 
                         (N126)? rf_reg_tmp[459] : 
                         (N97)? rf_reg_tmp[491] : 
                         (N99)? rf_reg_tmp[523] : 
                         (N101)? rf_reg_tmp[555] : 
                         (N103)? rf_reg_tmp[587] : 
                         (N105)? rf_reg_tmp[619] : 
                         (N107)? rf_reg_tmp[651] : 
                         (N109)? rf_reg_tmp[683] : 
                         (N111)? rf_reg_tmp[715] : 
                         (N113)? rf_reg_tmp[747] : 
                         (N115)? rf_reg_tmp[779] : 
                         (N117)? rf_reg_tmp[811] : 
                         (N119)? rf_reg_tmp[843] : 
                         (N121)? rf_reg_tmp[875] : 
                         (N123)? rf_reg_tmp[907] : 
                         (N125)? rf_reg_tmp[939] : 
                         (N127)? rf_reg_tmp[971] : 1'b0;
  assign rdata_a_o[10] = (N96)? 1'b0 : 
                         (N98)? rf_reg_tmp[10] : 
                         (N100)? rf_reg_tmp[42] : 
                         (N102)? rf_reg_tmp[74] : 
                         (N104)? rf_reg_tmp[106] : 
                         (N106)? rf_reg_tmp[138] : 
                         (N108)? rf_reg_tmp[170] : 
                         (N110)? rf_reg_tmp[202] : 
                         (N112)? rf_reg_tmp[234] : 
                         (N114)? rf_reg_tmp[266] : 
                         (N116)? rf_reg_tmp[298] : 
                         (N118)? rf_reg_tmp[330] : 
                         (N120)? rf_reg_tmp[362] : 
                         (N122)? rf_reg_tmp[394] : 
                         (N124)? rf_reg_tmp[426] : 
                         (N126)? rf_reg_tmp[458] : 
                         (N97)? rf_reg_tmp[490] : 
                         (N99)? rf_reg_tmp[522] : 
                         (N101)? rf_reg_tmp[554] : 
                         (N103)? rf_reg_tmp[586] : 
                         (N105)? rf_reg_tmp[618] : 
                         (N107)? rf_reg_tmp[650] : 
                         (N109)? rf_reg_tmp[682] : 
                         (N111)? rf_reg_tmp[714] : 
                         (N113)? rf_reg_tmp[746] : 
                         (N115)? rf_reg_tmp[778] : 
                         (N117)? rf_reg_tmp[810] : 
                         (N119)? rf_reg_tmp[842] : 
                         (N121)? rf_reg_tmp[874] : 
                         (N123)? rf_reg_tmp[906] : 
                         (N125)? rf_reg_tmp[938] : 
                         (N127)? rf_reg_tmp[970] : 1'b0;
  assign rdata_a_o[9] = (N96)? 1'b0 : 
                        (N98)? rf_reg_tmp[9] : 
                        (N100)? rf_reg_tmp[41] : 
                        (N102)? rf_reg_tmp[73] : 
                        (N104)? rf_reg_tmp[105] : 
                        (N106)? rf_reg_tmp[137] : 
                        (N108)? rf_reg_tmp[169] : 
                        (N110)? rf_reg_tmp[201] : 
                        (N112)? rf_reg_tmp[233] : 
                        (N114)? rf_reg_tmp[265] : 
                        (N116)? rf_reg_tmp[297] : 
                        (N118)? rf_reg_tmp[329] : 
                        (N120)? rf_reg_tmp[361] : 
                        (N122)? rf_reg_tmp[393] : 
                        (N124)? rf_reg_tmp[425] : 
                        (N126)? rf_reg_tmp[457] : 
                        (N97)? rf_reg_tmp[489] : 
                        (N99)? rf_reg_tmp[521] : 
                        (N101)? rf_reg_tmp[553] : 
                        (N103)? rf_reg_tmp[585] : 
                        (N105)? rf_reg_tmp[617] : 
                        (N107)? rf_reg_tmp[649] : 
                        (N109)? rf_reg_tmp[681] : 
                        (N111)? rf_reg_tmp[713] : 
                        (N113)? rf_reg_tmp[745] : 
                        (N115)? rf_reg_tmp[777] : 
                        (N117)? rf_reg_tmp[809] : 
                        (N119)? rf_reg_tmp[841] : 
                        (N121)? rf_reg_tmp[873] : 
                        (N123)? rf_reg_tmp[905] : 
                        (N125)? rf_reg_tmp[937] : 
                        (N127)? rf_reg_tmp[969] : 1'b0;
  assign rdata_a_o[8] = (N96)? 1'b0 : 
                        (N98)? rf_reg_tmp[8] : 
                        (N100)? rf_reg_tmp[40] : 
                        (N102)? rf_reg_tmp[72] : 
                        (N104)? rf_reg_tmp[104] : 
                        (N106)? rf_reg_tmp[136] : 
                        (N108)? rf_reg_tmp[168] : 
                        (N110)? rf_reg_tmp[200] : 
                        (N112)? rf_reg_tmp[232] : 
                        (N114)? rf_reg_tmp[264] : 
                        (N116)? rf_reg_tmp[296] : 
                        (N118)? rf_reg_tmp[328] : 
                        (N120)? rf_reg_tmp[360] : 
                        (N122)? rf_reg_tmp[392] : 
                        (N124)? rf_reg_tmp[424] : 
                        (N126)? rf_reg_tmp[456] : 
                        (N97)? rf_reg_tmp[488] : 
                        (N99)? rf_reg_tmp[520] : 
                        (N101)? rf_reg_tmp[552] : 
                        (N103)? rf_reg_tmp[584] : 
                        (N105)? rf_reg_tmp[616] : 
                        (N107)? rf_reg_tmp[648] : 
                        (N109)? rf_reg_tmp[680] : 
                        (N111)? rf_reg_tmp[712] : 
                        (N113)? rf_reg_tmp[744] : 
                        (N115)? rf_reg_tmp[776] : 
                        (N117)? rf_reg_tmp[808] : 
                        (N119)? rf_reg_tmp[840] : 
                        (N121)? rf_reg_tmp[872] : 
                        (N123)? rf_reg_tmp[904] : 
                        (N125)? rf_reg_tmp[936] : 
                        (N127)? rf_reg_tmp[968] : 1'b0;
  assign rdata_a_o[7] = (N96)? 1'b0 : 
                        (N98)? rf_reg_tmp[7] : 
                        (N100)? rf_reg_tmp[39] : 
                        (N102)? rf_reg_tmp[71] : 
                        (N104)? rf_reg_tmp[103] : 
                        (N106)? rf_reg_tmp[135] : 
                        (N108)? rf_reg_tmp[167] : 
                        (N110)? rf_reg_tmp[199] : 
                        (N112)? rf_reg_tmp[231] : 
                        (N114)? rf_reg_tmp[263] : 
                        (N116)? rf_reg_tmp[295] : 
                        (N118)? rf_reg_tmp[327] : 
                        (N120)? rf_reg_tmp[359] : 
                        (N122)? rf_reg_tmp[391] : 
                        (N124)? rf_reg_tmp[423] : 
                        (N126)? rf_reg_tmp[455] : 
                        (N97)? rf_reg_tmp[487] : 
                        (N99)? rf_reg_tmp[519] : 
                        (N101)? rf_reg_tmp[551] : 
                        (N103)? rf_reg_tmp[583] : 
                        (N105)? rf_reg_tmp[615] : 
                        (N107)? rf_reg_tmp[647] : 
                        (N109)? rf_reg_tmp[679] : 
                        (N111)? rf_reg_tmp[711] : 
                        (N113)? rf_reg_tmp[743] : 
                        (N115)? rf_reg_tmp[775] : 
                        (N117)? rf_reg_tmp[807] : 
                        (N119)? rf_reg_tmp[839] : 
                        (N121)? rf_reg_tmp[871] : 
                        (N123)? rf_reg_tmp[903] : 
                        (N125)? rf_reg_tmp[935] : 
                        (N127)? rf_reg_tmp[967] : 1'b0;
  assign rdata_a_o[6] = (N96)? 1'b0 : 
                        (N98)? rf_reg_tmp[6] : 
                        (N100)? rf_reg_tmp[38] : 
                        (N102)? rf_reg_tmp[70] : 
                        (N104)? rf_reg_tmp[102] : 
                        (N106)? rf_reg_tmp[134] : 
                        (N108)? rf_reg_tmp[166] : 
                        (N110)? rf_reg_tmp[198] : 
                        (N112)? rf_reg_tmp[230] : 
                        (N114)? rf_reg_tmp[262] : 
                        (N116)? rf_reg_tmp[294] : 
                        (N118)? rf_reg_tmp[326] : 
                        (N120)? rf_reg_tmp[358] : 
                        (N122)? rf_reg_tmp[390] : 
                        (N124)? rf_reg_tmp[422] : 
                        (N126)? rf_reg_tmp[454] : 
                        (N97)? rf_reg_tmp[486] : 
                        (N99)? rf_reg_tmp[518] : 
                        (N101)? rf_reg_tmp[550] : 
                        (N103)? rf_reg_tmp[582] : 
                        (N105)? rf_reg_tmp[614] : 
                        (N107)? rf_reg_tmp[646] : 
                        (N109)? rf_reg_tmp[678] : 
                        (N111)? rf_reg_tmp[710] : 
                        (N113)? rf_reg_tmp[742] : 
                        (N115)? rf_reg_tmp[774] : 
                        (N117)? rf_reg_tmp[806] : 
                        (N119)? rf_reg_tmp[838] : 
                        (N121)? rf_reg_tmp[870] : 
                        (N123)? rf_reg_tmp[902] : 
                        (N125)? rf_reg_tmp[934] : 
                        (N127)? rf_reg_tmp[966] : 1'b0;
  assign rdata_a_o[5] = (N96)? 1'b0 : 
                        (N98)? rf_reg_tmp[5] : 
                        (N100)? rf_reg_tmp[37] : 
                        (N102)? rf_reg_tmp[69] : 
                        (N104)? rf_reg_tmp[101] : 
                        (N106)? rf_reg_tmp[133] : 
                        (N108)? rf_reg_tmp[165] : 
                        (N110)? rf_reg_tmp[197] : 
                        (N112)? rf_reg_tmp[229] : 
                        (N114)? rf_reg_tmp[261] : 
                        (N116)? rf_reg_tmp[293] : 
                        (N118)? rf_reg_tmp[325] : 
                        (N120)? rf_reg_tmp[357] : 
                        (N122)? rf_reg_tmp[389] : 
                        (N124)? rf_reg_tmp[421] : 
                        (N126)? rf_reg_tmp[453] : 
                        (N97)? rf_reg_tmp[485] : 
                        (N99)? rf_reg_tmp[517] : 
                        (N101)? rf_reg_tmp[549] : 
                        (N103)? rf_reg_tmp[581] : 
                        (N105)? rf_reg_tmp[613] : 
                        (N107)? rf_reg_tmp[645] : 
                        (N109)? rf_reg_tmp[677] : 
                        (N111)? rf_reg_tmp[709] : 
                        (N113)? rf_reg_tmp[741] : 
                        (N115)? rf_reg_tmp[773] : 
                        (N117)? rf_reg_tmp[805] : 
                        (N119)? rf_reg_tmp[837] : 
                        (N121)? rf_reg_tmp[869] : 
                        (N123)? rf_reg_tmp[901] : 
                        (N125)? rf_reg_tmp[933] : 
                        (N127)? rf_reg_tmp[965] : 1'b0;
  assign rdata_a_o[4] = (N96)? 1'b0 : 
                        (N98)? rf_reg_tmp[4] : 
                        (N100)? rf_reg_tmp[36] : 
                        (N102)? rf_reg_tmp[68] : 
                        (N104)? rf_reg_tmp[100] : 
                        (N106)? rf_reg_tmp[132] : 
                        (N108)? rf_reg_tmp[164] : 
                        (N110)? rf_reg_tmp[196] : 
                        (N112)? rf_reg_tmp[228] : 
                        (N114)? rf_reg_tmp[260] : 
                        (N116)? rf_reg_tmp[292] : 
                        (N118)? rf_reg_tmp[324] : 
                        (N120)? rf_reg_tmp[356] : 
                        (N122)? rf_reg_tmp[388] : 
                        (N124)? rf_reg_tmp[420] : 
                        (N126)? rf_reg_tmp[452] : 
                        (N97)? rf_reg_tmp[484] : 
                        (N99)? rf_reg_tmp[516] : 
                        (N101)? rf_reg_tmp[548] : 
                        (N103)? rf_reg_tmp[580] : 
                        (N105)? rf_reg_tmp[612] : 
                        (N107)? rf_reg_tmp[644] : 
                        (N109)? rf_reg_tmp[676] : 
                        (N111)? rf_reg_tmp[708] : 
                        (N113)? rf_reg_tmp[740] : 
                        (N115)? rf_reg_tmp[772] : 
                        (N117)? rf_reg_tmp[804] : 
                        (N119)? rf_reg_tmp[836] : 
                        (N121)? rf_reg_tmp[868] : 
                        (N123)? rf_reg_tmp[900] : 
                        (N125)? rf_reg_tmp[932] : 
                        (N127)? rf_reg_tmp[964] : 1'b0;
  assign rdata_a_o[3] = (N96)? 1'b0 : 
                        (N98)? rf_reg_tmp[3] : 
                        (N100)? rf_reg_tmp[35] : 
                        (N102)? rf_reg_tmp[67] : 
                        (N104)? rf_reg_tmp[99] : 
                        (N106)? rf_reg_tmp[131] : 
                        (N108)? rf_reg_tmp[163] : 
                        (N110)? rf_reg_tmp[195] : 
                        (N112)? rf_reg_tmp[227] : 
                        (N114)? rf_reg_tmp[259] : 
                        (N116)? rf_reg_tmp[291] : 
                        (N118)? rf_reg_tmp[323] : 
                        (N120)? rf_reg_tmp[355] : 
                        (N122)? rf_reg_tmp[387] : 
                        (N124)? rf_reg_tmp[419] : 
                        (N126)? rf_reg_tmp[451] : 
                        (N97)? rf_reg_tmp[483] : 
                        (N99)? rf_reg_tmp[515] : 
                        (N101)? rf_reg_tmp[547] : 
                        (N103)? rf_reg_tmp[579] : 
                        (N105)? rf_reg_tmp[611] : 
                        (N107)? rf_reg_tmp[643] : 
                        (N109)? rf_reg_tmp[675] : 
                        (N111)? rf_reg_tmp[707] : 
                        (N113)? rf_reg_tmp[739] : 
                        (N115)? rf_reg_tmp[771] : 
                        (N117)? rf_reg_tmp[803] : 
                        (N119)? rf_reg_tmp[835] : 
                        (N121)? rf_reg_tmp[867] : 
                        (N123)? rf_reg_tmp[899] : 
                        (N125)? rf_reg_tmp[931] : 
                        (N127)? rf_reg_tmp[963] : 1'b0;
  assign rdata_a_o[2] = (N96)? 1'b0 : 
                        (N98)? rf_reg_tmp[2] : 
                        (N100)? rf_reg_tmp[34] : 
                        (N102)? rf_reg_tmp[66] : 
                        (N104)? rf_reg_tmp[98] : 
                        (N106)? rf_reg_tmp[130] : 
                        (N108)? rf_reg_tmp[162] : 
                        (N110)? rf_reg_tmp[194] : 
                        (N112)? rf_reg_tmp[226] : 
                        (N114)? rf_reg_tmp[258] : 
                        (N116)? rf_reg_tmp[290] : 
                        (N118)? rf_reg_tmp[322] : 
                        (N120)? rf_reg_tmp[354] : 
                        (N122)? rf_reg_tmp[386] : 
                        (N124)? rf_reg_tmp[418] : 
                        (N126)? rf_reg_tmp[450] : 
                        (N97)? rf_reg_tmp[482] : 
                        (N99)? rf_reg_tmp[514] : 
                        (N101)? rf_reg_tmp[546] : 
                        (N103)? rf_reg_tmp[578] : 
                        (N105)? rf_reg_tmp[610] : 
                        (N107)? rf_reg_tmp[642] : 
                        (N109)? rf_reg_tmp[674] : 
                        (N111)? rf_reg_tmp[706] : 
                        (N113)? rf_reg_tmp[738] : 
                        (N115)? rf_reg_tmp[770] : 
                        (N117)? rf_reg_tmp[802] : 
                        (N119)? rf_reg_tmp[834] : 
                        (N121)? rf_reg_tmp[866] : 
                        (N123)? rf_reg_tmp[898] : 
                        (N125)? rf_reg_tmp[930] : 
                        (N127)? rf_reg_tmp[962] : 1'b0;
  assign rdata_a_o[1] = (N96)? 1'b0 : 
                        (N98)? rf_reg_tmp[1] : 
                        (N100)? rf_reg_tmp[33] : 
                        (N102)? rf_reg_tmp[65] : 
                        (N104)? rf_reg_tmp[97] : 
                        (N106)? rf_reg_tmp[129] : 
                        (N108)? rf_reg_tmp[161] : 
                        (N110)? rf_reg_tmp[193] : 
                        (N112)? rf_reg_tmp[225] : 
                        (N114)? rf_reg_tmp[257] : 
                        (N116)? rf_reg_tmp[289] : 
                        (N118)? rf_reg_tmp[321] : 
                        (N120)? rf_reg_tmp[353] : 
                        (N122)? rf_reg_tmp[385] : 
                        (N124)? rf_reg_tmp[417] : 
                        (N126)? rf_reg_tmp[449] : 
                        (N97)? rf_reg_tmp[481] : 
                        (N99)? rf_reg_tmp[513] : 
                        (N101)? rf_reg_tmp[545] : 
                        (N103)? rf_reg_tmp[577] : 
                        (N105)? rf_reg_tmp[609] : 
                        (N107)? rf_reg_tmp[641] : 
                        (N109)? rf_reg_tmp[673] : 
                        (N111)? rf_reg_tmp[705] : 
                        (N113)? rf_reg_tmp[737] : 
                        (N115)? rf_reg_tmp[769] : 
                        (N117)? rf_reg_tmp[801] : 
                        (N119)? rf_reg_tmp[833] : 
                        (N121)? rf_reg_tmp[865] : 
                        (N123)? rf_reg_tmp[897] : 
                        (N125)? rf_reg_tmp[929] : 
                        (N127)? rf_reg_tmp[961] : 1'b0;
  assign rdata_a_o[0] = (N96)? 1'b0 : 
                        (N98)? rf_reg_tmp[0] : 
                        (N100)? rf_reg_tmp[32] : 
                        (N102)? rf_reg_tmp[64] : 
                        (N104)? rf_reg_tmp[96] : 
                        (N106)? rf_reg_tmp[128] : 
                        (N108)? rf_reg_tmp[160] : 
                        (N110)? rf_reg_tmp[192] : 
                        (N112)? rf_reg_tmp[224] : 
                        (N114)? rf_reg_tmp[256] : 
                        (N116)? rf_reg_tmp[288] : 
                        (N118)? rf_reg_tmp[320] : 
                        (N120)? rf_reg_tmp[352] : 
                        (N122)? rf_reg_tmp[384] : 
                        (N124)? rf_reg_tmp[416] : 
                        (N126)? rf_reg_tmp[448] : 
                        (N97)? rf_reg_tmp[480] : 
                        (N99)? rf_reg_tmp[512] : 
                        (N101)? rf_reg_tmp[544] : 
                        (N103)? rf_reg_tmp[576] : 
                        (N105)? rf_reg_tmp[608] : 
                        (N107)? rf_reg_tmp[640] : 
                        (N109)? rf_reg_tmp[672] : 
                        (N111)? rf_reg_tmp[704] : 
                        (N113)? rf_reg_tmp[736] : 
                        (N115)? rf_reg_tmp[768] : 
                        (N117)? rf_reg_tmp[800] : 
                        (N119)? rf_reg_tmp[832] : 
                        (N121)? rf_reg_tmp[864] : 
                        (N123)? rf_reg_tmp[896] : 
                        (N125)? rf_reg_tmp[928] : 
                        (N127)? rf_reg_tmp[960] : 1'b0;
  assign rdata_b_o[31] = (N161)? 1'b0 : 
                         (N163)? rf_reg_tmp[31] : 
                         (N165)? rf_reg_tmp[63] : 
                         (N167)? rf_reg_tmp[95] : 
                         (N169)? rf_reg_tmp[127] : 
                         (N171)? rf_reg_tmp[159] : 
                         (N173)? rf_reg_tmp[191] : 
                         (N175)? rf_reg_tmp[223] : 
                         (N177)? rf_reg_tmp[255] : 
                         (N179)? rf_reg_tmp[287] : 
                         (N181)? rf_reg_tmp[319] : 
                         (N183)? rf_reg_tmp[351] : 
                         (N185)? rf_reg_tmp[383] : 
                         (N187)? rf_reg_tmp[415] : 
                         (N189)? rf_reg_tmp[447] : 
                         (N191)? rf_reg_tmp[479] : 
                         (N162)? rf_reg_tmp[511] : 
                         (N164)? rf_reg_tmp[543] : 
                         (N166)? rf_reg_tmp[575] : 
                         (N168)? rf_reg_tmp[607] : 
                         (N170)? rf_reg_tmp[639] : 
                         (N172)? rf_reg_tmp[671] : 
                         (N174)? rf_reg_tmp[703] : 
                         (N176)? rf_reg_tmp[735] : 
                         (N178)? rf_reg_tmp[767] : 
                         (N180)? rf_reg_tmp[799] : 
                         (N182)? rf_reg_tmp[831] : 
                         (N184)? rf_reg_tmp[863] : 
                         (N186)? rf_reg_tmp[895] : 
                         (N188)? rf_reg_tmp[927] : 
                         (N190)? rf_reg_tmp[959] : 
                         (N192)? rf_reg_tmp[991] : 1'b0;
  assign rdata_b_o[30] = (N161)? 1'b0 : 
                         (N163)? rf_reg_tmp[30] : 
                         (N165)? rf_reg_tmp[62] : 
                         (N167)? rf_reg_tmp[94] : 
                         (N169)? rf_reg_tmp[126] : 
                         (N171)? rf_reg_tmp[158] : 
                         (N173)? rf_reg_tmp[190] : 
                         (N175)? rf_reg_tmp[222] : 
                         (N177)? rf_reg_tmp[254] : 
                         (N179)? rf_reg_tmp[286] : 
                         (N181)? rf_reg_tmp[318] : 
                         (N183)? rf_reg_tmp[350] : 
                         (N185)? rf_reg_tmp[382] : 
                         (N187)? rf_reg_tmp[414] : 
                         (N189)? rf_reg_tmp[446] : 
                         (N191)? rf_reg_tmp[478] : 
                         (N162)? rf_reg_tmp[510] : 
                         (N164)? rf_reg_tmp[542] : 
                         (N166)? rf_reg_tmp[574] : 
                         (N168)? rf_reg_tmp[606] : 
                         (N170)? rf_reg_tmp[638] : 
                         (N172)? rf_reg_tmp[670] : 
                         (N174)? rf_reg_tmp[702] : 
                         (N176)? rf_reg_tmp[734] : 
                         (N178)? rf_reg_tmp[766] : 
                         (N180)? rf_reg_tmp[798] : 
                         (N182)? rf_reg_tmp[830] : 
                         (N184)? rf_reg_tmp[862] : 
                         (N186)? rf_reg_tmp[894] : 
                         (N188)? rf_reg_tmp[926] : 
                         (N190)? rf_reg_tmp[958] : 
                         (N192)? rf_reg_tmp[990] : 1'b0;
  assign rdata_b_o[29] = (N161)? 1'b0 : 
                         (N163)? rf_reg_tmp[29] : 
                         (N165)? rf_reg_tmp[61] : 
                         (N167)? rf_reg_tmp[93] : 
                         (N169)? rf_reg_tmp[125] : 
                         (N171)? rf_reg_tmp[157] : 
                         (N173)? rf_reg_tmp[189] : 
                         (N175)? rf_reg_tmp[221] : 
                         (N177)? rf_reg_tmp[253] : 
                         (N179)? rf_reg_tmp[285] : 
                         (N181)? rf_reg_tmp[317] : 
                         (N183)? rf_reg_tmp[349] : 
                         (N185)? rf_reg_tmp[381] : 
                         (N187)? rf_reg_tmp[413] : 
                         (N189)? rf_reg_tmp[445] : 
                         (N191)? rf_reg_tmp[477] : 
                         (N162)? rf_reg_tmp[509] : 
                         (N164)? rf_reg_tmp[541] : 
                         (N166)? rf_reg_tmp[573] : 
                         (N168)? rf_reg_tmp[605] : 
                         (N170)? rf_reg_tmp[637] : 
                         (N172)? rf_reg_tmp[669] : 
                         (N174)? rf_reg_tmp[701] : 
                         (N176)? rf_reg_tmp[733] : 
                         (N178)? rf_reg_tmp[765] : 
                         (N180)? rf_reg_tmp[797] : 
                         (N182)? rf_reg_tmp[829] : 
                         (N184)? rf_reg_tmp[861] : 
                         (N186)? rf_reg_tmp[893] : 
                         (N188)? rf_reg_tmp[925] : 
                         (N190)? rf_reg_tmp[957] : 
                         (N192)? rf_reg_tmp[989] : 1'b0;
  assign rdata_b_o[28] = (N161)? 1'b0 : 
                         (N163)? rf_reg_tmp[28] : 
                         (N165)? rf_reg_tmp[60] : 
                         (N167)? rf_reg_tmp[92] : 
                         (N169)? rf_reg_tmp[124] : 
                         (N171)? rf_reg_tmp[156] : 
                         (N173)? rf_reg_tmp[188] : 
                         (N175)? rf_reg_tmp[220] : 
                         (N177)? rf_reg_tmp[252] : 
                         (N179)? rf_reg_tmp[284] : 
                         (N181)? rf_reg_tmp[316] : 
                         (N183)? rf_reg_tmp[348] : 
                         (N185)? rf_reg_tmp[380] : 
                         (N187)? rf_reg_tmp[412] : 
                         (N189)? rf_reg_tmp[444] : 
                         (N191)? rf_reg_tmp[476] : 
                         (N162)? rf_reg_tmp[508] : 
                         (N164)? rf_reg_tmp[540] : 
                         (N166)? rf_reg_tmp[572] : 
                         (N168)? rf_reg_tmp[604] : 
                         (N170)? rf_reg_tmp[636] : 
                         (N172)? rf_reg_tmp[668] : 
                         (N174)? rf_reg_tmp[700] : 
                         (N176)? rf_reg_tmp[732] : 
                         (N178)? rf_reg_tmp[764] : 
                         (N180)? rf_reg_tmp[796] : 
                         (N182)? rf_reg_tmp[828] : 
                         (N184)? rf_reg_tmp[860] : 
                         (N186)? rf_reg_tmp[892] : 
                         (N188)? rf_reg_tmp[924] : 
                         (N190)? rf_reg_tmp[956] : 
                         (N192)? rf_reg_tmp[988] : 1'b0;
  assign rdata_b_o[27] = (N161)? 1'b0 : 
                         (N163)? rf_reg_tmp[27] : 
                         (N165)? rf_reg_tmp[59] : 
                         (N167)? rf_reg_tmp[91] : 
                         (N169)? rf_reg_tmp[123] : 
                         (N171)? rf_reg_tmp[155] : 
                         (N173)? rf_reg_tmp[187] : 
                         (N175)? rf_reg_tmp[219] : 
                         (N177)? rf_reg_tmp[251] : 
                         (N179)? rf_reg_tmp[283] : 
                         (N181)? rf_reg_tmp[315] : 
                         (N183)? rf_reg_tmp[347] : 
                         (N185)? rf_reg_tmp[379] : 
                         (N187)? rf_reg_tmp[411] : 
                         (N189)? rf_reg_tmp[443] : 
                         (N191)? rf_reg_tmp[475] : 
                         (N162)? rf_reg_tmp[507] : 
                         (N164)? rf_reg_tmp[539] : 
                         (N166)? rf_reg_tmp[571] : 
                         (N168)? rf_reg_tmp[603] : 
                         (N170)? rf_reg_tmp[635] : 
                         (N172)? rf_reg_tmp[667] : 
                         (N174)? rf_reg_tmp[699] : 
                         (N176)? rf_reg_tmp[731] : 
                         (N178)? rf_reg_tmp[763] : 
                         (N180)? rf_reg_tmp[795] : 
                         (N182)? rf_reg_tmp[827] : 
                         (N184)? rf_reg_tmp[859] : 
                         (N186)? rf_reg_tmp[891] : 
                         (N188)? rf_reg_tmp[923] : 
                         (N190)? rf_reg_tmp[955] : 
                         (N192)? rf_reg_tmp[987] : 1'b0;
  assign rdata_b_o[26] = (N161)? 1'b0 : 
                         (N163)? rf_reg_tmp[26] : 
                         (N165)? rf_reg_tmp[58] : 
                         (N167)? rf_reg_tmp[90] : 
                         (N169)? rf_reg_tmp[122] : 
                         (N171)? rf_reg_tmp[154] : 
                         (N173)? rf_reg_tmp[186] : 
                         (N175)? rf_reg_tmp[218] : 
                         (N177)? rf_reg_tmp[250] : 
                         (N179)? rf_reg_tmp[282] : 
                         (N181)? rf_reg_tmp[314] : 
                         (N183)? rf_reg_tmp[346] : 
                         (N185)? rf_reg_tmp[378] : 
                         (N187)? rf_reg_tmp[410] : 
                         (N189)? rf_reg_tmp[442] : 
                         (N191)? rf_reg_tmp[474] : 
                         (N162)? rf_reg_tmp[506] : 
                         (N164)? rf_reg_tmp[538] : 
                         (N166)? rf_reg_tmp[570] : 
                         (N168)? rf_reg_tmp[602] : 
                         (N170)? rf_reg_tmp[634] : 
                         (N172)? rf_reg_tmp[666] : 
                         (N174)? rf_reg_tmp[698] : 
                         (N176)? rf_reg_tmp[730] : 
                         (N178)? rf_reg_tmp[762] : 
                         (N180)? rf_reg_tmp[794] : 
                         (N182)? rf_reg_tmp[826] : 
                         (N184)? rf_reg_tmp[858] : 
                         (N186)? rf_reg_tmp[890] : 
                         (N188)? rf_reg_tmp[922] : 
                         (N190)? rf_reg_tmp[954] : 
                         (N192)? rf_reg_tmp[986] : 1'b0;
  assign rdata_b_o[25] = (N161)? 1'b0 : 
                         (N163)? rf_reg_tmp[25] : 
                         (N165)? rf_reg_tmp[57] : 
                         (N167)? rf_reg_tmp[89] : 
                         (N169)? rf_reg_tmp[121] : 
                         (N171)? rf_reg_tmp[153] : 
                         (N173)? rf_reg_tmp[185] : 
                         (N175)? rf_reg_tmp[217] : 
                         (N177)? rf_reg_tmp[249] : 
                         (N179)? rf_reg_tmp[281] : 
                         (N181)? rf_reg_tmp[313] : 
                         (N183)? rf_reg_tmp[345] : 
                         (N185)? rf_reg_tmp[377] : 
                         (N187)? rf_reg_tmp[409] : 
                         (N189)? rf_reg_tmp[441] : 
                         (N191)? rf_reg_tmp[473] : 
                         (N162)? rf_reg_tmp[505] : 
                         (N164)? rf_reg_tmp[537] : 
                         (N166)? rf_reg_tmp[569] : 
                         (N168)? rf_reg_tmp[601] : 
                         (N170)? rf_reg_tmp[633] : 
                         (N172)? rf_reg_tmp[665] : 
                         (N174)? rf_reg_tmp[697] : 
                         (N176)? rf_reg_tmp[729] : 
                         (N178)? rf_reg_tmp[761] : 
                         (N180)? rf_reg_tmp[793] : 
                         (N182)? rf_reg_tmp[825] : 
                         (N184)? rf_reg_tmp[857] : 
                         (N186)? rf_reg_tmp[889] : 
                         (N188)? rf_reg_tmp[921] : 
                         (N190)? rf_reg_tmp[953] : 
                         (N192)? rf_reg_tmp[985] : 1'b0;
  assign rdata_b_o[24] = (N161)? 1'b0 : 
                         (N163)? rf_reg_tmp[24] : 
                         (N165)? rf_reg_tmp[56] : 
                         (N167)? rf_reg_tmp[88] : 
                         (N169)? rf_reg_tmp[120] : 
                         (N171)? rf_reg_tmp[152] : 
                         (N173)? rf_reg_tmp[184] : 
                         (N175)? rf_reg_tmp[216] : 
                         (N177)? rf_reg_tmp[248] : 
                         (N179)? rf_reg_tmp[280] : 
                         (N181)? rf_reg_tmp[312] : 
                         (N183)? rf_reg_tmp[344] : 
                         (N185)? rf_reg_tmp[376] : 
                         (N187)? rf_reg_tmp[408] : 
                         (N189)? rf_reg_tmp[440] : 
                         (N191)? rf_reg_tmp[472] : 
                         (N162)? rf_reg_tmp[504] : 
                         (N164)? rf_reg_tmp[536] : 
                         (N166)? rf_reg_tmp[568] : 
                         (N168)? rf_reg_tmp[600] : 
                         (N170)? rf_reg_tmp[632] : 
                         (N172)? rf_reg_tmp[664] : 
                         (N174)? rf_reg_tmp[696] : 
                         (N176)? rf_reg_tmp[728] : 
                         (N178)? rf_reg_tmp[760] : 
                         (N180)? rf_reg_tmp[792] : 
                         (N182)? rf_reg_tmp[824] : 
                         (N184)? rf_reg_tmp[856] : 
                         (N186)? rf_reg_tmp[888] : 
                         (N188)? rf_reg_tmp[920] : 
                         (N190)? rf_reg_tmp[952] : 
                         (N192)? rf_reg_tmp[984] : 1'b0;
  assign rdata_b_o[23] = (N161)? 1'b0 : 
                         (N163)? rf_reg_tmp[23] : 
                         (N165)? rf_reg_tmp[55] : 
                         (N167)? rf_reg_tmp[87] : 
                         (N169)? rf_reg_tmp[119] : 
                         (N171)? rf_reg_tmp[151] : 
                         (N173)? rf_reg_tmp[183] : 
                         (N175)? rf_reg_tmp[215] : 
                         (N177)? rf_reg_tmp[247] : 
                         (N179)? rf_reg_tmp[279] : 
                         (N181)? rf_reg_tmp[311] : 
                         (N183)? rf_reg_tmp[343] : 
                         (N185)? rf_reg_tmp[375] : 
                         (N187)? rf_reg_tmp[407] : 
                         (N189)? rf_reg_tmp[439] : 
                         (N191)? rf_reg_tmp[471] : 
                         (N162)? rf_reg_tmp[503] : 
                         (N164)? rf_reg_tmp[535] : 
                         (N166)? rf_reg_tmp[567] : 
                         (N168)? rf_reg_tmp[599] : 
                         (N170)? rf_reg_tmp[631] : 
                         (N172)? rf_reg_tmp[663] : 
                         (N174)? rf_reg_tmp[695] : 
                         (N176)? rf_reg_tmp[727] : 
                         (N178)? rf_reg_tmp[759] : 
                         (N180)? rf_reg_tmp[791] : 
                         (N182)? rf_reg_tmp[823] : 
                         (N184)? rf_reg_tmp[855] : 
                         (N186)? rf_reg_tmp[887] : 
                         (N188)? rf_reg_tmp[919] : 
                         (N190)? rf_reg_tmp[951] : 
                         (N192)? rf_reg_tmp[983] : 1'b0;
  assign rdata_b_o[22] = (N161)? 1'b0 : 
                         (N163)? rf_reg_tmp[22] : 
                         (N165)? rf_reg_tmp[54] : 
                         (N167)? rf_reg_tmp[86] : 
                         (N169)? rf_reg_tmp[118] : 
                         (N171)? rf_reg_tmp[150] : 
                         (N173)? rf_reg_tmp[182] : 
                         (N175)? rf_reg_tmp[214] : 
                         (N177)? rf_reg_tmp[246] : 
                         (N179)? rf_reg_tmp[278] : 
                         (N181)? rf_reg_tmp[310] : 
                         (N183)? rf_reg_tmp[342] : 
                         (N185)? rf_reg_tmp[374] : 
                         (N187)? rf_reg_tmp[406] : 
                         (N189)? rf_reg_tmp[438] : 
                         (N191)? rf_reg_tmp[470] : 
                         (N162)? rf_reg_tmp[502] : 
                         (N164)? rf_reg_tmp[534] : 
                         (N166)? rf_reg_tmp[566] : 
                         (N168)? rf_reg_tmp[598] : 
                         (N170)? rf_reg_tmp[630] : 
                         (N172)? rf_reg_tmp[662] : 
                         (N174)? rf_reg_tmp[694] : 
                         (N176)? rf_reg_tmp[726] : 
                         (N178)? rf_reg_tmp[758] : 
                         (N180)? rf_reg_tmp[790] : 
                         (N182)? rf_reg_tmp[822] : 
                         (N184)? rf_reg_tmp[854] : 
                         (N186)? rf_reg_tmp[886] : 
                         (N188)? rf_reg_tmp[918] : 
                         (N190)? rf_reg_tmp[950] : 
                         (N192)? rf_reg_tmp[982] : 1'b0;
  assign rdata_b_o[21] = (N161)? 1'b0 : 
                         (N163)? rf_reg_tmp[21] : 
                         (N165)? rf_reg_tmp[53] : 
                         (N167)? rf_reg_tmp[85] : 
                         (N169)? rf_reg_tmp[117] : 
                         (N171)? rf_reg_tmp[149] : 
                         (N173)? rf_reg_tmp[181] : 
                         (N175)? rf_reg_tmp[213] : 
                         (N177)? rf_reg_tmp[245] : 
                         (N179)? rf_reg_tmp[277] : 
                         (N181)? rf_reg_tmp[309] : 
                         (N183)? rf_reg_tmp[341] : 
                         (N185)? rf_reg_tmp[373] : 
                         (N187)? rf_reg_tmp[405] : 
                         (N189)? rf_reg_tmp[437] : 
                         (N191)? rf_reg_tmp[469] : 
                         (N162)? rf_reg_tmp[501] : 
                         (N164)? rf_reg_tmp[533] : 
                         (N166)? rf_reg_tmp[565] : 
                         (N168)? rf_reg_tmp[597] : 
                         (N170)? rf_reg_tmp[629] : 
                         (N172)? rf_reg_tmp[661] : 
                         (N174)? rf_reg_tmp[693] : 
                         (N176)? rf_reg_tmp[725] : 
                         (N178)? rf_reg_tmp[757] : 
                         (N180)? rf_reg_tmp[789] : 
                         (N182)? rf_reg_tmp[821] : 
                         (N184)? rf_reg_tmp[853] : 
                         (N186)? rf_reg_tmp[885] : 
                         (N188)? rf_reg_tmp[917] : 
                         (N190)? rf_reg_tmp[949] : 
                         (N192)? rf_reg_tmp[981] : 1'b0;
  assign rdata_b_o[20] = (N161)? 1'b0 : 
                         (N163)? rf_reg_tmp[20] : 
                         (N165)? rf_reg_tmp[52] : 
                         (N167)? rf_reg_tmp[84] : 
                         (N169)? rf_reg_tmp[116] : 
                         (N171)? rf_reg_tmp[148] : 
                         (N173)? rf_reg_tmp[180] : 
                         (N175)? rf_reg_tmp[212] : 
                         (N177)? rf_reg_tmp[244] : 
                         (N179)? rf_reg_tmp[276] : 
                         (N181)? rf_reg_tmp[308] : 
                         (N183)? rf_reg_tmp[340] : 
                         (N185)? rf_reg_tmp[372] : 
                         (N187)? rf_reg_tmp[404] : 
                         (N189)? rf_reg_tmp[436] : 
                         (N191)? rf_reg_tmp[468] : 
                         (N162)? rf_reg_tmp[500] : 
                         (N164)? rf_reg_tmp[532] : 
                         (N166)? rf_reg_tmp[564] : 
                         (N168)? rf_reg_tmp[596] : 
                         (N170)? rf_reg_tmp[628] : 
                         (N172)? rf_reg_tmp[660] : 
                         (N174)? rf_reg_tmp[692] : 
                         (N176)? rf_reg_tmp[724] : 
                         (N178)? rf_reg_tmp[756] : 
                         (N180)? rf_reg_tmp[788] : 
                         (N182)? rf_reg_tmp[820] : 
                         (N184)? rf_reg_tmp[852] : 
                         (N186)? rf_reg_tmp[884] : 
                         (N188)? rf_reg_tmp[916] : 
                         (N190)? rf_reg_tmp[948] : 
                         (N192)? rf_reg_tmp[980] : 1'b0;
  assign rdata_b_o[19] = (N161)? 1'b0 : 
                         (N163)? rf_reg_tmp[19] : 
                         (N165)? rf_reg_tmp[51] : 
                         (N167)? rf_reg_tmp[83] : 
                         (N169)? rf_reg_tmp[115] : 
                         (N171)? rf_reg_tmp[147] : 
                         (N173)? rf_reg_tmp[179] : 
                         (N175)? rf_reg_tmp[211] : 
                         (N177)? rf_reg_tmp[243] : 
                         (N179)? rf_reg_tmp[275] : 
                         (N181)? rf_reg_tmp[307] : 
                         (N183)? rf_reg_tmp[339] : 
                         (N185)? rf_reg_tmp[371] : 
                         (N187)? rf_reg_tmp[403] : 
                         (N189)? rf_reg_tmp[435] : 
                         (N191)? rf_reg_tmp[467] : 
                         (N162)? rf_reg_tmp[499] : 
                         (N164)? rf_reg_tmp[531] : 
                         (N166)? rf_reg_tmp[563] : 
                         (N168)? rf_reg_tmp[595] : 
                         (N170)? rf_reg_tmp[627] : 
                         (N172)? rf_reg_tmp[659] : 
                         (N174)? rf_reg_tmp[691] : 
                         (N176)? rf_reg_tmp[723] : 
                         (N178)? rf_reg_tmp[755] : 
                         (N180)? rf_reg_tmp[787] : 
                         (N182)? rf_reg_tmp[819] : 
                         (N184)? rf_reg_tmp[851] : 
                         (N186)? rf_reg_tmp[883] : 
                         (N188)? rf_reg_tmp[915] : 
                         (N190)? rf_reg_tmp[947] : 
                         (N192)? rf_reg_tmp[979] : 1'b0;
  assign rdata_b_o[18] = (N161)? 1'b0 : 
                         (N163)? rf_reg_tmp[18] : 
                         (N165)? rf_reg_tmp[50] : 
                         (N167)? rf_reg_tmp[82] : 
                         (N169)? rf_reg_tmp[114] : 
                         (N171)? rf_reg_tmp[146] : 
                         (N173)? rf_reg_tmp[178] : 
                         (N175)? rf_reg_tmp[210] : 
                         (N177)? rf_reg_tmp[242] : 
                         (N179)? rf_reg_tmp[274] : 
                         (N181)? rf_reg_tmp[306] : 
                         (N183)? rf_reg_tmp[338] : 
                         (N185)? rf_reg_tmp[370] : 
                         (N187)? rf_reg_tmp[402] : 
                         (N189)? rf_reg_tmp[434] : 
                         (N191)? rf_reg_tmp[466] : 
                         (N162)? rf_reg_tmp[498] : 
                         (N164)? rf_reg_tmp[530] : 
                         (N166)? rf_reg_tmp[562] : 
                         (N168)? rf_reg_tmp[594] : 
                         (N170)? rf_reg_tmp[626] : 
                         (N172)? rf_reg_tmp[658] : 
                         (N174)? rf_reg_tmp[690] : 
                         (N176)? rf_reg_tmp[722] : 
                         (N178)? rf_reg_tmp[754] : 
                         (N180)? rf_reg_tmp[786] : 
                         (N182)? rf_reg_tmp[818] : 
                         (N184)? rf_reg_tmp[850] : 
                         (N186)? rf_reg_tmp[882] : 
                         (N188)? rf_reg_tmp[914] : 
                         (N190)? rf_reg_tmp[946] : 
                         (N192)? rf_reg_tmp[978] : 1'b0;
  assign rdata_b_o[17] = (N161)? 1'b0 : 
                         (N163)? rf_reg_tmp[17] : 
                         (N165)? rf_reg_tmp[49] : 
                         (N167)? rf_reg_tmp[81] : 
                         (N169)? rf_reg_tmp[113] : 
                         (N171)? rf_reg_tmp[145] : 
                         (N173)? rf_reg_tmp[177] : 
                         (N175)? rf_reg_tmp[209] : 
                         (N177)? rf_reg_tmp[241] : 
                         (N179)? rf_reg_tmp[273] : 
                         (N181)? rf_reg_tmp[305] : 
                         (N183)? rf_reg_tmp[337] : 
                         (N185)? rf_reg_tmp[369] : 
                         (N187)? rf_reg_tmp[401] : 
                         (N189)? rf_reg_tmp[433] : 
                         (N191)? rf_reg_tmp[465] : 
                         (N162)? rf_reg_tmp[497] : 
                         (N164)? rf_reg_tmp[529] : 
                         (N166)? rf_reg_tmp[561] : 
                         (N168)? rf_reg_tmp[593] : 
                         (N170)? rf_reg_tmp[625] : 
                         (N172)? rf_reg_tmp[657] : 
                         (N174)? rf_reg_tmp[689] : 
                         (N176)? rf_reg_tmp[721] : 
                         (N178)? rf_reg_tmp[753] : 
                         (N180)? rf_reg_tmp[785] : 
                         (N182)? rf_reg_tmp[817] : 
                         (N184)? rf_reg_tmp[849] : 
                         (N186)? rf_reg_tmp[881] : 
                         (N188)? rf_reg_tmp[913] : 
                         (N190)? rf_reg_tmp[945] : 
                         (N192)? rf_reg_tmp[977] : 1'b0;
  assign rdata_b_o[16] = (N161)? 1'b0 : 
                         (N163)? rf_reg_tmp[16] : 
                         (N165)? rf_reg_tmp[48] : 
                         (N167)? rf_reg_tmp[80] : 
                         (N169)? rf_reg_tmp[112] : 
                         (N171)? rf_reg_tmp[144] : 
                         (N173)? rf_reg_tmp[176] : 
                         (N175)? rf_reg_tmp[208] : 
                         (N177)? rf_reg_tmp[240] : 
                         (N179)? rf_reg_tmp[272] : 
                         (N181)? rf_reg_tmp[304] : 
                         (N183)? rf_reg_tmp[336] : 
                         (N185)? rf_reg_tmp[368] : 
                         (N187)? rf_reg_tmp[400] : 
                         (N189)? rf_reg_tmp[432] : 
                         (N191)? rf_reg_tmp[464] : 
                         (N162)? rf_reg_tmp[496] : 
                         (N164)? rf_reg_tmp[528] : 
                         (N166)? rf_reg_tmp[560] : 
                         (N168)? rf_reg_tmp[592] : 
                         (N170)? rf_reg_tmp[624] : 
                         (N172)? rf_reg_tmp[656] : 
                         (N174)? rf_reg_tmp[688] : 
                         (N176)? rf_reg_tmp[720] : 
                         (N178)? rf_reg_tmp[752] : 
                         (N180)? rf_reg_tmp[784] : 
                         (N182)? rf_reg_tmp[816] : 
                         (N184)? rf_reg_tmp[848] : 
                         (N186)? rf_reg_tmp[880] : 
                         (N188)? rf_reg_tmp[912] : 
                         (N190)? rf_reg_tmp[944] : 
                         (N192)? rf_reg_tmp[976] : 1'b0;
  assign rdata_b_o[15] = (N161)? 1'b0 : 
                         (N163)? rf_reg_tmp[15] : 
                         (N165)? rf_reg_tmp[47] : 
                         (N167)? rf_reg_tmp[79] : 
                         (N169)? rf_reg_tmp[111] : 
                         (N171)? rf_reg_tmp[143] : 
                         (N173)? rf_reg_tmp[175] : 
                         (N175)? rf_reg_tmp[207] : 
                         (N177)? rf_reg_tmp[239] : 
                         (N179)? rf_reg_tmp[271] : 
                         (N181)? rf_reg_tmp[303] : 
                         (N183)? rf_reg_tmp[335] : 
                         (N185)? rf_reg_tmp[367] : 
                         (N187)? rf_reg_tmp[399] : 
                         (N189)? rf_reg_tmp[431] : 
                         (N191)? rf_reg_tmp[463] : 
                         (N162)? rf_reg_tmp[495] : 
                         (N164)? rf_reg_tmp[527] : 
                         (N166)? rf_reg_tmp[559] : 
                         (N168)? rf_reg_tmp[591] : 
                         (N170)? rf_reg_tmp[623] : 
                         (N172)? rf_reg_tmp[655] : 
                         (N174)? rf_reg_tmp[687] : 
                         (N176)? rf_reg_tmp[719] : 
                         (N178)? rf_reg_tmp[751] : 
                         (N180)? rf_reg_tmp[783] : 
                         (N182)? rf_reg_tmp[815] : 
                         (N184)? rf_reg_tmp[847] : 
                         (N186)? rf_reg_tmp[879] : 
                         (N188)? rf_reg_tmp[911] : 
                         (N190)? rf_reg_tmp[943] : 
                         (N192)? rf_reg_tmp[975] : 1'b0;
  assign rdata_b_o[14] = (N161)? 1'b0 : 
                         (N163)? rf_reg_tmp[14] : 
                         (N165)? rf_reg_tmp[46] : 
                         (N167)? rf_reg_tmp[78] : 
                         (N169)? rf_reg_tmp[110] : 
                         (N171)? rf_reg_tmp[142] : 
                         (N173)? rf_reg_tmp[174] : 
                         (N175)? rf_reg_tmp[206] : 
                         (N177)? rf_reg_tmp[238] : 
                         (N179)? rf_reg_tmp[270] : 
                         (N181)? rf_reg_tmp[302] : 
                         (N183)? rf_reg_tmp[334] : 
                         (N185)? rf_reg_tmp[366] : 
                         (N187)? rf_reg_tmp[398] : 
                         (N189)? rf_reg_tmp[430] : 
                         (N191)? rf_reg_tmp[462] : 
                         (N162)? rf_reg_tmp[494] : 
                         (N164)? rf_reg_tmp[526] : 
                         (N166)? rf_reg_tmp[558] : 
                         (N168)? rf_reg_tmp[590] : 
                         (N170)? rf_reg_tmp[622] : 
                         (N172)? rf_reg_tmp[654] : 
                         (N174)? rf_reg_tmp[686] : 
                         (N176)? rf_reg_tmp[718] : 
                         (N178)? rf_reg_tmp[750] : 
                         (N180)? rf_reg_tmp[782] : 
                         (N182)? rf_reg_tmp[814] : 
                         (N184)? rf_reg_tmp[846] : 
                         (N186)? rf_reg_tmp[878] : 
                         (N188)? rf_reg_tmp[910] : 
                         (N190)? rf_reg_tmp[942] : 
                         (N192)? rf_reg_tmp[974] : 1'b0;
  assign rdata_b_o[13] = (N161)? 1'b0 : 
                         (N163)? rf_reg_tmp[13] : 
                         (N165)? rf_reg_tmp[45] : 
                         (N167)? rf_reg_tmp[77] : 
                         (N169)? rf_reg_tmp[109] : 
                         (N171)? rf_reg_tmp[141] : 
                         (N173)? rf_reg_tmp[173] : 
                         (N175)? rf_reg_tmp[205] : 
                         (N177)? rf_reg_tmp[237] : 
                         (N179)? rf_reg_tmp[269] : 
                         (N181)? rf_reg_tmp[301] : 
                         (N183)? rf_reg_tmp[333] : 
                         (N185)? rf_reg_tmp[365] : 
                         (N187)? rf_reg_tmp[397] : 
                         (N189)? rf_reg_tmp[429] : 
                         (N191)? rf_reg_tmp[461] : 
                         (N162)? rf_reg_tmp[493] : 
                         (N164)? rf_reg_tmp[525] : 
                         (N166)? rf_reg_tmp[557] : 
                         (N168)? rf_reg_tmp[589] : 
                         (N170)? rf_reg_tmp[621] : 
                         (N172)? rf_reg_tmp[653] : 
                         (N174)? rf_reg_tmp[685] : 
                         (N176)? rf_reg_tmp[717] : 
                         (N178)? rf_reg_tmp[749] : 
                         (N180)? rf_reg_tmp[781] : 
                         (N182)? rf_reg_tmp[813] : 
                         (N184)? rf_reg_tmp[845] : 
                         (N186)? rf_reg_tmp[877] : 
                         (N188)? rf_reg_tmp[909] : 
                         (N190)? rf_reg_tmp[941] : 
                         (N192)? rf_reg_tmp[973] : 1'b0;
  assign rdata_b_o[12] = (N161)? 1'b0 : 
                         (N163)? rf_reg_tmp[12] : 
                         (N165)? rf_reg_tmp[44] : 
                         (N167)? rf_reg_tmp[76] : 
                         (N169)? rf_reg_tmp[108] : 
                         (N171)? rf_reg_tmp[140] : 
                         (N173)? rf_reg_tmp[172] : 
                         (N175)? rf_reg_tmp[204] : 
                         (N177)? rf_reg_tmp[236] : 
                         (N179)? rf_reg_tmp[268] : 
                         (N181)? rf_reg_tmp[300] : 
                         (N183)? rf_reg_tmp[332] : 
                         (N185)? rf_reg_tmp[364] : 
                         (N187)? rf_reg_tmp[396] : 
                         (N189)? rf_reg_tmp[428] : 
                         (N191)? rf_reg_tmp[460] : 
                         (N162)? rf_reg_tmp[492] : 
                         (N164)? rf_reg_tmp[524] : 
                         (N166)? rf_reg_tmp[556] : 
                         (N168)? rf_reg_tmp[588] : 
                         (N170)? rf_reg_tmp[620] : 
                         (N172)? rf_reg_tmp[652] : 
                         (N174)? rf_reg_tmp[684] : 
                         (N176)? rf_reg_tmp[716] : 
                         (N178)? rf_reg_tmp[748] : 
                         (N180)? rf_reg_tmp[780] : 
                         (N182)? rf_reg_tmp[812] : 
                         (N184)? rf_reg_tmp[844] : 
                         (N186)? rf_reg_tmp[876] : 
                         (N188)? rf_reg_tmp[908] : 
                         (N190)? rf_reg_tmp[940] : 
                         (N192)? rf_reg_tmp[972] : 1'b0;
  assign rdata_b_o[11] = (N161)? 1'b0 : 
                         (N163)? rf_reg_tmp[11] : 
                         (N165)? rf_reg_tmp[43] : 
                         (N167)? rf_reg_tmp[75] : 
                         (N169)? rf_reg_tmp[107] : 
                         (N171)? rf_reg_tmp[139] : 
                         (N173)? rf_reg_tmp[171] : 
                         (N175)? rf_reg_tmp[203] : 
                         (N177)? rf_reg_tmp[235] : 
                         (N179)? rf_reg_tmp[267] : 
                         (N181)? rf_reg_tmp[299] : 
                         (N183)? rf_reg_tmp[331] : 
                         (N185)? rf_reg_tmp[363] : 
                         (N187)? rf_reg_tmp[395] : 
                         (N189)? rf_reg_tmp[427] : 
                         (N191)? rf_reg_tmp[459] : 
                         (N162)? rf_reg_tmp[491] : 
                         (N164)? rf_reg_tmp[523] : 
                         (N166)? rf_reg_tmp[555] : 
                         (N168)? rf_reg_tmp[587] : 
                         (N170)? rf_reg_tmp[619] : 
                         (N172)? rf_reg_tmp[651] : 
                         (N174)? rf_reg_tmp[683] : 
                         (N176)? rf_reg_tmp[715] : 
                         (N178)? rf_reg_tmp[747] : 
                         (N180)? rf_reg_tmp[779] : 
                         (N182)? rf_reg_tmp[811] : 
                         (N184)? rf_reg_tmp[843] : 
                         (N186)? rf_reg_tmp[875] : 
                         (N188)? rf_reg_tmp[907] : 
                         (N190)? rf_reg_tmp[939] : 
                         (N192)? rf_reg_tmp[971] : 1'b0;
  assign rdata_b_o[10] = (N161)? 1'b0 : 
                         (N163)? rf_reg_tmp[10] : 
                         (N165)? rf_reg_tmp[42] : 
                         (N167)? rf_reg_tmp[74] : 
                         (N169)? rf_reg_tmp[106] : 
                         (N171)? rf_reg_tmp[138] : 
                         (N173)? rf_reg_tmp[170] : 
                         (N175)? rf_reg_tmp[202] : 
                         (N177)? rf_reg_tmp[234] : 
                         (N179)? rf_reg_tmp[266] : 
                         (N181)? rf_reg_tmp[298] : 
                         (N183)? rf_reg_tmp[330] : 
                         (N185)? rf_reg_tmp[362] : 
                         (N187)? rf_reg_tmp[394] : 
                         (N189)? rf_reg_tmp[426] : 
                         (N191)? rf_reg_tmp[458] : 
                         (N162)? rf_reg_tmp[490] : 
                         (N164)? rf_reg_tmp[522] : 
                         (N166)? rf_reg_tmp[554] : 
                         (N168)? rf_reg_tmp[586] : 
                         (N170)? rf_reg_tmp[618] : 
                         (N172)? rf_reg_tmp[650] : 
                         (N174)? rf_reg_tmp[682] : 
                         (N176)? rf_reg_tmp[714] : 
                         (N178)? rf_reg_tmp[746] : 
                         (N180)? rf_reg_tmp[778] : 
                         (N182)? rf_reg_tmp[810] : 
                         (N184)? rf_reg_tmp[842] : 
                         (N186)? rf_reg_tmp[874] : 
                         (N188)? rf_reg_tmp[906] : 
                         (N190)? rf_reg_tmp[938] : 
                         (N192)? rf_reg_tmp[970] : 1'b0;
  assign rdata_b_o[9] = (N161)? 1'b0 : 
                        (N163)? rf_reg_tmp[9] : 
                        (N165)? rf_reg_tmp[41] : 
                        (N167)? rf_reg_tmp[73] : 
                        (N169)? rf_reg_tmp[105] : 
                        (N171)? rf_reg_tmp[137] : 
                        (N173)? rf_reg_tmp[169] : 
                        (N175)? rf_reg_tmp[201] : 
                        (N177)? rf_reg_tmp[233] : 
                        (N179)? rf_reg_tmp[265] : 
                        (N181)? rf_reg_tmp[297] : 
                        (N183)? rf_reg_tmp[329] : 
                        (N185)? rf_reg_tmp[361] : 
                        (N187)? rf_reg_tmp[393] : 
                        (N189)? rf_reg_tmp[425] : 
                        (N191)? rf_reg_tmp[457] : 
                        (N162)? rf_reg_tmp[489] : 
                        (N164)? rf_reg_tmp[521] : 
                        (N166)? rf_reg_tmp[553] : 
                        (N168)? rf_reg_tmp[585] : 
                        (N170)? rf_reg_tmp[617] : 
                        (N172)? rf_reg_tmp[649] : 
                        (N174)? rf_reg_tmp[681] : 
                        (N176)? rf_reg_tmp[713] : 
                        (N178)? rf_reg_tmp[745] : 
                        (N180)? rf_reg_tmp[777] : 
                        (N182)? rf_reg_tmp[809] : 
                        (N184)? rf_reg_tmp[841] : 
                        (N186)? rf_reg_tmp[873] : 
                        (N188)? rf_reg_tmp[905] : 
                        (N190)? rf_reg_tmp[937] : 
                        (N192)? rf_reg_tmp[969] : 1'b0;
  assign rdata_b_o[8] = (N161)? 1'b0 : 
                        (N163)? rf_reg_tmp[8] : 
                        (N165)? rf_reg_tmp[40] : 
                        (N167)? rf_reg_tmp[72] : 
                        (N169)? rf_reg_tmp[104] : 
                        (N171)? rf_reg_tmp[136] : 
                        (N173)? rf_reg_tmp[168] : 
                        (N175)? rf_reg_tmp[200] : 
                        (N177)? rf_reg_tmp[232] : 
                        (N179)? rf_reg_tmp[264] : 
                        (N181)? rf_reg_tmp[296] : 
                        (N183)? rf_reg_tmp[328] : 
                        (N185)? rf_reg_tmp[360] : 
                        (N187)? rf_reg_tmp[392] : 
                        (N189)? rf_reg_tmp[424] : 
                        (N191)? rf_reg_tmp[456] : 
                        (N162)? rf_reg_tmp[488] : 
                        (N164)? rf_reg_tmp[520] : 
                        (N166)? rf_reg_tmp[552] : 
                        (N168)? rf_reg_tmp[584] : 
                        (N170)? rf_reg_tmp[616] : 
                        (N172)? rf_reg_tmp[648] : 
                        (N174)? rf_reg_tmp[680] : 
                        (N176)? rf_reg_tmp[712] : 
                        (N178)? rf_reg_tmp[744] : 
                        (N180)? rf_reg_tmp[776] : 
                        (N182)? rf_reg_tmp[808] : 
                        (N184)? rf_reg_tmp[840] : 
                        (N186)? rf_reg_tmp[872] : 
                        (N188)? rf_reg_tmp[904] : 
                        (N190)? rf_reg_tmp[936] : 
                        (N192)? rf_reg_tmp[968] : 1'b0;
  assign rdata_b_o[7] = (N161)? 1'b0 : 
                        (N163)? rf_reg_tmp[7] : 
                        (N165)? rf_reg_tmp[39] : 
                        (N167)? rf_reg_tmp[71] : 
                        (N169)? rf_reg_tmp[103] : 
                        (N171)? rf_reg_tmp[135] : 
                        (N173)? rf_reg_tmp[167] : 
                        (N175)? rf_reg_tmp[199] : 
                        (N177)? rf_reg_tmp[231] : 
                        (N179)? rf_reg_tmp[263] : 
                        (N181)? rf_reg_tmp[295] : 
                        (N183)? rf_reg_tmp[327] : 
                        (N185)? rf_reg_tmp[359] : 
                        (N187)? rf_reg_tmp[391] : 
                        (N189)? rf_reg_tmp[423] : 
                        (N191)? rf_reg_tmp[455] : 
                        (N162)? rf_reg_tmp[487] : 
                        (N164)? rf_reg_tmp[519] : 
                        (N166)? rf_reg_tmp[551] : 
                        (N168)? rf_reg_tmp[583] : 
                        (N170)? rf_reg_tmp[615] : 
                        (N172)? rf_reg_tmp[647] : 
                        (N174)? rf_reg_tmp[679] : 
                        (N176)? rf_reg_tmp[711] : 
                        (N178)? rf_reg_tmp[743] : 
                        (N180)? rf_reg_tmp[775] : 
                        (N182)? rf_reg_tmp[807] : 
                        (N184)? rf_reg_tmp[839] : 
                        (N186)? rf_reg_tmp[871] : 
                        (N188)? rf_reg_tmp[903] : 
                        (N190)? rf_reg_tmp[935] : 
                        (N192)? rf_reg_tmp[967] : 1'b0;
  assign rdata_b_o[6] = (N161)? 1'b0 : 
                        (N163)? rf_reg_tmp[6] : 
                        (N165)? rf_reg_tmp[38] : 
                        (N167)? rf_reg_tmp[70] : 
                        (N169)? rf_reg_tmp[102] : 
                        (N171)? rf_reg_tmp[134] : 
                        (N173)? rf_reg_tmp[166] : 
                        (N175)? rf_reg_tmp[198] : 
                        (N177)? rf_reg_tmp[230] : 
                        (N179)? rf_reg_tmp[262] : 
                        (N181)? rf_reg_tmp[294] : 
                        (N183)? rf_reg_tmp[326] : 
                        (N185)? rf_reg_tmp[358] : 
                        (N187)? rf_reg_tmp[390] : 
                        (N189)? rf_reg_tmp[422] : 
                        (N191)? rf_reg_tmp[454] : 
                        (N162)? rf_reg_tmp[486] : 
                        (N164)? rf_reg_tmp[518] : 
                        (N166)? rf_reg_tmp[550] : 
                        (N168)? rf_reg_tmp[582] : 
                        (N170)? rf_reg_tmp[614] : 
                        (N172)? rf_reg_tmp[646] : 
                        (N174)? rf_reg_tmp[678] : 
                        (N176)? rf_reg_tmp[710] : 
                        (N178)? rf_reg_tmp[742] : 
                        (N180)? rf_reg_tmp[774] : 
                        (N182)? rf_reg_tmp[806] : 
                        (N184)? rf_reg_tmp[838] : 
                        (N186)? rf_reg_tmp[870] : 
                        (N188)? rf_reg_tmp[902] : 
                        (N190)? rf_reg_tmp[934] : 
                        (N192)? rf_reg_tmp[966] : 1'b0;
  assign rdata_b_o[5] = (N161)? 1'b0 : 
                        (N163)? rf_reg_tmp[5] : 
                        (N165)? rf_reg_tmp[37] : 
                        (N167)? rf_reg_tmp[69] : 
                        (N169)? rf_reg_tmp[101] : 
                        (N171)? rf_reg_tmp[133] : 
                        (N173)? rf_reg_tmp[165] : 
                        (N175)? rf_reg_tmp[197] : 
                        (N177)? rf_reg_tmp[229] : 
                        (N179)? rf_reg_tmp[261] : 
                        (N181)? rf_reg_tmp[293] : 
                        (N183)? rf_reg_tmp[325] : 
                        (N185)? rf_reg_tmp[357] : 
                        (N187)? rf_reg_tmp[389] : 
                        (N189)? rf_reg_tmp[421] : 
                        (N191)? rf_reg_tmp[453] : 
                        (N162)? rf_reg_tmp[485] : 
                        (N164)? rf_reg_tmp[517] : 
                        (N166)? rf_reg_tmp[549] : 
                        (N168)? rf_reg_tmp[581] : 
                        (N170)? rf_reg_tmp[613] : 
                        (N172)? rf_reg_tmp[645] : 
                        (N174)? rf_reg_tmp[677] : 
                        (N176)? rf_reg_tmp[709] : 
                        (N178)? rf_reg_tmp[741] : 
                        (N180)? rf_reg_tmp[773] : 
                        (N182)? rf_reg_tmp[805] : 
                        (N184)? rf_reg_tmp[837] : 
                        (N186)? rf_reg_tmp[869] : 
                        (N188)? rf_reg_tmp[901] : 
                        (N190)? rf_reg_tmp[933] : 
                        (N192)? rf_reg_tmp[965] : 1'b0;
  assign rdata_b_o[4] = (N161)? 1'b0 : 
                        (N163)? rf_reg_tmp[4] : 
                        (N165)? rf_reg_tmp[36] : 
                        (N167)? rf_reg_tmp[68] : 
                        (N169)? rf_reg_tmp[100] : 
                        (N171)? rf_reg_tmp[132] : 
                        (N173)? rf_reg_tmp[164] : 
                        (N175)? rf_reg_tmp[196] : 
                        (N177)? rf_reg_tmp[228] : 
                        (N179)? rf_reg_tmp[260] : 
                        (N181)? rf_reg_tmp[292] : 
                        (N183)? rf_reg_tmp[324] : 
                        (N185)? rf_reg_tmp[356] : 
                        (N187)? rf_reg_tmp[388] : 
                        (N189)? rf_reg_tmp[420] : 
                        (N191)? rf_reg_tmp[452] : 
                        (N162)? rf_reg_tmp[484] : 
                        (N164)? rf_reg_tmp[516] : 
                        (N166)? rf_reg_tmp[548] : 
                        (N168)? rf_reg_tmp[580] : 
                        (N170)? rf_reg_tmp[612] : 
                        (N172)? rf_reg_tmp[644] : 
                        (N174)? rf_reg_tmp[676] : 
                        (N176)? rf_reg_tmp[708] : 
                        (N178)? rf_reg_tmp[740] : 
                        (N180)? rf_reg_tmp[772] : 
                        (N182)? rf_reg_tmp[804] : 
                        (N184)? rf_reg_tmp[836] : 
                        (N186)? rf_reg_tmp[868] : 
                        (N188)? rf_reg_tmp[900] : 
                        (N190)? rf_reg_tmp[932] : 
                        (N192)? rf_reg_tmp[964] : 1'b0;
  assign rdata_b_o[3] = (N161)? 1'b0 : 
                        (N163)? rf_reg_tmp[3] : 
                        (N165)? rf_reg_tmp[35] : 
                        (N167)? rf_reg_tmp[67] : 
                        (N169)? rf_reg_tmp[99] : 
                        (N171)? rf_reg_tmp[131] : 
                        (N173)? rf_reg_tmp[163] : 
                        (N175)? rf_reg_tmp[195] : 
                        (N177)? rf_reg_tmp[227] : 
                        (N179)? rf_reg_tmp[259] : 
                        (N181)? rf_reg_tmp[291] : 
                        (N183)? rf_reg_tmp[323] : 
                        (N185)? rf_reg_tmp[355] : 
                        (N187)? rf_reg_tmp[387] : 
                        (N189)? rf_reg_tmp[419] : 
                        (N191)? rf_reg_tmp[451] : 
                        (N162)? rf_reg_tmp[483] : 
                        (N164)? rf_reg_tmp[515] : 
                        (N166)? rf_reg_tmp[547] : 
                        (N168)? rf_reg_tmp[579] : 
                        (N170)? rf_reg_tmp[611] : 
                        (N172)? rf_reg_tmp[643] : 
                        (N174)? rf_reg_tmp[675] : 
                        (N176)? rf_reg_tmp[707] : 
                        (N178)? rf_reg_tmp[739] : 
                        (N180)? rf_reg_tmp[771] : 
                        (N182)? rf_reg_tmp[803] : 
                        (N184)? rf_reg_tmp[835] : 
                        (N186)? rf_reg_tmp[867] : 
                        (N188)? rf_reg_tmp[899] : 
                        (N190)? rf_reg_tmp[931] : 
                        (N192)? rf_reg_tmp[963] : 1'b0;
  assign rdata_b_o[2] = (N161)? 1'b0 : 
                        (N163)? rf_reg_tmp[2] : 
                        (N165)? rf_reg_tmp[34] : 
                        (N167)? rf_reg_tmp[66] : 
                        (N169)? rf_reg_tmp[98] : 
                        (N171)? rf_reg_tmp[130] : 
                        (N173)? rf_reg_tmp[162] : 
                        (N175)? rf_reg_tmp[194] : 
                        (N177)? rf_reg_tmp[226] : 
                        (N179)? rf_reg_tmp[258] : 
                        (N181)? rf_reg_tmp[290] : 
                        (N183)? rf_reg_tmp[322] : 
                        (N185)? rf_reg_tmp[354] : 
                        (N187)? rf_reg_tmp[386] : 
                        (N189)? rf_reg_tmp[418] : 
                        (N191)? rf_reg_tmp[450] : 
                        (N162)? rf_reg_tmp[482] : 
                        (N164)? rf_reg_tmp[514] : 
                        (N166)? rf_reg_tmp[546] : 
                        (N168)? rf_reg_tmp[578] : 
                        (N170)? rf_reg_tmp[610] : 
                        (N172)? rf_reg_tmp[642] : 
                        (N174)? rf_reg_tmp[674] : 
                        (N176)? rf_reg_tmp[706] : 
                        (N178)? rf_reg_tmp[738] : 
                        (N180)? rf_reg_tmp[770] : 
                        (N182)? rf_reg_tmp[802] : 
                        (N184)? rf_reg_tmp[834] : 
                        (N186)? rf_reg_tmp[866] : 
                        (N188)? rf_reg_tmp[898] : 
                        (N190)? rf_reg_tmp[930] : 
                        (N192)? rf_reg_tmp[962] : 1'b0;
  assign rdata_b_o[1] = (N161)? 1'b0 : 
                        (N163)? rf_reg_tmp[1] : 
                        (N165)? rf_reg_tmp[33] : 
                        (N167)? rf_reg_tmp[65] : 
                        (N169)? rf_reg_tmp[97] : 
                        (N171)? rf_reg_tmp[129] : 
                        (N173)? rf_reg_tmp[161] : 
                        (N175)? rf_reg_tmp[193] : 
                        (N177)? rf_reg_tmp[225] : 
                        (N179)? rf_reg_tmp[257] : 
                        (N181)? rf_reg_tmp[289] : 
                        (N183)? rf_reg_tmp[321] : 
                        (N185)? rf_reg_tmp[353] : 
                        (N187)? rf_reg_tmp[385] : 
                        (N189)? rf_reg_tmp[417] : 
                        (N191)? rf_reg_tmp[449] : 
                        (N162)? rf_reg_tmp[481] : 
                        (N164)? rf_reg_tmp[513] : 
                        (N166)? rf_reg_tmp[545] : 
                        (N168)? rf_reg_tmp[577] : 
                        (N170)? rf_reg_tmp[609] : 
                        (N172)? rf_reg_tmp[641] : 
                        (N174)? rf_reg_tmp[673] : 
                        (N176)? rf_reg_tmp[705] : 
                        (N178)? rf_reg_tmp[737] : 
                        (N180)? rf_reg_tmp[769] : 
                        (N182)? rf_reg_tmp[801] : 
                        (N184)? rf_reg_tmp[833] : 
                        (N186)? rf_reg_tmp[865] : 
                        (N188)? rf_reg_tmp[897] : 
                        (N190)? rf_reg_tmp[929] : 
                        (N192)? rf_reg_tmp[961] : 1'b0;
  assign rdata_b_o[0] = (N161)? 1'b0 : 
                        (N163)? rf_reg_tmp[0] : 
                        (N165)? rf_reg_tmp[32] : 
                        (N167)? rf_reg_tmp[64] : 
                        (N169)? rf_reg_tmp[96] : 
                        (N171)? rf_reg_tmp[128] : 
                        (N173)? rf_reg_tmp[160] : 
                        (N175)? rf_reg_tmp[192] : 
                        (N177)? rf_reg_tmp[224] : 
                        (N179)? rf_reg_tmp[256] : 
                        (N181)? rf_reg_tmp[288] : 
                        (N183)? rf_reg_tmp[320] : 
                        (N185)? rf_reg_tmp[352] : 
                        (N187)? rf_reg_tmp[384] : 
                        (N189)? rf_reg_tmp[416] : 
                        (N191)? rf_reg_tmp[448] : 
                        (N162)? rf_reg_tmp[480] : 
                        (N164)? rf_reg_tmp[512] : 
                        (N166)? rf_reg_tmp[544] : 
                        (N168)? rf_reg_tmp[576] : 
                        (N170)? rf_reg_tmp[608] : 
                        (N172)? rf_reg_tmp[640] : 
                        (N174)? rf_reg_tmp[672] : 
                        (N176)? rf_reg_tmp[704] : 
                        (N178)? rf_reg_tmp[736] : 
                        (N180)? rf_reg_tmp[768] : 
                        (N182)? rf_reg_tmp[800] : 
                        (N184)? rf_reg_tmp[832] : 
                        (N186)? rf_reg_tmp[864] : 
                        (N188)? rf_reg_tmp[896] : 
                        (N190)? rf_reg_tmp[928] : 
                        (N192)? rf_reg_tmp[960] : 1'b0;
  assign N193 = waddr_a_i[3] & waddr_a_i[4];
  assign N194 = waddr_a_i[2] & N193;
  assign N195 = waddr_a_i[1] & N194;
  assign N196 = waddr_a_i[0] & N195;
  assign N197 = ~waddr_a_i[4];
  assign N198 = ~waddr_a_i[3];
  assign N199 = ~waddr_a_i[2];
  assign N200 = ~waddr_a_i[1];
  assign N201 = N198 | N197;
  assign N202 = N199 | N201;
  assign N203 = N200 | N202;
  assign N204 = waddr_a_i[0] | N203;
  assign N205 = ~N204;
  assign N206 = ~waddr_a_i[0];
  assign N207 = waddr_a_i[1] | N202;
  assign N208 = N206 | N207;
  assign N209 = ~N208;
  assign N210 = waddr_a_i[0] | N207;
  assign N211 = ~N210;
  assign N212 = waddr_a_i[2] | N201;
  assign N213 = N200 | N212;
  assign N214 = N206 | N213;
  assign N215 = ~N214;
  assign N216 = waddr_a_i[0] | N213;
  assign N217 = ~N216;
  assign N218 = waddr_a_i[1] | N212;
  assign N219 = N206 | N218;
  assign N220 = ~N219;
  assign N221 = waddr_a_i[0] | N218;
  assign N222 = ~N221;
  assign N223 = waddr_a_i[3] | N197;
  assign N224 = N199 | N223;
  assign N225 = N200 | N224;
  assign N226 = N206 | N225;
  assign N227 = ~N226;
  assign N228 = waddr_a_i[0] | N225;
  assign N229 = ~N228;
  assign N230 = waddr_a_i[1] | N224;
  assign N231 = N206 | N230;
  assign N232 = ~N231;
  assign N233 = waddr_a_i[0] | N230;
  assign N234 = ~N233;
  assign N235 = waddr_a_i[2] | N223;
  assign N236 = N200 | N235;
  assign N237 = N206 | N236;
  assign N238 = ~N237;
  assign N239 = waddr_a_i[0] | N236;
  assign N240 = ~N239;
  assign N241 = waddr_a_i[1] | N235;
  assign N242 = N206 | N241;
  assign N243 = ~N242;
  assign N244 = waddr_a_i[0] | N241;
  assign N245 = ~N244;
  assign N246 = N198 | waddr_a_i[4];
  assign N247 = N199 | N246;
  assign N248 = N200 | N247;
  assign N249 = N206 | N248;
  assign N250 = ~N249;
  assign N251 = waddr_a_i[0] | N248;
  assign N252 = ~N251;
  assign N253 = waddr_a_i[1] | N247;
  assign N254 = N206 | N253;
  assign N255 = ~N254;
  assign N256 = waddr_a_i[0] | N253;
  assign N257 = ~N256;
  assign N258 = waddr_a_i[2] | N246;
  assign N259 = N200 | N258;
  assign N260 = N206 | N259;
  assign N261 = ~N260;
  assign N262 = waddr_a_i[0] | N259;
  assign N263 = ~N262;
  assign N264 = waddr_a_i[1] | N258;
  assign N265 = N206 | N264;
  assign N266 = ~N265;
  assign N267 = waddr_a_i[0] | N264;
  assign N268 = ~N267;
  assign N269 = waddr_a_i[3] | waddr_a_i[4];
  assign N270 = N199 | N269;
  assign N271 = N200 | N270;
  assign N272 = N206 | N271;
  assign N273 = ~N272;
  assign N274 = waddr_a_i[0] | N271;
  assign N275 = ~N274;
  assign N276 = waddr_a_i[1] | N270;
  assign N277 = N206 | N276;
  assign N278 = ~N277;
  assign N279 = waddr_a_i[0] | N276;
  assign N280 = ~N279;
  assign N281 = waddr_a_i[2] | N269;
  assign N282 = N200 | N281;
  assign N283 = N206 | N282;
  assign N284 = ~N283;
  assign N285 = waddr_a_i[0] | N282;
  assign N286 = ~N285;
  assign N287 = waddr_a_i[1] | N281;
  assign N288 = N206 | N287;
  assign N289 = ~N288;
  assign we_a_dec[1] = (N0)? we_a_i : 
                       (N1)? 1'b0 : 1'b0;
  assign N0 = N289;
  assign N1 = N288;
  assign we_a_dec[2] = (N2)? we_a_i : 
                       (N3)? 1'b0 : 1'b0;
  assign N2 = N286;
  assign N3 = N285;
  assign we_a_dec[3] = (N4)? we_a_i : 
                       (N5)? 1'b0 : 1'b0;
  assign N4 = N284;
  assign N5 = N283;
  assign we_a_dec[4] = (N6)? we_a_i : 
                       (N7)? 1'b0 : 1'b0;
  assign N6 = N280;
  assign N7 = N279;
  assign we_a_dec[5] = (N8)? we_a_i : 
                       (N9)? 1'b0 : 1'b0;
  assign N8 = N278;
  assign N9 = N277;
  assign we_a_dec[6] = (N10)? we_a_i : 
                       (N11)? 1'b0 : 1'b0;
  assign N10 = N275;
  assign N11 = N274;
  assign we_a_dec[7] = (N12)? we_a_i : 
                       (N13)? 1'b0 : 1'b0;
  assign N12 = N273;
  assign N13 = N272;
  assign we_a_dec[8] = (N14)? we_a_i : 
                       (N15)? 1'b0 : 1'b0;
  assign N14 = N268;
  assign N15 = N267;
  assign we_a_dec[9] = (N16)? we_a_i : 
                       (N17)? 1'b0 : 1'b0;
  assign N16 = N266;
  assign N17 = N265;
  assign we_a_dec[10] = (N18)? we_a_i : 
                        (N19)? 1'b0 : 1'b0;
  assign N18 = N263;
  assign N19 = N262;
  assign we_a_dec[11] = (N20)? we_a_i : 
                        (N21)? 1'b0 : 1'b0;
  assign N20 = N261;
  assign N21 = N260;
  assign we_a_dec[12] = (N22)? we_a_i : 
                        (N23)? 1'b0 : 1'b0;
  assign N22 = N257;
  assign N23 = N256;
  assign we_a_dec[13] = (N24)? we_a_i : 
                        (N25)? 1'b0 : 1'b0;
  assign N24 = N255;
  assign N25 = N254;
  assign we_a_dec[14] = (N26)? we_a_i : 
                        (N27)? 1'b0 : 1'b0;
  assign N26 = N252;
  assign N27 = N251;
  assign we_a_dec[15] = (N28)? we_a_i : 
                        (N29)? 1'b0 : 1'b0;
  assign N28 = N250;
  assign N29 = N249;
  assign we_a_dec[16] = (N30)? we_a_i : 
                        (N31)? 1'b0 : 1'b0;
  assign N30 = N245;
  assign N31 = N244;
  assign we_a_dec[17] = (N32)? we_a_i : 
                        (N33)? 1'b0 : 1'b0;
  assign N32 = N243;
  assign N33 = N242;
  assign we_a_dec[18] = (N34)? we_a_i : 
                        (N35)? 1'b0 : 1'b0;
  assign N34 = N240;
  assign N35 = N239;
  assign we_a_dec[19] = (N36)? we_a_i : 
                        (N37)? 1'b0 : 1'b0;
  assign N36 = N238;
  assign N37 = N237;
  assign we_a_dec[20] = (N38)? we_a_i : 
                        (N39)? 1'b0 : 1'b0;
  assign N38 = N234;
  assign N39 = N233;
  assign we_a_dec[21] = (N40)? we_a_i : 
                        (N41)? 1'b0 : 1'b0;
  assign N40 = N232;
  assign N41 = N231;
  assign we_a_dec[22] = (N42)? we_a_i : 
                        (N43)? 1'b0 : 1'b0;
  assign N42 = N229;
  assign N43 = N228;
  assign we_a_dec[23] = (N44)? we_a_i : 
                        (N45)? 1'b0 : 1'b0;
  assign N44 = N227;
  assign N45 = N226;
  assign we_a_dec[24] = (N46)? we_a_i : 
                        (N47)? 1'b0 : 1'b0;
  assign N46 = N222;
  assign N47 = N221;
  assign we_a_dec[25] = (N48)? we_a_i : 
                        (N49)? 1'b0 : 1'b0;
  assign N48 = N220;
  assign N49 = N219;
  assign we_a_dec[26] = (N50)? we_a_i : 
                        (N51)? 1'b0 : 1'b0;
  assign N50 = N217;
  assign N51 = N216;
  assign we_a_dec[27] = (N52)? we_a_i : 
                        (N53)? 1'b0 : 1'b0;
  assign N52 = N215;
  assign N53 = N214;
  assign we_a_dec[28] = (N54)? we_a_i : 
                        (N55)? 1'b0 : 1'b0;
  assign N54 = N211;
  assign N55 = N210;
  assign we_a_dec[29] = (N56)? we_a_i : 
                        (N57)? 1'b0 : 1'b0;
  assign N56 = N209;
  assign N57 = N208;
  assign we_a_dec[30] = (N58)? we_a_i : 
                        (N59)? 1'b0 : 1'b0;
  assign N58 = N205;
  assign N59 = N204;
  assign we_a_dec[31] = (N60)? we_a_i : 
                        (N61)? 1'b0 : 1'b0;
  assign N60 = N196;
  assign N61 = ~N196;
  assign N62 = ~rst_ni;
  assign N63 = ~raddr_a_i[0];
  assign N64 = ~raddr_a_i[1];
  assign N65 = N63 & N64;
  assign N66 = N63 & raddr_a_i[1];
  assign N67 = raddr_a_i[0] & N64;
  assign N68 = raddr_a_i[0] & raddr_a_i[1];
  assign N69 = ~raddr_a_i[2];
  assign N70 = N65 & N69;
  assign N71 = N65 & raddr_a_i[2];
  assign N72 = N67 & N69;
  assign N73 = N67 & raddr_a_i[2];
  assign N74 = N66 & N69;
  assign N75 = N66 & raddr_a_i[2];
  assign N76 = N68 & N69;
  assign N77 = N68 & raddr_a_i[2];
  assign N78 = ~raddr_a_i[3];
  assign N79 = N70 & N78;
  assign N80 = N70 & raddr_a_i[3];
  assign N81 = N72 & N78;
  assign N82 = N72 & raddr_a_i[3];
  assign N83 = N74 & N78;
  assign N84 = N74 & raddr_a_i[3];
  assign N85 = N76 & N78;
  assign N86 = N76 & raddr_a_i[3];
  assign N87 = N71 & N78;
  assign N88 = N71 & raddr_a_i[3];
  assign N89 = N73 & N78;
  assign N90 = N73 & raddr_a_i[3];
  assign N91 = N75 & N78;
  assign N92 = N75 & raddr_a_i[3];
  assign N93 = N77 & N78;
  assign N94 = N77 & raddr_a_i[3];
  assign N95 = ~raddr_a_i[4];
  assign N96 = N79 & N95;
  assign N97 = N79 & raddr_a_i[4];
  assign N98 = N81 & N95;
  assign N99 = N81 & raddr_a_i[4];
  assign N100 = N83 & N95;
  assign N101 = N83 & raddr_a_i[4];
  assign N102 = N85 & N95;
  assign N103 = N85 & raddr_a_i[4];
  assign N104 = N87 & N95;
  assign N105 = N87 & raddr_a_i[4];
  assign N106 = N89 & N95;
  assign N107 = N89 & raddr_a_i[4];
  assign N108 = N91 & N95;
  assign N109 = N91 & raddr_a_i[4];
  assign N110 = N93 & N95;
  assign N111 = N93 & raddr_a_i[4];
  assign N112 = N80 & N95;
  assign N113 = N80 & raddr_a_i[4];
  assign N114 = N82 & N95;
  assign N115 = N82 & raddr_a_i[4];
  assign N116 = N84 & N95;
  assign N117 = N84 & raddr_a_i[4];
  assign N118 = N86 & N95;
  assign N119 = N86 & raddr_a_i[4];
  assign N120 = N88 & N95;
  assign N121 = N88 & raddr_a_i[4];
  assign N122 = N90 & N95;
  assign N123 = N90 & raddr_a_i[4];
  assign N124 = N92 & N95;
  assign N125 = N92 & raddr_a_i[4];
  assign N126 = N94 & N95;
  assign N127 = N94 & raddr_a_i[4];
  assign N128 = ~raddr_b_i[0];
  assign N129 = ~raddr_b_i[1];
  assign N130 = N128 & N129;
  assign N131 = N128 & raddr_b_i[1];
  assign N132 = raddr_b_i[0] & N129;
  assign N133 = raddr_b_i[0] & raddr_b_i[1];
  assign N134 = ~raddr_b_i[2];
  assign N135 = N130 & N134;
  assign N136 = N130 & raddr_b_i[2];
  assign N137 = N132 & N134;
  assign N138 = N132 & raddr_b_i[2];
  assign N139 = N131 & N134;
  assign N140 = N131 & raddr_b_i[2];
  assign N141 = N133 & N134;
  assign N142 = N133 & raddr_b_i[2];
  assign N143 = ~raddr_b_i[3];
  assign N144 = N135 & N143;
  assign N145 = N135 & raddr_b_i[3];
  assign N146 = N137 & N143;
  assign N147 = N137 & raddr_b_i[3];
  assign N148 = N139 & N143;
  assign N149 = N139 & raddr_b_i[3];
  assign N150 = N141 & N143;
  assign N151 = N141 & raddr_b_i[3];
  assign N152 = N136 & N143;
  assign N153 = N136 & raddr_b_i[3];
  assign N154 = N138 & N143;
  assign N155 = N138 & raddr_b_i[3];
  assign N156 = N140 & N143;
  assign N157 = N140 & raddr_b_i[3];
  assign N158 = N142 & N143;
  assign N159 = N142 & raddr_b_i[3];
  assign N160 = ~raddr_b_i[4];
  assign N161 = N144 & N160;
  assign N162 = N144 & raddr_b_i[4];
  assign N163 = N146 & N160;
  assign N164 = N146 & raddr_b_i[4];
  assign N165 = N148 & N160;
  assign N166 = N148 & raddr_b_i[4];
  assign N167 = N150 & N160;
  assign N168 = N150 & raddr_b_i[4];
  assign N169 = N152 & N160;
  assign N170 = N152 & raddr_b_i[4];
  assign N171 = N154 & N160;
  assign N172 = N154 & raddr_b_i[4];
  assign N173 = N156 & N160;
  assign N174 = N156 & raddr_b_i[4];
  assign N175 = N158 & N160;
  assign N176 = N158 & raddr_b_i[4];
  assign N177 = N145 & N160;
  assign N178 = N145 & raddr_b_i[4];
  assign N179 = N147 & N160;
  assign N180 = N147 & raddr_b_i[4];
  assign N181 = N149 & N160;
  assign N182 = N149 & raddr_b_i[4];
  assign N183 = N151 & N160;
  assign N184 = N151 & raddr_b_i[4];
  assign N185 = N153 & N160;
  assign N186 = N153 & raddr_b_i[4];
  assign N187 = N155 & N160;
  assign N188 = N155 & raddr_b_i[4];
  assign N189 = N157 & N160;
  assign N190 = N157 & raddr_b_i[4];
  assign N191 = N159 & N160;
  assign N192 = N159 & raddr_b_i[4];

endmodule



module ibex_decoder_0_1
(
  illegal_insn_o,
  ebrk_insn_o,
  mret_insn_o,
  dret_insn_o,
  ecall_insn_o,
  wfi_insn_o,
  jump_set_o,
  instr_new_i,
  instr_rdata_i,
  illegal_c_insn_i,
  imm_a_mux_sel_o,
  imm_b_mux_sel_o,
  imm_i_type_o,
  imm_s_type_o,
  imm_b_type_o,
  imm_u_type_o,
  imm_j_type_o,
  zimm_rs1_type_o,
  regfile_wdata_sel_o,
  regfile_we_o,
  regfile_raddr_a_o,
  regfile_raddr_b_o,
  regfile_waddr_o,
  alu_operator_o,
  alu_op_a_mux_sel_o,
  alu_op_b_mux_sel_o,
  mult_en_o,
  div_en_o,
  multdiv_operator_o,
  multdiv_signed_mode_o,
  csr_access_o,
  csr_op_o,
  csr_status_o,
  data_req_o,
  data_we_o,
  data_type_o,
  data_sign_extension_o,
  data_reg_offset_o,
  jump_in_dec_o,
  branch_in_dec_o
);

  input [31:0] instr_rdata_i;
  output [2:0] imm_b_mux_sel_o;
  output [31:0] imm_i_type_o;
  output [31:0] imm_s_type_o;
  output [31:0] imm_b_type_o;
  output [31:0] imm_u_type_o;
  output [31:0] imm_j_type_o;
  output [31:0] zimm_rs1_type_o;
  output [1:0] regfile_wdata_sel_o;
  output [4:0] regfile_raddr_a_o;
  output [4:0] regfile_raddr_b_o;
  output [4:0] regfile_waddr_o;
  output [4:0] alu_operator_o;
  output [1:0] alu_op_a_mux_sel_o;
  output [1:0] multdiv_operator_o;
  output [1:0] multdiv_signed_mode_o;
  output [1:0] csr_op_o;
  output [1:0] data_type_o;
  output [1:0] data_reg_offset_o;
  input instr_new_i;
  input illegal_c_insn_i;
  output illegal_insn_o;
  output ebrk_insn_o;
  output mret_insn_o;
  output dret_insn_o;
  output ecall_insn_o;
  output wfi_insn_o;
  output jump_set_o;
  output imm_a_mux_sel_o;
  output regfile_we_o;
  output alu_op_b_mux_sel_o;
  output mult_en_o;
  output div_en_o;
  output csr_access_o;
  output csr_status_o;
  output data_req_o;
  output data_we_o;
  output data_sign_extension_o;
  output jump_in_dec_o;
  output branch_in_dec_o;
  wire [2:0] imm_b_mux_sel_o;
  wire [31:0] imm_i_type_o,imm_s_type_o,imm_b_type_o,imm_u_type_o,imm_j_type_o,
  zimm_rs1_type_o;
  wire [1:0] regfile_wdata_sel_o,alu_op_a_mux_sel_o,multdiv_operator_o,multdiv_signed_mode_o,
  csr_op_o,data_type_o,data_reg_offset_o,csr_op;
  wire [4:0] regfile_raddr_a_o,regfile_raddr_b_o,regfile_waddr_o,alu_operator_o;
  wire illegal_insn_o,ebrk_insn_o,mret_insn_o,dret_insn_o,ecall_insn_o,wfi_insn_o,
  jump_set_o,imm_a_mux_sel_o,regfile_we_o,alu_op_b_mux_sel_o,mult_en_o,div_en_o,
  csr_access_o,csr_status_o,data_req_o,data_we_o,data_sign_extension_o,jump_in_dec_o,
  branch_in_dec_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,
  N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,
  N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
  N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,
  N79,N80,N81,N82,regfile_we,illegal_insn,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,
  N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,
  N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,
  N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,
  N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,
  N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,
  N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,
  N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,
  N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,
  N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,
  N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,
  N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
  N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,
  N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,
  N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,
  N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,
  N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,
  N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,
  N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,
  N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,
  N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,
  N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,
  N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,
  N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,
  N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,
  N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,
  N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
  N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,
  N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,
  N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,
  N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
  N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,
  N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,
  N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,
  N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,
  N638,N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,
  N654,N655,N656,N657,N658;
  assign data_reg_offset_o[0] = 1'b0;
  assign data_reg_offset_o[1] = 1'b0;
  assign zimm_rs1_type_o[5] = 1'b0;
  assign zimm_rs1_type_o[6] = 1'b0;
  assign zimm_rs1_type_o[7] = 1'b0;
  assign zimm_rs1_type_o[8] = 1'b0;
  assign zimm_rs1_type_o[9] = 1'b0;
  assign zimm_rs1_type_o[10] = 1'b0;
  assign zimm_rs1_type_o[11] = 1'b0;
  assign zimm_rs1_type_o[12] = 1'b0;
  assign zimm_rs1_type_o[13] = 1'b0;
  assign zimm_rs1_type_o[14] = 1'b0;
  assign zimm_rs1_type_o[15] = 1'b0;
  assign zimm_rs1_type_o[16] = 1'b0;
  assign zimm_rs1_type_o[17] = 1'b0;
  assign zimm_rs1_type_o[18] = 1'b0;
  assign zimm_rs1_type_o[19] = 1'b0;
  assign zimm_rs1_type_o[20] = 1'b0;
  assign zimm_rs1_type_o[21] = 1'b0;
  assign zimm_rs1_type_o[22] = 1'b0;
  assign zimm_rs1_type_o[23] = 1'b0;
  assign zimm_rs1_type_o[24] = 1'b0;
  assign zimm_rs1_type_o[25] = 1'b0;
  assign zimm_rs1_type_o[26] = 1'b0;
  assign zimm_rs1_type_o[27] = 1'b0;
  assign zimm_rs1_type_o[28] = 1'b0;
  assign zimm_rs1_type_o[29] = 1'b0;
  assign zimm_rs1_type_o[30] = 1'b0;
  assign zimm_rs1_type_o[31] = 1'b0;
  assign imm_j_type_o[0] = 1'b0;
  assign imm_u_type_o[0] = 1'b0;
  assign imm_u_type_o[1] = 1'b0;
  assign imm_u_type_o[2] = 1'b0;
  assign imm_u_type_o[3] = 1'b0;
  assign imm_u_type_o[4] = 1'b0;
  assign imm_u_type_o[5] = 1'b0;
  assign imm_u_type_o[6] = 1'b0;
  assign imm_u_type_o[7] = 1'b0;
  assign imm_u_type_o[8] = 1'b0;
  assign imm_u_type_o[9] = 1'b0;
  assign imm_u_type_o[10] = 1'b0;
  assign imm_u_type_o[11] = 1'b0;
  assign imm_b_type_o[0] = 1'b0;
  assign imm_j_type_o[20] = instr_rdata_i[31];
  assign imm_j_type_o[21] = instr_rdata_i[31];
  assign imm_j_type_o[22] = instr_rdata_i[31];
  assign imm_j_type_o[23] = instr_rdata_i[31];
  assign imm_j_type_o[24] = instr_rdata_i[31];
  assign imm_j_type_o[25] = instr_rdata_i[31];
  assign imm_j_type_o[26] = instr_rdata_i[31];
  assign imm_j_type_o[27] = instr_rdata_i[31];
  assign imm_j_type_o[28] = instr_rdata_i[31];
  assign imm_j_type_o[29] = instr_rdata_i[31];
  assign imm_j_type_o[30] = instr_rdata_i[31];
  assign imm_j_type_o[31] = instr_rdata_i[31];
  assign imm_u_type_o[31] = instr_rdata_i[31];
  assign imm_b_type_o[12] = instr_rdata_i[31];
  assign imm_b_type_o[13] = instr_rdata_i[31];
  assign imm_b_type_o[14] = instr_rdata_i[31];
  assign imm_b_type_o[15] = instr_rdata_i[31];
  assign imm_b_type_o[16] = instr_rdata_i[31];
  assign imm_b_type_o[17] = instr_rdata_i[31];
  assign imm_b_type_o[18] = instr_rdata_i[31];
  assign imm_b_type_o[19] = instr_rdata_i[31];
  assign imm_b_type_o[20] = instr_rdata_i[31];
  assign imm_b_type_o[21] = instr_rdata_i[31];
  assign imm_b_type_o[22] = instr_rdata_i[31];
  assign imm_b_type_o[23] = instr_rdata_i[31];
  assign imm_b_type_o[24] = instr_rdata_i[31];
  assign imm_b_type_o[25] = instr_rdata_i[31];
  assign imm_b_type_o[26] = instr_rdata_i[31];
  assign imm_b_type_o[27] = instr_rdata_i[31];
  assign imm_b_type_o[28] = instr_rdata_i[31];
  assign imm_b_type_o[29] = instr_rdata_i[31];
  assign imm_b_type_o[30] = instr_rdata_i[31];
  assign imm_b_type_o[31] = instr_rdata_i[31];
  assign imm_s_type_o[11] = instr_rdata_i[31];
  assign imm_s_type_o[12] = instr_rdata_i[31];
  assign imm_s_type_o[13] = instr_rdata_i[31];
  assign imm_s_type_o[14] = instr_rdata_i[31];
  assign imm_s_type_o[15] = instr_rdata_i[31];
  assign imm_s_type_o[16] = instr_rdata_i[31];
  assign imm_s_type_o[17] = instr_rdata_i[31];
  assign imm_s_type_o[18] = instr_rdata_i[31];
  assign imm_s_type_o[19] = instr_rdata_i[31];
  assign imm_s_type_o[20] = instr_rdata_i[31];
  assign imm_s_type_o[21] = instr_rdata_i[31];
  assign imm_s_type_o[22] = instr_rdata_i[31];
  assign imm_s_type_o[23] = instr_rdata_i[31];
  assign imm_s_type_o[24] = instr_rdata_i[31];
  assign imm_s_type_o[25] = instr_rdata_i[31];
  assign imm_s_type_o[26] = instr_rdata_i[31];
  assign imm_s_type_o[27] = instr_rdata_i[31];
  assign imm_s_type_o[28] = instr_rdata_i[31];
  assign imm_s_type_o[29] = instr_rdata_i[31];
  assign imm_s_type_o[30] = instr_rdata_i[31];
  assign imm_s_type_o[31] = instr_rdata_i[31];
  assign imm_i_type_o[11] = instr_rdata_i[31];
  assign imm_i_type_o[12] = instr_rdata_i[31];
  assign imm_i_type_o[13] = instr_rdata_i[31];
  assign imm_i_type_o[14] = instr_rdata_i[31];
  assign imm_i_type_o[15] = instr_rdata_i[31];
  assign imm_i_type_o[16] = instr_rdata_i[31];
  assign imm_i_type_o[17] = instr_rdata_i[31];
  assign imm_i_type_o[18] = instr_rdata_i[31];
  assign imm_i_type_o[19] = instr_rdata_i[31];
  assign imm_i_type_o[20] = instr_rdata_i[31];
  assign imm_i_type_o[21] = instr_rdata_i[31];
  assign imm_i_type_o[22] = instr_rdata_i[31];
  assign imm_i_type_o[23] = instr_rdata_i[31];
  assign imm_i_type_o[24] = instr_rdata_i[31];
  assign imm_i_type_o[25] = instr_rdata_i[31];
  assign imm_i_type_o[26] = instr_rdata_i[31];
  assign imm_i_type_o[27] = instr_rdata_i[31];
  assign imm_i_type_o[28] = instr_rdata_i[31];
  assign imm_i_type_o[29] = instr_rdata_i[31];
  assign imm_i_type_o[30] = instr_rdata_i[31];
  assign imm_i_type_o[31] = instr_rdata_i[31];
  assign imm_j_type_o[10] = instr_rdata_i[30];
  assign imm_u_type_o[30] = instr_rdata_i[30];
  assign imm_b_type_o[10] = instr_rdata_i[30];
  assign imm_s_type_o[10] = instr_rdata_i[30];
  assign imm_i_type_o[10] = instr_rdata_i[30];
  assign imm_j_type_o[9] = instr_rdata_i[29];
  assign imm_u_type_o[29] = instr_rdata_i[29];
  assign imm_b_type_o[9] = instr_rdata_i[29];
  assign imm_s_type_o[9] = instr_rdata_i[29];
  assign imm_i_type_o[9] = instr_rdata_i[29];
  assign imm_j_type_o[8] = instr_rdata_i[28];
  assign imm_u_type_o[28] = instr_rdata_i[28];
  assign imm_b_type_o[8] = instr_rdata_i[28];
  assign imm_s_type_o[8] = instr_rdata_i[28];
  assign imm_i_type_o[8] = instr_rdata_i[28];
  assign imm_j_type_o[7] = instr_rdata_i[27];
  assign imm_u_type_o[27] = instr_rdata_i[27];
  assign imm_b_type_o[7] = instr_rdata_i[27];
  assign imm_s_type_o[7] = instr_rdata_i[27];
  assign imm_i_type_o[7] = instr_rdata_i[27];
  assign imm_j_type_o[6] = instr_rdata_i[26];
  assign imm_u_type_o[26] = instr_rdata_i[26];
  assign imm_b_type_o[6] = instr_rdata_i[26];
  assign imm_s_type_o[6] = instr_rdata_i[26];
  assign imm_i_type_o[6] = instr_rdata_i[26];
  assign imm_j_type_o[5] = instr_rdata_i[25];
  assign imm_u_type_o[25] = instr_rdata_i[25];
  assign imm_b_type_o[5] = instr_rdata_i[25];
  assign imm_s_type_o[5] = instr_rdata_i[25];
  assign imm_i_type_o[5] = instr_rdata_i[25];
  assign regfile_raddr_b_o[4] = instr_rdata_i[24];
  assign imm_j_type_o[4] = instr_rdata_i[24];
  assign imm_u_type_o[24] = instr_rdata_i[24];
  assign imm_i_type_o[4] = instr_rdata_i[24];
  assign regfile_raddr_b_o[3] = instr_rdata_i[23];
  assign imm_j_type_o[3] = instr_rdata_i[23];
  assign imm_u_type_o[23] = instr_rdata_i[23];
  assign imm_i_type_o[3] = instr_rdata_i[23];
  assign regfile_raddr_b_o[2] = instr_rdata_i[22];
  assign imm_j_type_o[2] = instr_rdata_i[22];
  assign imm_u_type_o[22] = instr_rdata_i[22];
  assign imm_i_type_o[2] = instr_rdata_i[22];
  assign regfile_raddr_b_o[1] = instr_rdata_i[21];
  assign imm_j_type_o[1] = instr_rdata_i[21];
  assign imm_u_type_o[21] = instr_rdata_i[21];
  assign imm_i_type_o[1] = instr_rdata_i[21];
  assign regfile_raddr_b_o[0] = instr_rdata_i[20];
  assign imm_j_type_o[11] = instr_rdata_i[20];
  assign imm_u_type_o[20] = instr_rdata_i[20];
  assign imm_i_type_o[0] = instr_rdata_i[20];
  assign regfile_waddr_o[4] = instr_rdata_i[11];
  assign imm_b_type_o[4] = instr_rdata_i[11];
  assign imm_s_type_o[4] = instr_rdata_i[11];
  assign regfile_waddr_o[3] = instr_rdata_i[10];
  assign imm_b_type_o[3] = instr_rdata_i[10];
  assign imm_s_type_o[3] = instr_rdata_i[10];
  assign regfile_waddr_o[2] = instr_rdata_i[9];
  assign imm_b_type_o[2] = instr_rdata_i[9];
  assign imm_s_type_o[2] = instr_rdata_i[9];
  assign regfile_waddr_o[1] = instr_rdata_i[8];
  assign imm_b_type_o[1] = instr_rdata_i[8];
  assign imm_s_type_o[1] = instr_rdata_i[8];
  assign regfile_waddr_o[0] = instr_rdata_i[7];
  assign imm_b_type_o[11] = instr_rdata_i[7];
  assign imm_s_type_o[0] = instr_rdata_i[7];
  assign regfile_raddr_a_o[4] = instr_rdata_i[19];
  assign zimm_rs1_type_o[4] = instr_rdata_i[19];
  assign imm_j_type_o[19] = instr_rdata_i[19];
  assign imm_u_type_o[19] = instr_rdata_i[19];
  assign regfile_raddr_a_o[3] = instr_rdata_i[18];
  assign zimm_rs1_type_o[3] = instr_rdata_i[18];
  assign imm_j_type_o[18] = instr_rdata_i[18];
  assign imm_u_type_o[18] = instr_rdata_i[18];
  assign regfile_raddr_a_o[2] = instr_rdata_i[17];
  assign zimm_rs1_type_o[2] = instr_rdata_i[17];
  assign imm_j_type_o[17] = instr_rdata_i[17];
  assign imm_u_type_o[17] = instr_rdata_i[17];
  assign regfile_raddr_a_o[1] = instr_rdata_i[16];
  assign zimm_rs1_type_o[1] = instr_rdata_i[16];
  assign imm_j_type_o[16] = instr_rdata_i[16];
  assign imm_u_type_o[16] = instr_rdata_i[16];
  assign regfile_raddr_a_o[0] = instr_rdata_i[15];
  assign zimm_rs1_type_o[0] = instr_rdata_i[15];
  assign imm_j_type_o[15] = instr_rdata_i[15];
  assign imm_u_type_o[15] = instr_rdata_i[15];
  assign imm_j_type_o[14] = instr_rdata_i[14];
  assign imm_u_type_o[14] = instr_rdata_i[14];
  assign imm_j_type_o[13] = instr_rdata_i[13];
  assign imm_u_type_o[13] = instr_rdata_i[13];
  assign imm_j_type_o[12] = instr_rdata_i[12];
  assign imm_u_type_o[12] = instr_rdata_i[12];
  assign N83 = instr_rdata_i[1] & instr_rdata_i[0];
  assign N85 = N100 | N101;
  assign N86 = instr_rdata_i[4] | N103;
  assign N87 = N85 | N86;
  assign N88 = N87 | N104;
  assign N90 = instr_rdata_i[4] | instr_rdata_i[3];
  assign N91 = N85 | N90;
  assign N92 = N91 | N104;
  assign N94 = N91 | instr_rdata_i[2];
  assign N96 = instr_rdata_i[6] | N101;
  assign N97 = N96 | N90;
  assign N98 = N97 | instr_rdata_i[2];
  assign N105 = N100 & N101;
  assign N106 = N102 & N103;
  assign N107 = N105 & N106;
  assign N108 = N107 & N104;
  assign N109 = N102 | instr_rdata_i[3];
  assign N110 = N96 | N109;
  assign N111 = N110 | N104;
  assign N113 = instr_rdata_i[6] | instr_rdata_i[5];
  assign N114 = N113 | N109;
  assign N115 = N114 | N104;
  assign N117 = N114 | instr_rdata_i[2];
  assign N119 = N110 | instr_rdata_i[2];
  assign N121 = N113 | N86;
  assign N122 = N121 | N104;
  assign N124 = N85 | N109;
  assign N125 = N124 | instr_rdata_i[2];
  assign N127 = instr_rdata_i[4] & instr_rdata_i[3];
  assign N128 = N100 & instr_rdata_i[5];
  assign N129 = N128 & instr_rdata_i[3];
  assign N130 = instr_rdata_i[6] & N101;
  assign N131 = N130 & instr_rdata_i[3];
  assign N132 = instr_rdata_i[6] & instr_rdata_i[4];
  assign N133 = N132 & instr_rdata_i[2];
  assign N134 = N100 & N102;
  assign N135 = N103 & instr_rdata_i[2];
  assign N136 = N134 & N135;
  assign N137 = N101 & N102;
  assign N138 = N137 & N135;
  assign N139 = instr_rdata_i[3] & N104;
  assign N140 = N130 & N104;
  assign N143 = N142 & N603;
  assign N144 = N143 & N604;
  assign N145 = instr_rdata_i[14] | instr_rdata_i[13];
  assign N146 = N145 | N604;
  assign N148 = N142 | instr_rdata_i[13];
  assign N149 = N148 | instr_rdata_i[12];
  assign N151 = N142 | instr_rdata_i[13];
  assign N152 = N151 | N604;
  assign N154 = N142 | N603;
  assign N155 = N154 | instr_rdata_i[12];
  assign N157 = instr_rdata_i[14] & instr_rdata_i[13];
  assign N158 = N157 & instr_rdata_i[12];
  assign N159 = instr_rdata_i[14] | N603;
  assign N173 = N603 & N604;
  assign N174 = instr_rdata_i[13] | N604;
  assign N176 = N603 | instr_rdata_i[12];
  assign N178 = instr_rdata_i[13] & instr_rdata_i[12];
  assign N180 = N603 & N604;
  assign N181 = instr_rdata_i[13] | N604;
  assign N186 = N184 & N548;
  assign N187 = N185 & N549;
  assign N188 = N186 & N187;
  assign N190 = N547 & N533;
  assign N191 = N190 & N534;
  assign N192 = N547 | instr_rdata_i[29];
  assign N193 = N192 | instr_rdata_i[28];
  assign N195 = instr_rdata_i[30] | instr_rdata_i[29];
  assign N196 = N195 | N534;
  assign N197 = N547 | instr_rdata_i[29];
  assign N198 = N197 | N534;
  assign N200 = instr_rdata_i[30] | N533;
  assign N201 = N200 | instr_rdata_i[28];
  assign N203 = instr_rdata_i[29] & instr_rdata_i[28];
  assign N204 = instr_rdata_i[30] & instr_rdata_i[29];
  assign N221 = N218 & N219;
  assign N222 = N221 & N220;
  assign N223 = instr_rdata_i[14] | N219;
  assign N224 = N223 | instr_rdata_i[12];
  assign N226 = instr_rdata_i[14] | N219;
  assign N227 = N226 | N220;
  assign N229 = N218 | instr_rdata_i[13];
  assign N230 = N229 | instr_rdata_i[12];
  assign N232 = N218 | N219;
  assign N233 = N232 | instr_rdata_i[12];
  assign N235 = instr_rdata_i[14] & instr_rdata_i[13];
  assign N236 = N235 & instr_rdata_i[12];
  assign N237 = instr_rdata_i[14] | instr_rdata_i[13];
  assign N238 = N237 | N220;
  assign N240 = N218 | instr_rdata_i[13];
  assign N241 = N240 | N220;
  assign N255 = N533 & N534;
  assign N256 = N548 & N185;
  assign N257 = N255 & N256;
  assign N259 = N547 & N549;
  assign N260 = N142 & N603;
  assign N261 = N259 & N260;
  assign N262 = N261 & N604;
  assign N263 = N547 | instr_rdata_i[25];
  assign N264 = instr_rdata_i[14] | instr_rdata_i[13];
  assign N265 = N263 | N264;
  assign N266 = N265 | instr_rdata_i[12];
  assign N268 = instr_rdata_i[30] | instr_rdata_i[25];
  assign N269 = instr_rdata_i[14] | N603;
  assign N270 = N268 | N269;
  assign N271 = N270 | instr_rdata_i[12];
  assign N273 = instr_rdata_i[30] | instr_rdata_i[25];
  assign N274 = instr_rdata_i[14] | N603;
  assign N275 = N273 | N274;
  assign N276 = N275 | N604;
  assign N278 = instr_rdata_i[30] | instr_rdata_i[25];
  assign N279 = N142 | instr_rdata_i[13];
  assign N280 = N278 | N279;
  assign N281 = N280 | instr_rdata_i[12];
  assign N283 = instr_rdata_i[30] | instr_rdata_i[25];
  assign N284 = N142 | N603;
  assign N285 = N283 | N284;
  assign N286 = N285 | instr_rdata_i[12];
  assign N288 = instr_rdata_i[30] | instr_rdata_i[25];
  assign N289 = N142 | N603;
  assign N290 = N288 | N289;
  assign N291 = N290 | N604;
  assign N293 = instr_rdata_i[30] | instr_rdata_i[25];
  assign N294 = instr_rdata_i[14] | instr_rdata_i[13];
  assign N295 = N293 | N294;
  assign N296 = N295 | N604;
  assign N298 = instr_rdata_i[30] | instr_rdata_i[25];
  assign N299 = N142 | instr_rdata_i[13];
  assign N300 = N298 | N299;
  assign N301 = N300 | N604;
  assign N303 = N547 | instr_rdata_i[25];
  assign N304 = N142 | instr_rdata_i[13];
  assign N305 = N303 | N304;
  assign N306 = N305 | N604;
  assign N308 = instr_rdata_i[30] | N549;
  assign N309 = instr_rdata_i[14] | instr_rdata_i[13];
  assign N310 = N308 | N309;
  assign N311 = N310 | instr_rdata_i[12];
  assign N313 = instr_rdata_i[30] | N549;
  assign N314 = instr_rdata_i[14] | instr_rdata_i[13];
  assign N315 = N313 | N314;
  assign N316 = N315 | N604;
  assign N318 = instr_rdata_i[30] | N549;
  assign N319 = instr_rdata_i[14] | N603;
  assign N320 = N318 | N319;
  assign N321 = N320 | instr_rdata_i[12];
  assign N323 = instr_rdata_i[30] | N549;
  assign N324 = instr_rdata_i[14] | N603;
  assign N325 = N323 | N324;
  assign N326 = N325 | N604;
  assign N328 = instr_rdata_i[30] | N549;
  assign N329 = N142 | instr_rdata_i[13];
  assign N330 = N328 | N329;
  assign N331 = N330 | instr_rdata_i[12];
  assign N333 = instr_rdata_i[30] | N549;
  assign N334 = N142 | instr_rdata_i[13];
  assign N335 = N333 | N334;
  assign N336 = N335 | N604;
  assign N338 = instr_rdata_i[30] | N549;
  assign N339 = N142 | N603;
  assign N340 = N338 | N339;
  assign N341 = N340 | instr_rdata_i[12];
  assign N343 = instr_rdata_i[30] | N549;
  assign N344 = N142 | N603;
  assign N345 = N343 | N344;
  assign N346 = N345 | N604;
  assign N348 = instr_rdata_i[30] & N142;
  assign N349 = N348 & instr_rdata_i[12];
  assign N350 = instr_rdata_i[30] & instr_rdata_i[13];
  assign N351 = instr_rdata_i[30] & instr_rdata_i[14];
  assign N352 = N351 & N604;
  assign N353 = instr_rdata_i[30] & instr_rdata_i[25];
  assign N385 = N184 & N185;
  assign N386 = N385 & N384;
  assign N389 = N547 & N533;
  assign N390 = N534 & N548;
  assign N391 = N549 & N550;
  assign N392 = N388 & N576;
  assign N393 = N389 & N390;
  assign N394 = N391 & N392;
  assign N395 = N393 & N394;
  assign N396 = N395 & N563;
  assign N397 = instr_rdata_i[30] | instr_rdata_i[29];
  assign N398 = instr_rdata_i[28] | instr_rdata_i[27];
  assign N399 = instr_rdata_i[25] | instr_rdata_i[24];
  assign N400 = instr_rdata_i[22] | instr_rdata_i[21];
  assign N401 = N397 | N398;
  assign N402 = N399 | N400;
  assign N403 = N401 | N402;
  assign N404 = N403 | N563;
  assign N406 = instr_rdata_i[30] | N533;
  assign N407 = N534 | instr_rdata_i[27];
  assign N408 = instr_rdata_i[25] | instr_rdata_i[24];
  assign N409 = instr_rdata_i[22] | N576;
  assign N410 = N406 | N407;
  assign N411 = N408 | N409;
  assign N412 = N410 | N411;
  assign N413 = N412 | instr_rdata_i[20];
  assign N415 = N547 | N533;
  assign N416 = N534 | N548;
  assign N417 = N549 | N550;
  assign N418 = instr_rdata_i[22] | N576;
  assign N419 = N415 | N416;
  assign N420 = N417 | N418;
  assign N421 = N419 | N420;
  assign N422 = N421 | instr_rdata_i[20];
  assign N424 = instr_rdata_i[30] | instr_rdata_i[29];
  assign N425 = N534 | instr_rdata_i[27];
  assign N426 = instr_rdata_i[25] | instr_rdata_i[24];
  assign N427 = N388 | instr_rdata_i[21];
  assign N428 = N424 | N425;
  assign N429 = N426 | N427;
  assign N430 = N428 | N429;
  assign N431 = N430 | N563;
  assign N453 = instr_rdata_i[13] | N604;
  assign N455 = N603 | instr_rdata_i[12];
  assign N457 = instr_rdata_i[13] & instr_rdata_i[12];
  assign N458 = N603 & N604;
  assign N524 = ~csr_op[1];
  assign N525 = csr_op[0] | N524;
  assign N526 = ~N525;
  assign N527 = csr_op[0] & csr_op[1];
  assign N528 = instr_rdata_i[18] | instr_rdata_i[19];
  assign N529 = instr_rdata_i[17] | N528;
  assign N530 = instr_rdata_i[16] | N529;
  assign N531 = instr_rdata_i[15] | N530;
  assign N532 = ~N531;
  assign N533 = ~instr_rdata_i[29];
  assign N534 = ~instr_rdata_i[28];
  assign N535 = instr_rdata_i[30] | instr_rdata_i[31];
  assign N536 = N533 | N535;
  assign N537 = N534 | N536;
  assign N538 = instr_rdata_i[27] | N537;
  assign N539 = instr_rdata_i[26] | N538;
  assign N540 = instr_rdata_i[25] | N539;
  assign N541 = instr_rdata_i[24] | N540;
  assign N542 = instr_rdata_i[23] | N541;
  assign N543 = instr_rdata_i[22] | N542;
  assign N544 = instr_rdata_i[21] | N543;
  assign N545 = instr_rdata_i[20] | N544;
  assign N546 = ~N545;
  assign N547 = ~instr_rdata_i[30];
  assign N548 = ~instr_rdata_i[27];
  assign N549 = ~instr_rdata_i[25];
  assign N550 = ~instr_rdata_i[24];
  assign N551 = N547 | instr_rdata_i[31];
  assign N552 = N533 | N551;
  assign N553 = N534 | N552;
  assign N554 = N548 | N553;
  assign N555 = instr_rdata_i[26] | N554;
  assign N556 = N549 | N555;
  assign N557 = N550 | N556;
  assign N558 = instr_rdata_i[23] | N557;
  assign N559 = instr_rdata_i[22] | N558;
  assign N560 = instr_rdata_i[21] | N559;
  assign N561 = instr_rdata_i[20] | N560;
  assign N562 = ~N561;
  assign N563 = ~instr_rdata_i[20];
  assign N564 = N547 | instr_rdata_i[31];
  assign N565 = N533 | N564;
  assign N566 = N534 | N565;
  assign N567 = N548 | N566;
  assign N568 = instr_rdata_i[26] | N567;
  assign N569 = N549 | N568;
  assign N570 = N550 | N569;
  assign N571 = instr_rdata_i[23] | N570;
  assign N572 = instr_rdata_i[22] | N571;
  assign N573 = instr_rdata_i[21] | N572;
  assign N574 = N563 | N573;
  assign N575 = ~N574;
  assign N576 = ~instr_rdata_i[21];
  assign N577 = N547 | instr_rdata_i[31];
  assign N578 = N533 | N577;
  assign N579 = N534 | N578;
  assign N580 = N548 | N579;
  assign N581 = instr_rdata_i[26] | N580;
  assign N582 = N549 | N581;
  assign N583 = N550 | N582;
  assign N584 = instr_rdata_i[23] | N583;
  assign N585 = instr_rdata_i[22] | N584;
  assign N586 = N576 | N585;
  assign N587 = instr_rdata_i[20] | N586;
  assign N588 = ~N587;
  assign N589 = N547 | instr_rdata_i[31];
  assign N590 = N533 | N589;
  assign N591 = N534 | N590;
  assign N592 = N548 | N591;
  assign N593 = instr_rdata_i[26] | N592;
  assign N594 = N549 | N593;
  assign N595 = N550 | N594;
  assign N596 = instr_rdata_i[23] | N595;
  assign N597 = instr_rdata_i[22] | N596;
  assign N598 = N576 | N597;
  assign N599 = N563 | N598;
  assign N600 = ~N599;
  assign N601 = instr_rdata_i[13] | instr_rdata_i[14];
  assign N602 = instr_rdata_i[12] | N601;
  assign N603 = ~instr_rdata_i[13];
  assign N604 = ~instr_rdata_i[12];
  assign N605 = N603 | instr_rdata_i[14];
  assign N606 = N604 | N605;
  assign N607 = ~N606;
  assign N608 = instr_rdata_i[13] | instr_rdata_i[14];
  assign N609 = instr_rdata_i[12] | N608;
  assign N610 = instr_rdata_i[13] & instr_rdata_i[14];
  assign N611 = instr_rdata_i[12] & N610;
  assign N612 = instr_rdata_i[30] | instr_rdata_i[31];
  assign N613 = instr_rdata_i[29] | N612;
  assign N614 = instr_rdata_i[28] | N613;
  assign N615 = instr_rdata_i[27] | N614;
  assign N616 = instr_rdata_i[26] | N615;
  assign N617 = instr_rdata_i[25] | N616;
  assign N618 = N547 | instr_rdata_i[31];
  assign N619 = instr_rdata_i[29] | N618;
  assign N620 = instr_rdata_i[28] | N619;
  assign N621 = instr_rdata_i[27] | N620;
  assign N622 = instr_rdata_i[26] | N621;
  assign N623 = instr_rdata_i[25] | N622;
  assign N624 = ~N623;
  assign N625 = instr_rdata_i[30] | instr_rdata_i[31];
  assign N626 = instr_rdata_i[29] | N625;
  assign N627 = instr_rdata_i[28] | N626;
  assign N628 = instr_rdata_i[27] | N627;
  assign N629 = instr_rdata_i[26] | N628;
  assign N630 = instr_rdata_i[25] | N629;
  assign N631 = ~N630;
  assign N632 = instr_rdata_i[13] | instr_rdata_i[14];
  assign N633 = instr_rdata_i[12] | N632;
  assign N634 = ~N633;
  assign csr_op_o = (N0)? { 1'b0, 1'b0 } : 
                    (N82)? csr_op : 1'b0;
  assign N0 = N81;
  assign { N165, N164, N163, N162, N161 } = (N1)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                            (N2)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                            (N3)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                            (N4)? { 1'b0, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                                            (N5)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b1 } : 
                                            (N6)? { 1'b0, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                            (N7)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 1'b0;
  assign N1 = N144;
  assign N2 = N147;
  assign N3 = N150;
  assign N4 = N153;
  assign N5 = N156;
  assign N6 = N158;
  assign N7 = N160;
  assign N166 = (N1)? 1'b0 : 
                (N2)? 1'b0 : 
                (N3)? 1'b0 : 
                (N4)? 1'b0 : 
                (N5)? 1'b0 : 
                (N6)? 1'b0 : 
                (N7)? 1'b1 : 1'b0;
  assign { N172, N171, N170, N169, N168 } = (N8)? { N165, N164, N163, N162, N161 } : 
                                            (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = instr_new_i;
  assign N9 = N167;
  assign N179 = (N10)? instr_rdata_i[14] : 
                (N11)? instr_rdata_i[14] : 
                (N12)? instr_rdata_i[14] : 
                (N13)? 1'b1 : 1'b0;
  assign N10 = N173;
  assign N11 = N175;
  assign N12 = N177;
  assign N13 = N178;
  assign { N207, N206 } = (N14)? { 1'b1, 1'b0 } : 
                          (N15)? { 1'b0, 1'b1 } : 
                          (N16)? { 1'b0, 1'b0 } : 
                          (N17)? { N180, N182 } : 1'b0;
  assign N14 = N194;
  assign N15 = N199;
  assign N16 = N202;
  assign N17 = N205;
  assign N208 = (N14)? 1'b0 : 
                (N15)? 1'b0 : 
                (N16)? 1'b0 : 
                (N17)? 1'b1 : 1'b0;
  assign { N210, N209 } = (N18)? { N207, N206 } : 
                          (N189)? { N180, N182 } : 1'b0;
  assign N18 = N188;
  assign N211 = (N18)? N208 : 
                (N189)? 1'b1 : 1'b0;
  assign N212 = ~N611;
  assign N213 = (N19)? N547 : 
                (N183)? N142 : 1'b0;
  assign N19 = N611;
  assign N214 = (N19)? N211 : 
                (N183)? 1'b0 : 1'b0;
  assign { N216, N215 } = (N19)? { N210, N209 } : 
                          (N183)? { N180, N182 } : 1'b0;
  assign N217 = (N20)? 1'b1 : 
                (N21)? N214 : 1'b0;
  assign N20 = N607;
  assign N21 = N606;
  assign N245 = (N22)? 1'b0 : 
                (N23)? 1'b1 : 
                (N24)? 1'b1 : 1'b0;
  assign N22 = N631;
  assign N23 = N630;
  assign N24 = 1'b0;
  assign { N248, N247, N246 } = (N22)? { 1'b0, 1'b1, 1'b1 } : 
                                (N25)? { 1'b0, 1'b1, 1'b0 } : 
                                (N244)? { 1'b1, 1'b0, 1'b1 } : 1'b0;
  assign N25 = N624;
  assign { N252, N251, N250, N249 } = (N26)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N225)? { 1'b1, 1'b0, 1'b1, 1'b0 } : 
                                      (N228)? { 1'b1, 1'b0, 1'b1, 1'b1 } : 
                                      (N231)? { 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                      (N234)? { 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                      (N27)? { 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                      (N239)? { 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                      (N242)? { N248, N247, N246, N245 } : 1'b0;
  assign N26 = N222;
  assign N27 = N236;
  assign N253 = (N26)? 1'b0 : 
                (N225)? 1'b0 : 
                (N228)? 1'b0 : 
                (N231)? 1'b0 : 
                (N234)? 1'b0 : 
                (N27)? 1'b0 : 
                (N239)? N617 : 
                (N242)? N248 : 1'b0;
  assign { N358, N357, N356, N355 } = (N28)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N29)? { 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                      (N30)? { 1'b1, 1'b0, 1'b1, 1'b0 } : 
                                      (N31)? { 1'b1, 1'b0, 1'b1, 1'b1 } : 
                                      (N32)? { 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                      (N33)? { 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                      (N34)? { 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                      (N35)? { 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                      (N36)? { 1'b0, 1'b1, 1'b1, 1'b0 } : 
                                      (N37)? { 1'b0, 1'b1, 1'b0, 1'b1 } : 
                                      (N38)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N39)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N40)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N41)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N42)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N43)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N44)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N45)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N46)? { 1'b1, 1'b0, 1'b1, 1'b1 } : 1'b0;
  assign N28 = N262;
  assign N29 = N267;
  assign N30 = N272;
  assign N31 = N277;
  assign N32 = N282;
  assign N33 = N287;
  assign N34 = N292;
  assign N35 = N297;
  assign N36 = N302;
  assign N37 = N307;
  assign N38 = N312;
  assign N39 = N317;
  assign N40 = N322;
  assign N41 = N327;
  assign N42 = N332;
  assign N43 = N337;
  assign N44 = N342;
  assign N45 = N347;
  assign N46 = N354;
  assign { N360, N359 } = (N28)? { 1'b0, 1'b0 } : 
                          (N29)? { 1'b0, 1'b0 } : 
                          (N30)? { 1'b0, 1'b0 } : 
                          (N31)? { 1'b0, 1'b0 } : 
                          (N32)? { 1'b0, 1'b0 } : 
                          (N33)? { 1'b0, 1'b0 } : 
                          (N34)? { 1'b0, 1'b0 } : 
                          (N35)? { 1'b0, 1'b0 } : 
                          (N36)? { 1'b0, 1'b0 } : 
                          (N37)? { 1'b0, 1'b0 } : 
                          (N38)? { 1'b0, 1'b0 } : 
                          (N39)? { 1'b0, 1'b1 } : 
                          (N40)? { 1'b0, 1'b1 } : 
                          (N41)? { 1'b0, 1'b1 } : 
                          (N42)? { 1'b1, 1'b0 } : 
                          (N43)? { 1'b1, 1'b0 } : 
                          (N44)? { 1'b1, 1'b1 } : 
                          (N45)? { 1'b1, 1'b1 } : 
                          (N46)? { 1'b0, 1'b0 } : 1'b0;
  assign N361 = (N28)? 1'b0 : 
                (N29)? 1'b0 : 
                (N30)? 1'b0 : 
                (N31)? 1'b0 : 
                (N32)? 1'b0 : 
                (N33)? 1'b0 : 
                (N34)? 1'b0 : 
                (N35)? 1'b0 : 
                (N36)? 1'b0 : 
                (N37)? 1'b0 : 
                (N38)? 1'b1 : 
                (N39)? 1'b1 : 
                (N40)? 1'b1 : 
                (N41)? 1'b1 : 
                (N42)? 1'b0 : 
                (N43)? 1'b0 : 
                (N44)? 1'b0 : 
                (N45)? 1'b0 : 
                (N46)? 1'b0 : 1'b0;
  assign { N363, N362 } = (N28)? { 1'b0, 1'b0 } : 
                          (N29)? { 1'b0, 1'b0 } : 
                          (N30)? { 1'b0, 1'b0 } : 
                          (N31)? { 1'b0, 1'b0 } : 
                          (N32)? { 1'b0, 1'b0 } : 
                          (N33)? { 1'b0, 1'b0 } : 
                          (N34)? { 1'b0, 1'b0 } : 
                          (N35)? { 1'b0, 1'b0 } : 
                          (N36)? { 1'b0, 1'b0 } : 
                          (N37)? { 1'b0, 1'b0 } : 
                          (N38)? { 1'b0, 1'b0 } : 
                          (N39)? { 1'b1, 1'b1 } : 
                          (N40)? { 1'b0, 1'b1 } : 
                          (N41)? { 1'b0, 1'b0 } : 
                          (N42)? { 1'b1, 1'b1 } : 
                          (N43)? { 1'b0, 1'b0 } : 
                          (N44)? { 1'b1, 1'b1 } : 
                          (N45)? { 1'b0, 1'b0 } : 
                          (N46)? { 1'b0, 1'b0 } : 1'b0;
  assign N364 = (N47)? N354 : 
                (N258)? 1'b1 : 1'b0;
  assign N47 = N257;
  assign { N368, N367, N366, N365 } = (N47)? { N358, N357, N356, N355 } : 
                                      (N258)? { 1'b1, 1'b0, 1'b1, 1'b1 } : 1'b0;
  assign { N370, N369 } = (N47)? { N360, N359 } : 
                          (N258)? { 1'b0, 1'b0 } : 1'b0;
  assign N371 = (N47)? N361 : 
                (N258)? 1'b0 : 1'b0;
  assign { N373, N372 } = (N47)? { N363, N362 } : 
                          (N258)? { 1'b0, 1'b0 } : 1'b0;
  assign N374 = (N48)? 1'b1 : 
                (N254)? N364 : 1'b0;
  assign N48 = instr_rdata_i[31];
  assign { N376, N375 } = (N48)? { 1'b0, 1'b0 } : 
                          (N254)? { N373, N372 } : 1'b0;
  assign { N380, N379, N378, N377 } = (N48)? { 1'b1, 1'b0, 1'b1, 1'b1 } : 
                                      (N254)? { N368, N367, N366, N365 } : 1'b0;
  assign { N382, N381 } = (N48)? { 1'b0, 1'b0 } : 
                          (N254)? { N370, N369 } : 1'b0;
  assign N383 = (N48)? 1'b0 : 
                (N254)? N371 : 1'b0;
  assign N438 = (N49)? 1'b1 : 
                (N50)? 1'b0 : 
                (N51)? 1'b0 : 
                (N52)? 1'b0 : 
                (N53)? 1'b0 : 
                (N437)? 1'b0 : 1'b0;
  assign N49 = N396;
  assign N50 = N405;
  assign N51 = N414;
  assign N52 = N423;
  assign N53 = N432;
  assign N439 = (N49)? 1'b0 : 
                (N50)? 1'b1 : 
                (N51)? 1'b0 : 
                (N52)? 1'b0 : 
                (N53)? 1'b0 : 
                (N437)? 1'b0 : 1'b0;
  assign N440 = (N49)? 1'b0 : 
                (N50)? 1'b0 : 
                (N51)? 1'b1 : 
                (N52)? 1'b0 : 
                (N53)? 1'b0 : 
                (N437)? 1'b0 : 1'b0;
  assign N441 = (N49)? 1'b0 : 
                (N50)? 1'b0 : 
                (N51)? 1'b0 : 
                (N52)? 1'b1 : 
                (N53)? 1'b0 : 
                (N437)? 1'b0 : 1'b0;
  assign N442 = (N49)? 1'b0 : 
                (N50)? 1'b0 : 
                (N51)? 1'b0 : 
                (N52)? 1'b0 : 
                (N53)? 1'b1 : 
                (N437)? 1'b0 : 1'b0;
  assign N443 = (N49)? 1'b0 : 
                (N50)? 1'b0 : 
                (N51)? 1'b0 : 
                (N52)? 1'b0 : 
                (N53)? 1'b0 : 
                (N437)? 1'b1 : 1'b0;
  assign N444 = (N54)? N442 : 
                (N387)? 1'b0 : 1'b0;
  assign N54 = N386;
  assign N445 = (N54)? N443 : 
                (N387)? 1'b1 : 1'b0;
  assign N446 = (N54)? N438 : 
                (N387)? 1'b0 : 1'b0;
  assign N447 = (N54)? N439 : 
                (N387)? 1'b0 : 1'b0;
  assign N448 = (N54)? N440 : 
                (N387)? 1'b0 : 1'b0;
  assign N449 = (N54)? N441 : 
                (N387)? 1'b0 : 1'b0;
  assign N452 = (N55)? 1'b1 : 
                (N451)? N445 : 1'b0;
  assign N55 = N450;
  assign { N460, N459 } = (N56)? { 1'b0, 1'b1 } : 
                          (N57)? { 1'b1, 1'b0 } : 
                          (N58)? { 1'b1, 1'b1 } : 
                          (N59)? { 1'b0, 1'b0 } : 1'b0;
  assign N56 = N454;
  assign N57 = N456;
  assign N58 = N457;
  assign N59 = N458;
  assign N461 = (N56)? 1'b0 : 
                (N57)? 1'b0 : 
                (N58)? 1'b0 : 
                (N59)? 1'b1 : 1'b0;
  assign N464 = (N60)? N463 : 
                (N61)? 1'b0 : 1'b0;
  assign N60 = N462;
  assign N61 = N461;
  assign N465 = (N62)? 1'b0 : 
                (N63)? instr_rdata_i[14] : 1'b0;
  assign N62 = N634;
  assign N63 = N633;
  assign N466 = (N62)? N449 : 
                (N63)? 1'b0 : 1'b0;
  assign N467 = (N62)? N444 : 
                (N63)? 1'b0 : 1'b0;
  assign N468 = (N62)? N452 : 
                (N63)? N461 : 1'b0;
  assign N469 = (N62)? N446 : 
                (N63)? 1'b0 : 1'b0;
  assign N470 = (N62)? N447 : 
                (N63)? 1'b0 : 1'b0;
  assign N471 = (N62)? N448 : 
                (N63)? 1'b0 : 1'b0;
  assign { N473, N472 } = (N62)? { 1'b0, 1'b0 } : 
                          (N63)? { N460, N459 } : 1'b0;
  assign N474 = (N62)? 1'b0 : 
                (N63)? N464 : 1'b0;
  assign N475 = (N64)? 1'b1 : 
                (N65)? 1'b1 : 
                (N66)? 1'b0 : 
                (N67)? 1'b0 : 
                (N68)? 1'b0 : 
                (N69)? 1'b0 : 
                (N70)? 1'b0 : 
                (N71)? 1'b0 : 
                (N72)? 1'b0 : 
                (N73)? 1'b0 : 
                (N74)? 1'b0 : 
                (N75)? 1'b0 : 1'b0;
  assign N64 = N89;
  assign N65 = N93;
  assign N66 = N95;
  assign N67 = N99;
  assign N68 = N108;
  assign N69 = N112;
  assign N70 = N116;
  assign N71 = N118;
  assign N72 = N120;
  assign N73 = N123;
  assign N74 = N126;
  assign N75 = N141;
  assign N476 = (N64)? instr_new_i : 
                (N65)? instr_new_i : 
                (N66)? 1'b0 : 
                (N67)? 1'b0 : 
                (N68)? 1'b0 : 
                (N69)? 1'b0 : 
                (N70)? 1'b0 : 
                (N71)? 1'b0 : 
                (N72)? 1'b0 : 
                (N73)? 1'b0 : 
                (N74)? 1'b0 : 
                (N75)? 1'b0 : 1'b0;
  assign { N478, N477 } = (N64)? { 1'b1, 1'b0 } : 
                          (N65)? { N167, 1'b0 } : 
                          (N66)? { N167, 1'b0 } : 
                          (N67)? { 1'b0, 1'b0 } : 
                          (N68)? { 1'b0, 1'b0 } : 
                          (N69)? { 1'b1, 1'b1 } : 
                          (N70)? { 1'b1, 1'b0 } : 
                          (N71)? { 1'b0, 1'b0 } : 
                          (N72)? { 1'b0, 1'b0 } : 
                          (N73)? { N609, N609 } : 
                          (N74)? { N465, N465 } : 
                          (N75)? { 1'b1, 1'b1 } : 1'b0;
  assign N479 = (N64)? 1'b1 : 
                (N65)? 1'b1 : 
                (N66)? N167 : 
                (N67)? N142 : 
                (N68)? N212 : 
                (N69)? 1'b1 : 
                (N70)? 1'b1 : 
                (N71)? 1'b1 : 
                (N72)? 1'b0 : 
                (N73)? 1'b1 : 
                (N74)? 1'b1 : 
                (N75)? 1'b1 : 1'b0;
  assign { N482, N481, N480 } = (N64)? { 1'b1, 1'b0, N167 } : 
                                (N65)? { N167, 1'b0, N167 } : 
                                (N66)? { 1'b0, N167, 1'b0 } : 
                                (N67)? { 1'b0, 1'b0, N142 } : 
                                (N68)? { 1'b0, 1'b0, 1'b0 } : 
                                (N69)? { 1'b0, 1'b1, 1'b1 } : 
                                (N70)? { 1'b0, 1'b1, 1'b1 } : 
                                (N71)? { 1'b0, 1'b0, 1'b0 } : 
                                (N72)? { 1'b0, 1'b0, 1'b0 } : 
                                (N73)? { 1'b0, 1'b0, 1'b0 } : 
                                (N74)? { 1'b0, 1'b0, 1'b0 } : 
                                (N75)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N488, N485, N484, N483 } = (N64)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N65)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N66)? { N172, N170, N169, N168 } : 
                                      (N67)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N68)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N69)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N70)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N71)? { N252, N251, N250, N249 } : 
                                      (N72)? { N380, N379, N378, N377 } : 
                                      (N73)? { N609, 1'b0, N609, N609 } : 
                                      (N74)? { 1'b1, 1'b0, 1'b1, 1'b1 } : 
                                      (N75)? { 1'b1, 1'b0, 1'b1, 1'b1 } : 1'b0;
  assign N487 = (N66)? N171 : 
                (N486)? 1'b0 : 1'b0;
  assign N489 = (N64)? N167 : 
                (N65)? N167 : 
                (N66)? 1'b0 : 
                (N67)? 1'b0 : 
                (N68)? 1'b1 : 
                (N69)? 1'b1 : 
                (N70)? 1'b1 : 
                (N71)? 1'b1 : 
                (N72)? 1'b1 : 
                (N73)? 1'b0 : 
                (N74)? N633 : 
                (N75)? 1'b0 : 1'b0;
  assign N490 = (N64)? 1'b0 : 
                (N65)? N602 : 
                (N66)? N166 : 
                (N67)? N179 : 
                (N68)? N217 : 
                (N69)? 1'b0 : 
                (N70)? 1'b0 : 
                (N71)? N253 : 
                (N72)? N374 : 
                (N73)? N609 : 
                (N74)? N468 : 
                (N75)? 1'b1 : 1'b0;
  assign N491 = (N64)? 1'b0 : 
                (N65)? 1'b0 : 
                (N66)? 1'b1 : 
                (N67)? 1'b0 : 
                (N68)? 1'b0 : 
                (N69)? 1'b0 : 
                (N70)? 1'b0 : 
                (N71)? 1'b0 : 
                (N72)? 1'b0 : 
                (N73)? 1'b0 : 
                (N74)? 1'b0 : 
                (N75)? 1'b0 : 1'b0;
  assign N492 = (N64)? 1'b0 : 
                (N65)? 1'b0 : 
                (N66)? 1'b0 : 
                (N67)? 1'b1 : 
                (N68)? 1'b1 : 
                (N69)? 1'b0 : 
                (N70)? 1'b0 : 
                (N71)? 1'b0 : 
                (N72)? 1'b0 : 
                (N73)? 1'b0 : 
                (N74)? 1'b0 : 
                (N75)? 1'b0 : 1'b0;
  assign N493 = (N64)? 1'b0 : 
                (N65)? 1'b0 : 
                (N66)? 1'b0 : 
                (N67)? 1'b1 : 
                (N68)? 1'b0 : 
                (N69)? 1'b0 : 
                (N70)? 1'b0 : 
                (N71)? 1'b0 : 
                (N72)? 1'b0 : 
                (N73)? 1'b0 : 
                (N74)? 1'b0 : 
                (N75)? 1'b0 : 1'b0;
  assign { N495, N494 } = (N64)? { 1'b0, 1'b0 } : 
                          (N65)? { 1'b0, 1'b0 } : 
                          (N66)? { 1'b0, 1'b0 } : 
                          (N67)? { N173, N175 } : 
                          (N68)? { N216, N215 } : 
                          (N69)? { 1'b0, 1'b0 } : 
                          (N70)? { 1'b0, 1'b0 } : 
                          (N71)? { 1'b0, 1'b0 } : 
                          (N72)? { 1'b0, 1'b0 } : 
                          (N73)? { 1'b0, 1'b0 } : 
                          (N74)? { 1'b0, 1'b0 } : 
                          (N75)? { 1'b0, 1'b0 } : 1'b0;
  assign { N497, N496 } = (N64)? { 1'b0, 1'b1 } : 
                          (N65)? { 1'b0, 1'b1 } : 
                          (N66)? { 1'b0, 1'b1 } : 
                          (N67)? { 1'b0, 1'b1 } : 
                          (N68)? { 1'b0, 1'b0 } : 
                          (N69)? { 1'b0, 1'b1 } : 
                          (N70)? { 1'b0, 1'b1 } : 
                          (N71)? { 1'b0, 1'b1 } : 
                          (N72)? { 1'b0, 1'b1 } : 
                          (N73)? { 1'b0, 1'b1 } : 
                          (N74)? { N633, N634 } : 
                          (N75)? { 1'b0, 1'b1 } : 1'b0;
  assign N498 = (N64)? 1'b0 : 
                (N65)? 1'b0 : 
                (N66)? 1'b0 : 
                (N67)? 1'b0 : 
                (N68)? N213 : 
                (N69)? 1'b0 : 
                (N70)? 1'b0 : 
                (N71)? 1'b0 : 
                (N72)? 1'b0 : 
                (N73)? 1'b0 : 
                (N74)? 1'b0 : 
                (N75)? 1'b0 : 1'b0;
  assign N499 = (N64)? 1'b1 : 
                (N65)? 1'b1 : 
                (N66)? 1'b1 : 
                (N67)? 1'b1 : 
                (N68)? 1'b1 : 
                (N69)? 1'b1 : 
                (N70)? 1'b1 : 
                (N71)? 1'b1 : 
                (N72)? 1'b1 : 
                (N73)? 1'b1 : 
                (N74)? N634 : 
                (N75)? 1'b1 : 1'b0;
  assign { N501, N500 } = (N64)? { 1'b0, 1'b0 } : 
                          (N65)? { 1'b0, 1'b0 } : 
                          (N66)? { 1'b0, 1'b0 } : 
                          (N67)? { 1'b0, 1'b0 } : 
                          (N68)? { 1'b0, 1'b0 } : 
                          (N69)? { 1'b0, 1'b0 } : 
                          (N70)? { 1'b0, 1'b0 } : 
                          (N71)? { 1'b0, 1'b0 } : 
                          (N72)? { N376, N375 } : 
                          (N73)? { 1'b0, 1'b0 } : 
                          (N74)? { 1'b0, 1'b0 } : 
                          (N75)? { 1'b0, 1'b0 } : 1'b0;
  assign { N503, N502 } = (N64)? { 1'b0, 1'b0 } : 
                          (N65)? { 1'b0, 1'b0 } : 
                          (N66)? { 1'b0, 1'b0 } : 
                          (N67)? { 1'b0, 1'b0 } : 
                          (N68)? { 1'b0, 1'b0 } : 
                          (N69)? { 1'b0, 1'b0 } : 
                          (N70)? { 1'b0, 1'b0 } : 
                          (N71)? { 1'b0, 1'b0 } : 
                          (N72)? { N382, N381 } : 
                          (N73)? { 1'b0, 1'b0 } : 
                          (N74)? { 1'b0, 1'b0 } : 
                          (N75)? { 1'b0, 1'b0 } : 1'b0;
  assign N504 = (N64)? 1'b0 : 
                (N65)? 1'b0 : 
                (N66)? 1'b0 : 
                (N67)? 1'b0 : 
                (N68)? 1'b0 : 
                (N69)? 1'b0 : 
                (N70)? 1'b0 : 
                (N71)? 1'b0 : 
                (N72)? N383 : 
                (N73)? 1'b0 : 
                (N74)? 1'b0 : 
                (N75)? 1'b0 : 1'b0;
  assign N505 = (N64)? 1'b0 : 
                (N65)? 1'b0 : 
                (N66)? 1'b0 : 
                (N67)? 1'b0 : 
                (N68)? 1'b0 : 
                (N69)? 1'b0 : 
                (N70)? 1'b0 : 
                (N71)? 1'b0 : 
                (N72)? 1'b0 : 
                (N73)? 1'b0 : 
                (N74)? N474 : 
                (N75)? 1'b0 : 1'b0;
  assign N506 = (N64)? 1'b0 : 
                (N65)? 1'b0 : 
                (N66)? 1'b0 : 
                (N67)? 1'b0 : 
                (N68)? 1'b0 : 
                (N69)? 1'b0 : 
                (N70)? 1'b0 : 
                (N71)? 1'b0 : 
                (N72)? 1'b0 : 
                (N73)? 1'b0 : 
                (N74)? N466 : 
                (N75)? 1'b0 : 1'b0;
  assign N507 = (N64)? 1'b0 : 
                (N65)? 1'b0 : 
                (N66)? 1'b0 : 
                (N67)? 1'b0 : 
                (N68)? 1'b0 : 
                (N69)? 1'b0 : 
                (N70)? 1'b0 : 
                (N71)? 1'b0 : 
                (N72)? 1'b0 : 
                (N73)? 1'b0 : 
                (N74)? N467 : 
                (N75)? 1'b0 : 1'b0;
  assign N508 = (N64)? 1'b0 : 
                (N65)? 1'b0 : 
                (N66)? 1'b0 : 
                (N67)? 1'b0 : 
                (N68)? 1'b0 : 
                (N69)? 1'b0 : 
                (N70)? 1'b0 : 
                (N71)? 1'b0 : 
                (N72)? 1'b0 : 
                (N73)? 1'b0 : 
                (N74)? N469 : 
                (N75)? 1'b0 : 1'b0;
  assign N509 = (N64)? 1'b0 : 
                (N65)? 1'b0 : 
                (N66)? 1'b0 : 
                (N67)? 1'b0 : 
                (N68)? 1'b0 : 
                (N69)? 1'b0 : 
                (N70)? 1'b0 : 
                (N71)? 1'b0 : 
                (N72)? 1'b0 : 
                (N73)? 1'b0 : 
                (N74)? N470 : 
                (N75)? 1'b0 : 1'b0;
  assign N510 = (N64)? 1'b0 : 
                (N65)? 1'b0 : 
                (N66)? 1'b0 : 
                (N67)? 1'b0 : 
                (N68)? 1'b0 : 
                (N69)? 1'b0 : 
                (N70)? 1'b0 : 
                (N71)? 1'b0 : 
                (N72)? 1'b0 : 
                (N73)? 1'b0 : 
                (N74)? N471 : 
                (N75)? 1'b0 : 1'b0;
  assign { N512, N511 } = (N64)? { 1'b0, 1'b0 } : 
                          (N65)? { 1'b0, 1'b0 } : 
                          (N66)? { 1'b0, 1'b0 } : 
                          (N67)? { 1'b0, 1'b0 } : 
                          (N68)? { 1'b0, 1'b0 } : 
                          (N69)? { 1'b0, 1'b0 } : 
                          (N70)? { 1'b0, 1'b0 } : 
                          (N71)? { 1'b0, 1'b0 } : 
                          (N72)? { 1'b0, 1'b0 } : 
                          (N73)? { 1'b0, 1'b0 } : 
                          (N74)? { N473, N472 } : 
                          (N75)? { 1'b0, 1'b0 } : 1'b0;
  assign N513 = (N76)? N497 : 
                (N84)? 1'b0 : 1'b0;
  assign N76 = N83;
  assign csr_op = (N76)? { N512, N511 } : 
                  (N84)? { 1'b0, 1'b0 } : 1'b0;
  assign N514 = (N76)? N475 : 
                (N84)? 1'b0 : 1'b0;
  assign jump_set_o = (N76)? N476 : 
                      (N84)? 1'b0 : 1'b0;
  assign alu_op_a_mux_sel_o = (N76)? { N478, N477 } : 
                              (N84)? { 1'b1, 1'b1 } : 1'b0;
  assign alu_op_b_mux_sel_o = (N76)? N479 : 
                              (N84)? 1'b1 : 1'b0;
  assign imm_b_mux_sel_o = (N76)? { N482, N481, N480 } : 
                           (N84)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign alu_operator_o = (N76)? { N488, N487, N485, N484, N483 } : 
                          (N84)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 1'b0;
  assign N515 = (N76)? N489 : 
                (N84)? 1'b0 : 1'b0;
  assign N516 = (N76)? N490 : 
                (N84)? 1'b1 : 1'b0;
  assign N517 = (N76)? N491 : 
                (N84)? 1'b0 : 1'b0;
  assign N518 = (N76)? N492 : 
                (N84)? 1'b0 : 1'b0;
  assign N519 = (N76)? N493 : 
                (N84)? 1'b0 : 1'b0;
  assign data_type_o = (N76)? { N495, N494 } : 
                       (N84)? { 1'b0, 1'b0 } : 1'b0;
  assign regfile_wdata_sel_o = (N76)? { N497, N496 } : 
                               (N84)? { 1'b0, 1'b1 } : 1'b0;
  assign data_sign_extension_o = (N76)? N498 : 
                                 (N84)? 1'b0 : 1'b0;
  assign imm_a_mux_sel_o = (N76)? N499 : 
                           (N84)? 1'b1 : 1'b0;
  assign multdiv_signed_mode_o = (N76)? { N501, N500 } : 
                                 (N84)? { 1'b0, 1'b0 } : 1'b0;
  assign N520 = (N76)? N503 : 
                (N84)? 1'b0 : 1'b0;
  assign multdiv_operator_o = (N76)? { N503, N502 } : 
                              (N84)? { 1'b0, 1'b0 } : 1'b0;
  assign N521 = (N76)? N504 : 
                (N84)? 1'b0 : 1'b0;
  assign csr_status_o = (N76)? N505 : 
                        (N84)? 1'b0 : 1'b0;
  assign dret_insn_o = (N76)? N506 : 
                       (N84)? 1'b0 : 1'b0;
  assign wfi_insn_o = (N76)? N507 : 
                      (N84)? 1'b0 : 1'b0;
  assign ecall_insn_o = (N76)? N508 : 
                        (N84)? 1'b0 : 1'b0;
  assign ebrk_insn_o = (N76)? N509 : 
                       (N84)? 1'b0 : 1'b0;
  assign mret_insn_o = (N76)? N510 : 
                       (N84)? 1'b0 : 1'b0;
  assign illegal_insn = (N77)? 1'b1 : 
                        (N78)? N516 : 1'b0;
  assign N77 = illegal_c_insn_i;
  assign N78 = N522;
  assign regfile_we = (N79)? 1'b0 : 
                      (N80)? N515 : 1'b0;
  assign N79 = illegal_insn;
  assign N80 = N523;
  assign data_req_o = (N79)? 1'b0 : 
                      (N80)? N518 : 1'b0;
  assign data_we_o = (N79)? 1'b0 : 
                     (N80)? N519 : 1'b0;
  assign mult_en_o = (N79)? 1'b0 : 
                     (N80)? N521 : 1'b0;
  assign div_en_o = (N79)? 1'b0 : 
                    (N80)? N520 : 1'b0;
  assign jump_in_dec_o = (N79)? 1'b0 : 
                         (N80)? N514 : 1'b0;
  assign branch_in_dec_o = (N79)? 1'b0 : 
                           (N80)? N517 : 1'b0;
  assign csr_access_o = (N79)? 1'b0 : 
                        (N80)? N513 : 1'b0;
  assign N81 = N635 & N532;
  assign N635 = N526 | N527;
  assign N82 = ~N81;
  assign N84 = ~N83;
  assign N89 = ~N88;
  assign N93 = ~N92;
  assign N95 = ~N94;
  assign N99 = ~N98;
  assign N100 = ~instr_rdata_i[6];
  assign N101 = ~instr_rdata_i[5];
  assign N102 = ~instr_rdata_i[4];
  assign N103 = ~instr_rdata_i[3];
  assign N104 = ~instr_rdata_i[2];
  assign N112 = ~N111;
  assign N116 = ~N115;
  assign N118 = ~N117;
  assign N120 = ~N119;
  assign N123 = ~N122;
  assign N126 = ~N125;
  assign N141 = N127 | N641;
  assign N641 = N129 | N640;
  assign N640 = N131 | N639;
  assign N639 = N133 | N638;
  assign N638 = N136 | N637;
  assign N637 = N138 | N636;
  assign N636 = N139 | N140;
  assign N142 = ~instr_rdata_i[14];
  assign N147 = ~N146;
  assign N150 = ~N149;
  assign N153 = ~N152;
  assign N156 = ~N155;
  assign N160 = ~N159;
  assign N167 = ~instr_new_i;
  assign N175 = ~N174;
  assign N177 = ~N176;
  assign N182 = ~N181;
  assign N183 = ~N611;
  assign N184 = ~instr_rdata_i[31];
  assign N185 = ~instr_rdata_i[26];
  assign N189 = ~N188;
  assign N194 = N191 | N642;
  assign N642 = ~N193;
  assign N199 = N643 | N644;
  assign N643 = ~N196;
  assign N644 = ~N198;
  assign N202 = ~N201;
  assign N205 = N203 | N204;
  assign N218 = ~instr_rdata_i[14];
  assign N219 = ~instr_rdata_i[13];
  assign N220 = ~instr_rdata_i[12];
  assign N225 = ~N224;
  assign N228 = ~N227;
  assign N231 = ~N230;
  assign N234 = ~N233;
  assign N239 = ~N238;
  assign N242 = ~N241;
  assign N243 = N624 | N631;
  assign N244 = ~N243;
  assign N254 = ~instr_rdata_i[31];
  assign N258 = ~N257;
  assign N267 = ~N266;
  assign N272 = ~N271;
  assign N277 = ~N276;
  assign N282 = ~N281;
  assign N287 = ~N286;
  assign N292 = ~N291;
  assign N297 = ~N296;
  assign N302 = ~N301;
  assign N307 = ~N306;
  assign N312 = ~N311;
  assign N317 = ~N316;
  assign N322 = ~N321;
  assign N327 = ~N326;
  assign N332 = ~N331;
  assign N337 = ~N336;
  assign N342 = ~N341;
  assign N347 = ~N346;
  assign N354 = N349 | N646;
  assign N646 = N350 | N645;
  assign N645 = N352 | N353;
  assign N384 = ~instr_rdata_i[23];
  assign N387 = ~N386;
  assign N388 = ~instr_rdata_i[22];
  assign N405 = ~N404;
  assign N414 = ~N413;
  assign N423 = ~N422;
  assign N432 = ~N431;
  assign N433 = N405 | N396;
  assign N434 = N414 | N433;
  assign N435 = N423 | N434;
  assign N436 = N432 | N435;
  assign N437 = ~N436;
  assign N450 = N650 | N654;
  assign N650 = N649 | instr_rdata_i[15];
  assign N649 = N648 | instr_rdata_i[16];
  assign N648 = N647 | instr_rdata_i[17];
  assign N647 = instr_rdata_i[19] | instr_rdata_i[18];
  assign N654 = N653 | instr_rdata_i[7];
  assign N653 = N652 | instr_rdata_i[8];
  assign N652 = N651 | instr_rdata_i[9];
  assign N651 = instr_rdata_i[11] | instr_rdata_i[10];
  assign N451 = ~N450;
  assign N454 = ~N453;
  assign N456 = ~N455;
  assign N462 = ~N461;
  assign N463 = N657 | N600;
  assign N657 = N656 | N588;
  assign N656 = N655 | N575;
  assign N655 = N546 | N562;
  assign N486 = N94;
  assign N522 = ~illegal_c_insn_i;
  assign N523 = ~illegal_insn;
  assign illegal_insn_o = illegal_insn | 1'b0;
  assign regfile_we_o = regfile_we & N658;
  assign N658 = ~1'b0;

endmodule



module ibex_controller
(
  clk_i,
  rst_ni,
  fetch_enable_i,
  ctrl_busy_o,
  first_fetch_o,
  illegal_insn_i,
  ecall_insn_i,
  mret_insn_i,
  dret_insn_i,
  wfi_insn_i,
  ebrk_insn_i,
  csr_status_i,
  instr_valid_i,
  instr_i,
  instr_compressed_i,
  instr_is_compressed_i,
  instr_valid_clear_o,
  id_in_ready_o,
  instr_req_o,
  pc_set_o,
  pc_mux_o,
  exc_pc_mux_o,
  lsu_addr_last_i,
  load_err_i,
  store_err_i,
  branch_set_i,
  jump_set_i,
  irq_i,
  irq_req_ctrl_i,
  irq_id_ctrl_i,
  m_IE_i,
  irq_ack_o,
  irq_id_o,
  exc_cause_o,
  exc_ack_o,
  exc_kill_o,
  debug_req_i,
  debug_cause_o,
  debug_csr_save_o,
  debug_single_step_i,
  debug_ebreakm_i,
  csr_save_if_o,
  csr_save_id_o,
  csr_restore_mret_id_o,
  csr_restore_dret_id_o,
  csr_save_cause_o,
  csr_mtval_o,
  stall_lsu_i,
  stall_multdiv_i,
  stall_jump_i,
  stall_branch_i,
  perf_jump_o,
  perf_tbranch_o
);

  input [31:0] instr_i;
  input [15:0] instr_compressed_i;
  output [2:0] pc_mux_o;
  output [1:0] exc_pc_mux_o;
  input [31:0] lsu_addr_last_i;
  input [4:0] irq_id_ctrl_i;
  output [4:0] irq_id_o;
  output [5:0] exc_cause_o;
  output [2:0] debug_cause_o;
  output [31:0] csr_mtval_o;
  input clk_i;
  input rst_ni;
  input fetch_enable_i;
  input illegal_insn_i;
  input ecall_insn_i;
  input mret_insn_i;
  input dret_insn_i;
  input wfi_insn_i;
  input ebrk_insn_i;
  input csr_status_i;
  input instr_valid_i;
  input instr_is_compressed_i;
  input load_err_i;
  input store_err_i;
  input branch_set_i;
  input jump_set_i;
  input irq_i;
  input irq_req_ctrl_i;
  input m_IE_i;
  input debug_req_i;
  input debug_single_step_i;
  input debug_ebreakm_i;
  input stall_lsu_i;
  input stall_multdiv_i;
  input stall_jump_i;
  input stall_branch_i;
  output ctrl_busy_o;
  output first_fetch_o;
  output instr_valid_clear_o;
  output id_in_ready_o;
  output instr_req_o;
  output pc_set_o;
  output irq_ack_o;
  output exc_ack_o;
  output exc_kill_o;
  output debug_csr_save_o;
  output csr_save_if_o;
  output csr_save_id_o;
  output csr_restore_mret_id_o;
  output csr_restore_dret_id_o;
  output csr_save_cause_o;
  output perf_jump_o;
  output perf_tbranch_o;
  wire [2:0] pc_mux_o,debug_cause_o;
  wire [1:0] exc_pc_mux_o;
  wire [4:0] irq_id_o;
  wire [5:0] exc_cause_o;
  wire [31:0] csr_mtval_o;
  wire ctrl_busy_o,first_fetch_o,instr_valid_clear_o,id_in_ready_o,instr_req_o,
  pc_set_o,irq_ack_o,exc_ack_o,exc_kill_o,debug_csr_save_o,csr_save_if_o,csr_save_id_o,
  csr_restore_mret_id_o,csr_restore_dret_id_o,csr_save_cause_o,perf_jump_o,
  perf_tbranch_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,
  N21,N22,exc_ack_o,exc_req,exc_req_lsu,special_req,enter_debug_mode,handle_irq,
  stall,N23,N24,N25,halt_if,halt_id,debug_mode_d,N26,N27,N28,N29,N30,N31,N32,N33,N34,
  N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,
  N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,
  N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,
  N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,
  N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,
  N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,
  N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,
  N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,
  N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,
  N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,
  N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,
  N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,
  N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,
  N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,
  N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,
  N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,
  N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,
  N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,
  N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
  N352,N353,N354,N355;
  wire [3:0] ctrl_fsm_ns;
  reg load_err_q,store_err_q,debug_mode_q;
  reg [3:0] ctrl_fsm_cs;
  assign exc_kill_o = 1'b0;
  assign irq_id_o[4] = irq_id_ctrl_i[4];
  assign irq_id_o[3] = irq_id_ctrl_i[3];
  assign irq_id_o[2] = irq_id_ctrl_i[2];
  assign irq_id_o[1] = irq_id_ctrl_i[1];
  assign irq_id_o[0] = irq_id_ctrl_i[0];
  assign irq_ack_o = exc_ack_o;
  assign N30 = N26 & N27;
  assign N31 = N28 & N29;
  assign N32 = N30 & N31;
  assign N33 = ctrl_fsm_cs[3] | ctrl_fsm_cs[2];
  assign N34 = ctrl_fsm_cs[1] | N29;
  assign N35 = N33 | N34;
  assign N37 = ctrl_fsm_cs[3] | ctrl_fsm_cs[2];
  assign N38 = N28 | ctrl_fsm_cs[0];
  assign N39 = N37 | N38;
  assign N41 = ctrl_fsm_cs[3] | ctrl_fsm_cs[2];
  assign N42 = N28 | N29;
  assign N43 = N41 | N42;
  assign N45 = ctrl_fsm_cs[3] | N27;
  assign N46 = ctrl_fsm_cs[1] | ctrl_fsm_cs[0];
  assign N47 = N45 | N46;
  assign N49 = ctrl_fsm_cs[3] | N27;
  assign N50 = ctrl_fsm_cs[1] | N29;
  assign N51 = N49 | N50;
  assign N53 = ctrl_fsm_cs[3] | N27;
  assign N54 = N28 | N29;
  assign N55 = N53 | N54;
  assign N57 = N26 | ctrl_fsm_cs[2];
  assign N58 = ctrl_fsm_cs[1] | ctrl_fsm_cs[0];
  assign N59 = N57 | N58;
  assign N61 = N26 | ctrl_fsm_cs[2];
  assign N62 = ctrl_fsm_cs[1] | N29;
  assign N63 = N61 | N62;
  assign N65 = ctrl_fsm_cs[3] | N27;
  assign N66 = N28 | ctrl_fsm_cs[0];
  assign N67 = N65 | N66;
  assign N69 = ctrl_fsm_cs[3] & ctrl_fsm_cs[1];
  assign N70 = ctrl_fsm_cs[3] & ctrl_fsm_cs[2];

  always @(posedge clk_i or posedge N319) begin
    if(N319) begin
      load_err_q <= 1'b0;
    end else if(1'b1) begin
      load_err_q <= load_err_i;
    end 
  end


  always @(posedge clk_i or posedge N319) begin
    if(N319) begin
      store_err_q <= 1'b0;
    end else if(1'b1) begin
      store_err_q <= store_err_i;
    end 
  end


  always @(posedge clk_i or posedge N319) begin
    if(N319) begin
      ctrl_fsm_cs[3] <= 1'b0;
    end else if(N323) begin
      ctrl_fsm_cs[3] <= ctrl_fsm_ns[3];
    end 
  end


  always @(posedge clk_i or posedge N319) begin
    if(N319) begin
      ctrl_fsm_cs[2] <= 1'b0;
    end else if(N323) begin
      ctrl_fsm_cs[2] <= ctrl_fsm_ns[2];
    end 
  end


  always @(posedge clk_i or posedge N319) begin
    if(N319) begin
      ctrl_fsm_cs[1] <= 1'b0;
    end else if(N323) begin
      ctrl_fsm_cs[1] <= ctrl_fsm_ns[1];
    end 
  end


  always @(posedge clk_i or posedge N319) begin
    if(N319) begin
      ctrl_fsm_cs[0] <= 1'b0;
    end else if(N323) begin
      ctrl_fsm_cs[0] <= ctrl_fsm_ns[0];
    end 
  end


  always @(posedge clk_i or posedge N319) begin
    if(N319) begin
      debug_mode_q <= 1'b0;
    end else if(N341) begin
      debug_mode_q <= debug_mode_d;
    end 
  end

  assign { N79, N78, N77, N76 } = (N0)? { 1'b0, 1'b1, 1'b0, 1'b1 } : 
                                  (N1)? ctrl_fsm_cs : 1'b0;
  assign N0 = id_in_ready_o;
  assign N1 = N75;
  assign { N84, N83, N82, N81 } = (N2)? { 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                  (N3)? { N79, N78, N77, N76 } : 1'b0;
  assign N2 = handle_irq;
  assign N3 = N80;
  assign { N89, N88, N87, N86 } = (N4)? { 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                  (N5)? { N84, N83, N82, N81 } : 1'b0;
  assign N4 = enter_debug_mode;
  assign N5 = N85;
  assign N90 = (N4)? 1'b1 : 
               (N5)? handle_irq : 1'b0;
  assign N96 = (N6)? 1'b1 : 
               (N95)? 1'b0 : 
               (N7)? 1'b0 : 1'b0;
  assign N6 = N92;
  assign N7 = 1'b0;
  assign N97 = (N6)? branch_set_i : 
               (N95)? 1'b0 : 
               (N7)? 1'b0 : 1'b0;
  assign N98 = (N6)? jump_set_i : 
               (N95)? 1'b0 : 
               (N7)? 1'b0 : 1'b0;
  assign { N102, N101, N100, N99 } = (N6)? ctrl_fsm_cs : 
                                     (N299)? { 1'b0, 1'b1, 1'b1, 1'b0 } : 
                                     (N94)? ctrl_fsm_cs : 1'b0;
  assign N103 = (N6)? 1'b0 : 
                (N299)? 1'b1 : 
                (N94)? 1'b0 : 1'b0;
  assign N106 = (N8)? 1'b1 : 
                (N105)? N103 : 1'b0;
  assign N8 = N104;
  assign { N113, N112, N111, N110 } = (N9)? { 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                      (N109)? { N102, N101, N100, N99 } : 1'b0;
  assign N9 = N108;
  assign N114 = (N10)? 1'b1 : 
                (N107)? N106 : 1'b0;
  assign N10 = N25;
  assign { N118, N117, N116, N115 } = (N10)? { N113, N112, N111, N110 } : 
                                      (N107)? { N102, N101, N100, N99 } : 1'b0;
  assign N119 = (N11)? N103 : 
                (N12)? 1'b0 : 1'b0;
  assign N11 = instr_valid_i;
  assign N12 = N91;
  assign N120 = (N11)? N96 : 
                (N12)? 1'b0 : 1'b0;
  assign N121 = (N11)? N97 : 
                (N12)? 1'b0 : 1'b0;
  assign N122 = (N11)? N98 : 
                (N12)? 1'b0 : 1'b0;
  assign { N126, N125, N124, N123 } = (N11)? { N118, N117, N116, N115 } : 
                                      (N12)? ctrl_fsm_cs : 1'b0;
  assign N127 = (N11)? N114 : 
                (N12)? 1'b0 : 1'b0;
  assign { N135, N134, N133, N132 } = (N4)? { 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                      (N301)? { 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                      (N131)? { N126, N125, N124, N123 } : 1'b0;
  assign N136 = (N4)? 1'b1 : 
                (N301)? 1'b1 : 
                (N131)? N127 : 1'b0;
  assign N137 = (N4)? 1'b1 : 
                (N301)? 1'b1 : 
                (N131)? N119 : 1'b0;
  assign N138 = (N13)? N137 : 
                (N129)? N119 : 1'b0;
  assign N13 = N128;
  assign { N142, N141, N140, N139 } = (N13)? { N135, N134, N133, N132 } : 
                                      (N129)? { N126, N125, N124, N123 } : 1'b0;
  assign N143 = (N13)? N136 : 
                (N129)? N127 : 1'b0;
  assign N147 = ~N144;
  assign { N150, N149, N148 } = (N14)? { debug_single_step_i, N146, N146 } : 
                                (N145)? { 1'b0, 1'b0, 1'b1 } : 1'b0;
  assign N14 = N144;
  assign N153 = (N15)? N152 : 
                (N16)? 1'b0 : 1'b0;
  assign N15 = ebrk_insn_i;
  assign N16 = N151;
  assign { N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165 } = (N17)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, instr_compressed_i } : 
                                                                                                                                                                                                              (N18)? instr_i : 1'b0;
  assign N17 = instr_is_compressed_i;
  assign N18 = N164;
  assign N199 = (N19)? 1'b0 : 
                (N318)? 1'b0 : 
                (N198)? 1'b1 : 1'b0;
  assign N19 = debug_mode_q;
  assign N200 = (N19)? 1'b1 : 
                (N318)? 1'b1 : 
                (N198)? 1'b0 : 1'b0;
  assign { N204, N201 } = (N20)? { 1'b0, 1'b0 } : 
                          (N205)? { 1'b0, 1'b1 } : 
                          (N310)? { 1'b0, N199 } : 
                          (N313)? { 1'b1, 1'b1 } : 
                          (N316)? { 1'b1, 1'b1 } : 
                          (N163)? { 1'b0, 1'b0 } : 1'b0;
  assign N20 = illegal_insn_i;
  assign N203 = (N20)? 1'b1 : 
                (N205)? 1'b1 : 
                (N310)? N199 : 
                (N313)? 1'b1 : 
                (N202)? 1'b0 : 
                (N7)? 1'b0 : 1'b0;
  assign { N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206 } = (N20)? { N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165 } : 
                                                                                                                                                                                                              (N205)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                              (N310)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                              (N313)? lsu_addr_last_i : 
                                                                                                                                                                                                              (N316)? lsu_addr_last_i : 
                                                                                                                                                                                                              (N163)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N239 = (N20)? 1'b1 : 
                (N205)? 1'b1 : 
                (N310)? N199 : 
                (N238)? 1'b1 : 
                (N7)? 1'b1 : 
                (N7)? 1'b1 : 1'b0;
  assign N240 = (N20)? 1'b0 : 
                (N205)? 1'b0 : 
                (N310)? N200 : 
                (N238)? 1'b0 : 
                (N7)? 1'b0 : 
                (N7)? 1'b0 : 1'b0;
  assign N242 = (N21)? N239 : 
                (N243)? 1'b1 : 
                (N246)? 1'b1 : 
                (N241)? 1'b0 : 
                (N7)? 1'b0 : 1'b0;
  assign N21 = N154;
  assign N245 = (N21)? 1'b1 : 
                (N243)? 1'b1 : 
                (N244)? 1'b0 : 
                (N7)? 1'b0 : 
                (N7)? 1'b0 : 1'b0;
  assign { N249, N248 } = (N21)? { debug_mode_q, debug_mode_q } : 
                          (N247)? { 1'b0, 1'b1 } : 
                          (N7)? { 1'b0, 1'b1 } : 
                          (N7)? { 1'b0, 1'b1 } : 
                          (N7)? { 1'b0, 1'b1 } : 1'b0;
  assign N250 = (N21)? N239 : 
                (N247)? 1'b0 : 
                (N7)? 1'b0 : 
                (N7)? 1'b0 : 
                (N7)? 1'b0 : 1'b0;
  assign { N253, N252, N251 } = (N21)? { N239, 1'b0, 1'b1 } : 
                                (N243)? { 1'b1, 1'b0, 1'b1 } : 
                                (N246)? { 1'b1, 1'b0, 1'b1 } : 
                                (N306)? { 1'b0, 1'b1, 1'b0 } : 
                                (N158)? { 1'b1, 1'b0, 1'b1 } : 1'b0;
  assign N254 = (N21)? N240 : 
                (N247)? 1'b0 : 
                (N7)? 1'b0 : 
                (N7)? 1'b0 : 
                (N7)? 1'b0 : 1'b0;
  assign { N258, N257, N256, N255 } = (N21)? { N205, N204, N203, N201 } : 
                                      (N247)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N7)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N7)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N7)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259 } = (N21)? { N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206 } : 
                                                                                                                                                                                                              (N247)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                              (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                              (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                              (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N291 = (N21)? 1'b0 : 
                (N243)? 1'b1 : 
                (N244)? 1'b0 : 
                (N7)? 1'b0 : 
                (N7)? 1'b0 : 1'b0;
  assign N292 = (N21)? 1'b0 : 
                (N243)? 1'b0 : 
                (N246)? 1'b1 : 
                (N241)? 1'b0 : 
                (N7)? 1'b0 : 1'b0;
  assign N293 = (N10)? 1'b0 : 
                (N107)? N242 : 1'b0;
  assign { N297, N296, N295, N294 } = (N10)? { 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                      (N107)? { N254, N253, N252, N251 } : 1'b0;
  assign instr_req_o = (N22)? 1'b0 : 
                       (N36)? 1'b1 : 
                       (N40)? 1'b0 : 
                       (N44)? 1'b0 : 
                       (N48)? 1'b1 : 
                       (N52)? 1'b1 : 
                       (N56)? 1'b1 : 
                       (N60)? 1'b1 : 
                       (N64)? 1'b1 : 
                       (N68)? 1'b1 : 
                       (N71)? 1'b0 : 1'b0;
  assign N22 = N32;
  assign pc_mux_o[1:0] = (N22)? { 1'b0, 1'b0 } : 
                         (N36)? { 1'b0, 1'b0 } : 
                         (N40)? { 1'b0, 1'b0 } : 
                         (N44)? { 1'b0, 1'b0 } : 
                         (N48)? { 1'b0, 1'b0 } : 
                         (N52)? { 1'b0, N120 } : 
                         (N56)? { 1'b1, 1'b0 } : 
                         (N60)? { N144, 1'b0 } : 
                         (N64)? { ebrk_insn_i, 1'b0 } : 
                         (N68)? { N245, N243 } : 
                         (N71)? { 1'b0, 1'b0 } : 1'b0;
  assign pc_mux_o[2] = (N68)? N246 : 
                       (N298)? 1'b0 : 1'b0;
  assign pc_set_o = (N22)? 1'b1 : 
                    (N36)? 1'b1 : 
                    (N40)? 1'b0 : 
                    (N44)? 1'b0 : 
                    (N48)? 1'b0 : 
                    (N52)? N120 : 
                    (N56)? 1'b1 : 
                    (N60)? N144 : 
                    (N64)? ebrk_insn_i : 
                    (N68)? N293 : 
                    (N71)? 1'b0 : 1'b0;
  assign ctrl_fsm_ns[0] = (N22)? 1'b1 : 
                          (N36)? 1'b0 : 
                          (N40)? 1'b1 : 
                          (N44)? 1'b0 : 
                          (N48)? N86 : 
                          (N52)? N139 : 
                          (N56)? 1'b1 : 
                          (N60)? 1'b1 : 
                          (N64)? 1'b1 : 
                          (N68)? N294 : 1'b0;
  assign ctrl_fsm_ns[3:1] = (N22)? { 1'b0, 1'b0, 1'b0 } : 
                            (N36)? { 1'b0, 1'b1, 1'b0 } : 
                            (N40)? { 1'b0, 1'b0, 1'b1 } : 
                            (N44)? { 1'b0, 1'b1, 1'b0 } : 
                            (N48)? { N89, N88, N87 } : 
                            (N52)? { N142, N141, N140 } : 
                            (N56)? { 1'b0, 1'b1, 1'b0 } : 
                            (N60)? { 1'b0, 1'b1, 1'b0 } : 
                            (N64)? { 1'b0, 1'b1, 1'b0 } : 
                            (N68)? { N297, N296, N295 } : 
                            (N71)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign ctrl_busy_o = (N22)? 1'b1 : 
                       (N36)? 1'b1 : 
                       (N40)? 1'b0 : 
                       (N44)? 1'b0 : 
                       (N48)? 1'b1 : 
                       (N52)? 1'b1 : 
                       (N56)? 1'b1 : 
                       (N60)? 1'b1 : 
                       (N64)? 1'b1 : 
                       (N68)? 1'b1 : 
                       (N71)? 1'b1 : 1'b0;
  assign halt_if = (N22)? 1'b0 : 
                   (N36)? 1'b0 : 
                   (N40)? 1'b1 : 
                   (N44)? 1'b1 : 
                   (N48)? N90 : 
                   (N52)? N143 : 
                   (N56)? 1'b0 : 
                   (N60)? 1'b0 : 
                   (N64)? 1'b0 : 
                   (N68)? 1'b1 : 
                   (N71)? 1'b0 : 1'b0;
  assign halt_id = (N22)? 1'b0 : 
                   (N36)? 1'b0 : 
                   (N40)? 1'b1 : 
                   (N44)? 1'b1 : 
                   (N48)? N90 : 
                   (N52)? N138 : 
                   (N56)? 1'b0 : 
                   (N60)? 1'b0 : 
                   (N64)? 1'b0 : 
                   (N68)? 1'b1 : 
                   (N71)? 1'b0 : 1'b0;
  assign first_fetch_o = (N22)? 1'b0 : 
                         (N36)? 1'b0 : 
                         (N40)? 1'b0 : 
                         (N44)? 1'b0 : 
                         (N48)? 1'b1 : 
                         (N52)? 1'b0 : 
                         (N56)? 1'b0 : 
                         (N60)? 1'b0 : 
                         (N64)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N71)? 1'b0 : 1'b0;
  assign perf_tbranch_o = (N22)? 1'b0 : 
                          (N36)? 1'b0 : 
                          (N40)? 1'b0 : 
                          (N44)? 1'b0 : 
                          (N48)? 1'b0 : 
                          (N52)? N121 : 
                          (N56)? 1'b0 : 
                          (N60)? 1'b0 : 
                          (N64)? 1'b0 : 
                          (N68)? 1'b0 : 
                          (N71)? 1'b0 : 1'b0;
  assign perf_jump_o = (N22)? 1'b0 : 
                       (N36)? 1'b0 : 
                       (N40)? 1'b0 : 
                       (N44)? 1'b0 : 
                       (N48)? 1'b0 : 
                       (N52)? N122 : 
                       (N56)? 1'b0 : 
                       (N60)? 1'b0 : 
                       (N64)? 1'b0 : 
                       (N68)? 1'b0 : 
                       (N71)? 1'b0 : 1'b0;
  assign exc_pc_mux_o = (N22)? { 1'b0, 1'b1 } : 
                        (N36)? { 1'b0, 1'b1 } : 
                        (N40)? { 1'b0, 1'b1 } : 
                        (N44)? { 1'b0, 1'b1 } : 
                        (N48)? { 1'b0, 1'b1 } : 
                        (N52)? { 1'b0, 1'b1 } : 
                        (N56)? { 1'b0, 1'b1 } : 
                        (N60)? { N144, N147 } : 
                        (N64)? { ebrk_insn_i, N151 } : 
                        (N68)? { N249, N248 } : 
                        (N71)? { 1'b0, 1'b1 } : 1'b0;
  assign exc_cause_o = (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N36)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N40)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N44)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N48)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N52)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N56)? { 1'b1, irq_id_ctrl_i } : 
                       (N60)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N64)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N68)? { 1'b0, 1'b0, N258, N257, N256, N255 } : 
                       (N71)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign csr_save_cause_o = (N22)? 1'b0 : 
                            (N36)? 1'b0 : 
                            (N40)? 1'b0 : 
                            (N44)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N56)? 1'b1 : 
                            (N60)? N144 : 
                            (N64)? N153 : 
                            (N68)? N250 : 
                            (N71)? 1'b0 : 1'b0;
  assign csr_save_if_o = (N22)? 1'b0 : 
                         (N36)? 1'b0 : 
                         (N40)? 1'b0 : 
                         (N44)? 1'b0 : 
                         (N48)? 1'b0 : 
                         (N52)? 1'b0 : 
                         (N56)? 1'b1 : 
                         (N60)? N144 : 
                         (N64)? 1'b0 : 
                         (N68)? 1'b0 : 
                         (N71)? 1'b0 : 1'b0;
  assign exc_ack_o = (N22)? 1'b0 : 
                     (N36)? 1'b0 : 
                     (N40)? 1'b0 : 
                     (N44)? 1'b0 : 
                     (N48)? 1'b0 : 
                     (N52)? 1'b0 : 
                     (N56)? 1'b1 : 
                     (N60)? 1'b0 : 
                     (N64)? 1'b0 : 
                     (N68)? 1'b0 : 
                     (N71)? 1'b0 : 1'b0;
  assign debug_mode_d = (N60)? 1'b1 : 
                        (N64)? 1'b1 : 
                        (N68)? 1'b0 : 1'b0;
  assign debug_csr_save_o = (N22)? 1'b0 : 
                            (N36)? 1'b0 : 
                            (N40)? 1'b0 : 
                            (N44)? 1'b0 : 
                            (N48)? 1'b0 : 
                            (N52)? 1'b0 : 
                            (N56)? 1'b0 : 
                            (N60)? N144 : 
                            (N64)? N153 : 
                            (N68)? 1'b0 : 
                            (N71)? 1'b0 : 1'b0;
  assign debug_cause_o = (N22)? { 1'b0, 1'b0, 1'b1 } : 
                         (N36)? { 1'b0, 1'b0, 1'b1 } : 
                         (N40)? { 1'b0, 1'b0, 1'b1 } : 
                         (N44)? { 1'b0, 1'b0, 1'b1 } : 
                         (N48)? { 1'b0, 1'b0, 1'b1 } : 
                         (N52)? { 1'b0, 1'b0, 1'b1 } : 
                         (N56)? { 1'b0, 1'b0, 1'b1 } : 
                         (N60)? { N150, N149, N148 } : 
                         (N64)? { 1'b0, 1'b0, 1'b1 } : 
                         (N68)? { 1'b0, 1'b0, 1'b1 } : 
                         (N71)? { 1'b0, 1'b0, 1'b1 } : 1'b0;
  assign csr_save_id_o = (N22)? 1'b0 : 
                         (N36)? 1'b0 : 
                         (N40)? 1'b0 : 
                         (N44)? 1'b0 : 
                         (N48)? 1'b0 : 
                         (N52)? 1'b0 : 
                         (N56)? 1'b0 : 
                         (N60)? 1'b0 : 
                         (N64)? N153 : 
                         (N68)? N250 : 
                         (N71)? 1'b0 : 1'b0;
  assign csr_mtval_o = (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N36)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N40)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N44)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N48)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N52)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N56)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N60)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N64)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                       (N68)? { N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259 } : 
                       (N71)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign csr_restore_mret_id_o = (N22)? 1'b0 : 
                                 (N36)? 1'b0 : 
                                 (N40)? 1'b0 : 
                                 (N44)? 1'b0 : 
                                 (N48)? 1'b0 : 
                                 (N52)? 1'b0 : 
                                 (N56)? 1'b0 : 
                                 (N60)? 1'b0 : 
                                 (N64)? 1'b0 : 
                                 (N68)? N291 : 
                                 (N71)? 1'b0 : 1'b0;
  assign csr_restore_dret_id_o = (N22)? 1'b0 : 
                                 (N36)? 1'b0 : 
                                 (N40)? 1'b0 : 
                                 (N44)? 1'b0 : 
                                 (N48)? 1'b0 : 
                                 (N52)? 1'b0 : 
                                 (N56)? 1'b0 : 
                                 (N60)? 1'b0 : 
                                 (N64)? 1'b0 : 
                                 (N68)? N292 : 
                                 (N71)? 1'b0 : 1'b0;
  assign exc_req = N342 | illegal_insn_i;
  assign N342 = ecall_insn_i | ebrk_insn_i;
  assign exc_req_lsu = store_err_i | load_err_i;
  assign special_req = N346 | exc_req_lsu;
  assign N346 = N345 | exc_req;
  assign N345 = N344 | csr_status_i;
  assign N344 = N343 | wfi_insn_i;
  assign N343 = mret_insn_i | dret_insn_i;
  assign enter_debug_mode = debug_req_i & N347;
  assign N347 = ~debug_mode_q;
  assign handle_irq = N348 & N347;
  assign N348 = irq_req_ctrl_i & m_IE_i;
  assign N23 = ~special_req;
  assign N24 = ~stall;
  assign N25 = debug_single_step_i & N347;
  assign N26 = ~ctrl_fsm_cs[3];
  assign N27 = ~ctrl_fsm_cs[2];
  assign N28 = ~ctrl_fsm_cs[1];
  assign N29 = ~ctrl_fsm_cs[0];
  assign N36 = ~N35;
  assign N40 = ~N39;
  assign N44 = ~N43;
  assign N48 = ~N47;
  assign N52 = ~N51;
  assign N56 = ~N55;
  assign N60 = ~N59;
  assign N64 = ~N63;
  assign N68 = ~N67;
  assign N71 = N69 | N70;
  assign N72 = ~fetch_enable_i;
  assign N73 = N350 | debug_single_step_i;
  assign N350 = N349 | debug_mode_q;
  assign N349 = irq_i | debug_req_i;
  assign N74 = ~N73;
  assign N75 = ~id_in_ready_o;
  assign N80 = ~handle_irq;
  assign N85 = ~enter_debug_mode;
  assign N91 = ~instr_valid_i;
  assign N92 = branch_set_i | jump_set_i;
  assign N93 = special_req | N92;
  assign N94 = ~N93;
  assign N95 = ~N92;
  assign N104 = N351 & stall;
  assign N351 = enter_debug_mode | handle_irq;
  assign N105 = ~N104;
  assign N107 = ~N25;
  assign N108 = N23 & N24;
  assign N109 = ~N108;
  assign N128 = N24 & N23;
  assign N129 = ~N128;
  assign N130 = handle_irq | enter_debug_mode;
  assign N131 = ~N130;
  assign N144 = debug_single_step_i | debug_req_i;
  assign N145 = ~N144;
  assign N146 = ~debug_single_step_i;
  assign N151 = ~ebrk_insn_i;
  assign N152 = debug_ebreakm_i & N347;
  assign N154 = N352 | load_err_q;
  assign N352 = exc_req | store_err_q;
  assign N155 = mret_insn_i | N154;
  assign N156 = dret_insn_i | N155;
  assign N157 = wfi_insn_i | N156;
  assign N158 = ~N157;
  assign N159 = ecall_insn_i | illegal_insn_i;
  assign N160 = ebrk_insn_i | N159;
  assign N161 = store_err_q | N160;
  assign N162 = load_err_q | N161;
  assign N163 = ~N162;
  assign N164 = ~instr_is_compressed_i;
  assign N197 = debug_ebreakm_i | debug_mode_q;
  assign N198 = ~N197;
  assign N202 = ~N161;
  assign N238 = ~N160;
  assign N241 = ~N156;
  assign N244 = ~N155;
  assign N247 = ~N154;
  assign N298 = N67;
  assign N299 = special_req & N95;
  assign N300 = ~enter_debug_mode;
  assign N301 = handle_irq & N300;
  assign N243 = mret_insn_i & N247;
  assign N302 = ~mret_insn_i;
  assign N303 = N247 & N302;
  assign N246 = dret_insn_i & N303;
  assign N304 = ~dret_insn_i;
  assign N305 = N303 & N304;
  assign N306 = wfi_insn_i & N305;
  assign N307 = ~illegal_insn_i;
  assign N205 = ecall_insn_i & N307;
  assign N308 = ~ecall_insn_i;
  assign N309 = N307 & N308;
  assign N310 = ebrk_insn_i & N309;
  assign N311 = ~ebrk_insn_i;
  assign N312 = N309 & N311;
  assign N313 = store_err_q & N312;
  assign N314 = ~store_err_q;
  assign N315 = N312 & N314;
  assign N316 = load_err_q & N315;
  assign N317 = ~debug_mode_q;
  assign N318 = debug_ebreakm_i & N317;
  assign stall = N354 | stall_branch_i;
  assign N354 = N353 | stall_jump_i;
  assign N353 = stall_lsu_i | stall_multdiv_i;
  assign id_in_ready_o = N24 & N355;
  assign N355 = ~halt_if;
  assign instr_valid_clear_o = N24 | halt_id;
  assign N319 = ~rst_ni;
  assign N320 = N72 & N32;
  assign N321 = N74 & N44;
  assign N322 = N320 | N321;
  assign N323 = ~N322;
  assign N324 = N32 | N36;
  assign N325 = N324 | N40;
  assign N326 = N325 | N44;
  assign N327 = N326 | N48;
  assign N328 = N327 | N52;
  assign N329 = N328 | N56;
  assign N330 = N145 & N60;
  assign N331 = N329 | N330;
  assign N332 = N151 & N64;
  assign N333 = N331 | N332;
  assign N334 = N154 & N68;
  assign N335 = N333 | N334;
  assign N336 = N243 & N68;
  assign N337 = N335 | N336;
  assign N338 = N241 & N68;
  assign N339 = N337 | N338;
  assign N340 = N339 | N71;
  assign N341 = ~N340;

endmodule



module ibex_int_controller
(
  clk_i,
  rst_ni,
  irq_req_ctrl_o,
  irq_id_ctrl_o,
  ctrl_ack_i,
  ctrl_kill_i,
  irq_i,
  irq_id_i,
  m_IE_i
);

  output [4:0] irq_id_ctrl_o;
  input [4:0] irq_id_i;
  input clk_i;
  input rst_ni;
  input ctrl_ack_i;
  input ctrl_kill_i;
  input irq_i;
  input m_IE_i;
  output irq_req_ctrl_o;
  wire irq_req_ctrl_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,
  N18,N19,N20,N21,N22,N23,N24,N25,N26;
  wire [1:0] exc_ctrl_ns;
  reg [1:0] exc_ctrl_cs;
  reg [4:0] irq_id_ctrl_o;

  always @(posedge clk_i or posedge N4) begin
    if(N4) begin
      exc_ctrl_cs[1] <= 1'b0;
    end else if(N20) begin
      exc_ctrl_cs[1] <= exc_ctrl_ns[1];
    end 
  end


  always @(posedge clk_i or posedge N4) begin
    if(N4) begin
      exc_ctrl_cs[0] <= 1'b0;
    end else if(N20) begin
      exc_ctrl_cs[0] <= exc_ctrl_ns[0];
    end 
  end


  always @(posedge clk_i or posedge N4) begin
    if(N4) begin
      irq_id_ctrl_o[4] <= 1'b0;
    end else if(N24) begin
      irq_id_ctrl_o[4] <= irq_id_i[4];
    end 
  end


  always @(posedge clk_i or posedge N4) begin
    if(N4) begin
      irq_id_ctrl_o[3] <= 1'b0;
    end else if(N24) begin
      irq_id_ctrl_o[3] <= irq_id_i[3];
    end 
  end


  always @(posedge clk_i or posedge N4) begin
    if(N4) begin
      irq_id_ctrl_o[2] <= 1'b0;
    end else if(N24) begin
      irq_id_ctrl_o[2] <= irq_id_i[2];
    end 
  end


  always @(posedge clk_i or posedge N4) begin
    if(N4) begin
      irq_id_ctrl_o[1] <= 1'b0;
    end else if(N24) begin
      irq_id_ctrl_o[1] <= irq_id_i[1];
    end 
  end


  always @(posedge clk_i or posedge N4) begin
    if(N4) begin
      irq_id_ctrl_o[0] <= 1'b0;
    end else if(N24) begin
      irq_id_ctrl_o[0] <= irq_id_i[0];
    end 
  end

  assign N7 = N5 & N6;
  assign N8 = exc_ctrl_cs[1] | N6;
  assign N10 = N5 | exc_ctrl_cs[0];
  assign N12 = exc_ctrl_cs[1] & exc_ctrl_cs[0];
  assign N25 = ~exc_ctrl_cs[0];
  assign N26 = N25 | exc_ctrl_cs[1];
  assign irq_req_ctrl_o = ~N26;
  assign { N18, N17 } = (N0)? { 1'b1, 1'b0 } : 
                        (N1)? { 1'b0, 1'b0 } : 
                        (N16)? { 1'b0, 1'b1 } : 1'b0;
  assign N0 = ctrl_ack_i;
  assign N1 = ctrl_kill_i;
  assign exc_ctrl_ns[0] = (N2)? 1'b1 : 
                          (N9)? N17 : 
                          (N11)? 1'b0 : 1'b0;
  assign N2 = N7;
  assign exc_ctrl_ns[1] = (N2)? 1'b0 : 
                          (N9)? N18 : 
                          (N11)? 1'b0 : 
                          (N3)? 1'b0 : 1'b0;
  assign N3 = N12;
  assign N4 = ~rst_ni;
  assign N5 = ~exc_ctrl_cs[1];
  assign N6 = ~exc_ctrl_cs[0];
  assign N9 = ~N8;
  assign N11 = ~N10;
  assign N13 = m_IE_i & irq_i;
  assign N14 = ~N13;
  assign N15 = ctrl_kill_i | ctrl_ack_i;
  assign N16 = ~N15;
  assign N19 = N14 & N7;
  assign N20 = ~N19;
  assign N21 = N19 | N9;
  assign N22 = N21 | N11;
  assign N23 = N22 | N12;
  assign N24 = ~N23;

endmodule



module ibex_id_stage_0_1
(
  clk_i,
  rst_ni,
  test_en_i,
  fetch_enable_i,
  ctrl_busy_o,
  core_ctrl_firstfetch_o,
  illegal_insn_o,
  instr_valid_i,
  instr_new_i,
  instr_rdata_i,
  instr_rdata_c_i,
  instr_is_compressed_i,
  instr_req_o,
  instr_valid_clear_o,
  id_in_ready_o,
  branch_decision_i,
  pc_set_o,
  pc_mux_o,
  exc_pc_mux_o,
  illegal_c_insn_i,
  pc_id_i,
  ex_valid_i,
  lsu_valid_i,
  alu_operator_ex_o,
  alu_operand_a_ex_o,
  alu_operand_b_ex_o,
  mult_en_ex_o,
  div_en_ex_o,
  multdiv_operator_ex_o,
  multdiv_signed_mode_ex_o,
  multdiv_operand_a_ex_o,
  multdiv_operand_b_ex_o,
  csr_access_o,
  csr_op_o,
  csr_save_if_o,
  csr_save_id_o,
  csr_restore_mret_id_o,
  csr_restore_dret_id_o,
  csr_save_cause_o,
  csr_mtval_o,
  illegal_csr_insn_i,
  data_req_ex_o,
  data_we_ex_o,
  data_type_ex_o,
  data_sign_ext_ex_o,
  data_reg_offset_ex_o,
  data_wdata_ex_o,
  lsu_addr_incr_req_i,
  lsu_addr_last_i,
  irq_i,
  irq_id_i,
  m_irq_enable_i,
  irq_ack_o,
  irq_id_o,
  exc_cause_o,
  lsu_load_err_i,
  lsu_store_err_i,
  debug_cause_o,
  debug_csr_save_o,
  debug_req_i,
  debug_single_step_i,
  debug_ebreakm_i,
  regfile_wdata_lsu_i,
  regfile_wdata_ex_i,
  csr_rdata_i,
  perf_jump_o,
  perf_branch_o,
  perf_tbranch_o,
  instr_ret_o,
  instr_ret_compressed_o
);

  input [31:0] instr_rdata_i;
  input [15:0] instr_rdata_c_i;
  output [2:0] pc_mux_o;
  output [1:0] exc_pc_mux_o;
  input [31:0] pc_id_i;
  output [4:0] alu_operator_ex_o;
  output [31:0] alu_operand_a_ex_o;
  output [31:0] alu_operand_b_ex_o;
  output [1:0] multdiv_operator_ex_o;
  output [1:0] multdiv_signed_mode_ex_o;
  output [31:0] multdiv_operand_a_ex_o;
  output [31:0] multdiv_operand_b_ex_o;
  output [1:0] csr_op_o;
  output [31:0] csr_mtval_o;
  output [1:0] data_type_ex_o;
  output [1:0] data_reg_offset_ex_o;
  output [31:0] data_wdata_ex_o;
  input [31:0] lsu_addr_last_i;
  input [4:0] irq_id_i;
  output [4:0] irq_id_o;
  output [5:0] exc_cause_o;
  output [2:0] debug_cause_o;
  input [31:0] regfile_wdata_lsu_i;
  input [31:0] regfile_wdata_ex_i;
  input [31:0] csr_rdata_i;
  input clk_i;
  input rst_ni;
  input test_en_i;
  input fetch_enable_i;
  input instr_valid_i;
  input instr_new_i;
  input instr_is_compressed_i;
  input branch_decision_i;
  input illegal_c_insn_i;
  input ex_valid_i;
  input lsu_valid_i;
  input illegal_csr_insn_i;
  input lsu_addr_incr_req_i;
  input irq_i;
  input m_irq_enable_i;
  input lsu_load_err_i;
  input lsu_store_err_i;
  input debug_req_i;
  input debug_single_step_i;
  input debug_ebreakm_i;
  output ctrl_busy_o;
  output core_ctrl_firstfetch_o;
  output illegal_insn_o;
  output instr_req_o;
  output instr_valid_clear_o;
  output id_in_ready_o;
  output pc_set_o;
  output mult_en_ex_o;
  output div_en_ex_o;
  output csr_access_o;
  output csr_save_if_o;
  output csr_save_id_o;
  output csr_restore_mret_id_o;
  output csr_restore_dret_id_o;
  output csr_save_cause_o;
  output data_req_ex_o;
  output data_we_ex_o;
  output data_sign_ext_ex_o;
  output irq_ack_o;
  output debug_csr_save_o;
  output perf_jump_o;
  output perf_branch_o;
  output perf_tbranch_o;
  output instr_ret_o;
  output instr_ret_compressed_o;
  wire [2:0] pc_mux_o,debug_cause_o,imm_b_mux_sel,imm_b_mux_sel_dec;
  wire [1:0] exc_pc_mux_o,multdiv_operator_ex_o,multdiv_signed_mode_ex_o,csr_op_o,
  data_type_ex_o,data_reg_offset_ex_o,alu_op_a_mux_sel,alu_op_a_mux_sel_dec,
  regfile_wdata_sel;
  wire [4:0] alu_operator_ex_o,irq_id_o,regfile_raddr_a,regfile_raddr_b,regfile_waddr,
  irq_id_ctrl;
  wire [31:0] alu_operand_a_ex_o,alu_operand_b_ex_o,multdiv_operand_a_ex_o,
  multdiv_operand_b_ex_o,csr_mtval_o,data_wdata_ex_o,imm_a,zimm_rs1_type,imm_b,imm_i_type,imm_s_type,
  imm_b_type,imm_u_type,imm_j_type,regfile_wdata;
  wire [5:0] exc_cause_o;
  wire ctrl_busy_o,core_ctrl_firstfetch_o,illegal_insn_o,instr_req_o,
  instr_valid_clear_o,id_in_ready_o,pc_set_o,mult_en_ex_o,div_en_ex_o,csr_access_o,csr_save_if_o,
  csr_save_id_o,csr_restore_mret_id_o,csr_restore_dret_id_o,csr_save_cause_o,
  data_req_ex_o,data_we_ex_o,data_sign_ext_ex_o,irq_ack_o,debug_csr_save_o,perf_jump_o,
  perf_branch_o,perf_tbranch_o,instr_ret_o,instr_ret_compressed_o,N0,N1,N2,N3,N4,N5,
  N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,
  N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,alu_op_b_mux_sel,
  alu_op_b_mux_sel_dec,N43,imm_a_mux_sel,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,
  N54,N55,N56,N57,N58,N59,N60,N61,instr_executing,N62,data_req_dec,multdiv_en_dec,
  N63,N64,N65,regfile_we,regfile_we_wb,regfile_we_dec,N66,N67,N68,illegal_insn_dec,
  ebrk_insn,mret_insn_dec,dret_insn_dec,ecall_insn_dec,wfi_insn_dec,jump_set,
  mult_en_dec,div_en_dec,csr_status,jump_in_dec,branch_in_dec,irq_req_ctrl,exc_ack,
  exc_kill,stall_lsu,stall_multdiv,stall_jump,stall_branch,N69,id_wb_fsm_ns,
  branch_set_n,instr_multicycle_done_n,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,
  N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111;
  reg branch_set_q,instr_multicycle_done_q,id_wb_fsm_cs;
  assign multdiv_operand_b_ex_o[31] = data_wdata_ex_o[31];
  assign multdiv_operand_b_ex_o[30] = data_wdata_ex_o[30];
  assign multdiv_operand_b_ex_o[29] = data_wdata_ex_o[29];
  assign multdiv_operand_b_ex_o[28] = data_wdata_ex_o[28];
  assign multdiv_operand_b_ex_o[27] = data_wdata_ex_o[27];
  assign multdiv_operand_b_ex_o[26] = data_wdata_ex_o[26];
  assign multdiv_operand_b_ex_o[25] = data_wdata_ex_o[25];
  assign multdiv_operand_b_ex_o[24] = data_wdata_ex_o[24];
  assign multdiv_operand_b_ex_o[23] = data_wdata_ex_o[23];
  assign multdiv_operand_b_ex_o[22] = data_wdata_ex_o[22];
  assign multdiv_operand_b_ex_o[21] = data_wdata_ex_o[21];
  assign multdiv_operand_b_ex_o[20] = data_wdata_ex_o[20];
  assign multdiv_operand_b_ex_o[19] = data_wdata_ex_o[19];
  assign multdiv_operand_b_ex_o[18] = data_wdata_ex_o[18];
  assign multdiv_operand_b_ex_o[17] = data_wdata_ex_o[17];
  assign multdiv_operand_b_ex_o[16] = data_wdata_ex_o[16];
  assign multdiv_operand_b_ex_o[15] = data_wdata_ex_o[15];
  assign multdiv_operand_b_ex_o[14] = data_wdata_ex_o[14];
  assign multdiv_operand_b_ex_o[13] = data_wdata_ex_o[13];
  assign multdiv_operand_b_ex_o[12] = data_wdata_ex_o[12];
  assign multdiv_operand_b_ex_o[11] = data_wdata_ex_o[11];
  assign multdiv_operand_b_ex_o[10] = data_wdata_ex_o[10];
  assign multdiv_operand_b_ex_o[9] = data_wdata_ex_o[9];
  assign multdiv_operand_b_ex_o[8] = data_wdata_ex_o[8];
  assign multdiv_operand_b_ex_o[7] = data_wdata_ex_o[7];
  assign multdiv_operand_b_ex_o[6] = data_wdata_ex_o[6];
  assign multdiv_operand_b_ex_o[5] = data_wdata_ex_o[5];
  assign multdiv_operand_b_ex_o[4] = data_wdata_ex_o[4];
  assign multdiv_operand_b_ex_o[3] = data_wdata_ex_o[3];
  assign multdiv_operand_b_ex_o[2] = data_wdata_ex_o[2];
  assign multdiv_operand_b_ex_o[1] = data_wdata_ex_o[1];
  assign multdiv_operand_b_ex_o[0] = data_wdata_ex_o[0];
  assign N46 = N44 & N45;
  assign N47 = alu_op_a_mux_sel[1] | N45;
  assign N49 = N44 | alu_op_a_mux_sel[0];
  assign N51 = alu_op_a_mux_sel[1] & alu_op_a_mux_sel[0];

  ibex_register_file_0
  registers_i
  (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .test_en_i(test_en_i),
    .raddr_a_i(regfile_raddr_a),
    .rdata_a_o(multdiv_operand_a_ex_o),
    .raddr_b_i(regfile_raddr_b),
    .rdata_b_o(data_wdata_ex_o),
    .waddr_a_i(regfile_waddr),
    .wdata_a_i(regfile_wdata),
    .we_a_i(regfile_we)
  );


  ibex_decoder_0_1
  decoder_i
  (
    .illegal_insn_o(illegal_insn_dec),
    .ebrk_insn_o(ebrk_insn),
    .mret_insn_o(mret_insn_dec),
    .dret_insn_o(dret_insn_dec),
    .ecall_insn_o(ecall_insn_dec),
    .wfi_insn_o(wfi_insn_dec),
    .jump_set_o(jump_set),
    .instr_new_i(instr_new_i),
    .instr_rdata_i(instr_rdata_i),
    .illegal_c_insn_i(illegal_c_insn_i),
    .imm_a_mux_sel_o(imm_a_mux_sel),
    .imm_b_mux_sel_o(imm_b_mux_sel_dec),
    .imm_i_type_o(imm_i_type),
    .imm_s_type_o(imm_s_type),
    .imm_b_type_o(imm_b_type),
    .imm_u_type_o(imm_u_type),
    .imm_j_type_o(imm_j_type),
    .zimm_rs1_type_o(zimm_rs1_type),
    .regfile_wdata_sel_o(regfile_wdata_sel),
    .regfile_we_o(regfile_we_dec),
    .regfile_raddr_a_o(regfile_raddr_a),
    .regfile_raddr_b_o(regfile_raddr_b),
    .regfile_waddr_o(regfile_waddr),
    .alu_operator_o(alu_operator_ex_o),
    .alu_op_a_mux_sel_o(alu_op_a_mux_sel_dec),
    .alu_op_b_mux_sel_o(alu_op_b_mux_sel_dec),
    .mult_en_o(mult_en_dec),
    .div_en_o(div_en_dec),
    .multdiv_operator_o(multdiv_operator_ex_o),
    .multdiv_signed_mode_o(multdiv_signed_mode_ex_o),
    .csr_access_o(csr_access_o),
    .csr_op_o(csr_op_o),
    .csr_status_o(csr_status),
    .data_req_o(data_req_dec),
    .data_we_o(data_we_ex_o),
    .data_type_o(data_type_ex_o),
    .data_sign_extension_o(data_sign_ext_ex_o),
    .data_reg_offset_o(data_reg_offset_ex_o),
    .jump_in_dec_o(jump_in_dec),
    .branch_in_dec_o(branch_in_dec)
  );


  ibex_controller
  controller_i
  (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .fetch_enable_i(fetch_enable_i),
    .ctrl_busy_o(ctrl_busy_o),
    .first_fetch_o(core_ctrl_firstfetch_o),
    .illegal_insn_i(illegal_insn_o),
    .ecall_insn_i(ecall_insn_dec),
    .mret_insn_i(mret_insn_dec),
    .dret_insn_i(dret_insn_dec),
    .wfi_insn_i(wfi_insn_dec),
    .ebrk_insn_i(ebrk_insn),
    .csr_status_i(csr_status),
    .instr_valid_i(instr_valid_i),
    .instr_i(instr_rdata_i),
    .instr_compressed_i(instr_rdata_c_i),
    .instr_is_compressed_i(instr_is_compressed_i),
    .instr_valid_clear_o(instr_valid_clear_o),
    .id_in_ready_o(id_in_ready_o),
    .instr_req_o(instr_req_o),
    .pc_set_o(pc_set_o),
    .pc_mux_o(pc_mux_o),
    .exc_pc_mux_o(exc_pc_mux_o),
    .lsu_addr_last_i(lsu_addr_last_i),
    .load_err_i(lsu_load_err_i),
    .store_err_i(lsu_store_err_i),
    .branch_set_i(branch_set_q),
    .jump_set_i(jump_set),
    .irq_i(irq_i),
    .irq_req_ctrl_i(irq_req_ctrl),
    .irq_id_ctrl_i(irq_id_ctrl),
    .m_IE_i(m_irq_enable_i),
    .irq_ack_o(irq_ack_o),
    .irq_id_o(irq_id_o),
    .exc_cause_o(exc_cause_o),
    .exc_ack_o(exc_ack),
    .exc_kill_o(exc_kill),
    .debug_req_i(debug_req_i),
    .debug_cause_o(debug_cause_o),
    .debug_csr_save_o(debug_csr_save_o),
    .debug_single_step_i(debug_single_step_i),
    .debug_ebreakm_i(debug_ebreakm_i),
    .csr_save_if_o(csr_save_if_o),
    .csr_save_id_o(csr_save_id_o),
    .csr_restore_mret_id_o(csr_restore_mret_id_o),
    .csr_restore_dret_id_o(csr_restore_dret_id_o),
    .csr_save_cause_o(csr_save_cause_o),
    .csr_mtval_o(csr_mtval_o),
    .stall_lsu_i(stall_lsu),
    .stall_multdiv_i(stall_multdiv),
    .stall_jump_i(stall_jump),
    .stall_branch_i(stall_branch),
    .perf_jump_o(perf_jump_o),
    .perf_tbranch_o(perf_tbranch_o)
  );


  ibex_int_controller
  int_controller_i
  (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .irq_req_ctrl_o(irq_req_ctrl),
    .irq_id_ctrl_o(irq_id_ctrl),
    .ctrl_ack_i(exc_ack),
    .ctrl_kill_i(exc_kill),
    .irq_i(irq_i),
    .irq_id_i(irq_id_i),
    .m_IE_i(m_irq_enable_i)
  );


  always @(posedge clk_i or posedge N69) begin
    if(N69) begin
      branch_set_q <= 1'b0;
    end else if(1'b1) begin
      branch_set_q <= branch_set_n;
    end 
  end


  always @(posedge clk_i or posedge N69) begin
    if(N69) begin
      instr_multicycle_done_q <= 1'b0;
    end else if(N105) begin
      instr_multicycle_done_q <= instr_multicycle_done_n;
    end 
  end


  always @(posedge clk_i or posedge N69) begin
    if(N69) begin
      id_wb_fsm_cs <= 1'b0;
    end else if(N105) begin
      id_wb_fsm_cs <= id_wb_fsm_ns;
    end 
  end

  assign N106 = ~imm_a_mux_sel;
  assign N52 = N0 & N1 & N2;
  assign N0 = ~imm_b_mux_sel[0];
  assign N1 = ~imm_b_mux_sel[2];
  assign N2 = ~imm_b_mux_sel[1];
  assign N53 = imm_b_mux_sel[0] & N3 & N4;
  assign N3 = ~imm_b_mux_sel[2];
  assign N4 = ~imm_b_mux_sel[1];
  assign N54 = N5 & N6 & imm_b_mux_sel[1];
  assign N5 = ~imm_b_mux_sel[0];
  assign N6 = ~imm_b_mux_sel[2];
  assign N55 = imm_b_mux_sel[0] & imm_b_mux_sel[1];
  assign N56 = N7 & imm_b_mux_sel[2] & N8;
  assign N7 = ~imm_b_mux_sel[0];
  assign N8 = ~imm_b_mux_sel[1];
  assign N57 = imm_b_mux_sel[0] & imm_b_mux_sel[2];
  assign N58 = imm_b_mux_sel[2] & imm_b_mux_sel[1];
  assign N68 = N9 & N10;
  assign N9 = ~regfile_wdata_sel[1];
  assign N10 = ~regfile_wdata_sel[0];
  assign alu_op_a_mux_sel = (N11)? { 1'b0, 1'b1 } : 
                            (N12)? alu_op_a_mux_sel_dec : 1'b0;
  assign N11 = lsu_addr_incr_req_i;
  assign N12 = N43;
  assign alu_op_b_mux_sel = (N11)? 1'b1 : 
                            (N12)? alu_op_b_mux_sel_dec : 1'b0;
  assign imm_b_mux_sel = (N11)? { 1'b1, 1'b1, 1'b0 } : 
                         (N12)? imm_b_mux_sel_dec : 1'b0;
  assign imm_a = (N13)? zimm_rs1_type : 
                 (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = N106;
  assign N14 = imm_a_mux_sel;
  assign alu_operand_a_ex_o = (N15)? multdiv_operand_a_ex_o : 
                              (N16)? lsu_addr_last_i : 
                              (N17)? pc_id_i : 
                              (N18)? imm_a : 1'b0;
  assign N15 = N46;
  assign N16 = N48;
  assign N17 = N50;
  assign N18 = N51;
  assign imm_b = (N19)? imm_i_type : 
                 (N20)? imm_s_type : 
                 (N21)? imm_b_type : 
                 (N22)? imm_u_type : 
                 (N23)? imm_j_type : 
                 (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N59, N60, 1'b0 } : 
                 (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 1'b0;
  assign N19 = N52;
  assign N20 = N53;
  assign N21 = N54;
  assign N22 = N55;
  assign N23 = N56;
  assign N24 = N57;
  assign N25 = N58;
  assign alu_operand_b_ex_o = (N26)? imm_b : 
                              (N27)? data_wdata_ex_o : 1'b0;
  assign N26 = alu_op_b_mux_sel;
  assign N27 = N61;
  assign regfile_we = (N28)? 1'b0 : 
                      (N67)? regfile_we_wb : 
                      (N65)? regfile_we_dec : 1'b0;
  assign N28 = N62;
  assign regfile_wdata = (N29)? regfile_wdata_ex_i : 
                         (N30)? regfile_wdata_lsu_i : 
                         (N31)? csr_rdata_i : 1'b0;
  assign N29 = regfile_wdata_sel[0];
  assign N30 = N68;
  assign N31 = regfile_wdata_sel[1];
  assign data_req_ex_o = (N32)? data_req_dec : 
                         (N33)? 1'b0 : 1'b0;
  assign N32 = instr_executing;
  assign N33 = N107;
  assign mult_en_ex_o = (N32)? mult_en_dec : 
                        (N33)? 1'b0 : 1'b0;
  assign div_en_ex_o = (N32)? div_en_dec : 
                       (N33)? 1'b0 : 1'b0;
  assign N78 = (N34)? 1'b1 : 
               (N35)? 1'b1 : 
               (N36)? branch_decision_i : 
               (N37)? 1'b1 : 
               (N77)? id_wb_fsm_cs : 1'b0;
  assign N34 = data_req_dec;
  assign N35 = multdiv_en_dec;
  assign N36 = branch_in_dec;
  assign N37 = jump_in_dec;
  assign N80 = (N34)? 1'b1 : 
               (N79)? 1'b0 : 
               (N38)? 1'b0 : 
               (N38)? 1'b0 : 
               (N38)? 1'b0 : 1'b0;
  assign N38 = 1'b0;
  assign N81 = (N34)? 1'b0 : 
               (N35)? 1'b0 : 
               (N36)? N70 : 
               (N37)? 1'b0 : 
               (N77)? instr_multicycle_done_q : 1'b0;
  assign N83 = (N34)? 1'b0 : 
               (N35)? 1'b1 : 
               (N82)? 1'b0 : 
               (N38)? 1'b0 : 
               (N38)? 1'b0 : 1'b0;
  assign N85 = (N34)? 1'b0 : 
               (N35)? 1'b0 : 
               (N36)? branch_decision_i : 
               (N84)? 1'b0 : 
               (N38)? 1'b0 : 1'b0;
  assign N86 = (N34)? 1'b0 : 
               (N35)? 1'b0 : 
               (N36)? 1'b1 : 
               (N84)? 1'b0 : 
               (N38)? 1'b0 : 1'b0;
  assign N87 = (N34)? 1'b0 : 
               (N35)? 1'b0 : 
               (N36)? N70 : 
               (N37)? 1'b0 : 
               (N77)? 1'b1 : 1'b0;
  assign N88 = (N34)? 1'b0 : 
               (N35)? 1'b0 : 
               (N36)? 1'b0 : 
               (N37)? 1'b1 : 
               (N77)? 1'b0 : 1'b0;
  assign N89 = (N39)? N88 : 
               (N40)? 1'b0 : 1'b0;
  assign N39 = N73;
  assign N40 = N72;
  assign N90 = (N39)? N80 : 
               (N40)? 1'b0 : 1'b0;
  assign N91 = (N39)? N83 : 
               (N40)? 1'b0 : 1'b0;
  assign N92 = (N39)? N85 : 
               (N40)? 1'b0 : 1'b0;
  assign N93 = (N39)? N86 : 
               (N40)? 1'b0 : 1'b0;
  assign N94 = (N39)? N87 : 
               (N40)? 1'b0 : 1'b0;
  assign N97 = (N41)? 1'b0 : 
               (N96)? id_wb_fsm_cs : 1'b0;
  assign N41 = N95;
  assign N98 = (N41)? 1'b1 : 
               (N96)? instr_multicycle_done_q : 1'b0;
  assign N99 = (N41)? regfile_we_dec : 
               (N96)? 1'b0 : 1'b0;
  assign N100 = (N41)? 1'b0 : 
                (N96)? data_req_dec : 1'b0;
  assign N101 = (N41)? 1'b0 : 
                (N96)? multdiv_en_dec : 1'b0;
  assign N102 = (N41)? 1'b0 : 
                (N96)? branch_in_dec : 1'b0;
  assign N103 = (N41)? 1'b0 : 
                (N96)? jump_in_dec : 1'b0;
  assign instr_ret_o = (N71)? N94 : 
                       (N42)? N95 : 1'b0;
  assign N42 = id_wb_fsm_cs;
  assign stall_jump = (N71)? N89 : 
                      (N42)? N103 : 1'b0;
  assign id_wb_fsm_ns = (N71)? N78 : 
                        (N42)? N97 : 1'b0;
  assign stall_lsu = (N71)? N90 : 
                     (N42)? N100 : 1'b0;
  assign instr_multicycle_done_n = (N71)? N81 : 
                                   (N42)? N98 : 1'b0;
  assign stall_multdiv = (N71)? N91 : 
                         (N42)? N101 : 1'b0;
  assign stall_branch = (N71)? N92 : 
                        (N42)? N102 : 1'b0;
  assign branch_set_n = (N71)? N92 : 
                        (N42)? 1'b0 : 1'b0;
  assign perf_branch_o = (N71)? N93 : 
                         (N42)? 1'b0 : 1'b0;
  assign regfile_we_wb = (N71)? 1'b0 : 
                         (N42)? N99 : 1'b0;
  assign N43 = ~lsu_addr_incr_req_i;
  assign N44 = ~alu_op_a_mux_sel[1];
  assign N45 = ~alu_op_a_mux_sel[0];
  assign N48 = ~N47;
  assign N50 = ~N49;
  assign N59 = ~instr_is_compressed_i;
  assign N60 = instr_is_compressed_i;
  assign N61 = ~alu_op_b_mux_sel;
  assign N62 = illegal_csr_insn_i | N107;
  assign N107 = ~instr_executing;
  assign N63 = data_req_dec | multdiv_en_dec;
  assign N64 = N63 | N62;
  assign N65 = ~N64;
  assign N66 = ~N62;
  assign N67 = N63 & N66;
  assign illegal_insn_o = illegal_insn_dec | illegal_csr_insn_i;
  assign instr_executing = instr_new_i | N108;
  assign N108 = ~instr_multicycle_done_q;
  assign N69 = ~rst_ni;
  assign multdiv_en_dec = mult_en_dec | div_en_dec;
  assign N70 = ~branch_decision_i;
  assign N71 = ~id_wb_fsm_cs;
  assign N72 = ~instr_new_i;
  assign N73 = instr_new_i;
  assign N74 = multdiv_en_dec | data_req_dec;
  assign N75 = branch_in_dec | N74;
  assign N76 = jump_in_dec | N75;
  assign N77 = ~N76;
  assign N79 = ~data_req_dec;
  assign N82 = ~N74;
  assign N84 = ~N75;
  assign N95 = N109 | N111;
  assign N109 = data_req_dec & lsu_valid_i;
  assign N111 = N110 & ex_valid_i;
  assign N110 = ~data_req_dec;
  assign N96 = ~N95;
  assign instr_ret_compressed_o = instr_ret_o & instr_is_compressed_i;
  assign N104 = N72 & N71;
  assign N105 = ~N104;

endmodule



module ibex_alu
(
  operator_i,
  operand_a_i,
  operand_b_i,
  multdiv_operand_a_i,
  multdiv_operand_b_i,
  multdiv_en_i,
  adder_result_o,
  adder_result_ext_o,
  result_o,
  comparison_result_o,
  is_equal_result_o
);

  input [4:0] operator_i;
  input [31:0] operand_a_i;
  input [31:0] operand_b_i;
  input [32:0] multdiv_operand_a_i;
  input [32:0] multdiv_operand_b_i;
  output [31:0] adder_result_o;
  output [33:0] adder_result_ext_o;
  output [31:0] result_o;
  input multdiv_en_i;
  output comparison_result_o;
  output is_equal_result_o;
  wire [31:0] adder_result_o,result_o,shift_op_a,shift_right_result_signed,shift_result;
  wire [33:0] adder_result_ext_o;
  wire comparison_result_o,is_equal_result_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,
  N13,N14,N15,N16,N17,N18,N19,N20,N21,cmp_signed,N22,is_greater_equal,N23,N24,N25,
  N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,
  N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,
  N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,
  N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,
  N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,
  N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,
  N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,
  N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,
  N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,
  N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,
  N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,
  N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,
  N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,
  N248,N249,N250,N251,N252,SV2V_UNCONNECTED_1;
  wire [32:0] adder_in_a,operand_b_neg,adder_in_b;
  wire [32:32] shift_op_a_32;
  assign adder_result_o[31] = adder_result_ext_o[32];
  assign adder_result_o[30] = adder_result_ext_o[31];
  assign adder_result_o[29] = adder_result_ext_o[30];
  assign adder_result_o[28] = adder_result_ext_o[29];
  assign adder_result_o[27] = adder_result_ext_o[28];
  assign adder_result_o[26] = adder_result_ext_o[27];
  assign adder_result_o[25] = adder_result_ext_o[26];
  assign adder_result_o[24] = adder_result_ext_o[25];
  assign adder_result_o[23] = adder_result_ext_o[24];
  assign adder_result_o[22] = adder_result_ext_o[23];
  assign adder_result_o[21] = adder_result_ext_o[22];
  assign adder_result_o[20] = adder_result_ext_o[21];
  assign adder_result_o[19] = adder_result_ext_o[20];
  assign adder_result_o[18] = adder_result_ext_o[19];
  assign adder_result_o[17] = adder_result_ext_o[18];
  assign adder_result_o[16] = adder_result_ext_o[17];
  assign adder_result_o[15] = adder_result_ext_o[16];
  assign adder_result_o[14] = adder_result_ext_o[15];
  assign adder_result_o[13] = adder_result_ext_o[14];
  assign adder_result_o[12] = adder_result_ext_o[13];
  assign adder_result_o[11] = adder_result_ext_o[12];
  assign adder_result_o[10] = adder_result_ext_o[11];
  assign adder_result_o[9] = adder_result_ext_o[10];
  assign adder_result_o[8] = adder_result_ext_o[9];
  assign adder_result_o[7] = adder_result_ext_o[8];
  assign adder_result_o[6] = adder_result_ext_o[7];
  assign adder_result_o[5] = adder_result_ext_o[6];
  assign adder_result_o[4] = adder_result_ext_o[5];
  assign adder_result_o[3] = adder_result_ext_o[4];
  assign adder_result_o[2] = adder_result_ext_o[3];
  assign adder_result_o[1] = adder_result_ext_o[2];
  assign adder_result_o[0] = adder_result_ext_o[1];
  assign { SV2V_UNCONNECTED_1, shift_right_result_signed } = $signed({ shift_op_a_32[32:32], shift_op_a }) >>> operand_b_i[4:0];
  assign is_equal_result_o = adder_result_ext_o[32:1] == 1'b0;
  assign N30 = N33 & operator_i[2];
  assign N31 = N30 & operator_i[1];
  assign N34 = N32 & N33;
  assign N38 = operator_i[4] | operator_i[3];
  assign N39 = N186 | operator_i[1];
  assign N40 = N38 | N39;
  assign N41 = N40 | operator_i[0];
  assign N43 = operator_i[2] | N194;
  assign N44 = N38 | N43;
  assign N45 = N44 | N187;
  assign N47 = N44 | operator_i[0];
  assign N49 = N186 & N194;
  assign N50 = N34 & N49;
  assign N51 = N50 & N187;
  assign N52 = operator_i[2] | operator_i[1];
  assign N53 = N38 | N52;
  assign N54 = N53 | N187;
  assign N56 = N186 | N194;
  assign N57 = N38 | N56;
  assign N58 = N57 | N187;
  assign N59 = N57 | operator_i[0];
  assign N60 = N40 | N187;
  assign N62 = N32 | operator_i[3];
  assign N63 = N62 | N52;
  assign N64 = N63 | operator_i[0];
  assign N65 = N63 | N187;
  assign N66 = operator_i[4] | N33;
  assign N67 = N66 | N39;
  assign N68 = N67 | N187;
  assign N69 = N66 | N56;
  assign N70 = N69 | N187;
  assign N71 = N66 | N52;
  assign N72 = N71 | N187;
  assign N73 = N66 | N43;
  assign N74 = N73 | N187;
  assign N75 = N67 | operator_i[0];
  assign N76 = N69 | operator_i[0];
  assign N77 = N71 | operator_i[0];
  assign N78 = N73 | operator_i[0];
  assign N79 = N62 | N43;
  assign N80 = N79 | operator_i[0];
  assign N81 = N79 | N187;
  assign N82 = N62 | N39;
  assign N83 = N82 | operator_i[0];
  assign N84 = N82 | N187;
  assign N86 = operator_i[4] & operator_i[2];
  assign N87 = N86 & operator_i[1];
  assign N88 = operator_i[4] & operator_i[3];
  assign N186 = ~operator_i[2];
  assign N187 = ~operator_i[0];
  assign N188 = operator_i[3] | operator_i[4];
  assign N189 = N186 | N188;
  assign N190 = operator_i[1] | N189;
  assign N191 = N187 | N190;
  assign N192 = ~N191;
  assign N193 = ~adder_result_ext_o[32];
  assign N194 = ~operator_i[1];
  assign N195 = N194 | N189;
  assign N196 = N187 | N195;
  assign N197 = ~N196;
  assign N198 = ~N154;
  assign adder_result_ext_o = adder_in_a + adder_in_b;
  assign adder_in_a = (N0)? multdiv_operand_a_i : 
                      (N1)? { operand_a_i, 1'b1 } : 1'b0;
  assign N0 = multdiv_en_i;
  assign N1 = N21;
  assign adder_in_b = (N0)? multdiv_operand_b_i : 
                      (N1)? operand_b_neg : 1'b0;
  assign shift_op_a = (N2)? { operand_a_i[0:0], operand_a_i[1:1], operand_a_i[2:2], operand_a_i[3:3], operand_a_i[4:4], operand_a_i[5:5], operand_a_i[6:6], operand_a_i[7:7], operand_a_i[8:8], operand_a_i[9:9], operand_a_i[10:10], operand_a_i[11:11], operand_a_i[12:12], operand_a_i[13:13], operand_a_i[14:14], operand_a_i[15:15], operand_a_i[16:16], operand_a_i[17:17], operand_a_i[18:18], operand_a_i[19:19], operand_a_i[20:20], operand_a_i[21:21], operand_a_i[22:22], operand_a_i[23:23], operand_a_i[24:24], operand_a_i[25:25], operand_a_i[26:26], operand_a_i[27:27], operand_a_i[28:28], operand_a_i[29:29], operand_a_i[30:30], operand_a_i[31:31] } : 
                      (N3)? operand_a_i : 1'b0;
  assign N2 = N197;
  assign N3 = N196;
  assign shift_result = (N2)? { shift_right_result_signed[0:0], shift_right_result_signed[1:1], shift_right_result_signed[2:2], shift_right_result_signed[3:3], shift_right_result_signed[4:4], shift_right_result_signed[5:5], shift_right_result_signed[6:6], shift_right_result_signed[7:7], shift_right_result_signed[8:8], shift_right_result_signed[9:9], shift_right_result_signed[10:10], shift_right_result_signed[11:11], shift_right_result_signed[12:12], shift_right_result_signed[13:13], shift_right_result_signed[14:14], shift_right_result_signed[15:15], shift_right_result_signed[16:16], shift_right_result_signed[17:17], shift_right_result_signed[18:18], shift_right_result_signed[19:19], shift_right_result_signed[20:20], shift_right_result_signed[21:21], shift_right_result_signed[22:22], shift_right_result_signed[23:23], shift_right_result_signed[24:24], shift_right_result_signed[25:25], shift_right_result_signed[26:26], shift_right_result_signed[27:27], shift_right_result_signed[28:28], shift_right_result_signed[29:29], shift_right_result_signed[30:30], shift_right_result_signed[31:31] } : 
                        (N3)? shift_right_result_signed : 1'b0;
  assign is_greater_equal = (N4)? N193 : 
                            (N5)? N23 : 1'b0;
  assign N4 = N198;
  assign N5 = N154;
  assign comparison_result_o = (N6)? is_equal_result_o : 
                               (N7)? N24 : 
                               (N8)? N36 : 
                               (N9)? is_greater_equal : 
                               (N10)? N25 : 
                               (N11)? N37 : 
                               (N12)? is_equal_result_o : 1'b0;
  assign N6 = N200;
  assign N7 = N202;
  assign N8 = N26;
  assign N9 = N27;
  assign N10 = N28;
  assign N11 = N29;
  assign N12 = N35;
  assign result_o = (N13)? { N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121 } : 
                    (N14)? { N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153 } : 
                    (N15)? { N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185 } : 
                    (N16)? adder_result_ext_o[32:1] : 
                    (N17)? shift_result : 
                    (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, comparison_result_o } : 
                    (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = N42;
  assign N14 = N46;
  assign N15 = N48;
  assign N16 = N55;
  assign N17 = N61;
  assign N18 = N85;
  assign N19 = N89;
  assign N20 = N225 | N226;
  assign N225 = N223 | N224;
  assign N223 = N221 | N222;
  assign N221 = N219 | N220;
  assign N219 = N217 | N218;
  assign N217 = N215 | N216;
  assign N215 = N213 | N214;
  assign N213 = N211 | N212;
  assign N211 = N209 | N210;
  assign N209 = N207 | N208;
  assign N207 = N205 | N206;
  assign N205 = N203 | N204;
  assign N203 = N201 | N202;
  assign N201 = N199 | N200;
  assign N199 = ~N54;
  assign N200 = ~N64;
  assign N202 = ~N65;
  assign N204 = ~N68;
  assign N206 = ~N70;
  assign N208 = ~N72;
  assign N210 = ~N74;
  assign N212 = ~N75;
  assign N214 = ~N76;
  assign N216 = ~N77;
  assign N218 = ~N78;
  assign N220 = ~N80;
  assign N222 = ~N81;
  assign N224 = ~N83;
  assign N226 = ~N84;
  assign operand_b_neg[0] = N20;
  assign N21 = ~multdiv_en_i;
  assign operand_b_neg[32] = operand_b_i[31] ^ operand_b_neg[0];
  assign operand_b_neg[31] = operand_b_i[30] ^ operand_b_neg[0];
  assign operand_b_neg[30] = operand_b_i[29] ^ operand_b_neg[0];
  assign operand_b_neg[29] = operand_b_i[28] ^ operand_b_neg[0];
  assign operand_b_neg[28] = operand_b_i[27] ^ operand_b_neg[0];
  assign operand_b_neg[27] = operand_b_i[26] ^ operand_b_neg[0];
  assign operand_b_neg[26] = operand_b_i[25] ^ operand_b_neg[0];
  assign operand_b_neg[25] = operand_b_i[24] ^ operand_b_neg[0];
  assign operand_b_neg[24] = operand_b_i[23] ^ operand_b_neg[0];
  assign operand_b_neg[23] = operand_b_i[22] ^ operand_b_neg[0];
  assign operand_b_neg[22] = operand_b_i[21] ^ operand_b_neg[0];
  assign operand_b_neg[21] = operand_b_i[20] ^ operand_b_neg[0];
  assign operand_b_neg[20] = operand_b_i[19] ^ operand_b_neg[0];
  assign operand_b_neg[19] = operand_b_i[18] ^ operand_b_neg[0];
  assign operand_b_neg[18] = operand_b_i[17] ^ operand_b_neg[0];
  assign operand_b_neg[17] = operand_b_i[16] ^ operand_b_neg[0];
  assign operand_b_neg[16] = operand_b_i[15] ^ operand_b_neg[0];
  assign operand_b_neg[15] = operand_b_i[14] ^ operand_b_neg[0];
  assign operand_b_neg[14] = operand_b_i[13] ^ operand_b_neg[0];
  assign operand_b_neg[13] = operand_b_i[12] ^ operand_b_neg[0];
  assign operand_b_neg[12] = operand_b_i[11] ^ operand_b_neg[0];
  assign operand_b_neg[11] = operand_b_i[10] ^ operand_b_neg[0];
  assign operand_b_neg[10] = operand_b_i[9] ^ operand_b_neg[0];
  assign operand_b_neg[9] = operand_b_i[8] ^ operand_b_neg[0];
  assign operand_b_neg[8] = operand_b_i[7] ^ operand_b_neg[0];
  assign operand_b_neg[7] = operand_b_i[6] ^ operand_b_neg[0];
  assign operand_b_neg[6] = operand_b_i[5] ^ operand_b_neg[0];
  assign operand_b_neg[5] = operand_b_i[4] ^ operand_b_neg[0];
  assign operand_b_neg[4] = operand_b_i[3] ^ operand_b_neg[0];
  assign operand_b_neg[3] = operand_b_i[2] ^ operand_b_neg[0];
  assign operand_b_neg[2] = operand_b_i[1] ^ operand_b_neg[0];
  assign operand_b_neg[1] = operand_b_i[0] ^ operand_b_neg[0];
  assign shift_op_a_32[32] = N192 & shift_op_a[31];
  assign N22 = N230 | N224;
  assign N230 = N229 | N220;
  assign N229 = N228 | N218;
  assign N228 = N227 | N216;
  assign N227 = N212 | N214;
  assign cmp_signed = N22;
  assign N23 = operand_a_i[31] ^ cmp_signed;
  assign N24 = ~is_equal_result_o;
  assign N25 = ~is_greater_equal;
  assign N26 = N212 | N204;
  assign N27 = N214 | N206;
  assign N28 = N232 | N222;
  assign N232 = N231 | N208;
  assign N231 = N216 | N220;
  assign N29 = N234 | N210;
  assign N234 = N233 | N218;
  assign N233 = N224 | N226;
  assign N32 = ~operator_i[4];
  assign N33 = ~operator_i[3];
  assign N35 = N87 | N236;
  assign N236 = N31 | N235;
  assign N235 = N88 | N34;
  assign N36 = is_greater_equal & N24;
  assign N37 = N25 | is_equal_result_o;
  assign N42 = ~N41;
  assign N46 = ~N45;
  assign N48 = ~N47;
  assign N55 = N51 | N199;
  assign N61 = N239 | N240;
  assign N239 = N237 | N238;
  assign N237 = ~N58;
  assign N238 = ~N59;
  assign N240 = ~N60;
  assign N85 = N252 | N226;
  assign N252 = N251 | N224;
  assign N251 = N250 | N222;
  assign N250 = N249 | N220;
  assign N249 = N248 | N218;
  assign N248 = N247 | N216;
  assign N247 = N246 | N214;
  assign N246 = N245 | N212;
  assign N245 = N244 | N210;
  assign N244 = N243 | N208;
  assign N243 = N242 | N206;
  assign N242 = N241 | N204;
  assign N241 = N200 | N202;
  assign N89 = N87 | N88;
  assign N90 = operand_a_i[31] & operand_b_i[31];
  assign N91 = operand_a_i[30] & operand_b_i[30];
  assign N92 = operand_a_i[29] & operand_b_i[29];
  assign N93 = operand_a_i[28] & operand_b_i[28];
  assign N94 = operand_a_i[27] & operand_b_i[27];
  assign N95 = operand_a_i[26] & operand_b_i[26];
  assign N96 = operand_a_i[25] & operand_b_i[25];
  assign N97 = operand_a_i[24] & operand_b_i[24];
  assign N98 = operand_a_i[23] & operand_b_i[23];
  assign N99 = operand_a_i[22] & operand_b_i[22];
  assign N100 = operand_a_i[21] & operand_b_i[21];
  assign N101 = operand_a_i[20] & operand_b_i[20];
  assign N102 = operand_a_i[19] & operand_b_i[19];
  assign N103 = operand_a_i[18] & operand_b_i[18];
  assign N104 = operand_a_i[17] & operand_b_i[17];
  assign N105 = operand_a_i[16] & operand_b_i[16];
  assign N106 = operand_a_i[15] & operand_b_i[15];
  assign N107 = operand_a_i[14] & operand_b_i[14];
  assign N108 = operand_a_i[13] & operand_b_i[13];
  assign N109 = operand_a_i[12] & operand_b_i[12];
  assign N110 = operand_a_i[11] & operand_b_i[11];
  assign N111 = operand_a_i[10] & operand_b_i[10];
  assign N112 = operand_a_i[9] & operand_b_i[9];
  assign N113 = operand_a_i[8] & operand_b_i[8];
  assign N114 = operand_a_i[7] & operand_b_i[7];
  assign N115 = operand_a_i[6] & operand_b_i[6];
  assign N116 = operand_a_i[5] & operand_b_i[5];
  assign N117 = operand_a_i[4] & operand_b_i[4];
  assign N118 = operand_a_i[3] & operand_b_i[3];
  assign N119 = operand_a_i[2] & operand_b_i[2];
  assign N120 = operand_a_i[1] & operand_b_i[1];
  assign N121 = operand_a_i[0] & operand_b_i[0];
  assign N122 = operand_a_i[31] | operand_b_i[31];
  assign N123 = operand_a_i[30] | operand_b_i[30];
  assign N124 = operand_a_i[29] | operand_b_i[29];
  assign N125 = operand_a_i[28] | operand_b_i[28];
  assign N126 = operand_a_i[27] | operand_b_i[27];
  assign N127 = operand_a_i[26] | operand_b_i[26];
  assign N128 = operand_a_i[25] | operand_b_i[25];
  assign N129 = operand_a_i[24] | operand_b_i[24];
  assign N130 = operand_a_i[23] | operand_b_i[23];
  assign N131 = operand_a_i[22] | operand_b_i[22];
  assign N132 = operand_a_i[21] | operand_b_i[21];
  assign N133 = operand_a_i[20] | operand_b_i[20];
  assign N134 = operand_a_i[19] | operand_b_i[19];
  assign N135 = operand_a_i[18] | operand_b_i[18];
  assign N136 = operand_a_i[17] | operand_b_i[17];
  assign N137 = operand_a_i[16] | operand_b_i[16];
  assign N138 = operand_a_i[15] | operand_b_i[15];
  assign N139 = operand_a_i[14] | operand_b_i[14];
  assign N140 = operand_a_i[13] | operand_b_i[13];
  assign N141 = operand_a_i[12] | operand_b_i[12];
  assign N142 = operand_a_i[11] | operand_b_i[11];
  assign N143 = operand_a_i[10] | operand_b_i[10];
  assign N144 = operand_a_i[9] | operand_b_i[9];
  assign N145 = operand_a_i[8] | operand_b_i[8];
  assign N146 = operand_a_i[7] | operand_b_i[7];
  assign N147 = operand_a_i[6] | operand_b_i[6];
  assign N148 = operand_a_i[5] | operand_b_i[5];
  assign N149 = operand_a_i[4] | operand_b_i[4];
  assign N150 = operand_a_i[3] | operand_b_i[3];
  assign N151 = operand_a_i[2] | operand_b_i[2];
  assign N152 = operand_a_i[1] | operand_b_i[1];
  assign N153 = operand_a_i[0] | operand_b_i[0];
  assign N154 = operand_a_i[31] ^ operand_b_i[31];
  assign N155 = operand_a_i[30] ^ operand_b_i[30];
  assign N156 = operand_a_i[29] ^ operand_b_i[29];
  assign N157 = operand_a_i[28] ^ operand_b_i[28];
  assign N158 = operand_a_i[27] ^ operand_b_i[27];
  assign N159 = operand_a_i[26] ^ operand_b_i[26];
  assign N160 = operand_a_i[25] ^ operand_b_i[25];
  assign N161 = operand_a_i[24] ^ operand_b_i[24];
  assign N162 = operand_a_i[23] ^ operand_b_i[23];
  assign N163 = operand_a_i[22] ^ operand_b_i[22];
  assign N164 = operand_a_i[21] ^ operand_b_i[21];
  assign N165 = operand_a_i[20] ^ operand_b_i[20];
  assign N166 = operand_a_i[19] ^ operand_b_i[19];
  assign N167 = operand_a_i[18] ^ operand_b_i[18];
  assign N168 = operand_a_i[17] ^ operand_b_i[17];
  assign N169 = operand_a_i[16] ^ operand_b_i[16];
  assign N170 = operand_a_i[15] ^ operand_b_i[15];
  assign N171 = operand_a_i[14] ^ operand_b_i[14];
  assign N172 = operand_a_i[13] ^ operand_b_i[13];
  assign N173 = operand_a_i[12] ^ operand_b_i[12];
  assign N174 = operand_a_i[11] ^ operand_b_i[11];
  assign N175 = operand_a_i[10] ^ operand_b_i[10];
  assign N176 = operand_a_i[9] ^ operand_b_i[9];
  assign N177 = operand_a_i[8] ^ operand_b_i[8];
  assign N178 = operand_a_i[7] ^ operand_b_i[7];
  assign N179 = operand_a_i[6] ^ operand_b_i[6];
  assign N180 = operand_a_i[5] ^ operand_b_i[5];
  assign N181 = operand_a_i[4] ^ operand_b_i[4];
  assign N182 = operand_a_i[3] ^ operand_b_i[3];
  assign N183 = operand_a_i[2] ^ operand_b_i[2];
  assign N184 = operand_a_i[1] ^ operand_b_i[1];
  assign N185 = operand_a_i[0] ^ operand_b_i[0];

endmodule



module ibex_multdiv_fast
(
  clk_i,
  rst_ni,
  mult_en_i,
  div_en_i,
  operator_i,
  signed_mode_i,
  op_a_i,
  op_b_i,
  alu_adder_ext_i,
  alu_adder_i,
  equal_to_zero,
  alu_operand_a_o,
  alu_operand_b_o,
  multdiv_result_o,
  valid_o
);

  input [1:0] operator_i;
  input [1:0] signed_mode_i;
  input [31:0] op_a_i;
  input [31:0] op_b_i;
  input [33:0] alu_adder_ext_i;
  input [31:0] alu_adder_i;
  output [32:0] alu_operand_a_o;
  output [32:0] alu_operand_b_o;
  output [31:0] multdiv_result_o;
  input clk_i;
  input rst_ni;
  input mult_en_i;
  input div_en_i;
  input equal_to_zero;
  output valid_o;
  wire [32:0] alu_operand_a_o,alu_operand_b_o;
  wire [31:0] multdiv_result_o,op_quotient_n,next_remainder,one_shift,next_quotient;
  wire valid_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
  sign_a,sign_b,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,
  N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,
  is_greater_equal,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,
  N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,
  N126,div_sign_a,div_sign_b,div_change_sign,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,div_valid,
  N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,
  N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,
  N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,
  N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
  N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,
  N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,
  N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,
  N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,
  N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,
  N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,
  N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,
  N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,
  N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,
  N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,
  N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,
  N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,
  N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,
  N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,
  N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,
  N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,
  N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,
  N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,
  N548,N549,N550,N551,N552,N553,mult_valid,N554,N555,N556,N557,N558,N559,N560,N561,
  N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,
  N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
  N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,
  N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,
  N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,
  N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,
  N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,
  N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,
  N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,
  N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,
  N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732;
  wire [1:0] mult_state_n;
  wire [4:0] div_counter_n;
  wire [2:0] md_state_n;
  wire [33:0] mac_res_n,op_remainder_n,accum,mac_res_signed;
  wire [15:0] mult_op_a,mult_op_b;
  reg [31:0] op_numerator_q,op_quotient_q,op_denominator_q;
  reg [1:0] mult_state_q;
  reg [33:0] mac_res_q;
  reg [4:0] div_counter_q;
  reg [2:0] md_state_q;
  assign alu_operand_b_o[0] = 1'b1;
  assign alu_operand_a_o[0] = 1'b1;

  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[31] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[31] <= N286;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[30] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[30] <= N285;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[29] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[29] <= N284;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[28] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[28] <= N283;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[27] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[27] <= N282;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[26] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[26] <= N281;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[25] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[25] <= N280;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[24] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[24] <= N279;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[23] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[23] <= N278;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[22] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[22] <= N277;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[21] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[21] <= N276;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[20] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[20] <= N275;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[19] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[19] <= N274;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[18] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[18] <= N273;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[17] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[17] <= N272;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[16] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[16] <= N271;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[15] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[15] <= N270;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[14] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[14] <= N269;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[13] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[13] <= N268;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[12] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[12] <= N267;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[11] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[11] <= N266;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[10] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[10] <= N265;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[9] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[9] <= N264;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[8] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[8] <= N263;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[7] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[7] <= N262;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[6] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[6] <= N261;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[5] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[5] <= N260;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[4] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[4] <= N259;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[3] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[3] <= N258;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[2] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[2] <= N257;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[1] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[1] <= N256;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_numerator_q[0] <= 1'b0;
    end else if(N696) begin
      op_numerator_q[0] <= N255;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[31] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[31] <= op_quotient_n[31];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[30] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[30] <= op_quotient_n[30];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[29] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[29] <= op_quotient_n[29];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[28] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[28] <= op_quotient_n[28];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[27] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[27] <= op_quotient_n[27];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[26] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[26] <= op_quotient_n[26];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[25] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[25] <= op_quotient_n[25];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[24] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[24] <= op_quotient_n[24];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[23] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[23] <= op_quotient_n[23];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[22] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[22] <= op_quotient_n[22];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[21] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[21] <= op_quotient_n[21];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[20] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[20] <= op_quotient_n[20];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[19] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[19] <= op_quotient_n[19];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[18] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[18] <= op_quotient_n[18];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[17] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[17] <= op_quotient_n[17];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[16] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[16] <= op_quotient_n[16];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[15] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[15] <= op_quotient_n[15];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[14] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[14] <= op_quotient_n[14];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[13] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[13] <= op_quotient_n[13];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[12] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[12] <= op_quotient_n[12];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[11] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[11] <= op_quotient_n[11];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[10] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[10] <= op_quotient_n[10];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[9] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[9] <= op_quotient_n[9];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[8] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[8] <= op_quotient_n[8];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[7] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[7] <= op_quotient_n[7];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[6] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[6] <= op_quotient_n[6];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[5] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[5] <= op_quotient_n[5];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[4] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[4] <= op_quotient_n[4];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[3] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[3] <= op_quotient_n[3];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[2] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[2] <= op_quotient_n[2];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[1] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[1] <= op_quotient_n[1];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_quotient_q[0] <= 1'b0;
    end else if(N702) begin
      op_quotient_q[0] <= op_quotient_n[0];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mult_state_q[1] <= 1'b0;
    end else if(mult_en_i) begin
      mult_state_q[1] <= mult_state_n[1];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mult_state_q[0] <= 1'b0;
    end else if(mult_en_i) begin
      mult_state_q[0] <= mult_state_n[0];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[33] <= 1'b0;
    end else if(N709) begin
      mac_res_q[33] <= N57;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[32] <= 1'b0;
    end else if(N709) begin
      mac_res_q[32] <= N56;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[31] <= 1'b0;
    end else if(N709) begin
      mac_res_q[31] <= N55;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[30] <= 1'b0;
    end else if(N709) begin
      mac_res_q[30] <= N54;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[29] <= 1'b0;
    end else if(N709) begin
      mac_res_q[29] <= N53;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[28] <= 1'b0;
    end else if(N709) begin
      mac_res_q[28] <= N52;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[27] <= 1'b0;
    end else if(N709) begin
      mac_res_q[27] <= N51;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[26] <= 1'b0;
    end else if(N709) begin
      mac_res_q[26] <= N50;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[25] <= 1'b0;
    end else if(N709) begin
      mac_res_q[25] <= N49;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[24] <= 1'b0;
    end else if(N709) begin
      mac_res_q[24] <= N48;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[23] <= 1'b0;
    end else if(N709) begin
      mac_res_q[23] <= N47;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[22] <= 1'b0;
    end else if(N709) begin
      mac_res_q[22] <= N46;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[21] <= 1'b0;
    end else if(N709) begin
      mac_res_q[21] <= N45;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[20] <= 1'b0;
    end else if(N709) begin
      mac_res_q[20] <= N44;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[19] <= 1'b0;
    end else if(N709) begin
      mac_res_q[19] <= N43;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[18] <= 1'b0;
    end else if(N709) begin
      mac_res_q[18] <= N42;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[17] <= 1'b0;
    end else if(N709) begin
      mac_res_q[17] <= N41;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[16] <= 1'b0;
    end else if(N709) begin
      mac_res_q[16] <= N40;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[15] <= 1'b0;
    end else if(N709) begin
      mac_res_q[15] <= N39;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[14] <= 1'b0;
    end else if(N709) begin
      mac_res_q[14] <= N38;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[13] <= 1'b0;
    end else if(N709) begin
      mac_res_q[13] <= N37;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[12] <= 1'b0;
    end else if(N709) begin
      mac_res_q[12] <= N36;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[11] <= 1'b0;
    end else if(N709) begin
      mac_res_q[11] <= N35;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[10] <= 1'b0;
    end else if(N709) begin
      mac_res_q[10] <= N34;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[9] <= 1'b0;
    end else if(N709) begin
      mac_res_q[9] <= N33;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[8] <= 1'b0;
    end else if(N709) begin
      mac_res_q[8] <= N32;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[7] <= 1'b0;
    end else if(N709) begin
      mac_res_q[7] <= N31;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[6] <= 1'b0;
    end else if(N709) begin
      mac_res_q[6] <= N30;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[5] <= 1'b0;
    end else if(N709) begin
      mac_res_q[5] <= N29;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[4] <= 1'b0;
    end else if(N709) begin
      mac_res_q[4] <= N28;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[3] <= 1'b0;
    end else if(N709) begin
      mac_res_q[3] <= N27;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[2] <= 1'b0;
    end else if(N709) begin
      mac_res_q[2] <= N26;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[1] <= 1'b0;
    end else if(N709) begin
      mac_res_q[1] <= N25;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      mac_res_q[0] <= 1'b0;
    end else if(N709) begin
      mac_res_q[0] <= N24;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      div_counter_q[4] <= 1'b0;
    end else if(div_en_i) begin
      div_counter_q[4] <= div_counter_n[4];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      div_counter_q[3] <= 1'b0;
    end else if(div_en_i) begin
      div_counter_q[3] <= div_counter_n[3];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      div_counter_q[2] <= 1'b0;
    end else if(div_en_i) begin
      div_counter_q[2] <= div_counter_n[2];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      div_counter_q[1] <= 1'b0;
    end else if(div_en_i) begin
      div_counter_q[1] <= div_counter_n[1];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      div_counter_q[0] <= 1'b0;
    end else if(div_en_i) begin
      div_counter_q[0] <= div_counter_n[0];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      md_state_q[2] <= 1'b0;
    end else if(div_en_i) begin
      md_state_q[2] <= md_state_n[2];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      md_state_q[1] <= 1'b0;
    end else if(div_en_i) begin
      md_state_q[1] <= md_state_n[1];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      md_state_q[0] <= 1'b0;
    end else if(div_en_i) begin
      md_state_q[0] <= md_state_n[0];
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[31] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[31] <= N351;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[30] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[30] <= N350;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[29] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[29] <= N349;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[28] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[28] <= N348;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[27] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[27] <= N347;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[26] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[26] <= N346;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[25] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[25] <= N345;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[24] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[24] <= N344;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[23] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[23] <= N343;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[22] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[22] <= N342;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[21] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[21] <= N341;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[20] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[20] <= N340;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[19] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[19] <= N339;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[18] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[18] <= N338;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[17] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[17] <= N337;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[16] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[16] <= N336;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[15] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[15] <= N335;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[14] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[14] <= N334;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[13] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[13] <= N333;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[12] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[12] <= N332;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[11] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[11] <= N331;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[10] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[10] <= N330;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[9] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[9] <= N329;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[8] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[8] <= N328;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[7] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[7] <= N327;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[6] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[6] <= N326;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[5] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[5] <= N325;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[4] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[4] <= N324;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[3] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[3] <= N323;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[2] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[2] <= N322;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[1] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[1] <= N321;
    end 
  end


  always @(posedge clk_i or posedge N21) begin
    if(N21) begin
      op_denominator_q[0] <= 1'b0;
    end else if(N718) begin
      op_denominator_q[0] <= N320;
    end 
  end

  assign one_shift = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << div_counter_q;
  assign N199 = N196 & N197;
  assign N200 = N199 & N198;
  assign N201 = md_state_q[2] | md_state_q[1];
  assign N202 = N201 | N198;
  assign N204 = md_state_q[2] | N197;
  assign N205 = N204 | md_state_q[0];
  assign N207 = md_state_q[2] | N197;
  assign N208 = N207 | N198;
  assign N210 = N196 | md_state_q[1];
  assign N211 = N210 | md_state_q[0];
  assign N213 = N196 | md_state_q[1];
  assign N214 = N213 | N198;
  assign N216 = N196 | N197;
  assign N217 = N216 | md_state_q[0];
  assign N219 = md_state_q[2] & md_state_q[1];
  assign N220 = N219 & md_state_q[0];
  assign N417 = (N385)? op_numerator_q[0] : 
                (N387)? op_numerator_q[1] : 
                (N389)? op_numerator_q[2] : 
                (N391)? op_numerator_q[3] : 
                (N393)? op_numerator_q[4] : 
                (N395)? op_numerator_q[5] : 
                (N397)? op_numerator_q[6] : 
                (N399)? op_numerator_q[7] : 
                (N401)? op_numerator_q[8] : 
                (N403)? op_numerator_q[9] : 
                (N405)? op_numerator_q[10] : 
                (N407)? op_numerator_q[11] : 
                (N409)? op_numerator_q[12] : 
                (N411)? op_numerator_q[13] : 
                (N413)? op_numerator_q[14] : 
                (N415)? op_numerator_q[15] : 
                (N386)? op_numerator_q[16] : 
                (N388)? op_numerator_q[17] : 
                (N390)? op_numerator_q[18] : 
                (N392)? op_numerator_q[19] : 
                (N394)? op_numerator_q[20] : 
                (N396)? op_numerator_q[21] : 
                (N398)? op_numerator_q[22] : 
                (N400)? op_numerator_q[23] : 
                (N402)? op_numerator_q[24] : 
                (N404)? op_numerator_q[25] : 
                (N406)? op_numerator_q[26] : 
                (N408)? op_numerator_q[27] : 
                (N410)? op_numerator_q[28] : 
                (N412)? op_numerator_q[29] : 
                (N414)? op_numerator_q[30] : 
                (N416)? op_numerator_q[31] : 1'b0;
  assign N558 = N556 & N557;
  assign N559 = mult_state_q[1] | N557;
  assign N561 = N556 | mult_state_q[0];
  assign N563 = mult_state_q[1] & mult_state_q[0];
  assign N719 = operator_i[0] | operator_i[1];
  assign N720 = ~N719;
  assign N721 = ~operator_i[1];
  assign N722 = operator_i[0] | N721;
  assign N723 = ~N722;
  assign N724 = ~div_counter_q[0];
  assign N725 = div_counter_q[3] | div_counter_q[4];
  assign N726 = div_counter_q[2] | N725;
  assign N727 = div_counter_q[1] | N726;
  assign N728 = N724 | N727;
  assign N729 = ~N728;
  assign N730 = signed_mode_i[0] | signed_mode_i[1];
  assign N731 = ~alu_adder_ext_i[32];
  assign N732 = ~N126;
  assign { N195, N194, N193, N192, N191 } = div_counter_q - 1'b1;
  assign { N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59 } = $signed({ sign_a, mult_op_a }) * $signed({ sign_b, mult_op_b });
  assign mac_res_signed = $signed({ N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59 }) + $signed(accum);
  assign { N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24 } = (N0)? mac_res_n : 
                                                                                                                                                                                        (N1)? op_remainder_n : 1'b0;
  assign N0 = mult_en_i;
  assign N1 = div_en_i;
  assign multdiv_result_o = (N1)? mac_res_q[31:0] : 
                            (N2)? mac_res_n[31:0] : 1'b0;
  assign N2 = N58;
  assign next_remainder = (N3)? alu_adder_ext_i[32:1] : 
                          (N4)? mac_res_q[31:0] : 1'b0;
  assign N3 = is_greater_equal;
  assign N4 = N93;
  assign next_quotient = (N3)? { N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125 } : 
                         (N4)? op_quotient_q : 1'b0;
  assign is_greater_equal = (N5)? N731 : 
                            (N6)? mac_res_q[31] : 1'b0;
  assign N5 = N732;
  assign N6 = N126;
  assign { N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222 } = (N7)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N8)? op_a_i : 1'b0;
  assign N7 = N723;
  assign N8 = N722;
  assign { N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255 } = (N9)? alu_adder_i : 
                                                                                                                                                                                                              (N10)? op_a_i : 1'b0;
  assign N9 = div_sign_a;
  assign N10 = N254;
  assign { N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320 } = (N11)? alu_adder_i : 
                                                                                                                                                                                                              (N12)? op_b_i : 1'b0;
  assign N11 = div_sign_b;
  assign N12 = N319;
  assign { N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418 } = (N7)? next_quotient : 
                                                                                                                                                                                                              (N8)? next_remainder : 1'b0;
  assign { N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453 } = (N13)? { 1'b0, 1'b0, alu_adder_i } : 
                                                                                                                                                                                                                          (N14)? mac_res_q : 1'b0;
  assign N13 = div_change_sign;
  assign N14 = N452;
  assign { N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487 } = (N7)? { N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453 } : 
                                                                                                                                                                                                                          (N553)? { 1'b0, 1'b0, alu_adder_i } : 
                                                                                                                                                                                                                          (N451)? mac_res_q : 1'b0;
  assign md_state_n[0] = (N15)? N221 : 
                         (N203)? 1'b0 : 
                         (N206)? 1'b1 : 
                         (N209)? N728 : 
                         (N212)? 1'b1 : 
                         (N215)? 1'b0 : 
                         (N218)? 1'b0 : 1'b0;
  assign N15 = N200;
  assign md_state_n[2:1] = (N15)? { equal_to_zero, equal_to_zero } : 
                           (N203)? { 1'b0, 1'b1 } : 
                           (N206)? { 1'b0, 1'b1 } : 
                           (N209)? { N729, N728 } : 
                           (N212)? { 1'b1, 1'b0 } : 
                           (N215)? { 1'b1, 1'b1 } : 
                           (N218)? { 1'b0, 1'b0 } : 
                           (N16)? { 1'b0, 1'b0 } : 1'b0;
  assign N16 = N220;
  assign op_remainder_n = (N15)? { N723, N723, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222 } : 
                          (N206)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, op_numerator_q[31:31] } : 
                          (N209)? { 1'b0, next_remainder, N417 } : 
                          (N212)? { 1'b0, 1'b0, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418 } : 
                          (N215)? { N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487 } : 1'b0;
  assign alu_operand_a_o[32:1] = (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                 (N203)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                 (N206)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                 (N209)? mac_res_q[31:0] : 
                                 (N212)? mac_res_q[31:0] : 
                                 (N215)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                 (N218)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                 (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign alu_operand_b_o[32:1] = (N15)? { N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158 } : 
                                 (N203)? { N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315, N316, N317, N318 } : 
                                 (N206)? { N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158 } : 
                                 (N209)? { N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190 } : 
                                 (N212)? { N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190 } : 
                                 (N215)? { N521, N522, N523, N524, N525, N526, N527, N528, N529, N530, N531, N532, N533, N534, N535, N536, N537, N538, N539, N540, N541, N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552 } : 
                                 (N218)? { N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158 } : 
                                 (N16)? { N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158 } : 1'b0;
  assign div_counter_n = (N15)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                         (N203)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                         (N206)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                         (N209)? { N195, N194, N193, N192, N191 } : 
                         (N212)? { N195, N194, N193, N192, N191 } : 
                         (N215)? { N195, N194, N193, N192, N191 } : 
                         (N218)? { N195, N194, N193, N192, N191 } : 
                         (N16)? { N195, N194, N193, N192, N191 } : 1'b0;
  assign op_quotient_n = (N203)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N209)? next_quotient : 1'b0;
  assign div_valid = (N15)? 1'b0 : 
                     (N203)? 1'b0 : 
                     (N206)? 1'b0 : 
                     (N209)? 1'b0 : 
                     (N212)? 1'b0 : 
                     (N215)? 1'b0 : 
                     (N218)? 1'b1 : 
                     (N16)? 1'b0 : 1'b0;
  assign { N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564 } = (N17)? { 1'b0, 1'b0, mac_res_signed[15:0], mac_res_q[15:0] } : 
                                                                                                                                                                                                                          (N18)? mac_res_signed : 1'b0;
  assign N17 = N720;
  assign N18 = N719;
  assign { N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598 } = (N17)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mac_res_q[31:16] } : 
                                                                                                                                                                                                                          (N18)? mac_res_q : 1'b0;
  assign { N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632 } = (N17)? { 1'b0, 1'b0, mac_res_signed[15:0], mac_res_q[15:0] } : 
                                                                                                                                                                                                                          (N18)? mac_res_signed : 1'b0;
  assign mult_op_a = (N19)? op_a_i[15:0] : 
                     (N560)? op_a_i[15:0] : 
                     (N562)? op_a_i[31:16] : 
                     (N20)? op_a_i[31:16] : 1'b0;
  assign N19 = N558;
  assign N20 = N563;
  assign mult_op_b = (N19)? op_b_i[15:0] : 
                     (N560)? op_b_i[31:16] : 
                     (N562)? op_b_i[15:0] : 
                     (N20)? op_b_i[31:16] : 1'b0;
  assign sign_a = (N19)? 1'b0 : 
                  (N560)? 1'b0 : 
                  (N562)? N555 : 
                  (N20)? N555 : 1'b0;
  assign sign_b = (N19)? 1'b0 : 
                  (N560)? N554 : 
                  (N562)? 1'b0 : 
                  (N20)? N554 : 1'b0;
  assign accum = (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                 (N560)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mac_res_q[31:16] } : 
                 (N562)? { N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598 } : 
                 (N20)? { N666, N667, N668, N669, N670, N671, N672, N673, N674, N675, N676, N677, N678, N679, N680, N681, mac_res_q[33:16] } : 1'b0;
  assign mac_res_n = (N19)? mac_res_signed : 
                     (N560)? { N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564 } : 
                     (N562)? { N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632 } : 
                     (N20)? mac_res_signed : 1'b0;
  assign mult_state_n = (N19)? { 1'b0, 1'b1 } : 
                        (N560)? { 1'b1, 1'b0 } : 
                        (N562)? { N719, N719 } : 
                        (N20)? { 1'b0, 1'b0 } : 1'b0;
  assign mult_valid = (N19)? 1'b0 : 
                      (N560)? 1'b0 : 
                      (N562)? N720 : 
                      (N20)? 1'b1 : 1'b0;
  assign N21 = ~rst_ni;
  assign N22 = div_en_i | mult_en_i;
  assign N23 = ~N22;
  assign N58 = ~div_en_i;
  assign N93 = ~is_greater_equal;
  assign N94 = op_quotient_q[31] | one_shift[31];
  assign N95 = op_quotient_q[30] | one_shift[30];
  assign N96 = op_quotient_q[29] | one_shift[29];
  assign N97 = op_quotient_q[28] | one_shift[28];
  assign N98 = op_quotient_q[27] | one_shift[27];
  assign N99 = op_quotient_q[26] | one_shift[26];
  assign N100 = op_quotient_q[25] | one_shift[25];
  assign N101 = op_quotient_q[24] | one_shift[24];
  assign N102 = op_quotient_q[23] | one_shift[23];
  assign N103 = op_quotient_q[22] | one_shift[22];
  assign N104 = op_quotient_q[21] | one_shift[21];
  assign N105 = op_quotient_q[20] | one_shift[20];
  assign N106 = op_quotient_q[19] | one_shift[19];
  assign N107 = op_quotient_q[18] | one_shift[18];
  assign N108 = op_quotient_q[17] | one_shift[17];
  assign N109 = op_quotient_q[16] | one_shift[16];
  assign N110 = op_quotient_q[15] | one_shift[15];
  assign N111 = op_quotient_q[14] | one_shift[14];
  assign N112 = op_quotient_q[13] | one_shift[13];
  assign N113 = op_quotient_q[12] | one_shift[12];
  assign N114 = op_quotient_q[11] | one_shift[11];
  assign N115 = op_quotient_q[10] | one_shift[10];
  assign N116 = op_quotient_q[9] | one_shift[9];
  assign N117 = op_quotient_q[8] | one_shift[8];
  assign N118 = op_quotient_q[7] | one_shift[7];
  assign N119 = op_quotient_q[6] | one_shift[6];
  assign N120 = op_quotient_q[5] | one_shift[5];
  assign N121 = op_quotient_q[4] | one_shift[4];
  assign N122 = op_quotient_q[3] | one_shift[3];
  assign N123 = op_quotient_q[2] | one_shift[2];
  assign N124 = op_quotient_q[1] | one_shift[1];
  assign N125 = op_quotient_q[0] | one_shift[0];
  assign N126 = mac_res_q[31] ^ op_denominator_q[31];
  assign div_sign_a = op_a_i[31] & signed_mode_i[0];
  assign div_sign_b = op_b_i[31] & signed_mode_i[1];
  assign div_change_sign = div_sign_a ^ div_sign_b;
  assign N127 = ~op_b_i[31];
  assign N128 = ~op_b_i[30];
  assign N129 = ~op_b_i[29];
  assign N130 = ~op_b_i[28];
  assign N131 = ~op_b_i[27];
  assign N132 = ~op_b_i[26];
  assign N133 = ~op_b_i[25];
  assign N134 = ~op_b_i[24];
  assign N135 = ~op_b_i[23];
  assign N136 = ~op_b_i[22];
  assign N137 = ~op_b_i[21];
  assign N138 = ~op_b_i[20];
  assign N139 = ~op_b_i[19];
  assign N140 = ~op_b_i[18];
  assign N141 = ~op_b_i[17];
  assign N142 = ~op_b_i[16];
  assign N143 = ~op_b_i[15];
  assign N144 = ~op_b_i[14];
  assign N145 = ~op_b_i[13];
  assign N146 = ~op_b_i[12];
  assign N147 = ~op_b_i[11];
  assign N148 = ~op_b_i[10];
  assign N149 = ~op_b_i[9];
  assign N150 = ~op_b_i[8];
  assign N151 = ~op_b_i[7];
  assign N152 = ~op_b_i[6];
  assign N153 = ~op_b_i[5];
  assign N154 = ~op_b_i[4];
  assign N155 = ~op_b_i[3];
  assign N156 = ~op_b_i[2];
  assign N157 = ~op_b_i[1];
  assign N158 = ~op_b_i[0];
  assign N159 = ~op_denominator_q[31];
  assign N160 = ~op_denominator_q[30];
  assign N161 = ~op_denominator_q[29];
  assign N162 = ~op_denominator_q[28];
  assign N163 = ~op_denominator_q[27];
  assign N164 = ~op_denominator_q[26];
  assign N165 = ~op_denominator_q[25];
  assign N166 = ~op_denominator_q[24];
  assign N167 = ~op_denominator_q[23];
  assign N168 = ~op_denominator_q[22];
  assign N169 = ~op_denominator_q[21];
  assign N170 = ~op_denominator_q[20];
  assign N171 = ~op_denominator_q[19];
  assign N172 = ~op_denominator_q[18];
  assign N173 = ~op_denominator_q[17];
  assign N174 = ~op_denominator_q[16];
  assign N175 = ~op_denominator_q[15];
  assign N176 = ~op_denominator_q[14];
  assign N177 = ~op_denominator_q[13];
  assign N178 = ~op_denominator_q[12];
  assign N179 = ~op_denominator_q[11];
  assign N180 = ~op_denominator_q[10];
  assign N181 = ~op_denominator_q[9];
  assign N182 = ~op_denominator_q[8];
  assign N183 = ~op_denominator_q[7];
  assign N184 = ~op_denominator_q[6];
  assign N185 = ~op_denominator_q[5];
  assign N186 = ~op_denominator_q[4];
  assign N187 = ~op_denominator_q[3];
  assign N188 = ~op_denominator_q[2];
  assign N189 = ~op_denominator_q[1];
  assign N190 = ~op_denominator_q[0];
  assign N196 = ~md_state_q[2];
  assign N197 = ~md_state_q[1];
  assign N198 = ~md_state_q[0];
  assign N203 = ~N202;
  assign N206 = ~N205;
  assign N209 = ~N208;
  assign N212 = ~N211;
  assign N215 = ~N214;
  assign N218 = ~N217;
  assign N221 = ~equal_to_zero;
  assign N254 = ~div_sign_a;
  assign N287 = ~op_a_i[31];
  assign N288 = ~op_a_i[30];
  assign N289 = ~op_a_i[29];
  assign N290 = ~op_a_i[28];
  assign N291 = ~op_a_i[27];
  assign N292 = ~op_a_i[26];
  assign N293 = ~op_a_i[25];
  assign N294 = ~op_a_i[24];
  assign N295 = ~op_a_i[23];
  assign N296 = ~op_a_i[22];
  assign N297 = ~op_a_i[21];
  assign N298 = ~op_a_i[20];
  assign N299 = ~op_a_i[19];
  assign N300 = ~op_a_i[18];
  assign N301 = ~op_a_i[17];
  assign N302 = ~op_a_i[16];
  assign N303 = ~op_a_i[15];
  assign N304 = ~op_a_i[14];
  assign N305 = ~op_a_i[13];
  assign N306 = ~op_a_i[12];
  assign N307 = ~op_a_i[11];
  assign N308 = ~op_a_i[10];
  assign N309 = ~op_a_i[9];
  assign N310 = ~op_a_i[8];
  assign N311 = ~op_a_i[7];
  assign N312 = ~op_a_i[6];
  assign N313 = ~op_a_i[5];
  assign N314 = ~op_a_i[4];
  assign N315 = ~op_a_i[3];
  assign N316 = ~op_a_i[2];
  assign N317 = ~op_a_i[1];
  assign N318 = ~op_a_i[0];
  assign N319 = ~div_sign_b;
  assign N352 = ~N191;
  assign N353 = ~N192;
  assign N354 = N352 & N353;
  assign N355 = N352 & N192;
  assign N356 = N191 & N353;
  assign N357 = N191 & N192;
  assign N358 = ~N193;
  assign N359 = N354 & N358;
  assign N360 = N354 & N193;
  assign N361 = N356 & N358;
  assign N362 = N356 & N193;
  assign N363 = N355 & N358;
  assign N364 = N355 & N193;
  assign N365 = N357 & N358;
  assign N366 = N357 & N193;
  assign N367 = ~N194;
  assign N368 = N359 & N367;
  assign N369 = N359 & N194;
  assign N370 = N361 & N367;
  assign N371 = N361 & N194;
  assign N372 = N363 & N367;
  assign N373 = N363 & N194;
  assign N374 = N365 & N367;
  assign N375 = N365 & N194;
  assign N376 = N360 & N367;
  assign N377 = N360 & N194;
  assign N378 = N362 & N367;
  assign N379 = N362 & N194;
  assign N380 = N364 & N367;
  assign N381 = N364 & N194;
  assign N382 = N366 & N367;
  assign N383 = N366 & N194;
  assign N384 = ~N195;
  assign N385 = N368 & N384;
  assign N386 = N368 & N195;
  assign N387 = N370 & N384;
  assign N388 = N370 & N195;
  assign N389 = N372 & N384;
  assign N390 = N372 & N195;
  assign N391 = N374 & N384;
  assign N392 = N374 & N195;
  assign N393 = N376 & N384;
  assign N394 = N376 & N195;
  assign N395 = N378 & N384;
  assign N396 = N378 & N195;
  assign N397 = N380 & N384;
  assign N398 = N380 & N195;
  assign N399 = N382 & N384;
  assign N400 = N382 & N195;
  assign N401 = N369 & N384;
  assign N402 = N369 & N195;
  assign N403 = N371 & N384;
  assign N404 = N371 & N195;
  assign N405 = N373 & N384;
  assign N406 = N373 & N195;
  assign N407 = N375 & N384;
  assign N408 = N375 & N195;
  assign N409 = N377 & N384;
  assign N410 = N377 & N195;
  assign N411 = N379 & N384;
  assign N412 = N379 & N195;
  assign N413 = N381 & N384;
  assign N414 = N381 & N195;
  assign N415 = N383 & N384;
  assign N416 = N383 & N195;
  assign N450 = div_sign_a | N723;
  assign N451 = ~N450;
  assign N452 = ~div_change_sign;
  assign N521 = ~mac_res_q[31];
  assign N522 = ~mac_res_q[30];
  assign N523 = ~mac_res_q[29];
  assign N524 = ~mac_res_q[28];
  assign N525 = ~mac_res_q[27];
  assign N526 = ~mac_res_q[26];
  assign N527 = ~mac_res_q[25];
  assign N528 = ~mac_res_q[24];
  assign N529 = ~mac_res_q[23];
  assign N530 = ~mac_res_q[22];
  assign N531 = ~mac_res_q[21];
  assign N532 = ~mac_res_q[20];
  assign N533 = ~mac_res_q[19];
  assign N534 = ~mac_res_q[18];
  assign N535 = ~mac_res_q[17];
  assign N536 = ~mac_res_q[16];
  assign N537 = ~mac_res_q[15];
  assign N538 = ~mac_res_q[14];
  assign N539 = ~mac_res_q[13];
  assign N540 = ~mac_res_q[12];
  assign N541 = ~mac_res_q[11];
  assign N542 = ~mac_res_q[10];
  assign N543 = ~mac_res_q[9];
  assign N544 = ~mac_res_q[8];
  assign N545 = ~mac_res_q[7];
  assign N546 = ~mac_res_q[6];
  assign N547 = ~mac_res_q[5];
  assign N548 = ~mac_res_q[4];
  assign N549 = ~mac_res_q[3];
  assign N550 = ~mac_res_q[2];
  assign N551 = ~mac_res_q[1];
  assign N552 = ~mac_res_q[0];
  assign N553 = div_sign_a & N722;
  assign valid_o = mult_valid | div_valid;
  assign N554 = signed_mode_i[1] & op_b_i[31];
  assign N555 = signed_mode_i[0] & op_a_i[31];
  assign N556 = ~mult_state_q[1];
  assign N557 = ~mult_state_q[0];
  assign N560 = ~N559;
  assign N562 = ~N561;
  assign N666 = N730 & mac_res_q[33];
  assign N667 = N730 & mac_res_q[33];
  assign N668 = N730 & mac_res_q[33];
  assign N669 = N730 & mac_res_q[33];
  assign N670 = N730 & mac_res_q[33];
  assign N671 = N730 & mac_res_q[33];
  assign N672 = N730 & mac_res_q[33];
  assign N673 = N730 & mac_res_q[33];
  assign N674 = N730 & mac_res_q[33];
  assign N675 = N730 & mac_res_q[33];
  assign N676 = N730 & mac_res_q[33];
  assign N677 = N730 & mac_res_q[33];
  assign N678 = N730 & mac_res_q[33];
  assign N679 = N730 & mac_res_q[33];
  assign N680 = N730 & mac_res_q[33];
  assign N681 = N730 & mac_res_q[33];
  assign N682 = N200 & div_en_i;
  assign N683 = N206 & div_en_i;
  assign N684 = N682 | N683;
  assign N685 = N209 & div_en_i;
  assign N686 = N684 | N685;
  assign N687 = N212 & div_en_i;
  assign N688 = N686 | N687;
  assign N689 = N215 & div_en_i;
  assign N690 = N688 | N689;
  assign N691 = N218 & div_en_i;
  assign N692 = N690 | N691;
  assign N693 = N220 & div_en_i;
  assign N694 = N692 | N693;
  assign N695 = ~N694;
  assign N696 = div_en_i & N695;
  assign N697 = N684 | N687;
  assign N698 = N697 | N689;
  assign N699 = N698 | N691;
  assign N700 = N699 | N693;
  assign N701 = ~N700;
  assign N702 = div_en_i & N701;
  assign N703 = N203 & div_en_i;
  assign N704 = N218 & div_en_i;
  assign N705 = N703 | N704;
  assign N706 = N220 & div_en_i;
  assign N707 = N705 | N706;
  assign N708 = N707 | N23;
  assign N709 = ~N708;
  assign N710 = N203 & div_en_i;
  assign N711 = N682 | N710;
  assign N712 = N711 | N685;
  assign N713 = N712 | N687;
  assign N714 = N713 | N689;
  assign N715 = N714 | N691;
  assign N716 = N715 | N693;
  assign N717 = ~N716;
  assign N718 = div_en_i & N717;

endmodule



module ibex_ex_block_1
(
  clk_i,
  rst_ni,
  alu_operator_i,
  alu_operand_a_i,
  alu_operand_b_i,
  multdiv_operator_i,
  mult_en_i,
  div_en_i,
  multdiv_signed_mode_i,
  multdiv_operand_a_i,
  multdiv_operand_b_i,
  alu_adder_result_ex_o,
  regfile_wdata_ex_o,
  jump_target_o,
  branch_decision_o,
  ex_valid_o
);

  input [4:0] alu_operator_i;
  input [31:0] alu_operand_a_i;
  input [31:0] alu_operand_b_i;
  input [1:0] multdiv_operator_i;
  input [1:0] multdiv_signed_mode_i;
  input [31:0] multdiv_operand_a_i;
  input [31:0] multdiv_operand_b_i;
  output [31:0] alu_adder_result_ex_o;
  output [31:0] regfile_wdata_ex_o;
  output [31:0] jump_target_o;
  input clk_i;
  input rst_ni;
  input mult_en_i;
  input div_en_i;
  output branch_decision_o;
  output ex_valid_o;
  wire [31:0] alu_adder_result_ex_o,regfile_wdata_ex_o,jump_target_o,multdiv_result,
  alu_result;
  wire branch_decision_o,ex_valid_o,N0,N1,multdiv_en,N2,alu_is_equal_result,
  multdiv_valid;
  wire [32:0] multdiv_alu_operand_a,multdiv_alu_operand_b;
  wire [33:0] alu_adder_result_ext;
  assign alu_adder_result_ex_o[31] = jump_target_o[31];
  assign alu_adder_result_ex_o[30] = jump_target_o[30];
  assign alu_adder_result_ex_o[29] = jump_target_o[29];
  assign alu_adder_result_ex_o[28] = jump_target_o[28];
  assign alu_adder_result_ex_o[27] = jump_target_o[27];
  assign alu_adder_result_ex_o[26] = jump_target_o[26];
  assign alu_adder_result_ex_o[25] = jump_target_o[25];
  assign alu_adder_result_ex_o[24] = jump_target_o[24];
  assign alu_adder_result_ex_o[23] = jump_target_o[23];
  assign alu_adder_result_ex_o[22] = jump_target_o[22];
  assign alu_adder_result_ex_o[21] = jump_target_o[21];
  assign alu_adder_result_ex_o[20] = jump_target_o[20];
  assign alu_adder_result_ex_o[19] = jump_target_o[19];
  assign alu_adder_result_ex_o[18] = jump_target_o[18];
  assign alu_adder_result_ex_o[17] = jump_target_o[17];
  assign alu_adder_result_ex_o[16] = jump_target_o[16];
  assign alu_adder_result_ex_o[15] = jump_target_o[15];
  assign alu_adder_result_ex_o[14] = jump_target_o[14];
  assign alu_adder_result_ex_o[13] = jump_target_o[13];
  assign alu_adder_result_ex_o[12] = jump_target_o[12];
  assign alu_adder_result_ex_o[11] = jump_target_o[11];
  assign alu_adder_result_ex_o[10] = jump_target_o[10];
  assign alu_adder_result_ex_o[9] = jump_target_o[9];
  assign alu_adder_result_ex_o[8] = jump_target_o[8];
  assign alu_adder_result_ex_o[7] = jump_target_o[7];
  assign alu_adder_result_ex_o[6] = jump_target_o[6];
  assign alu_adder_result_ex_o[5] = jump_target_o[5];
  assign alu_adder_result_ex_o[4] = jump_target_o[4];
  assign alu_adder_result_ex_o[3] = jump_target_o[3];
  assign alu_adder_result_ex_o[2] = jump_target_o[2];
  assign alu_adder_result_ex_o[1] = jump_target_o[1];
  assign alu_adder_result_ex_o[0] = jump_target_o[0];

  ibex_alu
  alu_i
  (
    .operator_i(alu_operator_i),
    .operand_a_i(alu_operand_a_i),
    .operand_b_i(alu_operand_b_i),
    .multdiv_operand_a_i(multdiv_alu_operand_a),
    .multdiv_operand_b_i(multdiv_alu_operand_b),
    .multdiv_en_i(div_en_i),
    .adder_result_o(jump_target_o),
    .adder_result_ext_o(alu_adder_result_ext),
    .result_o(alu_result),
    .comparison_result_o(branch_decision_o),
    .is_equal_result_o(alu_is_equal_result)
  );


  ibex_multdiv_fast
  gen_multdiv_fast_multdiv_i
  (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .mult_en_i(mult_en_i),
    .div_en_i(div_en_i),
    .operator_i(multdiv_operator_i),
    .signed_mode_i(multdiv_signed_mode_i),
    .op_a_i(multdiv_operand_a_i),
    .op_b_i(multdiv_operand_b_i),
    .alu_adder_ext_i(alu_adder_result_ext),
    .alu_adder_i(jump_target_o),
    .equal_to_zero(alu_is_equal_result),
    .alu_operand_a_o(multdiv_alu_operand_a),
    .alu_operand_b_o(multdiv_alu_operand_b),
    .multdiv_result_o(multdiv_result),
    .valid_o(multdiv_valid)
  );

  assign regfile_wdata_ex_o = (N0)? multdiv_result : 
                              (N1)? alu_result : 1'b0;
  assign N0 = multdiv_en;
  assign N1 = N2;
  assign ex_valid_o = (N0)? multdiv_valid : 
                      (N1)? 1'b1 : 1'b0;
  assign multdiv_en = mult_en_i | div_en_i;
  assign N2 = ~multdiv_en;

endmodule



module ibex_load_store_unit
(
  clk_i,
  rst_ni,
  data_req_o,
  data_gnt_i,
  data_rvalid_i,
  data_err_i,
  data_addr_o,
  data_we_o,
  data_be_o,
  data_wdata_o,
  data_rdata_i,
  data_we_ex_i,
  data_type_ex_i,
  data_wdata_ex_i,
  data_reg_offset_ex_i,
  data_sign_ext_ex_i,
  data_rdata_ex_o,
  data_req_ex_i,
  adder_result_ex_i,
  addr_incr_req_o,
  addr_last_o,
  data_valid_o,
  load_err_o,
  store_err_o,
  busy_o
);

  output [31:0] data_addr_o;
  output [3:0] data_be_o;
  output [31:0] data_wdata_o;
  input [31:0] data_rdata_i;
  input [1:0] data_type_ex_i;
  input [31:0] data_wdata_ex_i;
  input [1:0] data_reg_offset_ex_i;
  output [31:0] data_rdata_ex_o;
  input [31:0] adder_result_ex_i;
  output [31:0] addr_last_o;
  input clk_i;
  input rst_ni;
  input data_gnt_i;
  input data_rvalid_i;
  input data_err_i;
  input data_we_ex_i;
  input data_sign_ext_ex_i;
  input data_req_ex_i;
  output data_req_o;
  output data_we_o;
  output addr_incr_req_o;
  output data_valid_o;
  output load_err_o;
  output store_err_o;
  output busy_o;
  wire [31:0] data_addr_o,data_wdata_o,data_rdata_ex_o,rdata_w_ext,rdata_h_ext,rdata_b_ext,
  addr_last_d;
  wire [3:0] data_be_o;
  wire data_req_o,data_we_o,addr_incr_req_o,data_valid_o,load_err_o,store_err_o,busy_o,
  N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  data_we_ex_i,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
  N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,
  N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,
  N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,
  N115,split_misaligned_access,handle_misaligned_d,N116,N117,N118,N119,N120,N121,
  N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,
  N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,
  N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,
  N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,
  N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196;
  wire [1:0] wdata_offset;
  wire [2:0] ls_fsm_ns;
  reg data_we_q,data_sign_ext_q,handle_misaligned_q;
  reg [31:8] rdata_q;
  reg [1:0] rdata_offset_q,data_type_q;
  reg [2:0] ls_fsm_cs;
  reg [31:0] addr_last_o;
  assign data_addr_o[0] = 1'b0;
  assign data_addr_o[1] = 1'b0;
  assign data_addr_o[31] = adder_result_ex_i[31];
  assign data_addr_o[30] = adder_result_ex_i[30];
  assign data_addr_o[29] = adder_result_ex_i[29];
  assign data_addr_o[28] = adder_result_ex_i[28];
  assign data_addr_o[27] = adder_result_ex_i[27];
  assign data_addr_o[26] = adder_result_ex_i[26];
  assign data_addr_o[25] = adder_result_ex_i[25];
  assign data_addr_o[24] = adder_result_ex_i[24];
  assign data_addr_o[23] = adder_result_ex_i[23];
  assign data_addr_o[22] = adder_result_ex_i[22];
  assign data_addr_o[21] = adder_result_ex_i[21];
  assign data_addr_o[20] = adder_result_ex_i[20];
  assign data_addr_o[19] = adder_result_ex_i[19];
  assign data_addr_o[18] = adder_result_ex_i[18];
  assign data_addr_o[17] = adder_result_ex_i[17];
  assign data_addr_o[16] = adder_result_ex_i[16];
  assign data_addr_o[15] = adder_result_ex_i[15];
  assign data_addr_o[14] = adder_result_ex_i[14];
  assign data_addr_o[13] = adder_result_ex_i[13];
  assign data_addr_o[12] = adder_result_ex_i[12];
  assign data_addr_o[11] = adder_result_ex_i[11];
  assign data_addr_o[10] = adder_result_ex_i[10];
  assign data_addr_o[9] = adder_result_ex_i[9];
  assign data_addr_o[8] = adder_result_ex_i[8];
  assign data_addr_o[7] = adder_result_ex_i[7];
  assign data_addr_o[6] = adder_result_ex_i[6];
  assign data_addr_o[5] = adder_result_ex_i[5];
  assign data_addr_o[4] = adder_result_ex_i[4];
  assign data_addr_o[3] = adder_result_ex_i[3];
  assign data_addr_o[2] = adder_result_ex_i[2];
  assign data_we_o = data_we_ex_i;
  assign N58 = N56 & N57;
  assign N59 = adder_result_ex_i[1] | N57;
  assign N61 = N56 | adder_result_ex_i[0];
  assign N63 = adder_result_ex_i[1] & adder_result_ex_i[0];
  assign N70 = N68 & N69;
  assign N71 = wdata_offset[1] | N69;
  assign N73 = N68 | wdata_offset[0];
  assign N75 = wdata_offset[1] & wdata_offset[0];

  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      data_we_q <= 1'b0;
    end else if(data_gnt_i) begin
      data_we_q <= data_we_ex_i;
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_q[31] <= 1'b0;
    end else if(N76) begin
      rdata_q[31] <= data_rdata_i[31];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_q[30] <= 1'b0;
    end else if(N76) begin
      rdata_q[30] <= data_rdata_i[30];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_q[29] <= 1'b0;
    end else if(N76) begin
      rdata_q[29] <= data_rdata_i[29];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_q[28] <= 1'b0;
    end else if(N76) begin
      rdata_q[28] <= data_rdata_i[28];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_q[27] <= 1'b0;
    end else if(N76) begin
      rdata_q[27] <= data_rdata_i[27];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_q[26] <= 1'b0;
    end else if(N76) begin
      rdata_q[26] <= data_rdata_i[26];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_q[25] <= 1'b0;
    end else if(N76) begin
      rdata_q[25] <= data_rdata_i[25];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_q[24] <= 1'b0;
    end else if(N76) begin
      rdata_q[24] <= data_rdata_i[24];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_q[23] <= 1'b0;
    end else if(N76) begin
      rdata_q[23] <= data_rdata_i[23];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_q[22] <= 1'b0;
    end else if(N76) begin
      rdata_q[22] <= data_rdata_i[22];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_q[21] <= 1'b0;
    end else if(N76) begin
      rdata_q[21] <= data_rdata_i[21];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_q[20] <= 1'b0;
    end else if(N76) begin
      rdata_q[20] <= data_rdata_i[20];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_q[19] <= 1'b0;
    end else if(N76) begin
      rdata_q[19] <= data_rdata_i[19];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_q[18] <= 1'b0;
    end else if(N76) begin
      rdata_q[18] <= data_rdata_i[18];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_q[17] <= 1'b0;
    end else if(N76) begin
      rdata_q[17] <= data_rdata_i[17];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_q[16] <= 1'b0;
    end else if(N76) begin
      rdata_q[16] <= data_rdata_i[16];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_q[15] <= 1'b0;
    end else if(N76) begin
      rdata_q[15] <= data_rdata_i[15];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_q[14] <= 1'b0;
    end else if(N76) begin
      rdata_q[14] <= data_rdata_i[14];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_q[13] <= 1'b0;
    end else if(N76) begin
      rdata_q[13] <= data_rdata_i[13];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_q[12] <= 1'b0;
    end else if(N76) begin
      rdata_q[12] <= data_rdata_i[12];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_q[11] <= 1'b0;
    end else if(N76) begin
      rdata_q[11] <= data_rdata_i[11];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_q[10] <= 1'b0;
    end else if(N76) begin
      rdata_q[10] <= data_rdata_i[10];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_q[9] <= 1'b0;
    end else if(N76) begin
      rdata_q[9] <= data_rdata_i[9];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_q[8] <= 1'b0;
    end else if(N76) begin
      rdata_q[8] <= data_rdata_i[8];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_offset_q[1] <= 1'b0;
    end else if(data_gnt_i) begin
      rdata_offset_q[1] <= adder_result_ex_i[1];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      rdata_offset_q[0] <= 1'b0;
    end else if(data_gnt_i) begin
      rdata_offset_q[0] <= adder_result_ex_i[0];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      data_type_q[1] <= 1'b0;
    end else if(data_gnt_i) begin
      data_type_q[1] <= data_type_ex_i[1];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      data_type_q[0] <= 1'b0;
    end else if(data_gnt_i) begin
      data_type_q[0] <= data_type_ex_i[0];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      data_sign_ext_q <= 1'b0;
    end else if(data_gnt_i) begin
      data_sign_ext_q <= data_sign_ext_ex_i;
    end 
  end

  assign N81 = N79 & N80;
  assign N82 = rdata_offset_q[1] | N80;
  assign N84 = N79 | rdata_offset_q[0];
  assign N86 = rdata_offset_q[1] & rdata_offset_q[0];
  assign N88 = N79 & N80;
  assign N89 = rdata_offset_q[1] | N80;
  assign N91 = N79 | rdata_offset_q[0];
  assign N93 = rdata_offset_q[1] & rdata_offset_q[0];
  assign N98 = N79 & N80;
  assign N99 = rdata_offset_q[1] | N80;
  assign N101 = N79 | rdata_offset_q[0];
  assign N103 = rdata_offset_q[1] & rdata_offset_q[0];
  assign N110 = N108 & N109;
  assign N111 = data_type_q[1] | N109;
  assign N113 = N108 | data_type_q[0];
  assign N114 = data_type_q[1] & data_type_q[0];
  assign N119 = N116 & N117;
  assign N120 = N119 & N118;
  assign N121 = ls_fsm_cs[2] | ls_fsm_cs[1];
  assign N122 = N121 | N118;
  assign N124 = ls_fsm_cs[2] | N117;
  assign N125 = N124 | ls_fsm_cs[0];
  assign N127 = ls_fsm_cs[2] | N117;
  assign N128 = N127 | N118;
  assign N130 = N116 | ls_fsm_cs[1];
  assign N131 = N130 | ls_fsm_cs[0];
  assign N133 = ls_fsm_cs[2] & ls_fsm_cs[0];
  assign N134 = ls_fsm_cs[2] & ls_fsm_cs[1];

  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      handle_misaligned_q <= 1'b0;
    end else if(N171) begin
      handle_misaligned_q <= handle_misaligned_d;
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      ls_fsm_cs[2] <= 1'b0;
    end else if(N175) begin
      ls_fsm_cs[2] <= ls_fsm_ns[2];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      ls_fsm_cs[1] <= 1'b0;
    end else if(N175) begin
      ls_fsm_cs[1] <= ls_fsm_ns[1];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      ls_fsm_cs[0] <= 1'b0;
    end else if(N175) begin
      ls_fsm_cs[0] <= ls_fsm_ns[0];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[31] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[31] <= addr_last_d[31];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[30] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[30] <= addr_last_d[30];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[29] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[29] <= addr_last_d[29];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[28] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[28] <= addr_last_d[28];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[27] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[27] <= addr_last_d[27];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[26] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[26] <= addr_last_d[26];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[25] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[25] <= addr_last_d[25];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[24] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[24] <= addr_last_d[24];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[23] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[23] <= addr_last_d[23];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[22] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[22] <= addr_last_d[22];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[21] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[21] <= addr_last_d[21];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[20] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[20] <= addr_last_d[20];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[19] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[19] <= addr_last_d[19];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[18] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[18] <= addr_last_d[18];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[17] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[17] <= addr_last_d[17];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[16] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[16] <= addr_last_d[16];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[15] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[15] <= addr_last_d[15];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[14] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[14] <= addr_last_d[14];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[13] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[13] <= addr_last_d[13];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[12] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[12] <= addr_last_d[12];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[11] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[11] <= addr_last_d[11];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[10] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[10] <= addr_last_d[10];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[9] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[9] <= addr_last_d[9];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[8] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[8] <= addr_last_d[8];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[7] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[7] <= addr_last_d[7];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[6] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[6] <= addr_last_d[6];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[5] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[5] <= addr_last_d[5];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[4] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[4] <= addr_last_d[4];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[3] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[3] <= addr_last_d[3];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[2] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[2] <= addr_last_d[2];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[1] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[1] <= addr_last_d[1];
    end 
  end


  always @(posedge clk_i or posedge N78) begin
    if(N78) begin
      addr_last_o[0] <= 1'b0;
    end else if(1'b1) begin
      addr_last_o[0] <= addr_last_d[0];
    end 
  end

  assign N176 = ~ls_fsm_cs[2];
  assign N177 = ls_fsm_cs[1] | N176;
  assign N178 = ls_fsm_cs[0] | N177;
  assign N179 = ~N178;
  assign N180 = data_type_ex_i[0] | data_type_ex_i[1];
  assign N181 = ~N180;
  assign N182 = adder_result_ex_i[0] | adder_result_ex_i[1];
  assign N183 = ~data_type_ex_i[0];
  assign N184 = N183 | data_type_ex_i[1];
  assign N185 = ~N184;
  assign N186 = adder_result_ex_i[0] & adder_result_ex_i[1];
  assign wdata_offset = adder_result_ex_i[1:0] - data_reg_offset_ex_i;
  assign N42 = N0 & N1;
  assign N0 = ~data_type_ex_i[1];
  assign N1 = ~data_type_ex_i[0];
  assign N43 = N2 & N3;
  assign N2 = ~data_type_ex_i[1];
  assign N3 = ~N42;
  assign { N45, N44 } = (N4)? { 1'b1, 1'b1 } : 
                        (N5)? { 1'b1, 1'b1 } : 
                        (N6)? { 1'b1, 1'b0 } : 
                        (N7)? { 1'b0, 1'b0 } : 1'b0;
  assign N4 = N58;
  assign N5 = N60;
  assign N6 = N62;
  assign N7 = N63;
  assign { N47, N46 } = (N4)? { 1'b0, 1'b0 } : 
                        (N5)? { 1'b0, 1'b1 } : 
                        (N6)? { 1'b1, 1'b1 } : 
                        (N7)? { 1'b1, 1'b1 } : 1'b0;
  assign { N50, N49, N48 } = (N8)? { N45, N44, N64 } : 
                             (N9)? { N67, N47, N46 } : 1'b0;
  assign N8 = N41;
  assign N9 = handle_misaligned_q;
  assign N51 = (N4)? 1'b0 : 
               (N5)? 1'b1 : 
               (N6)? 1'b1 : 
               (N7)? 1'b0 : 1'b0;
  assign { N55, N54, N53, N52 } = (N8)? { N47, N51, N44, N64 } : 
                                  (N9)? { 1'b0, 1'b0, 1'b0, 1'b1 } : 1'b0;
  assign { N67, N66, N65, N64 } = (N4)? { 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                  (N5)? { 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                  (N6)? { 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                  (N7)? { 1'b1, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign data_be_o = (N10)? { N41, N50, N49, N48 } : 
                     (N11)? { N55, N54, N53, N52 } : 
                     (N12)? { N67, N66, N65, N64 } : 1'b0;
  assign N10 = N42;
  assign N11 = N43;
  assign N12 = data_type_ex_i[1];
  assign data_wdata_o = (N13)? data_wdata_ex_i : 
                        (N14)? { data_wdata_ex_i[23:0], data_wdata_ex_i[31:24] } : 
                        (N15)? { data_wdata_ex_i[15:0], data_wdata_ex_i[31:16] } : 
                        (N16)? { data_wdata_ex_i[7:0], data_wdata_ex_i[31:8] } : 1'b0;
  assign N13 = N70;
  assign N14 = N72;
  assign N15 = N74;
  assign N16 = N75;
  assign rdata_w_ext = (N17)? data_rdata_i : 
                       (N18)? { data_rdata_i[7:0], rdata_q } : 
                       (N19)? { data_rdata_i[15:0], rdata_q[31:16] } : 
                       (N20)? { data_rdata_i[23:0], rdata_q[31:24] } : 1'b0;
  assign N17 = N81;
  assign N18 = N83;
  assign N19 = N85;
  assign N20 = N86;
  assign N94 = (N21)? 1'b0 : 
               (N22)? data_rdata_i[15] : 1'b0;
  assign N21 = N87;
  assign N22 = data_sign_ext_q;
  assign N95 = (N21)? 1'b0 : 
               (N22)? data_rdata_i[23] : 1'b0;
  assign N96 = (N21)? 1'b0 : 
               (N22)? data_rdata_i[31] : 1'b0;
  assign N97 = (N21)? 1'b0 : 
               (N22)? data_rdata_i[7] : 1'b0;
  assign rdata_h_ext = (N23)? { N94, N94, N94, N94, N94, N94, N94, N94, N94, N94, N94, N94, N94, N94, N94, N94, data_rdata_i[15:0] } : 
                       (N24)? { N95, N95, N95, N95, N95, N95, N95, N95, N95, N95, N95, N95, N95, N95, N95, N95, data_rdata_i[23:8] } : 
                       (N25)? { N96, N96, N96, N96, N96, N96, N96, N96, N96, N96, N96, N96, N96, N96, N96, N96, data_rdata_i[31:16] } : 
                       (N26)? { N97, N97, N97, N97, N97, N97, N97, N97, N97, N97, N97, N97, N97, N97, N97, N97, data_rdata_i[7:0], rdata_q[31:24] } : 1'b0;
  assign N23 = N88;
  assign N24 = N90;
  assign N25 = N92;
  assign N26 = N93;
  assign N104 = (N21)? 1'b0 : 
                (N22)? data_rdata_i[7] : 1'b0;
  assign N105 = (N21)? 1'b0 : 
                (N22)? data_rdata_i[15] : 1'b0;
  assign N106 = (N21)? 1'b0 : 
                (N22)? data_rdata_i[23] : 1'b0;
  assign N107 = (N21)? 1'b0 : 
                (N22)? data_rdata_i[31] : 1'b0;
  assign rdata_b_ext = (N27)? { N104, N104, N104, N104, N104, N104, N104, N104, N104, N104, N104, N104, N104, N104, N104, N104, N104, N104, N104, N104, N104, N104, N104, N104, data_rdata_i[7:0] } : 
                       (N28)? { N105, N105, N105, N105, N105, N105, N105, N105, N105, N105, N105, N105, N105, N105, N105, N105, N105, N105, N105, N105, N105, N105, N105, N105, data_rdata_i[15:8] } : 
                       (N29)? { N106, N106, N106, N106, N106, N106, N106, N106, N106, N106, N106, N106, N106, N106, N106, N106, N106, N106, N106, N106, N106, N106, N106, N106, data_rdata_i[23:16] } : 
                       (N30)? { N107, N107, N107, N107, N107, N107, N107, N107, N107, N107, N107, N107, N107, N107, N107, N107, N107, N107, N107, N107, N107, N107, N107, N107, data_rdata_i[31:24] } : 1'b0;
  assign N27 = N98;
  assign N28 = N100;
  assign N29 = N102;
  assign N30 = N103;
  assign data_rdata_ex_o = (N31)? rdata_w_ext : 
                           (N32)? rdata_h_ext : 
                           (N33)? rdata_b_ext : 1'b0;
  assign N31 = N110;
  assign N32 = N112;
  assign N33 = N115;
  assign { N143, N142, N141 } = (N34)? { N139, split_misaligned_access, 1'b0 } : 
                                (N153)? { 1'b0, 1'b0, 1'b1 } : 
                                (N138)? { 1'b0, 1'b1, 1'b1 } : 1'b0;
  assign N34 = data_gnt_i;
  assign { N146, N145 } = (N35)? { 1'b0, 1'b0 } : 
                          (N36)? { data_gnt_i, N77 } : 1'b0;
  assign N35 = data_err_i;
  assign N36 = N144;
  assign N147 = (N37)? N144 : 
                (N38)? 1'b0 : 1'b0;
  assign N37 = data_rvalid_i;
  assign N38 = N152;
  assign N148 = (N37)? data_err_i : 
                (N38)? 1'b0 : 1'b0;
  assign { N151, N150, N149 } = (N37)? { N146, N145, N145 } : 
                                (N38)? { 1'b0, 1'b1, 1'b0 } : 1'b0;
  assign handle_misaligned_d = (N39)? split_misaligned_access : 
                               (N123)? 1'b1 : 
                               (N126)? 1'b0 : 
                               (N132)? 1'b0 : 1'b0;
  assign N39 = N120;
  assign data_req_o = (N39)? data_req_ex_i : 
                      (N123)? 1'b1 : 
                      (N126)? N147 : 
                      (N129)? 1'b1 : 
                      (N132)? 1'b0 : 
                      (N135)? 1'b0 : 1'b0;
  assign ls_fsm_ns[0] = (N39)? N141 : 
                        (N123)? 1'b0 : 
                        (N126)? N149 : 
                        (N129)? 1'b0 : 
                        (N132)? 1'b0 : 1'b0;
  assign ls_fsm_ns[2:1] = (N39)? { N143, N142 } : 
                          (N123)? { 1'b0, 1'b1 } : 
                          (N126)? { N151, N150 } : 
                          (N129)? { 1'b1, 1'b0 } : 
                          (N132)? { N152, 1'b0 } : 
                          (N135)? { 1'b0, 1'b0 } : 1'b0;
  assign addr_incr_req_o = (N39)? 1'b0 : 
                           (N123)? 1'b0 : 
                           (N126)? 1'b1 : 
                           (N129)? handle_misaligned_q : 
                           (N132)? 1'b0 : 
                           (N135)? 1'b0 : 1'b0;
  assign data_valid_o = (N39)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N126)? N148 : 
                        (N129)? 1'b0 : 
                        (N132)? data_rvalid_i : 
                        (N135)? 1'b0 : 1'b0;
  assign addr_last_d = (N40)? adder_result_ex_i : 
                       (N155)? addr_last_o : 1'b0;
  assign N40 = N154;
  assign N41 = ~handle_misaligned_q;
  assign N56 = ~adder_result_ex_i[1];
  assign N57 = ~adder_result_ex_i[0];
  assign N60 = ~N59;
  assign N62 = ~N61;
  assign N68 = ~wdata_offset[1];
  assign N69 = ~wdata_offset[0];
  assign N72 = ~N71;
  assign N74 = ~N73;
  assign N76 = N188 & handle_misaligned_q;
  assign N188 = data_rvalid_i & N187;
  assign N187 = ~data_we_q;
  assign N77 = ~data_gnt_i;
  assign N78 = ~rst_ni;
  assign N79 = ~rdata_offset_q[1];
  assign N80 = ~rdata_offset_q[0];
  assign N83 = ~N82;
  assign N85 = ~N84;
  assign N87 = ~data_sign_ext_q;
  assign N90 = ~N89;
  assign N92 = ~N91;
  assign N100 = ~N99;
  assign N102 = ~N101;
  assign N108 = ~data_type_q[1];
  assign N109 = ~data_type_q[0];
  assign N112 = ~N111;
  assign N115 = N189 | N114;
  assign N189 = ~N113;
  assign split_misaligned_access = N190 | N191;
  assign N190 = N181 & N182;
  assign N191 = N185 & N186;
  assign N116 = ~ls_fsm_cs[2];
  assign N117 = ~ls_fsm_cs[1];
  assign N118 = ~ls_fsm_cs[0];
  assign N123 = ~N122;
  assign N126 = ~N125;
  assign N129 = ~N128;
  assign N132 = ~N131;
  assign N135 = N133 | N134;
  assign N136 = ~data_req_ex_i;
  assign N137 = split_misaligned_access | data_gnt_i;
  assign N138 = ~N137;
  assign N139 = ~split_misaligned_access;
  assign N140 = ~data_gnt_i;
  assign N144 = ~data_err_i;
  assign N152 = ~data_rvalid_i;
  assign N153 = split_misaligned_access & N140;
  assign N154 = N192 & N194;
  assign N192 = data_req_o & data_gnt_i;
  assign N194 = ~N193;
  assign N193 = load_err_o | store_err_o;
  assign N155 = ~N154;
  assign load_err_o = N195 & N187;
  assign N195 = data_err_i & data_rvalid_i;
  assign store_err_o = N196 & data_we_q;
  assign N196 = data_err_i & data_rvalid_i;
  assign busy_o = N179 | data_req_o;
  assign N156 = data_req_ex_i & N120;
  assign N157 = N140 & N156;
  assign N158 = N136 & N120;
  assign N159 = N157 | N158;
  assign N160 = N77 & N123;
  assign N161 = N159 | N160;
  assign N162 = data_rvalid_i & N126;
  assign N163 = N144 & N162;
  assign N164 = N161 | N163;
  assign N165 = N152 & N126;
  assign N166 = N164 | N165;
  assign N167 = N166 | N129;
  assign N168 = N152 & N132;
  assign N169 = N167 | N168;
  assign N170 = N169 | N135;
  assign N171 = ~N170;
  assign N172 = N158 | N160;
  assign N173 = N77 & N129;
  assign N174 = N172 | N173;
  assign N175 = ~N174;

endmodule



module ibex_cs_registers_00000000_00000028_0_1
(
  clk_i,
  rst_ni,
  core_id_i,
  cluster_id_i,
  csr_access_i,
  csr_addr_i,
  csr_wdata_i,
  csr_op_i,
  csr_rdata_o,
  m_irq_enable_o,
  csr_mepc_o,
  debug_cause_i,
  debug_csr_save_i,
  csr_depc_o,
  debug_single_step_o,
  debug_ebreakm_o,
  pc_if_i,
  pc_id_i,
  csr_save_if_i,
  csr_save_id_i,
  csr_restore_mret_i,
  csr_restore_dret_i,
  csr_save_cause_i,
  csr_mtvec_i,
  csr_mcause_i,
  csr_mtval_i,
  illegal_csr_insn_o,
  instr_new_id_i,
  instr_ret_i,
  instr_ret_compressed_i,
  imiss_i,
  pc_set_i,
  jump_i,
  branch_i,
  branch_taken_i,
  mem_load_i,
  mem_store_i,
  lsu_busy_i
);

  input [3:0] core_id_i;
  input [5:0] cluster_id_i;
  input [11:0] csr_addr_i;
  input [31:0] csr_wdata_i;
  input [1:0] csr_op_i;
  output [31:0] csr_rdata_o;
  output [31:0] csr_mepc_o;
  input [2:0] debug_cause_i;
  output [31:0] csr_depc_o;
  input [31:0] pc_if_i;
  input [31:0] pc_id_i;
  input [31:0] csr_mtvec_i;
  input [5:0] csr_mcause_i;
  input [31:0] csr_mtval_i;
  input clk_i;
  input rst_ni;
  input csr_access_i;
  input debug_csr_save_i;
  input csr_save_if_i;
  input csr_save_id_i;
  input csr_restore_mret_i;
  input csr_restore_dret_i;
  input csr_save_cause_i;
  input instr_new_id_i;
  input instr_ret_i;
  input instr_ret_compressed_i;
  input imiss_i;
  input pc_set_i;
  input jump_i;
  input branch_i;
  input branch_taken_i;
  input mem_load_i;
  input mem_store_i;
  input lsu_busy_i;
  output m_irq_enable_o;
  output debug_single_step_o;
  output debug_ebreakm_o;
  output illegal_csr_insn_o;
  wire [31:0] csr_rdata_o,mcountinhibit,csr_wdata_int,mscratch_d,mepc_d,mtval_d,dcsr_d,depc_d,
  dscratch0_d,dscratch1_d,mhpmcounter_we,mhpmcounterh_we;
  wire illegal_csr_insn_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,
  N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,
  N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,
  N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,
  N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,
  N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,
  N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,
  N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,
  N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,
  N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,
  N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
  N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,csr_wreq,
  illegal_csr_write,illegal_csr,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,
  N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,
  N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,
  N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,
  N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,
  N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,
  N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,
  N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,
  N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,
  N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,
  N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,
  N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,
  N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,csr_we_int,
  mstatus_d_mie_,mstatus_d_mpie_,mcountinhibit_we,N407,N408,N409,N410,N411,N412,N413,
  N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,
  N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,
  N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,
  N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,
  N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,
  N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
  N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,
  N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,
  N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,
  N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
  N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,
  N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,
  N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,
  N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,
  N638,N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,
  N654,N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,
  N670,N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,
  N686,N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,
  N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,
  N718,N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
  N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,
  N750,N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,
  N766,N767,N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,
  N782,N783,N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,
  N798,N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,
  N814,N815,N816,N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,
  N830,N831,N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,
  N846,N847,N848,N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,
  N862,N863,N864,N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,
  N878,N879,N880,N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,
  N894,N895,N896,N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,
  N910,N911,N912,N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,
  N926,N927,N928,N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,
  N942,N943,N944,N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,
  N958,N959,N960,N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,
  N974,N975,N976,N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,
  N990,N991,N992,N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,
  N1005,N1006,N1007,N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,
  N1018,N1019,N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,
  N1032,N1033,N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,
  N1045,N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,
  N1058,N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,
  N1072,N1073,N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,
  N1085,N1086,N1087,N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,
  N1098,N1099,N1100,N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,
  N1112,N1113,N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,
  N1125,N1126,N1127,N1128,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,
  N1138,N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,
  N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,
  N1165,N1166,N1167,N1168,N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,
  N1178,N1179,N1180,N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,
  N1192,N1193,N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,
  N1205,N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,
  N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,
  N1232,N1233,N1234,N1235,N1236,N1237,N1238,N1239,mcountinhibit_d_0,N1240,N1241,
  N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,N1251,N1252,N1253,N1254,
  N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,
  N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281,
  N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,N1291,N1292,N1293,N1294,
  N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,
  N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,N1318,N1319,N1320,N1321,
  N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,N1331,N1332,N1333,N1334,
  N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,
  N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,
  N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,N1371,N1372,N1373,N1374,
  N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,
  N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,
  N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,N1411,N1412,N1413,N1414,
  N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,
  N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441,
  N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,N1451,N1452,N1453,N1454,
  N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,
  N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,
  N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,N1491,N1492,N1493,N1494,
  N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,
  N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,N1518,N1519,N1520,N1521,
  N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534,
  N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,
  N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561,
  N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,
  N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,
  N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1601,
  N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,N1611,N1612,N1613,N1614,
  N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624,N1625,N1626,N1627,N1628,
  N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,N1638,N1639,N1640,N1641,
  N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,N1651,N1652,N1653,N1654,
  N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,N1665,N1666,N1667,N1668,
  N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1681,
  N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,N1691,N1692,N1693,N1694,
  N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708,
  N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,N1718,N1719,N1720,N1721,
  N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730,N1731,N1732,N1733,N1734,
  N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744,N1745,N1746,N1747,N1748,
  N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757,N1758,N1759,N1760,N1761,
  N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1770,N1771,N1772,N1773,N1774,
  N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,N1784,N1785,N1786,N1787,N1788,
  N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1800,N1801,
  N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,N1810,N1811,N1812,N1813,N1814,
  N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1828,
  N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,N1838,N1839,N1840,N1841,
  N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,N1851,N1852,N1853,N1854,
  N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868,
  N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,N1878,N1879,N1880,N1881,
  N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,N1890,N1891,N1892,N1893,N1894,
  N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,N1904,N1905,N1906,N1907,N1908,
  N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,N1918,N1919,N1920,N1921,
  N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930,N1931,N1932,N1933,N1934,
  N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,N1945,N1946,N1947,N1948,
  N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,N1957,N1958,N1959,N1960,N1961,
  N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,N1970,N1971,N1972,N1973,N1974,
  N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,N1984,N1985,N1986,N1987,N1988,
  N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,N1998,N1999,N2000,N2001,
  N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,N2010,N2011,N2012,N2013,N2014,
  N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2028,
  N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,N2038,N2039,N2040,N2041,
  N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049,N2050,N2051,N2052,N2053,N2054,
  N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062,N2063,N2064,N2065,N2066,N2067,N2068,
  N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,N2077,N2078,N2079,N2080,N2081,
  N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2089,N2090,N2091,N2092,N2093,N2094,
  N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102,N2103,N2104,N2105,N2106,N2107,N2108,
  N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116,N2117,N2118,N2119,N2120,N2121,
  N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2129,N2130,N2131,N2132,N2133,N2134,
  N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148,
  N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156,N2157,N2158,N2159,N2160,N2161,
  N2162,N2163,N2164,N2165,N2166,N2167,N2168,N2169,N2170,N2171,N2172,N2173,N2174,
  N2175,N2176,N2177,N2178,N2179,N2180,N2181,N2182,N2183,N2184,N2185,N2186,N2187,N2188,
  N2189,N2190,N2191,N2192,N2193,N2194,N2195,N2196,N2197,N2198,N2199,N2200,N2201,
  N2202,N2203,N2204,N2205,N2206,N2207,N2208,N2209,N2210,N2211,N2212,N2213,N2214,
  N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222,N2223,N2224,N2225,N2226,N2227,N2228,
  N2229,N2230,N2231,N2232,N2233,N2234,N2235,N2236,N2237,N2238,N2239,N2240,N2241,
  N2242,N2243,N2244,N2245,N2246,N2247,N2248,N2249,N2250,N2251,N2252,N2253,N2254,
  N2255,N2256,N2257,N2258,N2259,N2260,N2261,N2262,N2263,N2264,N2265,N2266,N2267,N2268,
  N2269,N2270,N2271,N2272,N2273,N2274,N2275,N2276,N2277,N2278,N2279,N2280,N2281,
  N2282,N2283,N2284,N2285,N2286,N2287,N2288,N2289,N2290,N2291,N2292,N2293,N2294,
  N2295,N2296,N2297,N2298,N2299,N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,
  N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,N2318,N2319,N2320,N2321,
  N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,N2331,N2332,N2333,N2334,
  N2335,N2336,N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,N2345,N2346,N2347,N2348,
  N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,N2357,N2358,N2359,N2360,N2361,
  N2362,N2363,N2364,N2365,N2366,N2367,N2368,N2369,N2370,N2371,N2372,N2373,N2374,
  N2375,N2376,N2377,N2378,N2379,N2380,N2381,N2382,N2383,N2384,N2385,N2386,N2387,N2388,
  N2389,N2390,N2391,N2392,N2393,N2394,N2395,N2396,N2397,N2398,N2399,N2400,N2401,
  N2402,N2403,N2404,N2405,N2406,N2407,N2408,N2409,N2410,N2411,N2412,N2413,N2414,
  N2415,N2416,N2417,N2418,N2419,N2420,N2421,N2422,N2423,N2424,N2425,N2426,N2427,N2428,
  N2429,N2430,N2431,N2432,N2433,N2434,N2435,N2436,N2437,N2438,N2439,N2440,N2441,
  N2442,N2443,N2444,N2445,N2446,N2447,N2448,N2449,N2450,N2451,N2452,N2453,N2454,
  N2455,N2456,N2457,N2458,N2459,N2460,N2461,N2462,N2463,N2464,N2465,N2466,N2467,N2468,
  N2469,N2470,N2471,N2472,N2473,N2474,N2475,N2476,N2477,N2478,N2479,N2480,N2481,
  N2482,N2483,N2484,N2485,N2486,N2487,N2488,N2489,N2490,N2491,N2492,N2493,N2494,
  N2495,N2496,N2497,N2498,N2499,N2500,N2501,N2502,N2503,N2504,N2505,N2506,N2507,N2508,
  N2509,N2510,N2511,N2512,N2513,N2514,N2515,N2516,N2517,N2518,N2519,N2520,N2521,
  N2522,N2523,N2524,N2525,N2526,N2527,N2528,N2529,N2530,N2531,N2532,N2533,N2534,
  N2535,N2536,N2537,N2538,N2539,N2540,N2541,N2542,N2543,N2544,N2545,N2546,N2547,N2548,
  N2549,N2550,N2551,N2552,N2553,N2554,N2555,N2556,N2557,N2558,N2559,N2560,N2561,
  N2562,N2563,N2564,N2565,N2566,N2567,N2568,N2569,N2570,N2571,N2572,N2573,N2574,
  N2575,N2576,N2577,N2578,N2579,N2580,N2581,N2582,N2583,N2584,N2585,N2586,N2587,N2588,
  N2589,N2590,N2591,N2592,N2593,N2594,N2595,N2596,N2597,N2598,N2599,N2600,N2601,
  N2602,N2603,N2604,N2605,N2606,N2607,N2608,N2609,N2610,N2611,N2612,N2613,N2614,
  N2615,N2616,N2617,N2618,N2619,N2620,N2621,N2622,N2623,N2624,N2625,N2626,N2627,N2628,
  N2629,N2630,N2631,N2632,N2633,N2634,N2635,N2636,N2637,N2638,N2639,N2640,N2641,
  N2642,N2643,N2644,N2645,N2646,N2647,N2648,N2649,N2650,N2651,N2652,N2653,N2654,
  N2655,N2656,N2657,N2658,N2659,N2660,N2661,N2662,N2663,N2664,N2665,N2666,N2667,N2668,
  N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2677,N2678,N2679,N2680,N2681,
  N2682,N2683,N2684,N2685,N2686,N2687,N2688,N2689,N2690,N2691,N2692,N2693,N2694,
  N2695,N2696,N2697,N2698,N2699,N2700,N2701,N2702,N2703,N2704,N2705,N2706,N2707,N2708,
  N2709,N2710,N2711,N2712,N2713,N2714,N2715,N2716,N2717,N2718,N2719,N2720,N2721,
  N2722,N2723,N2724,N2725,N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,
  N2735,N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,N2746,N2747,N2748,
  N2749,N2750,N2751,N2752,N2753,N2754,N2755,N2756,N2757,N2758,N2759,N2760,N2761,
  N2762,N2763,N2764,N2765,N2766,N2767,N2768,N2769,N2770,N2771,N2772,N2773,N2774,
  N2775,N2776,N2777,N2778,N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2788,
  N2789,N2790,N2791,N2792,N2793,N2794,N2795,N2796,N2797,N2798,N2799,N2800,N2801,
  N2802,N2803,N2804,N2805,N2806,N2807,N2808,N2809,N2810,N2811,N2812,N2813,N2814,
  N2815,N2816,N2817,N2818,N2819,N2820,N2821,N2822,N2823,N2824,N2825,N2826,N2827,N2828,
  N2829,N2830,N2831,N2832,N2833,N2834,N2835,N2836,N2837,N2838,N2839,N2840,N2841,
  N2842,N2843,N2844,N2845,N2846,N2847,N2848,N2849,N2850,N2851,N2852,N2853,N2854,
  N2855,N2856,N2857,N2858,N2859,N2860,N2861,N2862,N2863,N2864,N2865,N2866,N2867,N2868,
  N2869,N2870,N2871,N2872,N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,
  N2882,N2883,N2884,N2885,N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2893,N2894,
  N2895,N2896,N2897,N2898,N2899,N2900,N2901,N2902,N2903,N2904,N2905,N2906,N2907,N2908,
  N2909,N2910,N2911,N2912,N2913,N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,
  N2922,N2923,N2924,N2925,N2926,N2927,N2928,N2929,N2930,N2931,N2932,N2933,N2934,
  N2935,N2936,N2937,N2938,N2939,N2940,N2941,N2942,N2943,N2944,N2945,N2946,N2947,N2948,
  N2949,N2950,N2951,N2952,N2953,N2954,N2955,N2956,N2957,N2958,N2959,N2960,N2961,
  N2962,N2963,N2964,N2965,N2966,N2967,N2968,N2969,N2970,N2971,N2972,N2973,N2974,
  N2975,N2976,N2977,N2978,N2979,N2980,N2981,N2982,N2983,N2984,N2985,N2986,N2987,N2988,
  N2989,N2990,N2991,N2992,N2993,N2994,N2995,N2996,N2997,N2998,N2999,N3000,N3001,
  N3002,N3003,N3004,N3005,N3006,N3007,N3008,N3009,N3010,N3011,N3012,N3013,N3014,
  N3015,N3016,N3017,N3018,N3019,N3020,N3021,N3022,N3023,N3024,N3025,N3026,N3027,N3028,
  N3029,N3030,N3031,N3032,N3033,N3034,N3035,N3036,N3037,N3038,N3039,N3040,N3041,
  N3042,N3043,N3044,N3045,N3046,N3047,N3048,N3049,N3050,N3051,N3052,N3053,N3054,
  N3055,N3056,N3057,N3058,N3059,N3060,N3061,N3062,N3063,N3064,N3065,N3066,N3067,N3068,
  N3069,N3070,N3071,N3072,N3073,N3074,N3075,N3076,N3077,N3078,N3079,N3080,N3081,
  N3082,N3083,N3084,N3085,N3086,N3087,N3088,N3089,N3090,N3091,N3092,N3093,N3094,
  N3095,N3096,N3097,N3098,N3099,N3100,N3101,N3102,N3103,N3104,N3105,N3106,N3107,N3108,
  N3109,N3110,N3111,N3112,N3113,N3114,N3115,N3116,N3117,N3118,N3119,N3120,N3121,
  N3122,N3123,N3124,N3125,N3126,N3127,N3128,N3129,N3130,N3131,N3132,N3133,N3134,
  N3135,N3136,N3137,N3138,N3139,N3140,N3141,N3142,N3143,N3144,N3145,N3146,N3147,N3148,
  N3149,N3150,N3151,N3152,N3153,N3154,N3155,N3156,N3157,N3158,N3159,N3160,N3161,
  N3162,N3163,N3164,N3165,N3166,N3167,N3168,N3169,N3170,N3171,N3172,N3173,N3174,
  N3175,N3176,N3177,N3178,N3179,N3180,N3181,N3182,N3183,N3184,N3185,N3186,N3187,N3188,
  N3189,N3190,N3191,N3192,N3193,N3194,N3195,N3196,N3197,N3198,N3199,N3200,N3201,
  N3202,N3203,N3204,N3205,N3206,N3207,N3208,N3209,N3210,N3211,N3212,N3213,N3214,
  N3215,N3216,N3217,N3218,N3219,N3220,N3221,N3222,N3223,N3224,N3225,N3226,N3227,N3228,
  N3229,N3230,N3231,N3232,N3233,N3234,N3235,N3236,N3237,N3238,N3239,N3240,N3241,
  N3242,N3243,N3244,N3245,N3246,N3247,N3248,N3249,N3250,N3251,N3252,N3253,N3254,
  N3255,N3256,N3257,N3258,N3259,N3260,N3261,N3262,N3263,N3264,N3265,N3266,N3267,N3268,
  N3269,N3270,N3271,N3272,N3273,N3274,N3275,N3276,N3277,N3278,N3279,N3280,N3281,
  N3282,N3283,N3284,N3285,N3286,N3287,N3288,N3289,N3290,N3291,N3292,N3293,N3294,
  N3295,N3296,N3297,N3298,N3299,N3300,N3301,N3302,N3303,N3304,N3305,N3306,N3307,N3308,
  N3309,N3310,N3311,N3312,N3313,N3314,N3315,N3316,N3317,N3318,N3319,N3320,N3321,
  N3322,N3323,N3324,N3325,N3326,N3327,N3328,N3329,N3330,N3331,N3332,N3333,N3334,
  N3335,N3336,N3337,N3338,N3339,N3340,N3341,N3342,N3343,N3344,N3345,N3346,N3347,N3348,
  N3349,N3350,N3351,N3352,N3353,N3354,N3355,N3356,N3357,N3358,N3359,N3360,N3361,
  N3362,N3363,N3364,N3365,N3366,N3367,N3368,N3369,N3370,N3371,N3372,N3373,N3374,
  N3375,N3376,N3377,N3378,N3379,N3380,N3381,N3382,N3383,N3384,N3385,N3386,N3387,N3388,
  N3389,N3390,N3391,N3392,N3393,N3394,N3395,N3396,N3397,N3398,N3399,N3400,N3401,
  N3402,N3403,N3404,N3405,N3406,N3407,N3408,N3409,N3410,N3411,N3412,N3413,N3414,
  N3415,N3416,N3417,N3418,N3419,N3420,N3421,N3422,N3423,N3424,N3425,N3426,N3427,N3428,
  N3429,N3430,N3431,N3432,N3433,N3434,N3435,N3436,N3437,N3438,N3439,N3440,N3441,
  N3442,N3443,N3444,N3445,N3446,N3447,N3448,N3449,N3450,N3451,N3452,N3453,N3454,
  N3455,N3456,N3457,N3458,N3459,N3460,N3461,N3462,N3463,N3464,N3465,N3466,N3467,N3468,
  N3469,N3470,N3471,N3472,N3473,N3474,N3475,N3476,N3477,N3478,N3479,N3480,N3481,
  N3482,N3483,N3484,N3485,N3486,N3487,N3488,N3489,N3490,N3491,N3492,N3493,N3494,
  N3495,N3496,N3497,N3498,N3499,N3500,N3501,N3502,N3503,N3504,N3505,N3506,N3507,N3508,
  N3509,N3510,N3511,N3512,N3513,N3514,N3515,N3516,N3517,N3518,N3519,N3520,N3521,
  N3522,N3523,N3524,N3525,N3526,N3527,N3528,N3529,N3530,N3531,N3532,N3533,N3534,
  N3535,N3536,N3537,N3538,N3539,N3540,N3541,N3542,N3543,N3544,N3545,N3546,N3547,N3548,
  N3549,N3550,N3551,N3552,N3553,N3554,N3555,N3556,N3557,N3558,N3559,N3560,N3561,
  N3562,N3563,N3564,N3565,N3566,N3567,N3568,N3569,N3570,N3571,N3572,N3573,N3574,
  N3575,N3576,N3577,N3578,N3579,N3580,N3581,N3582,N3583,N3584,N3585,N3586,N3587,N3588,
  N3589,N3590,N3591,N3592,N3593,N3594,N3595,N3596,N3597,N3598,N3599,N3600,N3601,
  N3602,N3603,N3604,N3605,N3606,N3607,N3608,N3609,N3610,N3611,N3612,N3613,N3614,
  N3615,N3616,N3617,N3618,N3619,N3620,N3621,N3622,N3623,N3624,N3625,N3626,N3627,N3628,
  N3629,N3630,N3631,N3632,N3633,N3634,N3635,N3636,N3637,N3638,N3639,N3640,N3641,
  N3642,N3643,N3644,N3645,N3646,N3647,N3648,N3649,N3650,N3651,N3652,N3653,N3654,
  N3655,N3656,N3657,N3658,N3659,N3660,N3661,N3662,N3663,N3664,N3665,N3666,N3667,N3668,
  N3669,N3670,N3671,N3672,N3673,N3674,N3675,N3676,N3677,N3678,N3679,N3680,N3681,
  N3682,N3683,N3684,N3685,N3686,N3687,N3688,N3689,N3690,N3691,N3692,N3693,N3694,
  N3695,N3696,N3697,N3698,N3699,N3700,N3701,N3702,N3703,N3704,N3705,N3706,N3707,N3708,
  N3709,N3710,N3711,N3712,N3713,N3714,N3715,N3716,N3717,N3718,N3719,N3720,N3721,
  N3722,N3723,N3724,N3725,N3726,N3727,N3728,N3729,N3730,N3731,N3732,N3733,N3734,
  N3735,N3736,N3737,N3738,N3739,N3740,N3741,N3742,N3743,N3744,N3745,N3746,N3747,N3748,
  N3749,N3750,N3751,N3752,N3753,N3754,N3755,N3756,N3757,N3758,N3759,N3760,N3761,
  N3762,N3763,N3764,N3765,N3766,N3767,N3768,N3769,N3770,N3771,N3772,N3773,N3774,
  N3775,N3776,N3777,N3778,N3779,N3780,N3781,N3782,N3783,N3784,N3785,N3786,N3787,N3788,
  N3789,N3790,N3791,N3792,N3793,N3794,N3795,N3796,N3797,N3798,N3799,N3800,N3801,
  N3802,N3803,N3804,N3805,N3806,N3807,N3808,N3809,N3810,N3811,N3812,N3813,N3814,
  N3815,N3816,N3817,N3818,N3819,N3820,N3821,N3822,N3823,N3824,N3825,N3826,N3827,N3828,
  N3829,N3830,N3831,N3832,N3833,N3834,N3835,N3836,N3837,N3838,N3839,N3840,N3841,
  N3842,N3843,N3844,N3845,N3846,N3847,N3848,N3849,N3850,N3851,N3852,N3853,N3854,
  N3855,N3856,N3857,N3858,N3859,N3860,N3861,N3862,N3863,N3864,N3865,N3866,N3867,N3868,
  N3869,N3870,N3871,N3872,N3873,N3874,N3875,N3876,N3877,N3878,N3879,N3880,N3881,
  N3882,N3883,N3884,N3885,N3886,N3887,N3888,N3889,N3890,N3891,N3892,N3893,N3894,
  N3895,N3896,N3897,N3898,N3899,N3900,N3901,N3902,N3903,N3904,N3905,N3906,N3907,N3908,
  N3909,N3910,N3911,N3912,N3913,N3914,N3915,N3916,N3917,N3918,N3919,N3920,N3921,
  N3922,N3923,N3924,N3925,N3926,N3927,N3928,N3929,N3930,N3931,N3932,N3933,N3934,
  N3935,N3936,N3937,N3938,N3939,N3940,N3941,N3942,N3943,N3944,N3945,N3946,N3947,N3948,
  N3949,N3950,N3951,N3952,N3953,N3954,N3955,N3956,N3957,N3958,N3959,N3960,N3961,
  N3962,N3963,N3964,N3965,N3966,N3967,N3968,N3969,N3970,N3971,N3972,N3973,N3974,
  N3975,N3976,N3977,N3978,N3979,N3980,N3981,N3982,N3983,N3984,N3985,N3986,N3987,N3988,
  N3989,N3990,N3991,N3992,N3993,N3994,N3995,N3996,N3997,N3998,N3999,N4000,N4001,
  N4002,N4003,N4004,N4005,N4006,N4007,N4008,N4009,N4010,N4011,N4012,N4013,N4014,
  N4015,N4016,N4017,N4018,N4019,N4020,N4021,N4022,N4023,N4024,N4025,N4026,N4027,N4028,
  N4029,N4030,N4031,N4032,N4033,N4034,N4035,N4036,N4037,N4038,N4039,N4040,N4041,
  N4042,N4043,N4044,N4045,N4046,N4047,N4048,N4049,N4050,N4051,N4052,N4053,N4054,
  N4055,N4056,N4057,N4058,N4059,N4060,N4061,N4062,N4063,N4064,N4065,N4066,N4067,N4068,
  N4069,N4070,N4071,N4072,N4073,N4074,N4075,N4076,N4077,N4078,N4079,N4080,N4081,
  N4082,N4083,N4084,N4085,N4086,N4087,N4088,N4089,N4090,N4091,N4092,N4093,N4094,
  N4095,N4096,N4097,N4098,N4099,N4100,N4101,N4102,N4103,N4104,N4105,N4106,N4107,N4108,
  N4109,N4110,N4111,N4112,N4113,N4114,N4115,N4116,N4117,N4118,N4119,N4120,N4121,
  N4122,N4123,N4124,N4125,N4126,N4127,N4128,N4129,N4130,N4131,N4132,N4133,N4134,
  N4135,N4136,N4137,N4138,N4139,N4140,N4141,N4142,N4143,N4144,N4145,N4146,N4147,N4148,
  N4149,N4150,N4151,N4152,N4153,N4154,N4155,N4156,N4157,N4158,N4159,N4160,N4161,
  N4162,N4163,N4164,N4165,N4166,N4167,N4168,N4169,N4170,N4171,N4172,N4173,N4174,
  N4175,N4176,N4177,N4178,N4179,N4180,N4181,N4182,N4183,N4184,N4185,N4186,N4187,N4188,
  N4189,N4190,N4191,N4192,N4193,N4194,N4195,N4196,N4197,N4198,N4199,N4200,N4201,
  N4202,N4203,N4204,N4205,N4206,N4207,N4208,N4209,N4210,N4211,N4212,N4213,N4214,
  N4215,N4216,N4217,N4218,N4219,N4220,N4221,N4222,N4223,N4224,N4225,N4226,N4227,N4228,
  N4229,N4230,N4231,N4232,N4233,N4234,N4235,N4236,N4237,N4238,N4239,N4240,N4241,
  N4242,N4243,N4244,N4245,N4246,N4247,N4248,N4249,N4250,N4251,N4252,N4253,N4254,
  N4255,N4256,N4257,N4258,N4259,N4260,N4261,N4262,N4263,N4264,N4265,N4266,N4267,N4268,
  N4269,N4270,N4271,N4272,N4273,N4274,N4275,N4276,N4277,N4278,N4279,N4280,N4281,
  N4282,N4283,N4284,N4285,N4286,N4287,N4288,N4289,N4290,N4291,N4292,N4293,N4294,
  N4295,N4296,N4297,N4298,N4299,N4300,N4301,N4302,N4303,N4304,N4305,N4306,N4307,N4308,
  N4309,N4310,N4311,N4312,N4313,N4314,N4315,N4316,N4317,N4318,N4319,N4320,N4321,
  N4322,N4323,N4324,N4325,N4326,N4327,N4328,N4329,N4330,N4331,N4332,N4333,N4334,
  N4335,N4336,N4337,N4338,N4339,N4340,N4341,N4342,N4343,N4344,N4345,N4346,N4347,N4348,
  N4349,N4350,N4351,N4352,N4353,N4354,N4355,N4356,N4357,N4358,N4359,N4360,N4361,
  N4362,N4363,N4364,N4365,N4366,N4367,N4368,N4369,N4370,N4371,N4372,N4373,N4374,
  N4375,N4376,N4377,N4378,N4379,N4380,N4381,N4382,N4383,N4384,N4385,N4386,N4387,N4388,
  N4389,N4390,N4391,N4392,N4393,N4394,N4395,N4396,N4397,N4398,N4399,N4400,N4401,
  N4402,N4403,N4404,N4405,N4406,N4407,N4408,N4409,N4410,N4411,N4412,N4413,N4414,
  N4415,N4416,N4417,N4418,N4419,N4420,N4421,N4422,N4423,N4424,N4425,N4426,N4427,N4428,
  N4429,N4430,N4431,N4432,N4433,N4434,N4435,N4436,N4437,N4438,N4439,N4440,N4441,
  N4442,N4443,N4444,N4445,N4446,N4447,N4448,N4449,N4450,N4451,N4452,N4453,N4454,
  N4455,N4456,N4457,N4458,N4459,N4460,N4461,N4462,N4463,N4464,N4465,N4466,N4467,N4468,
  N4469,N4470,N4471,N4472,N4473,N4474,N4475,N4476,N4477,N4478,N4479,N4480,N4481,
  N4482,N4483,N4484,N4485,N4486,N4487,N4488,N4489,N4490,N4491,N4492,N4493,N4494,
  N4495,N4496,N4497,N4498,N4499,N4500,N4501,N4502,N4503,N4504,N4505,N4506,N4507,N4508,
  N4509,N4510,N4511,N4512,N4513,N4514,N4515,N4516,N4517,N4518,N4519,N4520,N4521,
  N4522,N4523,N4524,N4525,N4526,N4527,N4528,N4529,N4530,N4531,N4532,N4533,N4534,
  N4535,N4536,N4537,N4538,N4539,N4540,N4541,N4542,N4543,N4544,N4545,N4546,N4547,N4548,
  N4549,N4550,N4551,N4552,N4553,N4554,N4555,N4556,N4557,N4558,N4559,N4560,N4561,
  N4562,N4563,N4564,N4565,N4566,N4567,N4568,N4569,N4570,N4571,N4572,N4573,N4574,
  N4575,N4576,N4577,N4578,N4579,N4580,N4581,N4582,N4583,N4584,N4585,N4586,N4587,N4588,
  N4589,N4590,N4591,N4592,N4593,N4594,N4595,N4596,N4597,N4598,N4599,N4600,N4601,
  N4602,N4603,N4604,N4605,N4606,N4607,N4608,N4609,N4610,N4611,N4612,N4613,N4614,
  N4615,N4616,N4617,N4618,N4619,N4620,N4621,N4622,N4623,N4624,N4625,N4626,N4627,N4628,
  N4629,N4630,N4631,N4632,N4633,N4634,N4635,N4636,N4637,N4638,N4639,N4640,N4641,
  N4642,N4643,N4644,N4645,N4646,N4647,N4648,N4649,N4650,N4651,N4652,N4653,N4654,
  N4655,N4656,N4657,N4658,N4659,N4660,N4661,N4662,N4663,N4664,N4665,N4666,N4667,N4668,
  N4669,N4670,N4671,N4672,N4673,N4674,N4675,N4676,N4677,N4678,N4679,N4680,N4681,
  N4682,N4683,N4684,N4685,N4686,N4687,N4688,N4689,N4690,N4691,N4692,N4693,N4694,
  N4695,N4696,N4697,N4698,N4699,N4700,N4701,N4702,N4703,N4704,N4705,N4706,N4707,N4708,
  N4709,N4710,N4711,N4712,N4713,N4714,N4715,N4716,N4717,N4718,N4719,N4720,N4721,
  N4722,N4723,N4724,N4725,N4726,N4727,N4728,N4729,N4730,N4731,N4732,N4733,N4734,
  N4735,N4736,N4737,N4738,N4739,N4740,N4741,N4742,N4743,N4744,N4745,N4746,N4747,N4748,
  N4749,N4750,N4751,N4752,N4753,N4754,N4755,N4756,N4757,N4758,N4759,N4760,N4761,
  N4762,N4763,N4764,N4765,N4766,N4767,N4768,N4769,N4770,N4771,N4772,N4773,N4774,
  N4775,N4776,N4777,N4778,N4779,N4780,N4781,N4782,N4783,N4784,N4785,N4786,N4787,N4788,
  N4789,N4790,N4791,N4792,N4793,N4794,N4795,N4796,N4797,N4798,N4799,N4800,N4801,
  N4802,N4803,N4804,N4805,N4806,N4807,N4808,N4809,N4810,N4811,N4812,N4813,N4814,
  N4815,N4816,N4817,N4818,N4819,N4820,N4821,N4822,N4823,N4824,N4825,N4826,N4827,N4828,
  N4829,N4830,N4831,N4832,N4833,N4834,N4835,N4836,N4837,N4838,N4839,N4840,N4841,
  N4842,N4843,N4844,N4845,N4846,N4847,N4848,N4849,N4850,N4851,N4852,N4853,N4854,
  N4855,N4856,N4857,N4858,N4859,N4860,N4861,N4862,N4863,N4864,N4865,N4866,N4867,N4868,
  N4869,N4870,N4871,N4872,N4873,N4874,N4875,N4876,N4877,N4878,N4879,N4880,N4881,
  N4882,N4883,N4884,N4885,N4886,N4887,N4888,N4889,N4890,N4891,N4892,N4893,N4894,
  N4895,N4896,N4897,N4898,N4899,N4900,N4901,N4902,N4903,N4904,N4905,N4906,N4907,N4908,
  N4909,N4910,N4911,N4912,N4913,N4914,N4915,N4916,N4917,N4918,N4919,N4920,N4921,
  N4922,N4923,N4924,N4925,N4926,N4927,N4928,N4929,N4930,N4931,N4932,N4933,N4934,
  N4935,N4936,N4937,N4938,N4939,N4940,N4941,N4942,N4943,N4944,N4945,N4946,N4947,N4948,
  N4949,N4950,N4951,N4952,N4953,N4954,N4955,N4956,N4957,N4958,N4959,N4960,N4961,
  N4962,N4963,N4964,N4965,N4966,N4967,N4968,N4969,N4970,N4971,N4972,N4973,N4974,
  N4975,N4976,N4977,N4978,N4979,N4980,N4981,N4982,N4983,N4984,N4985,N4986,N4987,N4988,
  N4989,N4990,N4991,N4992,N4993,N4994,N4995,N4996,N4997,N4998,N4999,N5000,N5001,
  N5002,N5003,N5004,N5005,N5006,N5007,N5008,N5009,N5010,N5011,N5012,N5013,N5014,
  N5015,N5016,N5017,N5018,N5019,N5020,N5021,N5022,N5023,N5024,N5025,N5026,N5027,N5028,
  N5029,N5030,N5031,N5032,N5033,N5034,N5035,N5036,N5037,N5038,N5039,N5040,N5041,
  N5042,N5043,N5044,N5045,N5046,N5047,N5048,N5049,N5050,N5051,N5052,N5053,N5054,
  N5055,N5056,N5057,N5058,N5059,N5060,N5061,N5062,N5063,N5064,N5065,N5066,N5067,N5068,
  N5069,N5070,N5071,N5072,N5073,N5074,N5075,N5076,N5077,N5078,N5079,N5080,N5081,
  N5082,N5083,N5084,N5085,N5086,N5087,N5088,N5089,N5090,N5091,N5092,N5093,N5094,
  N5095,N5096,N5097,N5098,N5099,N5100,N5101,N5102,N5103,N5104,N5105,N5106,N5107,N5108,
  N5109,N5110,N5111,N5112,N5113,N5114,N5115,N5116,N5117,N5118,N5119,N5120,N5121,
  N5122,N5123,N5124,N5125,N5126,N5127,N5128,N5129,N5130,N5131,N5132,N5133,N5134,
  N5135,N5136,N5137,N5138,N5139,N5140,N5141,N5142,N5143,N5144,N5145,N5146,N5147,N5148,
  N5149,N5150,N5151,N5152,N5153,N5154,N5155,N5156,N5157,N5158,N5159,N5160,N5161,
  N5162,N5163,N5164,N5165,N5166,N5167,N5168,N5169,N5170,N5171,N5172,N5173,N5174,
  N5175,N5176,N5177,N5178,N5179,N5180,N5181,N5182,N5183,N5184,N5185,N5186,N5187,N5188,
  N5189,N5190,N5191,N5192,N5193,N5194,N5195,N5196,N5197,N5198,N5199,N5200,N5201,
  N5202,N5203,N5204,N5205,N5206,N5207,N5208,N5209,N5210,N5211,N5212,N5213,N5214,
  N5215,N5216,N5217,N5218,N5219,N5220,N5221,N5222,N5223,N5224,N5225,N5226,N5227,N5228,
  N5229,N5230,N5231,N5232,N5233,N5234,N5235,N5236,N5237,N5238,N5239,N5240,N5241,
  N5242,N5243,N5244,N5245,N5246,N5247,N5248,N5249,N5250,N5251,N5252,N5253,N5254,
  N5255,N5256,N5257,N5258,N5259,N5260,N5261,N5262,N5263,N5264,N5265,N5266,N5267,N5268,
  N5269,N5270,N5271,N5272,N5273,N5274,N5275,N5276,N5277,N5278,N5279,N5280,N5281,
  N5282,N5283,N5284,N5285,N5286,N5287,N5288,N5289,N5290,N5291,N5292,N5293,N5294,
  N5295,N5296,N5297,N5298,N5299,N5300,N5301,N5302,N5303,N5304,N5305,N5306,N5307,N5308,
  N5309,N5310,N5311,N5312,N5313,N5314,N5315,N5316,N5317,N5318,N5319,N5320,N5321,
  N5322,N5323,N5324,N5325,N5326,N5327,N5328,N5329,N5330,N5331,N5332,N5333,N5334,
  N5335,N5336,N5337,N5338,N5339,N5340,N5341,N5342,N5343,N5344,N5345,N5346,N5347,N5348,
  N5349,N5350,N5351,N5352,N5353,N5354,N5355,N5356,N5357,N5358,N5359,N5360,N5361,
  N5362,N5363,N5364,N5365,N5366,N5367,N5368,N5369,N5370,N5371,N5372,N5373,N5374,
  N5375,N5376,N5377,N5378,N5379,N5380,N5381,N5382,N5383,N5384,N5385,N5386,N5387,N5388,
  N5389,N5390,N5391,N5392,N5393,N5394,N5395,N5396,N5397,N5398,N5399,N5400,N5401,
  N5402,N5403,N5404,N5405,N5406,N5407,N5408,N5409,N5410,N5411,N5412,N5413,N5414,
  N5415,N5416,N5417,N5418,N5419,N5420,N5421,N5422,N5423,N5424,N5425,N5426,N5427,N5428,
  N5429,N5430,N5431,N5432,N5433,N5434,N5435,N5436,N5437,N5438,N5439,N5440,N5441,
  N5442,N5443,N5444,N5445,N5446,N5447,N5448,N5449,N5450,N5451,N5452,N5453,N5454,
  N5455,N5456,N5457,N5458,N5459,N5460,N5461,N5462,N5463,N5464,N5465,N5466,N5467,N5468,
  N5469,N5470,N5471,N5472,N5473,N5474,N5475,N5476,N5477,N5478,N5479,N5480,N5481,
  N5482,N5483,N5484,N5485,N5486,N5487,N5488,N5489,N5490,N5491,N5492,N5493,N5494,
  N5495,N5496,N5497,N5498,N5499,N5500,N5501,N5502,N5503,N5504,N5505,N5506,N5507,N5508,
  N5509,N5510,N5511,N5512,N5513,N5514,N5515,N5516,N5517,N5518,N5519,N5520,N5521,
  N5522,N5523,N5524,N5525,N5526,N5527,N5528,N5529,N5530,N5531,N5532,N5533,N5534,
  N5535,N5536,N5537,N5538,N5539,N5540,N5541,N5542,N5543,N5544,N5545,N5546,N5547,N5548,
  N5549,N5550,N5551,N5552,N5553,N5554,N5555,N5556,N5557,N5558,N5559,N5560,N5561,
  N5562,N5563,N5564,N5565,N5566,N5567,N5568,N5569,N5570,N5571,N5572,N5573,N5574,
  N5575,N5576,N5577,N5578,N5579,N5580,N5581,N5582,N5583,N5584,N5585,N5586,N5587,N5588,
  N5589,N5590,N5591,N5592,N5593,N5594,N5595,N5596,N5597,N5598,N5599,N5600,N5601,
  N5602,N5603,N5604,N5605,N5606,N5607,N5608,N5609,N5610,N5611,N5612,N5613,N5614,
  N5615,N5616,N5617,N5618,N5619,N5620,N5621,N5622,N5623,N5624,N5625,N5626,N5627,N5628,
  N5629,N5630,N5631,N5632,N5633,N5634,N5635,N5636,N5637,N5638,N5639,N5640,N5641,
  N5642,N5643,N5644,N5645,N5646,N5647,N5648,N5649,N5650,N5651,N5652,N5653,N5654,
  N5655,N5656,N5657,N5658,N5659,N5660,N5661,N5662,N5663,N5664,N5665,N5666,N5667,N5668,
  N5669,N5670,N5671,N5672,N5673,N5674,N5675,N5676,N5677,N5678,N5679,N5680,N5681,
  N5682,N5683,N5684,N5685,N5686,N5687,N5688,N5689,N5690,N5691,N5692,N5693,N5694,
  N5695,N5696,N5697,N5698,N5699,N5700,N5701,N5702,N5703,N5704,N5705,N5706,N5707,N5708,
  N5709,N5710,N5711,N5712,N5713,N5714,N5715,N5716,N5717,N5718,N5719,N5720,N5721,
  N5722,N5723,N5724,N5725,N5726,N5727,N5728,N5729,N5730,N5731,N5732,N5733,N5734,
  N5735,N5736,N5737,N5738,N5739,N5740,N5741,N5742,N5743,N5744,N5745,N5746,N5747,N5748,
  N5749,N5750,N5751,N5752,N5753,N5754,N5755,N5756,N5757,N5758,N5759,N5760,N5761,
  N5762,N5763,N5764,N5765,N5766,N5767,N5768,N5769,N5770,N5771,N5772,N5773,N5774,
  N5775,N5776,N5777,N5778,N5779,N5780,N5781,N5782,N5783,N5784,N5785,N5786,N5787,N5788,
  N5789,N5790,N5791,N5792,N5793,N5794,N5795,N5796,N5797,N5798,N5799,N5800,N5801,
  N5802,N5803,N5804,N5805,N5806,N5807,N5808,N5809,N5810,N5811,N5812,N5813,N5814,
  N5815,N5816,N5817,N5818,N5819,N5820,N5821,N5822,N5823,N5824,N5825,N5826,N5827,N5828,
  N5829,N5830,N5831,N5832,N5833,N5834,N5835,N5836,N5837,N5838,N5839,N5840,N5841,
  N5842,N5843,N5844,N5845,N5846,N5847,N5848,N5849,N5850,N5851,N5852,N5853,N5854,
  N5855,N5856,N5857,N5858,N5859,N5860,N5861,N5862,N5863,N5864,N5865,N5866,N5867,N5868,
  N5869,N5870,N5871,N5872,N5873,N5874,N5875,N5876,N5877,N5878,N5879,N5880,N5881,
  N5882,N5883,N5884,N5885,N5886,N5887,N5888,N5889,N5890,N5891,N5892,N5893,N5894,
  N5895,N5896,N5897,N5898,N5899,N5900,N5901,N5902,N5903,N5904,N5905,N5906,N5907,N5908,
  N5909,N5910,N5911,N5912,N5913,N5914,N5915,N5916,N5917,N5918,N5919,N5920,N5921,
  N5922,N5923,N5924,N5925,N5926,N5927,N5928,N5929,N5930,N5931,N5932,N5933,N5934,
  N5935,N5936,N5937,N5938,N5939,N5940,N5941,N5942,N5943,N5944,N5945,N5946,N5947,N5948,
  N5949,N5950,N5951,N5952,N5953,N5954,N5955,N5956,N5957,N5958,N5959,N5960,N5961,
  N5962,N5963,N5964,N5965,N5966,N5967,N5968,N5969,N5970,N5971,N5972,N5973,N5974,
  N5975,N5976,N5977,N5978,N5979,N5980,N5981,N5982,N5983,N5984,N5985,N5986,N5987,N5988,
  N5989,N5990,N5991,N5992,N5993,N5994,N5995,N5996,N5997,N5998,N5999,N6000,N6001,
  N6002,N6003,N6004,N6005,N6006,N6007,N6008,N6009,N6010,N6011,N6012,N6013,N6014,
  N6015,N6016,N6017,N6018,N6019,N6020,N6021,N6022,N6023,N6024,N6025,N6026,N6027,N6028,
  N6029,N6030,N6031,N6032,N6033,N6034,N6035,N6036,N6037,N6038,N6039,N6040,N6041,
  N6042,N6043,N6044,N6045,N6046,N6047,N6048,N6049,N6050,N6051,N6052,N6053,N6054,
  N6055,N6056,N6057,N6058,N6059,N6060,N6061,N6062,N6063,N6064,N6065,N6066,N6067,N6068,
  N6069,N6070,N6071,N6072,N6073,N6074,N6075,N6076,N6077,N6078,N6079,N6080,N6081,
  N6082,N6083,N6084,N6085,N6086,N6087,N6088,N6089,N6090,N6091,N6092,N6093,N6094,
  N6095,N6096,N6097,N6098,N6099,N6100,N6101,N6102,N6103,N6104,N6105,N6106,N6107,N6108,
  N6109,N6110,N6111,N6112,N6113,N6114,N6115,N6116,N6117,N6118,N6119,N6120,N6121,
  N6122,N6123,N6124,N6125,N6126,N6127,N6128,N6129,N6130,N6131,N6132,N6133,N6134,
  N6135,N6136,N6137,N6138,N6139,N6140,N6141,N6142,N6143,N6144,N6145,N6146,N6147,N6148,
  N6149,N6150,N6151,N6152,N6153,N6154,N6155,N6156,N6157,N6158,N6159,N6160,N6161,
  N6162,N6163,N6164,N6165,N6166,N6167,N6168,N6169,N6170,N6171,N6172,N6173,N6174,
  N6175,N6176,N6177,N6178,N6179,N6180,N6181,N6182,N6183,N6184,N6185,N6186,N6187,N6188,
  N6189,N6190,N6191,N6192,N6193,N6194,N6195,N6196,N6197,N6198,N6199,N6200,N6201,
  N6202,N6203,N6204,N6205,N6206,N6207,N6208,N6209,N6210,N6211,N6212,N6213,N6214,
  N6215,N6216,N6217,N6218,N6219,N6220,N6221,N6222,N6223,N6224,N6225,N6226,N6227,N6228,
  N6229,N6230,N6231,N6232,N6233,N6234,N6235,N6236,N6237,N6238,N6239,N6240,N6241,
  N6242,N6243,N6244,N6245,N6246,N6247,N6248,N6249,N6250,N6251,N6252,N6253,N6254,
  N6255,N6256,N6257,N6258,N6259,N6260,N6261,N6262,N6263,N6264,N6265,N6266,N6267,N6268,
  N6269,N6270,N6271,N6272,N6273,N6274,N6275,N6276,N6277,N6278,N6279,N6280,N6281,
  N6282,N6283,N6284,N6285,N6286,N6287,N6288,N6289,N6290,N6291,N6292,N6293,N6294,
  N6295,N6296,N6297,N6298,N6299,N6300,N6301,N6302,N6303,N6304,N6305,N6306,N6307,N6308,
  N6309,N6310,N6311,N6312,N6313,N6314,N6315,N6316,N6317,N6318,N6319,N6320,N6321,
  N6322,N6323,N6324,N6325,N6326,N6327,N6328,N6329,N6330,N6331,N6332,N6333,N6334,
  N6335,N6336,N6337,N6338,N6339,N6340,N6341,N6342,N6343,N6344,N6345,N6346,N6347,N6348,
  N6349,N6350,N6351,N6352,N6353,N6354,N6355,N6356,N6357,N6358,N6359,N6360,N6361,
  N6362,N6363,N6364,N6365,N6366,N6367,N6368,N6369,N6370,N6371,N6372,N6373,N6374,
  N6375,N6376,N6377,N6378,N6379,N6380,N6381,N6382,N6383,N6384,N6385,N6386,N6387,N6388,
  N6389,N6390,N6391,N6392,N6393,N6394,N6395,N6396,N6397,N6398,N6399,N6400,N6401,
  N6402,N6403,N6404,N6405,N6406,N6407,N6408,N6409,N6410,N6411,N6412,N6413,N6414,
  N6415,N6416,N6417,N6418,N6419,N6420,N6421,N6422,N6423,N6424,N6425,N6426,N6427,N6428,
  N6429,N6430,N6431,N6432,N6433,N6434,N6435,N6436,N6437,N6438,N6439,N6440,N6441,
  N6442,N6443,N6444,N6445,N6446,N6447,N6448,N6449,N6450,N6451,N6452,N6453,N6454,
  N6455,N6456,N6457,N6458,N6459,N6460,N6461,N6462,N6463,N6464,N6465,N6466,N6467,N6468,
  N6469,N6470,N6471,N6472,N6473,N6474,N6475,N6476,N6477,N6478,N6479,N6480,N6481,
  N6482,N6483,N6484,N6485,N6486,N6487,N6488,N6489,N6490,N6491,N6492,N6493,N6494,
  N6495,N6496,N6497,N6498,N6499,N6500,N6501,N6502,N6503,N6504,N6505,N6506,N6507,N6508,
  N6509,N6510,N6511,N6512,N6513,N6514,N6515,N6516,N6517,N6518,N6519,N6520,N6521,
  N6522,N6523,N6524,N6525,N6526,N6527,N6528,N6529,N6530,N6531,N6532,N6533,N6534,
  N6535,N6536,N6537,N6538,N6539,N6540,N6541,N6542,N6543,N6544,N6545,N6546,N6547,N6548,
  N6549,N6550,N6551,N6552,N6553,N6554,N6555,N6556,N6557,N6558,N6559,N6560,N6561,
  N6562,N6563,N6564,N6565,N6566,N6567,N6568,N6569,N6570,N6571,N6572,N6573,N6574,
  N6575,N6576,N6577,N6578,N6579,N6580,N6581,N6582,N6583,N6584,N6585,N6586,N6587,N6588,
  N6589,N6590,N6591,N6592,N6593,N6594,N6595,N6596,N6597,N6598,N6599,N6600,N6601,
  N6602,N6603,N6604,N6605,N6606,N6607,N6608,N6609,N6610,N6611,N6612,N6613,N6614,
  N6615,N6616,N6617,N6618,N6619,N6620,N6621,N6622,N6623,N6624,N6625,N6626,N6627,N6628,
  N6629,N6630,N6631,N6632,N6633,N6634,N6635,N6636,N6637,N6638,N6639,N6640,N6641,
  N6642,N6643,N6644,N6645,N6646,N6647,N6648,N6649,N6650,N6651,N6652,N6653,N6654,
  N6655,N6656,N6657,N6658,N6659,N6660,N6661,N6662,N6663,N6664,N6665,N6666,N6667,N6668,
  N6669,N6670,N6671,N6672,N6673,N6674,N6675,N6676,N6677,N6678,N6679,N6680,N6681,
  N6682,N6683,N6684,N6685,N6686,N6687,N6688,N6689,N6690,N6691,N6692,N6693,N6694,
  N6695,N6696,N6697,N6698,N6699,N6700,N6701,N6702,N6703,N6704,N6705,N6706,N6707,N6708,
  N6709,N6710,N6711,N6712,N6713,N6714,N6715,N6716,N6717,N6718,N6719,N6720,N6721,
  N6722,N6723,N6724,N6725,N6726,N6727,N6728,N6729,N6730,N6731,N6732,N6733,N6734,
  N6735,N6736,N6737,N6738,N6739,N6740,N6741,N6742,N6743,N6744,N6745,N6746,N6747,N6748,
  N6749,N6750,N6751,N6752,N6753,N6754,N6755,N6756,N6757,N6758,N6759,N6760,N6761,
  N6762,N6763,N6764,N6765,N6766,N6767,N6768,N6769,N6770,N6771,N6772,N6773,N6774,
  N6775,N6776,N6777,N6778,N6779,N6780,N6781,N6782,N6783,N6784,N6785,N6786,N6787,N6788,
  N6789,N6790,N6791,N6792,N6793,N6794,N6795,N6796,N6797,N6798,N6799,N6800,N6801,
  N6802,N6803,N6804,N6805,N6806,N6807,N6808,N6809,N6810,N6811,N6812,N6813,N6814,
  N6815,N6816,N6817,N6818,N6819,N6820,N6821,N6822,N6823,N6824,N6825,N6826,N6827,N6828,
  N6829,N6830,N6831,N6832,N6833,N6834,N6835,N6836,N6837,N6838,N6839,N6840,N6841,
  N6842,N6843,N6844,N6845,N6846,N6847,N6848,N6849,N6850,N6851,N6852,N6853,N6854,
  N6855,N6856,N6857,N6858,N6859,N6860,N6861,N6862,N6863,N6864,N6865,N6866,N6867,N6868,
  N6869,N6870,N6871,N6872,N6873,N6874,N6875,N6876,N6877,N6878,N6879,N6880,N6881,
  N6882,N6883,N6884,N6885,N6886,N6887,N6888,N6889,N6890,N6891,N6892,N6893,N6894,
  N6895,N6896,N6897,N6898,N6899,N6900,N6901,N6902,N6903,N6904,N6905,N6906,N6907,N6908,
  N6909,N6910,N6911,N6912,N6913,N6914,N6915,N6916,N6917,N6918,N6919,N6920,N6921,
  N6922,N6923,N6924,N6925,N6926,N6927,N6928,N6929,N6930,N6931,N6932,N6933,N6934,
  N6935,N6936,N6937,N6938,N6939,N6940,N6941,N6942,N6943,N6944,N6945,N6946,N6947,N6948,
  N6949,N6950,N6951,N6952,N6953,N6954,N6955,N6956,N6957,N6958,N6959,N6960,N6961,
  N6962,N6963,N6964,N6965,N6966,N6967,N6968,N6969,N6970,N6971,N6972,N6973,N6974,
  N6975,N6976,N6977,N6978,N6979,N6980,N6981,N6982,N6983,N6984,N6985,N6986,N6987,N6988,
  N6989,N6990,N6991,N6992,N6993,N6994,N6995,N6996,N6997,N6998,N6999,N7000,N7001,
  N7002,N7003,N7004,N7005,N7006,N7007,N7008,N7009,N7010,N7011,N7012,N7013,N7014,
  N7015,N7016,N7017,N7018,N7019,N7020,N7021,N7022,N7023,N7024,N7025,N7026,N7027,N7028,
  N7029,N7030,N7031,N7032,N7033,N7034,N7035,N7036,N7037,N7038,N7039,N7040,N7041,
  N7042,N7043,N7044,N7045,N7046,N7047,N7048,N7049,N7050,N7051,N7052,N7053,N7054,
  N7055,N7056,N7057,N7058,N7059,N7060,N7061,N7062,N7063,N7064,N7065,N7066,N7067,N7068,
  N7069,N7070,N7071,N7072,N7073,N7074,N7075,N7076,N7077,N7078,N7079,N7080,N7081,
  N7082,N7083,N7084,N7085,N7086,N7087,N7088,N7089,N7090,N7091,N7092,N7093,N7094,
  N7095,N7096,N7097,N7098,N7099,N7100,N7101,N7102,N7103,N7104,N7105,N7106,N7107,N7108,
  N7109,N7110,N7111,N7112,N7113,N7114,N7115,N7116,N7117,N7118,N7119,N7120,N7121,
  N7122,N7123,N7124,N7125,N7126,N7127,N7128,N7129,N7130,N7131,N7132,N7133,N7134,
  N7135,N7136,N7137,N7138,N7139,N7140,N7141,N7142,N7143,N7144,N7145,N7146,N7147,N7148,
  N7149,N7150,N7151,N7152,N7153,N7154,N7155,N7156,N7157,N7158,N7159,N7160,N7161,
  N7162,N7163,N7164,N7165,N7166,N7167,N7168,N7169,N7170,N7171,N7172,N7173,N7174,
  N7175,N7176,N7177,N7178,N7179,N7180,N7181,N7182,N7183,N7184,N7185,N7186,N7187,N7188,
  N7189,N7190,N7191,N7192,N7193,N7194,N7195,N7196,N7197,N7198,N7199,N7200,N7201,
  N7202,N7203,N7204,N7205,N7206,N7207,N7208,N7209,N7210,N7211,N7212,N7213,N7214,
  N7215,N7216,N7217,N7218,N7219,N7220,N7221,N7222,N7223,N7224,N7225,N7226,N7227,N7228,
  N7229,N7230,N7231,N7232,N7233,N7234,N7235,N7236,N7237,N7238,N7239,N7240,N7241,
  N7242,N7243,N7244,N7245,N7246,N7247,N7248,N7249,N7250,N7251,N7252,N7253,N7254,
  N7255,N7256,N7257,N7258,N7259,N7260,N7261,N7262,N7263,N7264,N7265,N7266,N7267,N7268,
  N7269,N7270,N7271,N7272,N7273,N7274,N7275,N7276,N7277,N7278,N7279,N7280,N7281,
  N7282,N7283,N7284,N7285,N7286,N7287,N7288,N7289,N7290,N7291,N7292,N7293,N7294,
  N7295,N7296,N7297,N7298,N7299,N7300,N7301,N7302,N7303,N7304,N7305,N7306,N7307,N7308,
  N7309,N7310,N7311,N7312,N7313,N7314,N7315,N7316,N7317,N7318,N7319,N7320,N7321,
  N7322,N7323,N7324,N7325,N7326,N7327,N7328,N7329,N7330,N7331,N7332,N7333,N7334,
  N7335,N7336,N7337,N7338,N7339,N7340,N7341,N7342,N7343,N7344,N7345,N7346,N7347,N7348,
  N7349,N7350,N7351,N7352,N7353,N7354,N7355,N7356,N7357,N7358,N7359,N7360,N7361,
  N7362,N7363,N7364,N7365,N7366,N7367,N7368,N7369,N7370,N7371,N7372,N7373,N7374,
  N7375,N7376,N7377,N7378,N7379,N7380,N7381,N7382,N7383,N7384,N7385,N7386,N7387,N7388,
  N7389,N7390,N7391,N7392,N7393,N7394,N7395,N7396,N7397,N7398,N7399,N7400,N7401,
  N7402,N7403,N7404,N7405,N7406,N7407,N7408,N7409,N7410,N7411,N7412,N7413,N7414,
  N7415,N7416,N7417,N7418,N7419,N7420,N7421,N7422,N7423,N7424,N7425,N7426,N7427,N7428,
  N7429,N7430,N7431,N7432,N7433,N7434,N7435,N7436,N7437,N7438,N7439,N7440,N7441,
  N7442,N7443,N7444,N7445,N7446,N7447,N7448,N7449,N7450,N7451,N7452,N7453,N7454,
  N7455,N7456,N7457,N7458,N7459,N7460,N7461,N7462,N7463,N7464,N7465,N7466,N7467,N7468,
  N7469,N7470,N7471,N7472,N7473,N7474,N7475,N7476,N7477,N7478,N7479,N7480,N7481,
  N7482,N7483,N7484,N7485,N7486,N7487,N7488,N7489,N7490,N7491,N7492,N7493,N7494,
  N7495,N7496,N7497,N7498,N7499,N7500,N7501,N7502,N7503,N7504,N7505,N7506,N7507,N7508,
  N7509,N7510,N7511,N7512,N7513,N7514,N7515,N7516,N7517,N7518,N7519,N7520,N7521,
  N7522,N7523,N7524,N7525,N7526,N7527,N7528,N7529,N7530,N7531,N7532,N7533,N7534,
  N7535,N7536,N7537,N7538,N7539,N7540,N7541,N7542,N7543,N7544,N7545,N7546,N7547,N7548,
  N7549,N7550,N7551,N7552,N7553,N7554,N7555,N7556,N7557,N7558,N7559,N7560,N7561,
  N7562,N7563,N7564,N7565,N7566,N7567,N7568,N7569,N7570,N7571,N7572,N7573,N7574,
  N7575,N7576,N7577,N7578,N7579,N7580,N7581,N7582,N7583,N7584,N7585,N7586,N7587,N7588,
  N7589,N7590,N7591,N7592,N7593,N7594,N7595,N7596,N7597,N7598,N7599,N7600,N7601,
  N7602,N7603,N7604,N7605,N7606,N7607,N7608,N7609,N7610,N7611,N7612,N7613,N7614,
  N7615,N7616,N7617,N7618,N7619,N7620,N7621,N7622,N7623,N7624,N7625,N7626,N7627,N7628,
  N7629,N7630,N7631,N7632,N7633,N7634,N7635,N7636,N7637,N7638,N7639,N7640,N7641,
  N7642,N7643,N7644,N7645,N7646,N7647,N7648,N7649,N7650,N7651,N7652,N7653,N7654,
  N7655,N7656,N7657,N7658,N7659,N7660,N7661,N7662,N7663,N7664,N7665,N7666,N7667,N7668,
  N7669,N7670,N7671,N7672,N7673,N7674,N7675,N7676,N7677,N7678,N7679,N7680,N7681,
  N7682,N7683,N7684,N7685,N7686,N7687,N7688,N7689,N7690,N7691,N7692,N7693,N7694,
  N7695,N7696,N7697,N7698,N7699,N7700,N7701,N7702,N7703,N7704,N7705,N7706,N7707,N7708,
  N7709,N7710,N7711,N7712,N7713,N7714,N7715,N7716,N7717,N7718,N7719,N7720,N7721,
  N7722,N7723,N7724,N7725,N7726,N7727,N7728,N7729,N7730,N7731,N7732,N7733,N7734,
  N7735,N7736,N7737,N7738,N7739,N7740,N7741,N7742,N7743,N7744,N7745,N7746,N7747,N7748,
  N7749,N7750,N7751,N7752,N7753,N7754,N7755,N7756,N7757,N7758,N7759,N7760,N7761,
  N7762,N7763,N7764,N7765,N7766,N7767,N7768,N7769,N7770,N7771,N7772,N7773,N7774,
  N7775,N7776,N7777,N7778,N7779,N7780,N7781,N7782,N7783,N7784,N7785,N7786,N7787,N7788,
  N7789,N7790,N7791,N7792,N7793,N7794,N7795,N7796,N7797,N7798,N7799,N7800,N7801,
  N7802,N7803,N7804,N7805,N7806,N7807,N7808,N7809,N7810,N7811,N7812,N7813,N7814,
  N7815,N7816,N7817,N7818,N7819,N7820,N7821,N7822,N7823,N7824,N7825,N7826,N7827,N7828,
  N7829,N7830,N7831,N7832,N7833,N7834,N7835,N7836,N7837,N7838,N7839,N7840,N7841,
  N7842,N7843,N7844,N7845,N7846,N7847,N7848,N7849,N7850,N7851,N7852,N7853,N7854,
  N7855,N7856,N7857,N7858,N7859,N7860,N7861,N7862,N7863,N7864,N7865,N7866,N7867,N7868,
  N7869,N7870,N7871,N7872,N7873,N7874,N7875,N7876,N7877,N7878,N7879,N7880,N7881,
  N7882,N7883,N7884,N7885,N7886,N7887,N7888,N7889,N7890,N7891,N7892,N7893,N7894,
  N7895,N7896,N7897,N7898,N7899,N7900,N7901,N7902,N7903,N7904,N7905,N7906,N7907,N7908,
  N7909,N7910,N7911,N7912,N7913,N7914,N7915,N7916,N7917,N7918,N7919,N7920,N7921,
  N7922,N7923,N7924,N7925,N7926,N7927,N7928,N7929,N7930,N7931,N7932,N7933,N7934,
  N7935,N7936,N7937,N7938,N7939,N7940,N7941,N7942,N7943,N7944,N7945,N7946,N7947,N7948,
  N7949,N7950,N7951,N7952,N7953,N7954,N7955,N7956,N7957,N7958,N7959,N7960,N7961,
  N7962,N7963,N7964,N7965,N7966,N7967,N7968,N7969,N7970,N7971,N7972,N7973,N7974,
  N7975,N7976,N7977,N7978,N7979,N7980,N7981,N7982,N7983,N7984,N7985,N7986,N7987,N7988,
  N7989,N7990,N7991,N7992,N7993,N7994,N7995,N7996,N7997,N7998,N7999,N8000,N8001,
  N8002,N8003,N8004,N8005,N8006,N8007,N8008,N8009,N8010,N8011,N8012,N8013,N8014,
  N8015,N8016,N8017,N8018,N8019,N8020,N8021,N8022,N8023,N8024,N8025,N8026,N8027,N8028,
  N8029,N8030,N8031,N8032,N8033,N8034,N8035,N8036,N8037,N8038,N8039,N8040,N8041,
  N8042,N8043,N8044,N8045,N8046,N8047,N8048,N8049,N8050,N8051,N8052,N8053,N8054,
  N8055,N8056,N8057,N8058,N8059,N8060,N8061,N8062,N8063,N8064,N8065,N8066,N8067,N8068,
  N8069,N8070,N8071,N8072,N8073,N8074,N8075,N8076,N8077,N8078,N8079,N8080,N8081,
  N8082,N8083,N8084,N8085,N8086,N8087,N8088,N8089,N8090,N8091,N8092,N8093,N8094,
  N8095,N8096,N8097,N8098,N8099,N8100,N8101,N8102,N8103,N8104,N8105,N8106,N8107,N8108,
  N8109,N8110,N8111,N8112,N8113,N8114,N8115,N8116,N8117,N8118,N8119,N8120,N8121,
  N8122,N8123,N8124,N8125,N8126,N8127,N8128,N8129,N8130,N8131,N8132,N8133,N8134,
  N8135,N8136,N8137,N8138,N8139,N8140,N8141,N8142,N8143,N8144,N8145,N8146,N8147,N8148,
  N8149,N8150,N8151,N8152,N8153,N8154,N8155,N8156,N8157,N8158,N8159,N8160,N8161,
  N8162,N8163,N8164,N8165,N8166,N8167,N8168,N8169,N8170,N8171,N8172,N8173,N8174,
  N8175,N8176,N8177,N8178,N8179,N8180,N8181,N8182,N8183,N8184,N8185,N8186,N8187,N8188,
  N8189,N8190,N8191,N8192,N8193,N8194,N8195,N8196,N8197,N8198,N8199,N8200,N8201,
  N8202,N8203,N8204,N8205,N8206,N8207,N8208,N8209,N8210,N8211,N8212,N8213,N8214,
  N8215,N8216,N8217,N8218,N8219,N8220,N8221,N8222,N8223,N8224,N8225,N8226,N8227,N8228,
  N8229,N8230,N8231,N8232,N8233,N8234,N8235,N8236,N8237,N8238,N8239,N8240,N8241,
  N8242,N8243,N8244,N8245,N8246,N8247,N8248,N8249,N8250,N8251,N8252,N8253,N8254,
  N8255,N8256,N8257,N8258,N8259,N8260,N8261,N8262,N8263,N8264,N8265,N8266,N8267,N8268,
  N8269,N8270,N8271,N8272,N8273,N8274,N8275,N8276,N8277,N8278,N8279,N8280,N8281,
  N8282,N8283,N8284,N8285,N8286,N8287,N8288,N8289,N8290,N8291,N8292,N8293,N8294,
  N8295,N8296,N8297,N8298,N8299,N8300,N8301,N8302,N8303,N8304,N8305,N8306,N8307,N8308,
  N8309,N8310,N8311,N8312,N8313,N8314,N8315,N8316,N8317,N8318,N8319,N8320,N8321,
  N8322,N8323,N8324,N8325,N8326,N8327,N8328,N8329,N8330,N8331,N8332,N8333,N8334,
  N8335,N8336,N8337,N8338,N8339,N8340,N8341,N8342,N8343,N8344,N8345,N8346,N8347,N8348,
  N8349,N8350,N8351,N8352,N8353,N8354,N8355,N8356,N8357,N8358,N8359,N8360,N8361,
  N8362,N8363,N8364,N8365,N8366,N8367,N8368,N8369,N8370,N8371,N8372,N8373,N8374,
  N8375,N8376,N8377,N8378,N8379,N8380,N8381,N8382,N8383,N8384,N8385,N8386,N8387,N8388,
  N8389,N8390,N8391,N8392,N8393,N8394,N8395,N8396,N8397,N8398,N8399,N8400,N8401,
  N8402,N8403,N8404,N8405,N8406,N8407,N8408,N8409,N8410,N8411,N8412,N8413,N8414,
  N8415,N8416,N8417,N8418,N8419,N8420,N8421,N8422,N8423,N8424,N8425,N8426,N8427,N8428,
  N8429,N8430,N8431,N8432,N8433,N8434,N8435,N8436,N8437,N8438,N8439,N8440,N8441,
  N8442,N8443,N8444,N8445,N8446,N8447,N8448,N8449,N8450,N8451,N8452,N8453,N8454,
  N8455,N8456,N8457,N8458,N8459,N8460,N8461,N8462,N8463,N8464,N8465,N8466,N8467,N8468,
  N8469,N8470,N8471,N8472,N8473,N8474,N8475,N8476,N8477,N8478,N8479,N8480,N8481,
  N8482,N8483,N8484,N8485,N8486,N8487,N8488,N8489,N8490,N8491,N8492,N8493,N8494,
  N8495,N8496,N8497,N8498,N8499,N8500,N8501,N8502,N8503,N8504,N8505,N8506,N8507,N8508,
  N8509,N8510,N8511,N8512,N8513,N8514,N8515,N8516,N8517,N8518,N8519,N8520,N8521,
  N8522,N8523,N8524,N8525,N8526,N8527,N8528,N8529,N8530,N8531,N8532,N8533,N8534,
  N8535,N8536,N8537,N8538,N8539,N8540,N8541,N8542,N8543,N8544,N8545,N8546,N8547,N8548,
  N8549,N8550,N8551,N8552,N8553,N8554,N8555,N8556,N8557,N8558,N8559,N8560,N8561,
  N8562,N8563,N8564,N8565,N8566,N8567,N8568,N8569,N8570,N8571,N8572,N8573,N8574,
  N8575,N8576,N8577,N8578,N8579,N8580,N8581,N8582,N8583,N8584,N8585,N8586,N8587,N8588,
  N8589,N8590,N8591,N8592,N8593,N8594,N8595,N8596,N8597,N8598,N8599,N8600,N8601,
  N8602,N8603,N8604,N8605,N8606,N8607,N8608,N8609,N8610,N8611,N8612,N8613,N8614,
  N8615,N8616,N8617,N8618,N8619,N8620,N8621,N8622,N8623,N8624,N8625,N8626,N8627,N8628,
  N8629,N8630,N8631,N8632,N8633,N8634,N8635,N8636,N8637,N8638,N8639,N8640,N8641,
  N8642,N8643,N8644,N8645,N8646,N8647,N8648,N8649,N8650,N8651,N8652,N8653,N8654,
  N8655,N8656,N8657,N8658,N8659,N8660,N8661,N8662,N8663,N8664,N8665,N8666,N8667,N8668,
  N8669,N8670,N8671,N8672,N8673,N8674,N8675,N8676,N8677,N8678,N8679,N8680,N8681,
  N8682,N8683,N8684,N8685,N8686,N8687,N8688,N8689,N8690,N8691,N8692,N8693,N8694,
  N8695,N8696,N8697,N8698,N8699,N8700,N8701,N8702,N8703,N8704,N8705,N8706,N8707,N8708,
  N8709,N8710,N8711,N8712,N8713,N8714,N8715,N8716,N8717,N8718,N8719,N8720,N8721,
  N8722,N8723,N8724,N8725,N8726,N8727,N8728,N8729,N8730,N8731,N8732,N8733,N8734,
  N8735,N8736,N8737,N8738,N8739,N8740,N8741,N8742,N8743,N8744,N8745,N8746,N8747,N8748,
  N8749,N8750,N8751,N8752,N8753,N8754,N8755,N8756,N8757,N8758,N8759,N8760,N8761,
  N8762,N8763,N8764,N8765,N8766,N8767,N8768,N8769,N8770,N8771,N8772,N8773,N8774,
  N8775,N8776,N8777,N8778,N8779,N8780,N8781,N8782,N8783,N8784,N8785,N8786,N8787,N8788,
  N8789,N8790,N8791,N8792,N8793,N8794,N8795,N8796,N8797,N8798,N8799,N8800,N8801,
  N8802,N8803,N8804,N8805,N8806,N8807,N8808,N8809,N8810,N8811,N8812,N8813,N8814,
  N8815,N8816,N8817,N8818,N8819,N8820,N8821,N8822,N8823,N8824,N8825,N8826,N8827,N8828,
  N8829,N8830,N8831,N8832,N8833,N8834,N8835,N8836,N8837,N8838,N8839,N8840,N8841,
  N8842,N8843,N8844,N8845,N8846,N8847,N8848,N8849,N8850,N8851,N8852,N8853,N8854,
  N8855,N8856,N8857,N8858,N8859,N8860,N8861,N8862,N8863,N8864,N8865,N8866,N8867,N8868,
  N8869,N8870,N8871,N8872,N8873,N8874,N8875,N8876,N8877,N8878,N8879,N8880,N8881,
  N8882,N8883,N8884,N8885,N8886,N8887,N8888,N8889,N8890,N8891,N8892,N8893,N8894,
  N8895,N8896,N8897,N8898,N8899,N8900,N8901,N8902,N8903,N8904,N8905,N8906,N8907,N8908,
  N8909,N8910,N8911,N8912,N8913,N8914,N8915,N8916,N8917,N8918,N8919,N8920,N8921,
  N8922,N8923,N8924,N8925,N8926,N8927,N8928,N8929,N8930,N8931,N8932,N8933,N8934,
  N8935,N8936,N8937,N8938,N8939,N8940,N8941,N8942,N8943,N8944,N8945,N8946,N8947,N8948,
  N8949,N8950,N8951,N8952,N8953,N8954,N8955,N8956,N8957,N8958,N8959,N8960,N8961,
  N8962,N8963,N8964,N8965,N8966,N8967,N8968,N8969,N8970,N8971,N8972,N8973,N8974,
  N8975,N8976,N8977,N8978,N8979,N8980,N8981,N8982,N8983,N8984,N8985,N8986,N8987,N8988,
  N8989,N8990,N8991,N8992,N8993,N8994,N8995,N8996,N8997,N8998,N8999,N9000,N9001,
  N9002,N9003,N9004,N9005,N9006,N9007,N9008,N9009,N9010,N9011,N9012,N9013,N9014,
  N9015,N9016,N9017,N9018,N9019,N9020,N9021,N9022,N9023,N9024,N9025,N9026,N9027,N9028,
  N9029,N9030,N9031,N9032,N9033,N9034,N9035,N9036,N9037,N9038,N9039,N9040,N9041,
  N9042,N9043,N9044,N9045,N9046,N9047,N9048,N9049,N9050,N9051,N9052,N9053,N9054,
  N9055,N9056,N9057,N9058,N9059,N9060,N9061,N9062,N9063,N9064,N9065,N9066,N9067,N9068,
  N9069,N9070,N9071,N9072,N9073,N9074,N9075,N9076,N9077,N9078,N9079,N9080,N9081,
  N9082,N9083,N9084,N9085,N9086,N9087,N9088,N9089,N9090,N9091,N9092,N9093,N9094,
  N9095,N9096,N9097,N9098,N9099,N9100,N9101,N9102,N9103,N9104,N9105,N9106,N9107,N9108,
  N9109,N9110,N9111,N9112,N9113,N9114,N9115,N9116,N9117,N9118,N9119,N9120,N9121,
  N9122,N9123,N9124,N9125,N9126,N9127,N9128,N9129,N9130,N9131,N9132,N9133,N9134,
  N9135,N9136,N9137,N9138,N9139,N9140,N9141,N9142,N9143,N9144,N9145,N9146,N9147,N9148,
  N9149,N9150,N9151,N9152,N9153,N9154,N9155,N9156,N9157,N9158,N9159,N9160,N9161,
  N9162,N9163,N9164,N9165,N9166,N9167,N9168,N9169,N9170,N9171,N9172,N9173,N9174,
  N9175,N9176,N9177,N9178,N9179,N9180,N9181,N9182,N9183,N9184,N9185,N9186,N9187,N9188,
  N9189,N9190,N9191,N9192,N9193,N9194,N9195,N9196,N9197,N9198,N9199,N9200,N9201,
  N9202,N9203,N9204,N9205,N9206,N9207,N9208,N9209,N9210,N9211,N9212,N9213,N9214,
  N9215,N9216,N9217,N9218,N9219,N9220,N9221,N9222,N9223,N9224,N9225,N9226,N9227,N9228,
  N9229,N9230,N9231,N9232,N9233,N9234,N9235,N9236,N9237,N9238,N9239,N9240,N9241,
  N9242,N9243,N9244,N9245,N9246,N9247,N9248,N9249,N9250,N9251,N9252,N9253,N9254,
  N9255,N9256,N9257,N9258,N9259,N9260,N9261,N9262,N9263,N9264,N9265,N9266,N9267,N9268,
  N9269,N9270,N9271,N9272,N9273,N9274,N9275,N9276,N9277,N9278,N9279,N9280,N9281,
  N9282,N9283,N9284,N9285,N9286,N9287,N9288,N9289,N9290,N9291,N9292,N9293,N9294,
  N9295,N9296,N9297,N9298,N9299,N9300,N9301,N9302,N9303,N9304,N9305,N9306,N9307,N9308,
  N9309,N9310,N9311,N9312,N9313,N9314,N9315,N9316,N9317,N9318,N9319,N9320,N9321,
  N9322,N9323,N9324,N9325,N9326,N9327,N9328,N9329,N9330,N9331,N9332,N9333,N9334,
  N9335,N9336,N9337,N9338,N9339,N9340,N9341,N9342,N9343,N9344,N9345,N9346,N9347,N9348,
  N9349,N9350,N9351,N9352,N9353,N9354,N9355,N9356,N9357,N9358,N9359,N9360,N9361,
  N9362,N9363,N9364,N9365,N9366,N9367,N9368,N9369,N9370,N9371,N9372,N9373,N9374,
  N9375,N9376,N9377,N9378,N9379,N9380,N9381,N9382,N9383,N9384,N9385,N9386,N9387,N9388,
  N9389,N9390,N9391,N9392,N9393,N9394,N9395,N9396,N9397,N9398,N9399,N9400,N9401,
  N9402,N9403,N9404,N9405,N9406,N9407,N9408,N9409,N9410,N9411,N9412,N9413,N9414,
  N9415,N9416,N9417,N9418,N9419,N9420,N9421,N9422,N9423,N9424,N9425,N9426,N9427,N9428,
  N9429,N9430,N9431,N9432,N9433,N9434,N9435,N9436,N9437,N9438,N9439,N9440,N9441,
  N9442,N9443,N9444,N9445,N9446,N9447,N9448,N9449,N9450,N9451,N9452,N9453,N9454,
  N9455,N9456,N9457,N9458,N9459,N9460,N9461,N9462,N9463,N9464,N9465,N9466,N9467,N9468,
  N9469,N9470,N9471,N9472,N9473,N9474,N9475,N9476,N9477,N9478,N9479,N9480,N9481,
  N9482,N9483,N9484,N9485,N9486,N9487,N9488,N9489,N9490,N9491,N9492,N9493,N9494,
  N9495,N9496,N9497,N9498,N9499,N9500,N9501,N9502,N9503,N9504,N9505,N9506,N9507,N9508,
  N9509,N9510,N9511,N9512,N9513,N9514,N9515,N9516,N9517,N9518,N9519,N9520,N9521,
  N9522,N9523,N9524,N9525,N9526,N9527,N9528,N9529,N9530,N9531,N9532,N9533,N9534,
  N9535,N9536,N9537,N9538,N9539,N9540,N9541,N9542,N9543,N9544,N9545,N9546,N9547,N9548,
  N9549,N9550,N9551,N9552,N9553,N9554,N9555,N9556,N9557,N9558,N9559,N9560,N9561,
  N9562,N9563,N9564,N9565,N9566,N9567,N9568,N9569,N9570,N9571,N9572,N9573,N9574,
  N9575,N9576,N9577,N9578,N9579,N9580,N9581,N9582,N9583,N9584,N9585,N9586,N9587,N9588,
  N9589,N9590,N9591,N9592,N9593,N9594,N9595,N9596,N9597,N9598,N9599,N9600,N9601,
  N9602,N9603,N9604,N9605,N9606,N9607,N9608,N9609,N9610,N9611,N9612,N9613,N9614,
  N9615,N9616,N9617,N9618,N9619,N9620,N9621,N9622,N9623,N9624,N9625,N9626,N9627,N9628,
  N9629,N9630,N9631,N9632,N9633,N9634,N9635,N9636,N9637,N9638,N9639,N9640,N9641,
  N9642,N9643,N9644,N9645,N9646,N9647,N9648,N9649,N9650,N9651,N9652,N9653,N9654,
  N9655,N9656,N9657,N9658,N9659,N9660,N9661,N9662,N9663,N9664,N9665,N9666,N9667,N9668,
  N9669,N9670,N9671,N9672,N9673,N9674,N9675,N9676,N9677,N9678,N9679,N9680,N9681,
  N9682,N9683,N9684,N9685,N9686,N9687,N9688,N9689,N9690,N9691,N9692,N9693,N9694,
  N9695,N9696,N9697,N9698,N9699,N9700,N9701,N9702,N9703,N9704,N9705,N9706,N9707,N9708,
  N9709,N9710,N9711,N9712,N9713,N9714,N9715,N9716,N9717,N9718,N9719,N9720,N9721,
  N9722,N9723,N9724,N9725,N9726,N9727,N9728,N9729,N9730,N9731,N9732,N9733,N9734,
  N9735,N9736,N9737,N9738,N9739,N9740,N9741,N9742,N9743,N9744,N9745,N9746,N9747,N9748,
  N9749,N9750,N9751,N9752,N9753,N9754,N9755,N9756,N9757,N9758,N9759,N9760,N9761,
  N9762,N9763,N9764,N9765,N9766,N9767,N9768,N9769,N9770,N9771,N9772,N9773,N9774,
  N9775,N9776,N9777,N9778,N9779,N9780,N9781,N9782,N9783,N9784,N9785,N9786,N9787,N9788,
  N9789,N9790,N9791,N9792,N9793,N9794,N9795,N9796,N9797,N9798,N9799,N9800,N9801,
  N9802,N9803,N9804,N9805,N9806,N9807,N9808,N9809,N9810,N9811,N9812,N9813,N9814,
  N9815,N9816,N9817,N9818,N9819,N9820,N9821,N9822,N9823,N9824,N9825,N9826,N9827,N9828,
  N9829,N9830,N9831,N9832,N9833,N9834,N9835,N9836,N9837,N9838,N9839,N9840,N9841,
  N9842,N9843,N9844,N9845,N9846,N9847,N9848,N9849,N9850,N9851,N9852,N9853,N9854,
  N9855,N9856,N9857,N9858,N9859,N9860,N9861,N9862,N9863,N9864,N9865,N9866,N9867,N9868,
  N9869,N9870,N9871,N9872,N9873,N9874,N9875,N9876,N9877,N9878,N9879,N9880,N9881,
  N9882,N9883,N9884,N9885,N9886,N9887,N9888,N9889,N9890,N9891,N9892,N9893,N9894,
  N9895,N9896,N9897,N9898,N9899,N9900,N9901,N9902,N9903,N9904,N9905,N9906,N9907,N9908,
  N9909,N9910,N9911,N9912,N9913,N9914,N9915,N9916,N9917,N9918,N9919,N9920,N9921,
  N9922,N9923,N9924,N9925,N9926,N9927,N9928,N9929,N9930,N9931,N9932,N9933,N9934,
  N9935,N9936,N9937,N9938,N9939,N9940,N9941,N9942,N9943,N9944,N9945,N9946,N9947,N9948,
  N9949,N9950,N9951,N9952,N9953,N9954,N9955,N9956,N9957,N9958,N9959,N9960,N9961,
  N9962,N9963,N9964,N9965,N9966,N9967,N9968,N9969,N9970,N9971,N9972,N9973,N9974,
  N9975,N9976,N9977,N9978,N9979,N9980,N9981,N9982,N9983,N9984,N9985,N9986,N9987,N9988,
  N9989,N9990,N9991,N9992,N9993,N9994,N9995,N9996,N9997,N9998,N9999,N10000,N10001,
  N10002,N10003,N10004,N10005,N10006,N10007,N10008,N10009,N10010,N10011,N10012,
  N10013,N10014,N10015,N10016,N10017,N10018,N10019,N10020,N10021,N10022,N10023,N10024,
  N10025,N10026,N10027,N10028,N10029,N10030,N10031,N10032,N10033,N10034,N10035,
  N10036,N10037,N10038,N10039,N10040,N10041,N10042,N10043,N10044,N10045,N10046,
  N10047,N10048,N10049,N10050,N10051,N10052,N10053,N10054,N10055,N10056,N10057,N10058,
  N10059,N10060,N10061,N10062,N10063,N10064,N10065,N10066,N10067,N10068,N10069,
  N10070,N10071,N10072,N10073,N10074,N10075,N10076,N10077,N10078,N10079,N10080,N10081,
  N10082,N10083,N10084,N10085,N10086,N10087,N10088,N10089,N10090,N10091,N10092,
  N10093,N10094,N10095,N10096,N10097,N10098,N10099,N10100,N10101,N10102,N10103,N10104,
  N10105,N10106,N10107,N10108,N10109,N10110,N10111,N10112,N10113,N10114,N10115,
  N10116,N10117,N10118,N10119,N10120,N10121,N10122,N10123,N10124,N10125,N10126,
  N10127,N10128,N10129,N10130,N10131,N10132,N10133,N10134,N10135,N10136,N10137,N10138,
  N10139,N10140,N10141,N10142,N10143,N10144,N10145,N10146,N10147,N10148,N10149,
  N10150,N10151,N10152,N10153,N10154,N10155,N10156,N10157,N10158,N10159,N10160,N10161,
  N10162,N10163,N10164,N10165,N10166,N10167,N10168,N10169,N10170,N10171,N10172,
  N10173,N10174,N10175,N10176,N10177,N10178,N10179,N10180,N10181,N10182,N10183,N10184,
  N10185,N10186,N10187,N10188,N10189,N10190,N10191,N10192,N10193,N10194,N10195,
  N10196,N10197,N10198,N10199,N10200,N10201,N10202,N10203,N10204,N10205,N10206,
  N10207,N10208,N10209,N10210,N10211,N10212,N10213,N10214,N10215,N10216,N10217,N10218,
  N10219,N10220,N10221,N10222,N10223,N10224,N10225,N10226,N10227,N10228,N10229,
  N10230,N10231,N10232,N10233,N10234,N10235,N10236,N10237,N10238,N10239,N10240,N10241,
  N10242,N10243,N10244,N10245,N10246,N10247,N10248,N10249,N10250,N10251,N10252,
  N10253,N10254,N10255,N10256,N10257,N10258,N10259,N10260,N10261,N10262,N10263,N10264,
  N10265,N10266,N10267,N10268,N10269,N10270,N10271,N10272,N10273,N10274,N10275,
  N10276,N10277,N10278,N10279,N10280,N10281,N10282,N10283,N10284,N10285,N10286,
  N10287,N10288,N10289,N10290,N10291,N10292,N10293,N10294,N10295,N10296,N10297,N10298,
  N10299,N10300,N10301,N10302,N10303,N10304,N10305,N10306,N10307,N10308,N10309,
  N10310,N10311,N10312,N10313,N10314,N10315,N10316,N10317,N10318,N10319,N10320,N10321,
  N10322,N10323,N10324,N10325,N10326,N10327,N10328,N10329,N10330,N10331,N10332,
  N10333,N10334,N10335,N10336,N10337,N10338,N10339,N10340,N10341,N10342,N10343,N10344,
  N10345,N10346,N10347,N10348,N10349,N10350,N10351,N10352,N10353,N10354,N10355,
  N10356,N10357,N10358,N10359,N10360,N10361,N10362,N10363,N10364,N10365,N10366,
  N10367,N10368,N10369,N10370,N10371,N10372,N10373,N10374,N10375,N10376,N10377,N10378,
  N10379,N10380,N10381,N10382,N10383,N10384,N10385,N10386,N10387,N10388,N10389,
  N10390,N10391,N10392,N10393,N10394,N10395,N10396,N10397,N10398,N10399,N10400,N10401,
  N10402,N10403,N10404,N10405,N10406,N10407,N10408,N10409,N10410,N10411,N10412,
  N10413,N10414,N10415,N10416,N10417,N10418,N10419,N10420,N10421,N10422,N10423,N10424,
  N10425,N10426,N10427,N10428,N10429,N10430,N10431,N10432,N10433,N10434,N10435,
  N10436,N10437,N10438,N10439,N10440,N10441,N10442,N10443,N10444,N10445,N10446,
  N10447,N10448,N10449,N10450,N10451,N10452,N10453,N10454,N10455,N10456,N10457,N10458,
  N10459,N10460,N10461,N10462,N10463,N10464,N10465,N10466,N10467,N10468,N10469,
  N10470,N10471,N10472,N10473,N10474,N10475,N10476,N10477,N10478,N10479,N10480,N10481,
  N10482,N10483,N10484,N10485,N10486,N10487,N10488,N10489,N10490,N10491,N10492,
  N10493,N10494,N10495,N10496,N10497,N10498,N10499,N10500,N10501,N10502,N10503,N10504,
  N10505,N10506,N10507,N10508,N10509,N10510,N10511,N10512,N10513,N10514,N10515,
  N10516,N10517,N10518,N10519,N10520,N10521,N10522,N10523,N10524,N10525,N10526,
  N10527,N10528,N10529,N10530,N10531,N10532,N10533,N10534,N10535,N10536,N10537,N10538,
  N10539,N10540,N10541,N10542,N10543,N10544,N10545,N10546,N10547,N10548,N10549,
  N10550,N10551,N10552,N10553,N10554,N10555,N10556,N10557,N10558,N10559,N10560,N10561,
  N10562,N10563,N10564,N10565,N10566,N10567,N10568,N10569,N10570,N10571,N10572,
  N10573,N10574,N10575,N10576,N10577,N10578,N10579,N10580,N10581,N10582,N10583,N10584,
  N10585,N10586,N10587,N10588,N10589,N10590,N10591,N10592,N10593,N10594,N10595,
  N10596,N10597,N10598,N10599,N10600,N10601,N10602,N10603,N10604,N10605,N10606,
  N10607,N10608,N10609,N10610,N10611,N10612,N10613,N10614,N10615,N10616,N10617,N10618,
  N10619,N10620,N10621,N10622,N10623,N10624,N10625,N10626,N10627,N10628,N10629,
  N10630,N10631,N10632,N10633,N10634,N10635,N10636,N10637,N10638,N10639,N10640,N10641,
  N10642,N10643,N10644,N10645,N10646,N10647,N10648,N10649,N10650,N10651,N10652,
  N10653,N10654,N10655,N10656,N10657,N10658,N10659,N10660,N10661,N10662,N10663,N10664,
  N10665,N10666,N10667,N10668,N10669,N10670,N10671,N10672,N10673,N10674,N10675,
  N10676,N10677,N10678,N10679,N10680,N10681,N10682,N10683,N10684,N10685,N10686,
  N10687,N10688,N10689,N10690,N10691,N10692,N10693,N10694,N10695,N10696,N10697,N10698,
  N10699,N10700,N10701,N10702,N10703,N10704,N10705,N10706,N10707,N10708,N10709,
  N10710,N10711,N10712,N10713,N10714,N10715,N10716,N10717,N10718,N10719,N10720,N10721,
  N10722,N10723,N10724,N10725,N10726,N10727,N10728,N10729,N10730,N10731,N10732,
  N10733,N10734,N10735,N10736;
  wire [5:0] mcause_d;
  wire [31:2] mcountinhibit_d;
  wire [2047:0] mhpmcounter_d;
  reg [31:0] dscratch1_q,mscratch_q,csr_mepc_o,mtval_q,csr_depc_o,dscratch0_q,
  mcountinhibit_q;
  reg m_irq_enable_o,mstatus_q_mpie_,mstatus_q_mpp__1_,mstatus_q_mpp__0_,
  dcsr_q_xdebugver__3_,dcsr_q_xdebugver__2_,dcsr_q_xdebugver__1_,dcsr_q_xdebugver__0_,
  dcsr_q_zero2__11_,dcsr_q_zero2__10_,dcsr_q_zero2__9_,dcsr_q_zero2__8_,dcsr_q_zero2__7_,
  dcsr_q_zero2__6_,dcsr_q_zero2__5_,dcsr_q_zero2__4_,dcsr_q_zero2__3_,
  dcsr_q_zero2__2_,dcsr_q_zero2__1_,dcsr_q_zero2__0_,debug_ebreakm_o,dcsr_q_zero1_,
  dcsr_q_ebreaks_,dcsr_q_ebreaku_,dcsr_q_stepie_,dcsr_q_stopcount_,dcsr_q_stoptime_,
  dcsr_q_cause__2_,dcsr_q_cause__1_,dcsr_q_cause__0_,dcsr_q_zero0_,dcsr_q_mprven_,
  dcsr_q_nmip_,debug_single_step_o,dcsr_q_prv__1_,dcsr_q_prv__0_;
  reg [5:0] mcause_q;
  reg [2047:0] mhpmcounter_q;
  assign N206 = (N337)? mhpmcounter_q[2047] : 
                (N339)? mhpmcounter_q[1983] : 
                (N341)? mhpmcounter_q[1919] : 
                (N343)? mhpmcounter_q[1855] : 
                (N345)? mhpmcounter_q[1791] : 
                (N347)? mhpmcounter_q[1727] : 
                (N349)? mhpmcounter_q[1663] : 
                (N351)? mhpmcounter_q[1599] : 
                (N353)? mhpmcounter_q[1535] : 
                (N355)? mhpmcounter_q[1471] : 
                (N357)? mhpmcounter_q[1407] : 
                (N359)? mhpmcounter_q[1343] : 
                (N361)? mhpmcounter_q[1279] : 
                (N363)? mhpmcounter_q[1215] : 
                (N365)? mhpmcounter_q[1151] : 
                (N367)? mhpmcounter_q[1087] : 
                (N338)? mhpmcounter_q[1023] : 
                (N340)? mhpmcounter_q[959] : 
                (N342)? mhpmcounter_q[895] : 
                (N344)? mhpmcounter_q[831] : 
                (N346)? mhpmcounter_q[767] : 
                (N348)? mhpmcounter_q[703] : 
                (N350)? mhpmcounter_q[639] : 
                (N352)? mhpmcounter_q[575] : 
                (N354)? mhpmcounter_q[511] : 
                (N356)? mhpmcounter_q[447] : 
                (N358)? mhpmcounter_q[383] : 
                (N360)? mhpmcounter_q[319] : 
                (N362)? mhpmcounter_q[255] : 
                (N364)? mhpmcounter_q[191] : 
                (N366)? mhpmcounter_q[127] : 
                (N368)? mhpmcounter_q[63] : 1'b0;
  assign N207 = (N337)? mhpmcounter_q[2046] : 
                (N339)? mhpmcounter_q[1982] : 
                (N341)? mhpmcounter_q[1918] : 
                (N343)? mhpmcounter_q[1854] : 
                (N345)? mhpmcounter_q[1790] : 
                (N347)? mhpmcounter_q[1726] : 
                (N349)? mhpmcounter_q[1662] : 
                (N351)? mhpmcounter_q[1598] : 
                (N353)? mhpmcounter_q[1534] : 
                (N355)? mhpmcounter_q[1470] : 
                (N357)? mhpmcounter_q[1406] : 
                (N359)? mhpmcounter_q[1342] : 
                (N361)? mhpmcounter_q[1278] : 
                (N363)? mhpmcounter_q[1214] : 
                (N365)? mhpmcounter_q[1150] : 
                (N367)? mhpmcounter_q[1086] : 
                (N338)? mhpmcounter_q[1022] : 
                (N340)? mhpmcounter_q[958] : 
                (N342)? mhpmcounter_q[894] : 
                (N344)? mhpmcounter_q[830] : 
                (N346)? mhpmcounter_q[766] : 
                (N348)? mhpmcounter_q[702] : 
                (N350)? mhpmcounter_q[638] : 
                (N352)? mhpmcounter_q[574] : 
                (N354)? mhpmcounter_q[510] : 
                (N356)? mhpmcounter_q[446] : 
                (N358)? mhpmcounter_q[382] : 
                (N360)? mhpmcounter_q[318] : 
                (N362)? mhpmcounter_q[254] : 
                (N364)? mhpmcounter_q[190] : 
                (N366)? mhpmcounter_q[126] : 
                (N368)? mhpmcounter_q[62] : 1'b0;
  assign N208 = (N337)? mhpmcounter_q[2045] : 
                (N339)? mhpmcounter_q[1981] : 
                (N341)? mhpmcounter_q[1917] : 
                (N343)? mhpmcounter_q[1853] : 
                (N345)? mhpmcounter_q[1789] : 
                (N347)? mhpmcounter_q[1725] : 
                (N349)? mhpmcounter_q[1661] : 
                (N351)? mhpmcounter_q[1597] : 
                (N353)? mhpmcounter_q[1533] : 
                (N355)? mhpmcounter_q[1469] : 
                (N357)? mhpmcounter_q[1405] : 
                (N359)? mhpmcounter_q[1341] : 
                (N361)? mhpmcounter_q[1277] : 
                (N363)? mhpmcounter_q[1213] : 
                (N365)? mhpmcounter_q[1149] : 
                (N367)? mhpmcounter_q[1085] : 
                (N338)? mhpmcounter_q[1021] : 
                (N340)? mhpmcounter_q[957] : 
                (N342)? mhpmcounter_q[893] : 
                (N344)? mhpmcounter_q[829] : 
                (N346)? mhpmcounter_q[765] : 
                (N348)? mhpmcounter_q[701] : 
                (N350)? mhpmcounter_q[637] : 
                (N352)? mhpmcounter_q[573] : 
                (N354)? mhpmcounter_q[509] : 
                (N356)? mhpmcounter_q[445] : 
                (N358)? mhpmcounter_q[381] : 
                (N360)? mhpmcounter_q[317] : 
                (N362)? mhpmcounter_q[253] : 
                (N364)? mhpmcounter_q[189] : 
                (N366)? mhpmcounter_q[125] : 
                (N368)? mhpmcounter_q[61] : 1'b0;
  assign N209 = (N337)? mhpmcounter_q[2044] : 
                (N339)? mhpmcounter_q[1980] : 
                (N341)? mhpmcounter_q[1916] : 
                (N343)? mhpmcounter_q[1852] : 
                (N345)? mhpmcounter_q[1788] : 
                (N347)? mhpmcounter_q[1724] : 
                (N349)? mhpmcounter_q[1660] : 
                (N351)? mhpmcounter_q[1596] : 
                (N353)? mhpmcounter_q[1532] : 
                (N355)? mhpmcounter_q[1468] : 
                (N357)? mhpmcounter_q[1404] : 
                (N359)? mhpmcounter_q[1340] : 
                (N361)? mhpmcounter_q[1276] : 
                (N363)? mhpmcounter_q[1212] : 
                (N365)? mhpmcounter_q[1148] : 
                (N367)? mhpmcounter_q[1084] : 
                (N338)? mhpmcounter_q[1020] : 
                (N340)? mhpmcounter_q[956] : 
                (N342)? mhpmcounter_q[892] : 
                (N344)? mhpmcounter_q[828] : 
                (N346)? mhpmcounter_q[764] : 
                (N348)? mhpmcounter_q[700] : 
                (N350)? mhpmcounter_q[636] : 
                (N352)? mhpmcounter_q[572] : 
                (N354)? mhpmcounter_q[508] : 
                (N356)? mhpmcounter_q[444] : 
                (N358)? mhpmcounter_q[380] : 
                (N360)? mhpmcounter_q[316] : 
                (N362)? mhpmcounter_q[252] : 
                (N364)? mhpmcounter_q[188] : 
                (N366)? mhpmcounter_q[124] : 
                (N368)? mhpmcounter_q[60] : 1'b0;
  assign N210 = (N337)? mhpmcounter_q[2043] : 
                (N339)? mhpmcounter_q[1979] : 
                (N341)? mhpmcounter_q[1915] : 
                (N343)? mhpmcounter_q[1851] : 
                (N345)? mhpmcounter_q[1787] : 
                (N347)? mhpmcounter_q[1723] : 
                (N349)? mhpmcounter_q[1659] : 
                (N351)? mhpmcounter_q[1595] : 
                (N353)? mhpmcounter_q[1531] : 
                (N355)? mhpmcounter_q[1467] : 
                (N357)? mhpmcounter_q[1403] : 
                (N359)? mhpmcounter_q[1339] : 
                (N361)? mhpmcounter_q[1275] : 
                (N363)? mhpmcounter_q[1211] : 
                (N365)? mhpmcounter_q[1147] : 
                (N367)? mhpmcounter_q[1083] : 
                (N338)? mhpmcounter_q[1019] : 
                (N340)? mhpmcounter_q[955] : 
                (N342)? mhpmcounter_q[891] : 
                (N344)? mhpmcounter_q[827] : 
                (N346)? mhpmcounter_q[763] : 
                (N348)? mhpmcounter_q[699] : 
                (N350)? mhpmcounter_q[635] : 
                (N352)? mhpmcounter_q[571] : 
                (N354)? mhpmcounter_q[507] : 
                (N356)? mhpmcounter_q[443] : 
                (N358)? mhpmcounter_q[379] : 
                (N360)? mhpmcounter_q[315] : 
                (N362)? mhpmcounter_q[251] : 
                (N364)? mhpmcounter_q[187] : 
                (N366)? mhpmcounter_q[123] : 
                (N368)? mhpmcounter_q[59] : 1'b0;
  assign N211 = (N337)? mhpmcounter_q[2042] : 
                (N339)? mhpmcounter_q[1978] : 
                (N341)? mhpmcounter_q[1914] : 
                (N343)? mhpmcounter_q[1850] : 
                (N345)? mhpmcounter_q[1786] : 
                (N347)? mhpmcounter_q[1722] : 
                (N349)? mhpmcounter_q[1658] : 
                (N351)? mhpmcounter_q[1594] : 
                (N353)? mhpmcounter_q[1530] : 
                (N355)? mhpmcounter_q[1466] : 
                (N357)? mhpmcounter_q[1402] : 
                (N359)? mhpmcounter_q[1338] : 
                (N361)? mhpmcounter_q[1274] : 
                (N363)? mhpmcounter_q[1210] : 
                (N365)? mhpmcounter_q[1146] : 
                (N367)? mhpmcounter_q[1082] : 
                (N338)? mhpmcounter_q[1018] : 
                (N340)? mhpmcounter_q[954] : 
                (N342)? mhpmcounter_q[890] : 
                (N344)? mhpmcounter_q[826] : 
                (N346)? mhpmcounter_q[762] : 
                (N348)? mhpmcounter_q[698] : 
                (N350)? mhpmcounter_q[634] : 
                (N352)? mhpmcounter_q[570] : 
                (N354)? mhpmcounter_q[506] : 
                (N356)? mhpmcounter_q[442] : 
                (N358)? mhpmcounter_q[378] : 
                (N360)? mhpmcounter_q[314] : 
                (N362)? mhpmcounter_q[250] : 
                (N364)? mhpmcounter_q[186] : 
                (N366)? mhpmcounter_q[122] : 
                (N368)? mhpmcounter_q[58] : 1'b0;
  assign N212 = (N337)? mhpmcounter_q[2041] : 
                (N339)? mhpmcounter_q[1977] : 
                (N341)? mhpmcounter_q[1913] : 
                (N343)? mhpmcounter_q[1849] : 
                (N345)? mhpmcounter_q[1785] : 
                (N347)? mhpmcounter_q[1721] : 
                (N349)? mhpmcounter_q[1657] : 
                (N351)? mhpmcounter_q[1593] : 
                (N353)? mhpmcounter_q[1529] : 
                (N355)? mhpmcounter_q[1465] : 
                (N357)? mhpmcounter_q[1401] : 
                (N359)? mhpmcounter_q[1337] : 
                (N361)? mhpmcounter_q[1273] : 
                (N363)? mhpmcounter_q[1209] : 
                (N365)? mhpmcounter_q[1145] : 
                (N367)? mhpmcounter_q[1081] : 
                (N338)? mhpmcounter_q[1017] : 
                (N340)? mhpmcounter_q[953] : 
                (N342)? mhpmcounter_q[889] : 
                (N344)? mhpmcounter_q[825] : 
                (N346)? mhpmcounter_q[761] : 
                (N348)? mhpmcounter_q[697] : 
                (N350)? mhpmcounter_q[633] : 
                (N352)? mhpmcounter_q[569] : 
                (N354)? mhpmcounter_q[505] : 
                (N356)? mhpmcounter_q[441] : 
                (N358)? mhpmcounter_q[377] : 
                (N360)? mhpmcounter_q[313] : 
                (N362)? mhpmcounter_q[249] : 
                (N364)? mhpmcounter_q[185] : 
                (N366)? mhpmcounter_q[121] : 
                (N368)? mhpmcounter_q[57] : 1'b0;
  assign N213 = (N337)? mhpmcounter_q[2040] : 
                (N339)? mhpmcounter_q[1976] : 
                (N341)? mhpmcounter_q[1912] : 
                (N343)? mhpmcounter_q[1848] : 
                (N345)? mhpmcounter_q[1784] : 
                (N347)? mhpmcounter_q[1720] : 
                (N349)? mhpmcounter_q[1656] : 
                (N351)? mhpmcounter_q[1592] : 
                (N353)? mhpmcounter_q[1528] : 
                (N355)? mhpmcounter_q[1464] : 
                (N357)? mhpmcounter_q[1400] : 
                (N359)? mhpmcounter_q[1336] : 
                (N361)? mhpmcounter_q[1272] : 
                (N363)? mhpmcounter_q[1208] : 
                (N365)? mhpmcounter_q[1144] : 
                (N367)? mhpmcounter_q[1080] : 
                (N338)? mhpmcounter_q[1016] : 
                (N340)? mhpmcounter_q[952] : 
                (N342)? mhpmcounter_q[888] : 
                (N344)? mhpmcounter_q[824] : 
                (N346)? mhpmcounter_q[760] : 
                (N348)? mhpmcounter_q[696] : 
                (N350)? mhpmcounter_q[632] : 
                (N352)? mhpmcounter_q[568] : 
                (N354)? mhpmcounter_q[504] : 
                (N356)? mhpmcounter_q[440] : 
                (N358)? mhpmcounter_q[376] : 
                (N360)? mhpmcounter_q[312] : 
                (N362)? mhpmcounter_q[248] : 
                (N364)? mhpmcounter_q[184] : 
                (N366)? mhpmcounter_q[120] : 
                (N368)? mhpmcounter_q[56] : 1'b0;
  assign N214 = (N337)? mhpmcounter_q[2039] : 
                (N339)? mhpmcounter_q[1975] : 
                (N341)? mhpmcounter_q[1911] : 
                (N343)? mhpmcounter_q[1847] : 
                (N345)? mhpmcounter_q[1783] : 
                (N347)? mhpmcounter_q[1719] : 
                (N349)? mhpmcounter_q[1655] : 
                (N351)? mhpmcounter_q[1591] : 
                (N353)? mhpmcounter_q[1527] : 
                (N355)? mhpmcounter_q[1463] : 
                (N357)? mhpmcounter_q[1399] : 
                (N359)? mhpmcounter_q[1335] : 
                (N361)? mhpmcounter_q[1271] : 
                (N363)? mhpmcounter_q[1207] : 
                (N365)? mhpmcounter_q[1143] : 
                (N367)? mhpmcounter_q[1079] : 
                (N338)? mhpmcounter_q[1015] : 
                (N340)? mhpmcounter_q[951] : 
                (N342)? mhpmcounter_q[887] : 
                (N344)? mhpmcounter_q[823] : 
                (N346)? mhpmcounter_q[759] : 
                (N348)? mhpmcounter_q[695] : 
                (N350)? mhpmcounter_q[631] : 
                (N352)? mhpmcounter_q[567] : 
                (N354)? mhpmcounter_q[503] : 
                (N356)? mhpmcounter_q[439] : 
                (N358)? mhpmcounter_q[375] : 
                (N360)? mhpmcounter_q[311] : 
                (N362)? mhpmcounter_q[247] : 
                (N364)? mhpmcounter_q[183] : 
                (N366)? mhpmcounter_q[119] : 
                (N368)? mhpmcounter_q[55] : 1'b0;
  assign N215 = (N337)? mhpmcounter_q[2038] : 
                (N339)? mhpmcounter_q[1974] : 
                (N341)? mhpmcounter_q[1910] : 
                (N343)? mhpmcounter_q[1846] : 
                (N345)? mhpmcounter_q[1782] : 
                (N347)? mhpmcounter_q[1718] : 
                (N349)? mhpmcounter_q[1654] : 
                (N351)? mhpmcounter_q[1590] : 
                (N353)? mhpmcounter_q[1526] : 
                (N355)? mhpmcounter_q[1462] : 
                (N357)? mhpmcounter_q[1398] : 
                (N359)? mhpmcounter_q[1334] : 
                (N361)? mhpmcounter_q[1270] : 
                (N363)? mhpmcounter_q[1206] : 
                (N365)? mhpmcounter_q[1142] : 
                (N367)? mhpmcounter_q[1078] : 
                (N338)? mhpmcounter_q[1014] : 
                (N340)? mhpmcounter_q[950] : 
                (N342)? mhpmcounter_q[886] : 
                (N344)? mhpmcounter_q[822] : 
                (N346)? mhpmcounter_q[758] : 
                (N348)? mhpmcounter_q[694] : 
                (N350)? mhpmcounter_q[630] : 
                (N352)? mhpmcounter_q[566] : 
                (N354)? mhpmcounter_q[502] : 
                (N356)? mhpmcounter_q[438] : 
                (N358)? mhpmcounter_q[374] : 
                (N360)? mhpmcounter_q[310] : 
                (N362)? mhpmcounter_q[246] : 
                (N364)? mhpmcounter_q[182] : 
                (N366)? mhpmcounter_q[118] : 
                (N368)? mhpmcounter_q[54] : 1'b0;
  assign N216 = (N337)? mhpmcounter_q[2037] : 
                (N339)? mhpmcounter_q[1973] : 
                (N341)? mhpmcounter_q[1909] : 
                (N343)? mhpmcounter_q[1845] : 
                (N345)? mhpmcounter_q[1781] : 
                (N347)? mhpmcounter_q[1717] : 
                (N349)? mhpmcounter_q[1653] : 
                (N351)? mhpmcounter_q[1589] : 
                (N353)? mhpmcounter_q[1525] : 
                (N355)? mhpmcounter_q[1461] : 
                (N357)? mhpmcounter_q[1397] : 
                (N359)? mhpmcounter_q[1333] : 
                (N361)? mhpmcounter_q[1269] : 
                (N363)? mhpmcounter_q[1205] : 
                (N365)? mhpmcounter_q[1141] : 
                (N367)? mhpmcounter_q[1077] : 
                (N338)? mhpmcounter_q[1013] : 
                (N340)? mhpmcounter_q[949] : 
                (N342)? mhpmcounter_q[885] : 
                (N344)? mhpmcounter_q[821] : 
                (N346)? mhpmcounter_q[757] : 
                (N348)? mhpmcounter_q[693] : 
                (N350)? mhpmcounter_q[629] : 
                (N352)? mhpmcounter_q[565] : 
                (N354)? mhpmcounter_q[501] : 
                (N356)? mhpmcounter_q[437] : 
                (N358)? mhpmcounter_q[373] : 
                (N360)? mhpmcounter_q[309] : 
                (N362)? mhpmcounter_q[245] : 
                (N364)? mhpmcounter_q[181] : 
                (N366)? mhpmcounter_q[117] : 
                (N368)? mhpmcounter_q[53] : 1'b0;
  assign N217 = (N337)? mhpmcounter_q[2036] : 
                (N339)? mhpmcounter_q[1972] : 
                (N341)? mhpmcounter_q[1908] : 
                (N343)? mhpmcounter_q[1844] : 
                (N345)? mhpmcounter_q[1780] : 
                (N347)? mhpmcounter_q[1716] : 
                (N349)? mhpmcounter_q[1652] : 
                (N351)? mhpmcounter_q[1588] : 
                (N353)? mhpmcounter_q[1524] : 
                (N355)? mhpmcounter_q[1460] : 
                (N357)? mhpmcounter_q[1396] : 
                (N359)? mhpmcounter_q[1332] : 
                (N361)? mhpmcounter_q[1268] : 
                (N363)? mhpmcounter_q[1204] : 
                (N365)? mhpmcounter_q[1140] : 
                (N367)? mhpmcounter_q[1076] : 
                (N338)? mhpmcounter_q[1012] : 
                (N340)? mhpmcounter_q[948] : 
                (N342)? mhpmcounter_q[884] : 
                (N344)? mhpmcounter_q[820] : 
                (N346)? mhpmcounter_q[756] : 
                (N348)? mhpmcounter_q[692] : 
                (N350)? mhpmcounter_q[628] : 
                (N352)? mhpmcounter_q[564] : 
                (N354)? mhpmcounter_q[500] : 
                (N356)? mhpmcounter_q[436] : 
                (N358)? mhpmcounter_q[372] : 
                (N360)? mhpmcounter_q[308] : 
                (N362)? mhpmcounter_q[244] : 
                (N364)? mhpmcounter_q[180] : 
                (N366)? mhpmcounter_q[116] : 
                (N368)? mhpmcounter_q[52] : 1'b0;
  assign N218 = (N337)? mhpmcounter_q[2035] : 
                (N339)? mhpmcounter_q[1971] : 
                (N341)? mhpmcounter_q[1907] : 
                (N343)? mhpmcounter_q[1843] : 
                (N345)? mhpmcounter_q[1779] : 
                (N347)? mhpmcounter_q[1715] : 
                (N349)? mhpmcounter_q[1651] : 
                (N351)? mhpmcounter_q[1587] : 
                (N353)? mhpmcounter_q[1523] : 
                (N355)? mhpmcounter_q[1459] : 
                (N357)? mhpmcounter_q[1395] : 
                (N359)? mhpmcounter_q[1331] : 
                (N361)? mhpmcounter_q[1267] : 
                (N363)? mhpmcounter_q[1203] : 
                (N365)? mhpmcounter_q[1139] : 
                (N367)? mhpmcounter_q[1075] : 
                (N338)? mhpmcounter_q[1011] : 
                (N340)? mhpmcounter_q[947] : 
                (N342)? mhpmcounter_q[883] : 
                (N344)? mhpmcounter_q[819] : 
                (N346)? mhpmcounter_q[755] : 
                (N348)? mhpmcounter_q[691] : 
                (N350)? mhpmcounter_q[627] : 
                (N352)? mhpmcounter_q[563] : 
                (N354)? mhpmcounter_q[499] : 
                (N356)? mhpmcounter_q[435] : 
                (N358)? mhpmcounter_q[371] : 
                (N360)? mhpmcounter_q[307] : 
                (N362)? mhpmcounter_q[243] : 
                (N364)? mhpmcounter_q[179] : 
                (N366)? mhpmcounter_q[115] : 
                (N368)? mhpmcounter_q[51] : 1'b0;
  assign N219 = (N337)? mhpmcounter_q[2034] : 
                (N339)? mhpmcounter_q[1970] : 
                (N341)? mhpmcounter_q[1906] : 
                (N343)? mhpmcounter_q[1842] : 
                (N345)? mhpmcounter_q[1778] : 
                (N347)? mhpmcounter_q[1714] : 
                (N349)? mhpmcounter_q[1650] : 
                (N351)? mhpmcounter_q[1586] : 
                (N353)? mhpmcounter_q[1522] : 
                (N355)? mhpmcounter_q[1458] : 
                (N357)? mhpmcounter_q[1394] : 
                (N359)? mhpmcounter_q[1330] : 
                (N361)? mhpmcounter_q[1266] : 
                (N363)? mhpmcounter_q[1202] : 
                (N365)? mhpmcounter_q[1138] : 
                (N367)? mhpmcounter_q[1074] : 
                (N338)? mhpmcounter_q[1010] : 
                (N340)? mhpmcounter_q[946] : 
                (N342)? mhpmcounter_q[882] : 
                (N344)? mhpmcounter_q[818] : 
                (N346)? mhpmcounter_q[754] : 
                (N348)? mhpmcounter_q[690] : 
                (N350)? mhpmcounter_q[626] : 
                (N352)? mhpmcounter_q[562] : 
                (N354)? mhpmcounter_q[498] : 
                (N356)? mhpmcounter_q[434] : 
                (N358)? mhpmcounter_q[370] : 
                (N360)? mhpmcounter_q[306] : 
                (N362)? mhpmcounter_q[242] : 
                (N364)? mhpmcounter_q[178] : 
                (N366)? mhpmcounter_q[114] : 
                (N368)? mhpmcounter_q[50] : 1'b0;
  assign N220 = (N337)? mhpmcounter_q[2033] : 
                (N339)? mhpmcounter_q[1969] : 
                (N341)? mhpmcounter_q[1905] : 
                (N343)? mhpmcounter_q[1841] : 
                (N345)? mhpmcounter_q[1777] : 
                (N347)? mhpmcounter_q[1713] : 
                (N349)? mhpmcounter_q[1649] : 
                (N351)? mhpmcounter_q[1585] : 
                (N353)? mhpmcounter_q[1521] : 
                (N355)? mhpmcounter_q[1457] : 
                (N357)? mhpmcounter_q[1393] : 
                (N359)? mhpmcounter_q[1329] : 
                (N361)? mhpmcounter_q[1265] : 
                (N363)? mhpmcounter_q[1201] : 
                (N365)? mhpmcounter_q[1137] : 
                (N367)? mhpmcounter_q[1073] : 
                (N338)? mhpmcounter_q[1009] : 
                (N340)? mhpmcounter_q[945] : 
                (N342)? mhpmcounter_q[881] : 
                (N344)? mhpmcounter_q[817] : 
                (N346)? mhpmcounter_q[753] : 
                (N348)? mhpmcounter_q[689] : 
                (N350)? mhpmcounter_q[625] : 
                (N352)? mhpmcounter_q[561] : 
                (N354)? mhpmcounter_q[497] : 
                (N356)? mhpmcounter_q[433] : 
                (N358)? mhpmcounter_q[369] : 
                (N360)? mhpmcounter_q[305] : 
                (N362)? mhpmcounter_q[241] : 
                (N364)? mhpmcounter_q[177] : 
                (N366)? mhpmcounter_q[113] : 
                (N368)? mhpmcounter_q[49] : 1'b0;
  assign N221 = (N337)? mhpmcounter_q[2032] : 
                (N339)? mhpmcounter_q[1968] : 
                (N341)? mhpmcounter_q[1904] : 
                (N343)? mhpmcounter_q[1840] : 
                (N345)? mhpmcounter_q[1776] : 
                (N347)? mhpmcounter_q[1712] : 
                (N349)? mhpmcounter_q[1648] : 
                (N351)? mhpmcounter_q[1584] : 
                (N353)? mhpmcounter_q[1520] : 
                (N355)? mhpmcounter_q[1456] : 
                (N357)? mhpmcounter_q[1392] : 
                (N359)? mhpmcounter_q[1328] : 
                (N361)? mhpmcounter_q[1264] : 
                (N363)? mhpmcounter_q[1200] : 
                (N365)? mhpmcounter_q[1136] : 
                (N367)? mhpmcounter_q[1072] : 
                (N338)? mhpmcounter_q[1008] : 
                (N340)? mhpmcounter_q[944] : 
                (N342)? mhpmcounter_q[880] : 
                (N344)? mhpmcounter_q[816] : 
                (N346)? mhpmcounter_q[752] : 
                (N348)? mhpmcounter_q[688] : 
                (N350)? mhpmcounter_q[624] : 
                (N352)? mhpmcounter_q[560] : 
                (N354)? mhpmcounter_q[496] : 
                (N356)? mhpmcounter_q[432] : 
                (N358)? mhpmcounter_q[368] : 
                (N360)? mhpmcounter_q[304] : 
                (N362)? mhpmcounter_q[240] : 
                (N364)? mhpmcounter_q[176] : 
                (N366)? mhpmcounter_q[112] : 
                (N368)? mhpmcounter_q[48] : 1'b0;
  assign N222 = (N337)? mhpmcounter_q[2031] : 
                (N339)? mhpmcounter_q[1967] : 
                (N341)? mhpmcounter_q[1903] : 
                (N343)? mhpmcounter_q[1839] : 
                (N345)? mhpmcounter_q[1775] : 
                (N347)? mhpmcounter_q[1711] : 
                (N349)? mhpmcounter_q[1647] : 
                (N351)? mhpmcounter_q[1583] : 
                (N353)? mhpmcounter_q[1519] : 
                (N355)? mhpmcounter_q[1455] : 
                (N357)? mhpmcounter_q[1391] : 
                (N359)? mhpmcounter_q[1327] : 
                (N361)? mhpmcounter_q[1263] : 
                (N363)? mhpmcounter_q[1199] : 
                (N365)? mhpmcounter_q[1135] : 
                (N367)? mhpmcounter_q[1071] : 
                (N338)? mhpmcounter_q[1007] : 
                (N340)? mhpmcounter_q[943] : 
                (N342)? mhpmcounter_q[879] : 
                (N344)? mhpmcounter_q[815] : 
                (N346)? mhpmcounter_q[751] : 
                (N348)? mhpmcounter_q[687] : 
                (N350)? mhpmcounter_q[623] : 
                (N352)? mhpmcounter_q[559] : 
                (N354)? mhpmcounter_q[495] : 
                (N356)? mhpmcounter_q[431] : 
                (N358)? mhpmcounter_q[367] : 
                (N360)? mhpmcounter_q[303] : 
                (N362)? mhpmcounter_q[239] : 
                (N364)? mhpmcounter_q[175] : 
                (N366)? mhpmcounter_q[111] : 
                (N368)? mhpmcounter_q[47] : 1'b0;
  assign N223 = (N337)? mhpmcounter_q[2030] : 
                (N339)? mhpmcounter_q[1966] : 
                (N341)? mhpmcounter_q[1902] : 
                (N343)? mhpmcounter_q[1838] : 
                (N345)? mhpmcounter_q[1774] : 
                (N347)? mhpmcounter_q[1710] : 
                (N349)? mhpmcounter_q[1646] : 
                (N351)? mhpmcounter_q[1582] : 
                (N353)? mhpmcounter_q[1518] : 
                (N355)? mhpmcounter_q[1454] : 
                (N357)? mhpmcounter_q[1390] : 
                (N359)? mhpmcounter_q[1326] : 
                (N361)? mhpmcounter_q[1262] : 
                (N363)? mhpmcounter_q[1198] : 
                (N365)? mhpmcounter_q[1134] : 
                (N367)? mhpmcounter_q[1070] : 
                (N338)? mhpmcounter_q[1006] : 
                (N340)? mhpmcounter_q[942] : 
                (N342)? mhpmcounter_q[878] : 
                (N344)? mhpmcounter_q[814] : 
                (N346)? mhpmcounter_q[750] : 
                (N348)? mhpmcounter_q[686] : 
                (N350)? mhpmcounter_q[622] : 
                (N352)? mhpmcounter_q[558] : 
                (N354)? mhpmcounter_q[494] : 
                (N356)? mhpmcounter_q[430] : 
                (N358)? mhpmcounter_q[366] : 
                (N360)? mhpmcounter_q[302] : 
                (N362)? mhpmcounter_q[238] : 
                (N364)? mhpmcounter_q[174] : 
                (N366)? mhpmcounter_q[110] : 
                (N368)? mhpmcounter_q[46] : 1'b0;
  assign N224 = (N337)? mhpmcounter_q[2029] : 
                (N339)? mhpmcounter_q[1965] : 
                (N341)? mhpmcounter_q[1901] : 
                (N343)? mhpmcounter_q[1837] : 
                (N345)? mhpmcounter_q[1773] : 
                (N347)? mhpmcounter_q[1709] : 
                (N349)? mhpmcounter_q[1645] : 
                (N351)? mhpmcounter_q[1581] : 
                (N353)? mhpmcounter_q[1517] : 
                (N355)? mhpmcounter_q[1453] : 
                (N357)? mhpmcounter_q[1389] : 
                (N359)? mhpmcounter_q[1325] : 
                (N361)? mhpmcounter_q[1261] : 
                (N363)? mhpmcounter_q[1197] : 
                (N365)? mhpmcounter_q[1133] : 
                (N367)? mhpmcounter_q[1069] : 
                (N338)? mhpmcounter_q[1005] : 
                (N340)? mhpmcounter_q[941] : 
                (N342)? mhpmcounter_q[877] : 
                (N344)? mhpmcounter_q[813] : 
                (N346)? mhpmcounter_q[749] : 
                (N348)? mhpmcounter_q[685] : 
                (N350)? mhpmcounter_q[621] : 
                (N352)? mhpmcounter_q[557] : 
                (N354)? mhpmcounter_q[493] : 
                (N356)? mhpmcounter_q[429] : 
                (N358)? mhpmcounter_q[365] : 
                (N360)? mhpmcounter_q[301] : 
                (N362)? mhpmcounter_q[237] : 
                (N364)? mhpmcounter_q[173] : 
                (N366)? mhpmcounter_q[109] : 
                (N368)? mhpmcounter_q[45] : 1'b0;
  assign N225 = (N337)? mhpmcounter_q[2028] : 
                (N339)? mhpmcounter_q[1964] : 
                (N341)? mhpmcounter_q[1900] : 
                (N343)? mhpmcounter_q[1836] : 
                (N345)? mhpmcounter_q[1772] : 
                (N347)? mhpmcounter_q[1708] : 
                (N349)? mhpmcounter_q[1644] : 
                (N351)? mhpmcounter_q[1580] : 
                (N353)? mhpmcounter_q[1516] : 
                (N355)? mhpmcounter_q[1452] : 
                (N357)? mhpmcounter_q[1388] : 
                (N359)? mhpmcounter_q[1324] : 
                (N361)? mhpmcounter_q[1260] : 
                (N363)? mhpmcounter_q[1196] : 
                (N365)? mhpmcounter_q[1132] : 
                (N367)? mhpmcounter_q[1068] : 
                (N338)? mhpmcounter_q[1004] : 
                (N340)? mhpmcounter_q[940] : 
                (N342)? mhpmcounter_q[876] : 
                (N344)? mhpmcounter_q[812] : 
                (N346)? mhpmcounter_q[748] : 
                (N348)? mhpmcounter_q[684] : 
                (N350)? mhpmcounter_q[620] : 
                (N352)? mhpmcounter_q[556] : 
                (N354)? mhpmcounter_q[492] : 
                (N356)? mhpmcounter_q[428] : 
                (N358)? mhpmcounter_q[364] : 
                (N360)? mhpmcounter_q[300] : 
                (N362)? mhpmcounter_q[236] : 
                (N364)? mhpmcounter_q[172] : 
                (N366)? mhpmcounter_q[108] : 
                (N368)? mhpmcounter_q[44] : 1'b0;
  assign N226 = (N337)? mhpmcounter_q[2027] : 
                (N339)? mhpmcounter_q[1963] : 
                (N341)? mhpmcounter_q[1899] : 
                (N343)? mhpmcounter_q[1835] : 
                (N345)? mhpmcounter_q[1771] : 
                (N347)? mhpmcounter_q[1707] : 
                (N349)? mhpmcounter_q[1643] : 
                (N351)? mhpmcounter_q[1579] : 
                (N353)? mhpmcounter_q[1515] : 
                (N355)? mhpmcounter_q[1451] : 
                (N357)? mhpmcounter_q[1387] : 
                (N359)? mhpmcounter_q[1323] : 
                (N361)? mhpmcounter_q[1259] : 
                (N363)? mhpmcounter_q[1195] : 
                (N365)? mhpmcounter_q[1131] : 
                (N367)? mhpmcounter_q[1067] : 
                (N338)? mhpmcounter_q[1003] : 
                (N340)? mhpmcounter_q[939] : 
                (N342)? mhpmcounter_q[875] : 
                (N344)? mhpmcounter_q[811] : 
                (N346)? mhpmcounter_q[747] : 
                (N348)? mhpmcounter_q[683] : 
                (N350)? mhpmcounter_q[619] : 
                (N352)? mhpmcounter_q[555] : 
                (N354)? mhpmcounter_q[491] : 
                (N356)? mhpmcounter_q[427] : 
                (N358)? mhpmcounter_q[363] : 
                (N360)? mhpmcounter_q[299] : 
                (N362)? mhpmcounter_q[235] : 
                (N364)? mhpmcounter_q[171] : 
                (N366)? mhpmcounter_q[107] : 
                (N368)? mhpmcounter_q[43] : 1'b0;
  assign N227 = (N337)? mhpmcounter_q[2026] : 
                (N339)? mhpmcounter_q[1962] : 
                (N341)? mhpmcounter_q[1898] : 
                (N343)? mhpmcounter_q[1834] : 
                (N345)? mhpmcounter_q[1770] : 
                (N347)? mhpmcounter_q[1706] : 
                (N349)? mhpmcounter_q[1642] : 
                (N351)? mhpmcounter_q[1578] : 
                (N353)? mhpmcounter_q[1514] : 
                (N355)? mhpmcounter_q[1450] : 
                (N357)? mhpmcounter_q[1386] : 
                (N359)? mhpmcounter_q[1322] : 
                (N361)? mhpmcounter_q[1258] : 
                (N363)? mhpmcounter_q[1194] : 
                (N365)? mhpmcounter_q[1130] : 
                (N367)? mhpmcounter_q[1066] : 
                (N338)? mhpmcounter_q[1002] : 
                (N340)? mhpmcounter_q[938] : 
                (N342)? mhpmcounter_q[874] : 
                (N344)? mhpmcounter_q[810] : 
                (N346)? mhpmcounter_q[746] : 
                (N348)? mhpmcounter_q[682] : 
                (N350)? mhpmcounter_q[618] : 
                (N352)? mhpmcounter_q[554] : 
                (N354)? mhpmcounter_q[490] : 
                (N356)? mhpmcounter_q[426] : 
                (N358)? mhpmcounter_q[362] : 
                (N360)? mhpmcounter_q[298] : 
                (N362)? mhpmcounter_q[234] : 
                (N364)? mhpmcounter_q[170] : 
                (N366)? mhpmcounter_q[106] : 
                (N368)? mhpmcounter_q[42] : 1'b0;
  assign N228 = (N337)? mhpmcounter_q[2025] : 
                (N339)? mhpmcounter_q[1961] : 
                (N341)? mhpmcounter_q[1897] : 
                (N343)? mhpmcounter_q[1833] : 
                (N345)? mhpmcounter_q[1769] : 
                (N347)? mhpmcounter_q[1705] : 
                (N349)? mhpmcounter_q[1641] : 
                (N351)? mhpmcounter_q[1577] : 
                (N353)? mhpmcounter_q[1513] : 
                (N355)? mhpmcounter_q[1449] : 
                (N357)? mhpmcounter_q[1385] : 
                (N359)? mhpmcounter_q[1321] : 
                (N361)? mhpmcounter_q[1257] : 
                (N363)? mhpmcounter_q[1193] : 
                (N365)? mhpmcounter_q[1129] : 
                (N367)? mhpmcounter_q[1065] : 
                (N338)? mhpmcounter_q[1001] : 
                (N340)? mhpmcounter_q[937] : 
                (N342)? mhpmcounter_q[873] : 
                (N344)? mhpmcounter_q[809] : 
                (N346)? mhpmcounter_q[745] : 
                (N348)? mhpmcounter_q[681] : 
                (N350)? mhpmcounter_q[617] : 
                (N352)? mhpmcounter_q[553] : 
                (N354)? mhpmcounter_q[489] : 
                (N356)? mhpmcounter_q[425] : 
                (N358)? mhpmcounter_q[361] : 
                (N360)? mhpmcounter_q[297] : 
                (N362)? mhpmcounter_q[233] : 
                (N364)? mhpmcounter_q[169] : 
                (N366)? mhpmcounter_q[105] : 
                (N368)? mhpmcounter_q[41] : 1'b0;
  assign N229 = (N337)? mhpmcounter_q[2024] : 
                (N339)? mhpmcounter_q[1960] : 
                (N341)? mhpmcounter_q[1896] : 
                (N343)? mhpmcounter_q[1832] : 
                (N345)? mhpmcounter_q[1768] : 
                (N347)? mhpmcounter_q[1704] : 
                (N349)? mhpmcounter_q[1640] : 
                (N351)? mhpmcounter_q[1576] : 
                (N353)? mhpmcounter_q[1512] : 
                (N355)? mhpmcounter_q[1448] : 
                (N357)? mhpmcounter_q[1384] : 
                (N359)? mhpmcounter_q[1320] : 
                (N361)? mhpmcounter_q[1256] : 
                (N363)? mhpmcounter_q[1192] : 
                (N365)? mhpmcounter_q[1128] : 
                (N367)? mhpmcounter_q[1064] : 
                (N338)? mhpmcounter_q[1000] : 
                (N340)? mhpmcounter_q[936] : 
                (N342)? mhpmcounter_q[872] : 
                (N344)? mhpmcounter_q[808] : 
                (N346)? mhpmcounter_q[744] : 
                (N348)? mhpmcounter_q[680] : 
                (N350)? mhpmcounter_q[616] : 
                (N352)? mhpmcounter_q[552] : 
                (N354)? mhpmcounter_q[488] : 
                (N356)? mhpmcounter_q[424] : 
                (N358)? mhpmcounter_q[360] : 
                (N360)? mhpmcounter_q[296] : 
                (N362)? mhpmcounter_q[232] : 
                (N364)? mhpmcounter_q[168] : 
                (N366)? mhpmcounter_q[104] : 
                (N368)? mhpmcounter_q[40] : 1'b0;
  assign N230 = (N337)? mhpmcounter_q[2023] : 
                (N339)? mhpmcounter_q[1959] : 
                (N341)? mhpmcounter_q[1895] : 
                (N343)? mhpmcounter_q[1831] : 
                (N345)? mhpmcounter_q[1767] : 
                (N347)? mhpmcounter_q[1703] : 
                (N349)? mhpmcounter_q[1639] : 
                (N351)? mhpmcounter_q[1575] : 
                (N353)? mhpmcounter_q[1511] : 
                (N355)? mhpmcounter_q[1447] : 
                (N357)? mhpmcounter_q[1383] : 
                (N359)? mhpmcounter_q[1319] : 
                (N361)? mhpmcounter_q[1255] : 
                (N363)? mhpmcounter_q[1191] : 
                (N365)? mhpmcounter_q[1127] : 
                (N367)? mhpmcounter_q[1063] : 
                (N338)? mhpmcounter_q[999] : 
                (N340)? mhpmcounter_q[935] : 
                (N342)? mhpmcounter_q[871] : 
                (N344)? mhpmcounter_q[807] : 
                (N346)? mhpmcounter_q[743] : 
                (N348)? mhpmcounter_q[679] : 
                (N350)? mhpmcounter_q[615] : 
                (N352)? mhpmcounter_q[551] : 
                (N354)? mhpmcounter_q[487] : 
                (N356)? mhpmcounter_q[423] : 
                (N358)? mhpmcounter_q[359] : 
                (N360)? mhpmcounter_q[295] : 
                (N362)? mhpmcounter_q[231] : 
                (N364)? mhpmcounter_q[167] : 
                (N366)? mhpmcounter_q[103] : 
                (N368)? mhpmcounter_q[39] : 1'b0;
  assign N231 = (N337)? mhpmcounter_q[2022] : 
                (N339)? mhpmcounter_q[1958] : 
                (N341)? mhpmcounter_q[1894] : 
                (N343)? mhpmcounter_q[1830] : 
                (N345)? mhpmcounter_q[1766] : 
                (N347)? mhpmcounter_q[1702] : 
                (N349)? mhpmcounter_q[1638] : 
                (N351)? mhpmcounter_q[1574] : 
                (N353)? mhpmcounter_q[1510] : 
                (N355)? mhpmcounter_q[1446] : 
                (N357)? mhpmcounter_q[1382] : 
                (N359)? mhpmcounter_q[1318] : 
                (N361)? mhpmcounter_q[1254] : 
                (N363)? mhpmcounter_q[1190] : 
                (N365)? mhpmcounter_q[1126] : 
                (N367)? mhpmcounter_q[1062] : 
                (N338)? mhpmcounter_q[998] : 
                (N340)? mhpmcounter_q[934] : 
                (N342)? mhpmcounter_q[870] : 
                (N344)? mhpmcounter_q[806] : 
                (N346)? mhpmcounter_q[742] : 
                (N348)? mhpmcounter_q[678] : 
                (N350)? mhpmcounter_q[614] : 
                (N352)? mhpmcounter_q[550] : 
                (N354)? mhpmcounter_q[486] : 
                (N356)? mhpmcounter_q[422] : 
                (N358)? mhpmcounter_q[358] : 
                (N360)? mhpmcounter_q[294] : 
                (N362)? mhpmcounter_q[230] : 
                (N364)? mhpmcounter_q[166] : 
                (N366)? mhpmcounter_q[102] : 
                (N368)? mhpmcounter_q[38] : 1'b0;
  assign N232 = (N337)? mhpmcounter_q[2021] : 
                (N339)? mhpmcounter_q[1957] : 
                (N341)? mhpmcounter_q[1893] : 
                (N343)? mhpmcounter_q[1829] : 
                (N345)? mhpmcounter_q[1765] : 
                (N347)? mhpmcounter_q[1701] : 
                (N349)? mhpmcounter_q[1637] : 
                (N351)? mhpmcounter_q[1573] : 
                (N353)? mhpmcounter_q[1509] : 
                (N355)? mhpmcounter_q[1445] : 
                (N357)? mhpmcounter_q[1381] : 
                (N359)? mhpmcounter_q[1317] : 
                (N361)? mhpmcounter_q[1253] : 
                (N363)? mhpmcounter_q[1189] : 
                (N365)? mhpmcounter_q[1125] : 
                (N367)? mhpmcounter_q[1061] : 
                (N338)? mhpmcounter_q[997] : 
                (N340)? mhpmcounter_q[933] : 
                (N342)? mhpmcounter_q[869] : 
                (N344)? mhpmcounter_q[805] : 
                (N346)? mhpmcounter_q[741] : 
                (N348)? mhpmcounter_q[677] : 
                (N350)? mhpmcounter_q[613] : 
                (N352)? mhpmcounter_q[549] : 
                (N354)? mhpmcounter_q[485] : 
                (N356)? mhpmcounter_q[421] : 
                (N358)? mhpmcounter_q[357] : 
                (N360)? mhpmcounter_q[293] : 
                (N362)? mhpmcounter_q[229] : 
                (N364)? mhpmcounter_q[165] : 
                (N366)? mhpmcounter_q[101] : 
                (N368)? mhpmcounter_q[37] : 1'b0;
  assign N233 = (N337)? mhpmcounter_q[2020] : 
                (N339)? mhpmcounter_q[1956] : 
                (N341)? mhpmcounter_q[1892] : 
                (N343)? mhpmcounter_q[1828] : 
                (N345)? mhpmcounter_q[1764] : 
                (N347)? mhpmcounter_q[1700] : 
                (N349)? mhpmcounter_q[1636] : 
                (N351)? mhpmcounter_q[1572] : 
                (N353)? mhpmcounter_q[1508] : 
                (N355)? mhpmcounter_q[1444] : 
                (N357)? mhpmcounter_q[1380] : 
                (N359)? mhpmcounter_q[1316] : 
                (N361)? mhpmcounter_q[1252] : 
                (N363)? mhpmcounter_q[1188] : 
                (N365)? mhpmcounter_q[1124] : 
                (N367)? mhpmcounter_q[1060] : 
                (N338)? mhpmcounter_q[996] : 
                (N340)? mhpmcounter_q[932] : 
                (N342)? mhpmcounter_q[868] : 
                (N344)? mhpmcounter_q[804] : 
                (N346)? mhpmcounter_q[740] : 
                (N348)? mhpmcounter_q[676] : 
                (N350)? mhpmcounter_q[612] : 
                (N352)? mhpmcounter_q[548] : 
                (N354)? mhpmcounter_q[484] : 
                (N356)? mhpmcounter_q[420] : 
                (N358)? mhpmcounter_q[356] : 
                (N360)? mhpmcounter_q[292] : 
                (N362)? mhpmcounter_q[228] : 
                (N364)? mhpmcounter_q[164] : 
                (N366)? mhpmcounter_q[100] : 
                (N368)? mhpmcounter_q[36] : 1'b0;
  assign N234 = (N337)? mhpmcounter_q[2019] : 
                (N339)? mhpmcounter_q[1955] : 
                (N341)? mhpmcounter_q[1891] : 
                (N343)? mhpmcounter_q[1827] : 
                (N345)? mhpmcounter_q[1763] : 
                (N347)? mhpmcounter_q[1699] : 
                (N349)? mhpmcounter_q[1635] : 
                (N351)? mhpmcounter_q[1571] : 
                (N353)? mhpmcounter_q[1507] : 
                (N355)? mhpmcounter_q[1443] : 
                (N357)? mhpmcounter_q[1379] : 
                (N359)? mhpmcounter_q[1315] : 
                (N361)? mhpmcounter_q[1251] : 
                (N363)? mhpmcounter_q[1187] : 
                (N365)? mhpmcounter_q[1123] : 
                (N367)? mhpmcounter_q[1059] : 
                (N338)? mhpmcounter_q[995] : 
                (N340)? mhpmcounter_q[931] : 
                (N342)? mhpmcounter_q[867] : 
                (N344)? mhpmcounter_q[803] : 
                (N346)? mhpmcounter_q[739] : 
                (N348)? mhpmcounter_q[675] : 
                (N350)? mhpmcounter_q[611] : 
                (N352)? mhpmcounter_q[547] : 
                (N354)? mhpmcounter_q[483] : 
                (N356)? mhpmcounter_q[419] : 
                (N358)? mhpmcounter_q[355] : 
                (N360)? mhpmcounter_q[291] : 
                (N362)? mhpmcounter_q[227] : 
                (N364)? mhpmcounter_q[163] : 
                (N366)? mhpmcounter_q[99] : 
                (N368)? mhpmcounter_q[35] : 1'b0;
  assign N235 = (N337)? mhpmcounter_q[2018] : 
                (N339)? mhpmcounter_q[1954] : 
                (N341)? mhpmcounter_q[1890] : 
                (N343)? mhpmcounter_q[1826] : 
                (N345)? mhpmcounter_q[1762] : 
                (N347)? mhpmcounter_q[1698] : 
                (N349)? mhpmcounter_q[1634] : 
                (N351)? mhpmcounter_q[1570] : 
                (N353)? mhpmcounter_q[1506] : 
                (N355)? mhpmcounter_q[1442] : 
                (N357)? mhpmcounter_q[1378] : 
                (N359)? mhpmcounter_q[1314] : 
                (N361)? mhpmcounter_q[1250] : 
                (N363)? mhpmcounter_q[1186] : 
                (N365)? mhpmcounter_q[1122] : 
                (N367)? mhpmcounter_q[1058] : 
                (N338)? mhpmcounter_q[994] : 
                (N340)? mhpmcounter_q[930] : 
                (N342)? mhpmcounter_q[866] : 
                (N344)? mhpmcounter_q[802] : 
                (N346)? mhpmcounter_q[738] : 
                (N348)? mhpmcounter_q[674] : 
                (N350)? mhpmcounter_q[610] : 
                (N352)? mhpmcounter_q[546] : 
                (N354)? mhpmcounter_q[482] : 
                (N356)? mhpmcounter_q[418] : 
                (N358)? mhpmcounter_q[354] : 
                (N360)? mhpmcounter_q[290] : 
                (N362)? mhpmcounter_q[226] : 
                (N364)? mhpmcounter_q[162] : 
                (N366)? mhpmcounter_q[98] : 
                (N368)? mhpmcounter_q[34] : 1'b0;
  assign N236 = (N337)? mhpmcounter_q[2017] : 
                (N339)? mhpmcounter_q[1953] : 
                (N341)? mhpmcounter_q[1889] : 
                (N343)? mhpmcounter_q[1825] : 
                (N345)? mhpmcounter_q[1761] : 
                (N347)? mhpmcounter_q[1697] : 
                (N349)? mhpmcounter_q[1633] : 
                (N351)? mhpmcounter_q[1569] : 
                (N353)? mhpmcounter_q[1505] : 
                (N355)? mhpmcounter_q[1441] : 
                (N357)? mhpmcounter_q[1377] : 
                (N359)? mhpmcounter_q[1313] : 
                (N361)? mhpmcounter_q[1249] : 
                (N363)? mhpmcounter_q[1185] : 
                (N365)? mhpmcounter_q[1121] : 
                (N367)? mhpmcounter_q[1057] : 
                (N338)? mhpmcounter_q[993] : 
                (N340)? mhpmcounter_q[929] : 
                (N342)? mhpmcounter_q[865] : 
                (N344)? mhpmcounter_q[801] : 
                (N346)? mhpmcounter_q[737] : 
                (N348)? mhpmcounter_q[673] : 
                (N350)? mhpmcounter_q[609] : 
                (N352)? mhpmcounter_q[545] : 
                (N354)? mhpmcounter_q[481] : 
                (N356)? mhpmcounter_q[417] : 
                (N358)? mhpmcounter_q[353] : 
                (N360)? mhpmcounter_q[289] : 
                (N362)? mhpmcounter_q[225] : 
                (N364)? mhpmcounter_q[161] : 
                (N366)? mhpmcounter_q[97] : 
                (N368)? mhpmcounter_q[33] : 1'b0;
  assign N237 = (N337)? mhpmcounter_q[2016] : 
                (N339)? mhpmcounter_q[1952] : 
                (N341)? mhpmcounter_q[1888] : 
                (N343)? mhpmcounter_q[1824] : 
                (N345)? mhpmcounter_q[1760] : 
                (N347)? mhpmcounter_q[1696] : 
                (N349)? mhpmcounter_q[1632] : 
                (N351)? mhpmcounter_q[1568] : 
                (N353)? mhpmcounter_q[1504] : 
                (N355)? mhpmcounter_q[1440] : 
                (N357)? mhpmcounter_q[1376] : 
                (N359)? mhpmcounter_q[1312] : 
                (N361)? mhpmcounter_q[1248] : 
                (N363)? mhpmcounter_q[1184] : 
                (N365)? mhpmcounter_q[1120] : 
                (N367)? mhpmcounter_q[1056] : 
                (N338)? mhpmcounter_q[992] : 
                (N340)? mhpmcounter_q[928] : 
                (N342)? mhpmcounter_q[864] : 
                (N344)? mhpmcounter_q[800] : 
                (N346)? mhpmcounter_q[736] : 
                (N348)? mhpmcounter_q[672] : 
                (N350)? mhpmcounter_q[608] : 
                (N352)? mhpmcounter_q[544] : 
                (N354)? mhpmcounter_q[480] : 
                (N356)? mhpmcounter_q[416] : 
                (N358)? mhpmcounter_q[352] : 
                (N360)? mhpmcounter_q[288] : 
                (N362)? mhpmcounter_q[224] : 
                (N364)? mhpmcounter_q[160] : 
                (N366)? mhpmcounter_q[96] : 
                (N368)? mhpmcounter_q[32] : 1'b0;
  assign N238 = (N337)? mhpmcounter_q[2015] : 
                (N339)? mhpmcounter_q[1951] : 
                (N341)? mhpmcounter_q[1887] : 
                (N343)? mhpmcounter_q[1823] : 
                (N345)? mhpmcounter_q[1759] : 
                (N347)? mhpmcounter_q[1695] : 
                (N349)? mhpmcounter_q[1631] : 
                (N351)? mhpmcounter_q[1567] : 
                (N353)? mhpmcounter_q[1503] : 
                (N355)? mhpmcounter_q[1439] : 
                (N357)? mhpmcounter_q[1375] : 
                (N359)? mhpmcounter_q[1311] : 
                (N361)? mhpmcounter_q[1247] : 
                (N363)? mhpmcounter_q[1183] : 
                (N365)? mhpmcounter_q[1119] : 
                (N367)? mhpmcounter_q[1055] : 
                (N338)? mhpmcounter_q[991] : 
                (N340)? mhpmcounter_q[927] : 
                (N342)? mhpmcounter_q[863] : 
                (N344)? mhpmcounter_q[799] : 
                (N346)? mhpmcounter_q[735] : 
                (N348)? mhpmcounter_q[671] : 
                (N350)? mhpmcounter_q[607] : 
                (N352)? mhpmcounter_q[543] : 
                (N354)? mhpmcounter_q[479] : 
                (N356)? mhpmcounter_q[415] : 
                (N358)? mhpmcounter_q[351] : 
                (N360)? mhpmcounter_q[287] : 
                (N362)? mhpmcounter_q[223] : 
                (N364)? mhpmcounter_q[159] : 
                (N366)? mhpmcounter_q[95] : 
                (N368)? mhpmcounter_q[31] : 1'b0;
  assign N239 = (N337)? mhpmcounter_q[2014] : 
                (N339)? mhpmcounter_q[1950] : 
                (N341)? mhpmcounter_q[1886] : 
                (N343)? mhpmcounter_q[1822] : 
                (N345)? mhpmcounter_q[1758] : 
                (N347)? mhpmcounter_q[1694] : 
                (N349)? mhpmcounter_q[1630] : 
                (N351)? mhpmcounter_q[1566] : 
                (N353)? mhpmcounter_q[1502] : 
                (N355)? mhpmcounter_q[1438] : 
                (N357)? mhpmcounter_q[1374] : 
                (N359)? mhpmcounter_q[1310] : 
                (N361)? mhpmcounter_q[1246] : 
                (N363)? mhpmcounter_q[1182] : 
                (N365)? mhpmcounter_q[1118] : 
                (N367)? mhpmcounter_q[1054] : 
                (N338)? mhpmcounter_q[990] : 
                (N340)? mhpmcounter_q[926] : 
                (N342)? mhpmcounter_q[862] : 
                (N344)? mhpmcounter_q[798] : 
                (N346)? mhpmcounter_q[734] : 
                (N348)? mhpmcounter_q[670] : 
                (N350)? mhpmcounter_q[606] : 
                (N352)? mhpmcounter_q[542] : 
                (N354)? mhpmcounter_q[478] : 
                (N356)? mhpmcounter_q[414] : 
                (N358)? mhpmcounter_q[350] : 
                (N360)? mhpmcounter_q[286] : 
                (N362)? mhpmcounter_q[222] : 
                (N364)? mhpmcounter_q[158] : 
                (N366)? mhpmcounter_q[94] : 
                (N368)? mhpmcounter_q[30] : 1'b0;
  assign N240 = (N337)? mhpmcounter_q[2013] : 
                (N339)? mhpmcounter_q[1949] : 
                (N341)? mhpmcounter_q[1885] : 
                (N343)? mhpmcounter_q[1821] : 
                (N345)? mhpmcounter_q[1757] : 
                (N347)? mhpmcounter_q[1693] : 
                (N349)? mhpmcounter_q[1629] : 
                (N351)? mhpmcounter_q[1565] : 
                (N353)? mhpmcounter_q[1501] : 
                (N355)? mhpmcounter_q[1437] : 
                (N357)? mhpmcounter_q[1373] : 
                (N359)? mhpmcounter_q[1309] : 
                (N361)? mhpmcounter_q[1245] : 
                (N363)? mhpmcounter_q[1181] : 
                (N365)? mhpmcounter_q[1117] : 
                (N367)? mhpmcounter_q[1053] : 
                (N338)? mhpmcounter_q[989] : 
                (N340)? mhpmcounter_q[925] : 
                (N342)? mhpmcounter_q[861] : 
                (N344)? mhpmcounter_q[797] : 
                (N346)? mhpmcounter_q[733] : 
                (N348)? mhpmcounter_q[669] : 
                (N350)? mhpmcounter_q[605] : 
                (N352)? mhpmcounter_q[541] : 
                (N354)? mhpmcounter_q[477] : 
                (N356)? mhpmcounter_q[413] : 
                (N358)? mhpmcounter_q[349] : 
                (N360)? mhpmcounter_q[285] : 
                (N362)? mhpmcounter_q[221] : 
                (N364)? mhpmcounter_q[157] : 
                (N366)? mhpmcounter_q[93] : 
                (N368)? mhpmcounter_q[29] : 1'b0;
  assign N241 = (N337)? mhpmcounter_q[2012] : 
                (N339)? mhpmcounter_q[1948] : 
                (N341)? mhpmcounter_q[1884] : 
                (N343)? mhpmcounter_q[1820] : 
                (N345)? mhpmcounter_q[1756] : 
                (N347)? mhpmcounter_q[1692] : 
                (N349)? mhpmcounter_q[1628] : 
                (N351)? mhpmcounter_q[1564] : 
                (N353)? mhpmcounter_q[1500] : 
                (N355)? mhpmcounter_q[1436] : 
                (N357)? mhpmcounter_q[1372] : 
                (N359)? mhpmcounter_q[1308] : 
                (N361)? mhpmcounter_q[1244] : 
                (N363)? mhpmcounter_q[1180] : 
                (N365)? mhpmcounter_q[1116] : 
                (N367)? mhpmcounter_q[1052] : 
                (N338)? mhpmcounter_q[988] : 
                (N340)? mhpmcounter_q[924] : 
                (N342)? mhpmcounter_q[860] : 
                (N344)? mhpmcounter_q[796] : 
                (N346)? mhpmcounter_q[732] : 
                (N348)? mhpmcounter_q[668] : 
                (N350)? mhpmcounter_q[604] : 
                (N352)? mhpmcounter_q[540] : 
                (N354)? mhpmcounter_q[476] : 
                (N356)? mhpmcounter_q[412] : 
                (N358)? mhpmcounter_q[348] : 
                (N360)? mhpmcounter_q[284] : 
                (N362)? mhpmcounter_q[220] : 
                (N364)? mhpmcounter_q[156] : 
                (N366)? mhpmcounter_q[92] : 
                (N368)? mhpmcounter_q[28] : 1'b0;
  assign N242 = (N337)? mhpmcounter_q[2011] : 
                (N339)? mhpmcounter_q[1947] : 
                (N341)? mhpmcounter_q[1883] : 
                (N343)? mhpmcounter_q[1819] : 
                (N345)? mhpmcounter_q[1755] : 
                (N347)? mhpmcounter_q[1691] : 
                (N349)? mhpmcounter_q[1627] : 
                (N351)? mhpmcounter_q[1563] : 
                (N353)? mhpmcounter_q[1499] : 
                (N355)? mhpmcounter_q[1435] : 
                (N357)? mhpmcounter_q[1371] : 
                (N359)? mhpmcounter_q[1307] : 
                (N361)? mhpmcounter_q[1243] : 
                (N363)? mhpmcounter_q[1179] : 
                (N365)? mhpmcounter_q[1115] : 
                (N367)? mhpmcounter_q[1051] : 
                (N338)? mhpmcounter_q[987] : 
                (N340)? mhpmcounter_q[923] : 
                (N342)? mhpmcounter_q[859] : 
                (N344)? mhpmcounter_q[795] : 
                (N346)? mhpmcounter_q[731] : 
                (N348)? mhpmcounter_q[667] : 
                (N350)? mhpmcounter_q[603] : 
                (N352)? mhpmcounter_q[539] : 
                (N354)? mhpmcounter_q[475] : 
                (N356)? mhpmcounter_q[411] : 
                (N358)? mhpmcounter_q[347] : 
                (N360)? mhpmcounter_q[283] : 
                (N362)? mhpmcounter_q[219] : 
                (N364)? mhpmcounter_q[155] : 
                (N366)? mhpmcounter_q[91] : 
                (N368)? mhpmcounter_q[27] : 1'b0;
  assign N243 = (N337)? mhpmcounter_q[2010] : 
                (N339)? mhpmcounter_q[1946] : 
                (N341)? mhpmcounter_q[1882] : 
                (N343)? mhpmcounter_q[1818] : 
                (N345)? mhpmcounter_q[1754] : 
                (N347)? mhpmcounter_q[1690] : 
                (N349)? mhpmcounter_q[1626] : 
                (N351)? mhpmcounter_q[1562] : 
                (N353)? mhpmcounter_q[1498] : 
                (N355)? mhpmcounter_q[1434] : 
                (N357)? mhpmcounter_q[1370] : 
                (N359)? mhpmcounter_q[1306] : 
                (N361)? mhpmcounter_q[1242] : 
                (N363)? mhpmcounter_q[1178] : 
                (N365)? mhpmcounter_q[1114] : 
                (N367)? mhpmcounter_q[1050] : 
                (N338)? mhpmcounter_q[986] : 
                (N340)? mhpmcounter_q[922] : 
                (N342)? mhpmcounter_q[858] : 
                (N344)? mhpmcounter_q[794] : 
                (N346)? mhpmcounter_q[730] : 
                (N348)? mhpmcounter_q[666] : 
                (N350)? mhpmcounter_q[602] : 
                (N352)? mhpmcounter_q[538] : 
                (N354)? mhpmcounter_q[474] : 
                (N356)? mhpmcounter_q[410] : 
                (N358)? mhpmcounter_q[346] : 
                (N360)? mhpmcounter_q[282] : 
                (N362)? mhpmcounter_q[218] : 
                (N364)? mhpmcounter_q[154] : 
                (N366)? mhpmcounter_q[90] : 
                (N368)? mhpmcounter_q[26] : 1'b0;
  assign N244 = (N337)? mhpmcounter_q[2009] : 
                (N339)? mhpmcounter_q[1945] : 
                (N341)? mhpmcounter_q[1881] : 
                (N343)? mhpmcounter_q[1817] : 
                (N345)? mhpmcounter_q[1753] : 
                (N347)? mhpmcounter_q[1689] : 
                (N349)? mhpmcounter_q[1625] : 
                (N351)? mhpmcounter_q[1561] : 
                (N353)? mhpmcounter_q[1497] : 
                (N355)? mhpmcounter_q[1433] : 
                (N357)? mhpmcounter_q[1369] : 
                (N359)? mhpmcounter_q[1305] : 
                (N361)? mhpmcounter_q[1241] : 
                (N363)? mhpmcounter_q[1177] : 
                (N365)? mhpmcounter_q[1113] : 
                (N367)? mhpmcounter_q[1049] : 
                (N338)? mhpmcounter_q[985] : 
                (N340)? mhpmcounter_q[921] : 
                (N342)? mhpmcounter_q[857] : 
                (N344)? mhpmcounter_q[793] : 
                (N346)? mhpmcounter_q[729] : 
                (N348)? mhpmcounter_q[665] : 
                (N350)? mhpmcounter_q[601] : 
                (N352)? mhpmcounter_q[537] : 
                (N354)? mhpmcounter_q[473] : 
                (N356)? mhpmcounter_q[409] : 
                (N358)? mhpmcounter_q[345] : 
                (N360)? mhpmcounter_q[281] : 
                (N362)? mhpmcounter_q[217] : 
                (N364)? mhpmcounter_q[153] : 
                (N366)? mhpmcounter_q[89] : 
                (N368)? mhpmcounter_q[25] : 1'b0;
  assign N245 = (N337)? mhpmcounter_q[2008] : 
                (N339)? mhpmcounter_q[1944] : 
                (N341)? mhpmcounter_q[1880] : 
                (N343)? mhpmcounter_q[1816] : 
                (N345)? mhpmcounter_q[1752] : 
                (N347)? mhpmcounter_q[1688] : 
                (N349)? mhpmcounter_q[1624] : 
                (N351)? mhpmcounter_q[1560] : 
                (N353)? mhpmcounter_q[1496] : 
                (N355)? mhpmcounter_q[1432] : 
                (N357)? mhpmcounter_q[1368] : 
                (N359)? mhpmcounter_q[1304] : 
                (N361)? mhpmcounter_q[1240] : 
                (N363)? mhpmcounter_q[1176] : 
                (N365)? mhpmcounter_q[1112] : 
                (N367)? mhpmcounter_q[1048] : 
                (N338)? mhpmcounter_q[984] : 
                (N340)? mhpmcounter_q[920] : 
                (N342)? mhpmcounter_q[856] : 
                (N344)? mhpmcounter_q[792] : 
                (N346)? mhpmcounter_q[728] : 
                (N348)? mhpmcounter_q[664] : 
                (N350)? mhpmcounter_q[600] : 
                (N352)? mhpmcounter_q[536] : 
                (N354)? mhpmcounter_q[472] : 
                (N356)? mhpmcounter_q[408] : 
                (N358)? mhpmcounter_q[344] : 
                (N360)? mhpmcounter_q[280] : 
                (N362)? mhpmcounter_q[216] : 
                (N364)? mhpmcounter_q[152] : 
                (N366)? mhpmcounter_q[88] : 
                (N368)? mhpmcounter_q[24] : 1'b0;
  assign N246 = (N337)? mhpmcounter_q[2007] : 
                (N339)? mhpmcounter_q[1943] : 
                (N341)? mhpmcounter_q[1879] : 
                (N343)? mhpmcounter_q[1815] : 
                (N345)? mhpmcounter_q[1751] : 
                (N347)? mhpmcounter_q[1687] : 
                (N349)? mhpmcounter_q[1623] : 
                (N351)? mhpmcounter_q[1559] : 
                (N353)? mhpmcounter_q[1495] : 
                (N355)? mhpmcounter_q[1431] : 
                (N357)? mhpmcounter_q[1367] : 
                (N359)? mhpmcounter_q[1303] : 
                (N361)? mhpmcounter_q[1239] : 
                (N363)? mhpmcounter_q[1175] : 
                (N365)? mhpmcounter_q[1111] : 
                (N367)? mhpmcounter_q[1047] : 
                (N338)? mhpmcounter_q[983] : 
                (N340)? mhpmcounter_q[919] : 
                (N342)? mhpmcounter_q[855] : 
                (N344)? mhpmcounter_q[791] : 
                (N346)? mhpmcounter_q[727] : 
                (N348)? mhpmcounter_q[663] : 
                (N350)? mhpmcounter_q[599] : 
                (N352)? mhpmcounter_q[535] : 
                (N354)? mhpmcounter_q[471] : 
                (N356)? mhpmcounter_q[407] : 
                (N358)? mhpmcounter_q[343] : 
                (N360)? mhpmcounter_q[279] : 
                (N362)? mhpmcounter_q[215] : 
                (N364)? mhpmcounter_q[151] : 
                (N366)? mhpmcounter_q[87] : 
                (N368)? mhpmcounter_q[23] : 1'b0;
  assign N247 = (N337)? mhpmcounter_q[2006] : 
                (N339)? mhpmcounter_q[1942] : 
                (N341)? mhpmcounter_q[1878] : 
                (N343)? mhpmcounter_q[1814] : 
                (N345)? mhpmcounter_q[1750] : 
                (N347)? mhpmcounter_q[1686] : 
                (N349)? mhpmcounter_q[1622] : 
                (N351)? mhpmcounter_q[1558] : 
                (N353)? mhpmcounter_q[1494] : 
                (N355)? mhpmcounter_q[1430] : 
                (N357)? mhpmcounter_q[1366] : 
                (N359)? mhpmcounter_q[1302] : 
                (N361)? mhpmcounter_q[1238] : 
                (N363)? mhpmcounter_q[1174] : 
                (N365)? mhpmcounter_q[1110] : 
                (N367)? mhpmcounter_q[1046] : 
                (N338)? mhpmcounter_q[982] : 
                (N340)? mhpmcounter_q[918] : 
                (N342)? mhpmcounter_q[854] : 
                (N344)? mhpmcounter_q[790] : 
                (N346)? mhpmcounter_q[726] : 
                (N348)? mhpmcounter_q[662] : 
                (N350)? mhpmcounter_q[598] : 
                (N352)? mhpmcounter_q[534] : 
                (N354)? mhpmcounter_q[470] : 
                (N356)? mhpmcounter_q[406] : 
                (N358)? mhpmcounter_q[342] : 
                (N360)? mhpmcounter_q[278] : 
                (N362)? mhpmcounter_q[214] : 
                (N364)? mhpmcounter_q[150] : 
                (N366)? mhpmcounter_q[86] : 
                (N368)? mhpmcounter_q[22] : 1'b0;
  assign N248 = (N337)? mhpmcounter_q[2005] : 
                (N339)? mhpmcounter_q[1941] : 
                (N341)? mhpmcounter_q[1877] : 
                (N343)? mhpmcounter_q[1813] : 
                (N345)? mhpmcounter_q[1749] : 
                (N347)? mhpmcounter_q[1685] : 
                (N349)? mhpmcounter_q[1621] : 
                (N351)? mhpmcounter_q[1557] : 
                (N353)? mhpmcounter_q[1493] : 
                (N355)? mhpmcounter_q[1429] : 
                (N357)? mhpmcounter_q[1365] : 
                (N359)? mhpmcounter_q[1301] : 
                (N361)? mhpmcounter_q[1237] : 
                (N363)? mhpmcounter_q[1173] : 
                (N365)? mhpmcounter_q[1109] : 
                (N367)? mhpmcounter_q[1045] : 
                (N338)? mhpmcounter_q[981] : 
                (N340)? mhpmcounter_q[917] : 
                (N342)? mhpmcounter_q[853] : 
                (N344)? mhpmcounter_q[789] : 
                (N346)? mhpmcounter_q[725] : 
                (N348)? mhpmcounter_q[661] : 
                (N350)? mhpmcounter_q[597] : 
                (N352)? mhpmcounter_q[533] : 
                (N354)? mhpmcounter_q[469] : 
                (N356)? mhpmcounter_q[405] : 
                (N358)? mhpmcounter_q[341] : 
                (N360)? mhpmcounter_q[277] : 
                (N362)? mhpmcounter_q[213] : 
                (N364)? mhpmcounter_q[149] : 
                (N366)? mhpmcounter_q[85] : 
                (N368)? mhpmcounter_q[21] : 1'b0;
  assign N249 = (N337)? mhpmcounter_q[2004] : 
                (N339)? mhpmcounter_q[1940] : 
                (N341)? mhpmcounter_q[1876] : 
                (N343)? mhpmcounter_q[1812] : 
                (N345)? mhpmcounter_q[1748] : 
                (N347)? mhpmcounter_q[1684] : 
                (N349)? mhpmcounter_q[1620] : 
                (N351)? mhpmcounter_q[1556] : 
                (N353)? mhpmcounter_q[1492] : 
                (N355)? mhpmcounter_q[1428] : 
                (N357)? mhpmcounter_q[1364] : 
                (N359)? mhpmcounter_q[1300] : 
                (N361)? mhpmcounter_q[1236] : 
                (N363)? mhpmcounter_q[1172] : 
                (N365)? mhpmcounter_q[1108] : 
                (N367)? mhpmcounter_q[1044] : 
                (N338)? mhpmcounter_q[980] : 
                (N340)? mhpmcounter_q[916] : 
                (N342)? mhpmcounter_q[852] : 
                (N344)? mhpmcounter_q[788] : 
                (N346)? mhpmcounter_q[724] : 
                (N348)? mhpmcounter_q[660] : 
                (N350)? mhpmcounter_q[596] : 
                (N352)? mhpmcounter_q[532] : 
                (N354)? mhpmcounter_q[468] : 
                (N356)? mhpmcounter_q[404] : 
                (N358)? mhpmcounter_q[340] : 
                (N360)? mhpmcounter_q[276] : 
                (N362)? mhpmcounter_q[212] : 
                (N364)? mhpmcounter_q[148] : 
                (N366)? mhpmcounter_q[84] : 
                (N368)? mhpmcounter_q[20] : 1'b0;
  assign N250 = (N337)? mhpmcounter_q[2003] : 
                (N339)? mhpmcounter_q[1939] : 
                (N341)? mhpmcounter_q[1875] : 
                (N343)? mhpmcounter_q[1811] : 
                (N345)? mhpmcounter_q[1747] : 
                (N347)? mhpmcounter_q[1683] : 
                (N349)? mhpmcounter_q[1619] : 
                (N351)? mhpmcounter_q[1555] : 
                (N353)? mhpmcounter_q[1491] : 
                (N355)? mhpmcounter_q[1427] : 
                (N357)? mhpmcounter_q[1363] : 
                (N359)? mhpmcounter_q[1299] : 
                (N361)? mhpmcounter_q[1235] : 
                (N363)? mhpmcounter_q[1171] : 
                (N365)? mhpmcounter_q[1107] : 
                (N367)? mhpmcounter_q[1043] : 
                (N338)? mhpmcounter_q[979] : 
                (N340)? mhpmcounter_q[915] : 
                (N342)? mhpmcounter_q[851] : 
                (N344)? mhpmcounter_q[787] : 
                (N346)? mhpmcounter_q[723] : 
                (N348)? mhpmcounter_q[659] : 
                (N350)? mhpmcounter_q[595] : 
                (N352)? mhpmcounter_q[531] : 
                (N354)? mhpmcounter_q[467] : 
                (N356)? mhpmcounter_q[403] : 
                (N358)? mhpmcounter_q[339] : 
                (N360)? mhpmcounter_q[275] : 
                (N362)? mhpmcounter_q[211] : 
                (N364)? mhpmcounter_q[147] : 
                (N366)? mhpmcounter_q[83] : 
                (N368)? mhpmcounter_q[19] : 1'b0;
  assign N251 = (N337)? mhpmcounter_q[2002] : 
                (N339)? mhpmcounter_q[1938] : 
                (N341)? mhpmcounter_q[1874] : 
                (N343)? mhpmcounter_q[1810] : 
                (N345)? mhpmcounter_q[1746] : 
                (N347)? mhpmcounter_q[1682] : 
                (N349)? mhpmcounter_q[1618] : 
                (N351)? mhpmcounter_q[1554] : 
                (N353)? mhpmcounter_q[1490] : 
                (N355)? mhpmcounter_q[1426] : 
                (N357)? mhpmcounter_q[1362] : 
                (N359)? mhpmcounter_q[1298] : 
                (N361)? mhpmcounter_q[1234] : 
                (N363)? mhpmcounter_q[1170] : 
                (N365)? mhpmcounter_q[1106] : 
                (N367)? mhpmcounter_q[1042] : 
                (N338)? mhpmcounter_q[978] : 
                (N340)? mhpmcounter_q[914] : 
                (N342)? mhpmcounter_q[850] : 
                (N344)? mhpmcounter_q[786] : 
                (N346)? mhpmcounter_q[722] : 
                (N348)? mhpmcounter_q[658] : 
                (N350)? mhpmcounter_q[594] : 
                (N352)? mhpmcounter_q[530] : 
                (N354)? mhpmcounter_q[466] : 
                (N356)? mhpmcounter_q[402] : 
                (N358)? mhpmcounter_q[338] : 
                (N360)? mhpmcounter_q[274] : 
                (N362)? mhpmcounter_q[210] : 
                (N364)? mhpmcounter_q[146] : 
                (N366)? mhpmcounter_q[82] : 
                (N368)? mhpmcounter_q[18] : 1'b0;
  assign N252 = (N337)? mhpmcounter_q[2001] : 
                (N339)? mhpmcounter_q[1937] : 
                (N341)? mhpmcounter_q[1873] : 
                (N343)? mhpmcounter_q[1809] : 
                (N345)? mhpmcounter_q[1745] : 
                (N347)? mhpmcounter_q[1681] : 
                (N349)? mhpmcounter_q[1617] : 
                (N351)? mhpmcounter_q[1553] : 
                (N353)? mhpmcounter_q[1489] : 
                (N355)? mhpmcounter_q[1425] : 
                (N357)? mhpmcounter_q[1361] : 
                (N359)? mhpmcounter_q[1297] : 
                (N361)? mhpmcounter_q[1233] : 
                (N363)? mhpmcounter_q[1169] : 
                (N365)? mhpmcounter_q[1105] : 
                (N367)? mhpmcounter_q[1041] : 
                (N338)? mhpmcounter_q[977] : 
                (N340)? mhpmcounter_q[913] : 
                (N342)? mhpmcounter_q[849] : 
                (N344)? mhpmcounter_q[785] : 
                (N346)? mhpmcounter_q[721] : 
                (N348)? mhpmcounter_q[657] : 
                (N350)? mhpmcounter_q[593] : 
                (N352)? mhpmcounter_q[529] : 
                (N354)? mhpmcounter_q[465] : 
                (N356)? mhpmcounter_q[401] : 
                (N358)? mhpmcounter_q[337] : 
                (N360)? mhpmcounter_q[273] : 
                (N362)? mhpmcounter_q[209] : 
                (N364)? mhpmcounter_q[145] : 
                (N366)? mhpmcounter_q[81] : 
                (N368)? mhpmcounter_q[17] : 1'b0;
  assign N253 = (N337)? mhpmcounter_q[2000] : 
                (N339)? mhpmcounter_q[1936] : 
                (N341)? mhpmcounter_q[1872] : 
                (N343)? mhpmcounter_q[1808] : 
                (N345)? mhpmcounter_q[1744] : 
                (N347)? mhpmcounter_q[1680] : 
                (N349)? mhpmcounter_q[1616] : 
                (N351)? mhpmcounter_q[1552] : 
                (N353)? mhpmcounter_q[1488] : 
                (N355)? mhpmcounter_q[1424] : 
                (N357)? mhpmcounter_q[1360] : 
                (N359)? mhpmcounter_q[1296] : 
                (N361)? mhpmcounter_q[1232] : 
                (N363)? mhpmcounter_q[1168] : 
                (N365)? mhpmcounter_q[1104] : 
                (N367)? mhpmcounter_q[1040] : 
                (N338)? mhpmcounter_q[976] : 
                (N340)? mhpmcounter_q[912] : 
                (N342)? mhpmcounter_q[848] : 
                (N344)? mhpmcounter_q[784] : 
                (N346)? mhpmcounter_q[720] : 
                (N348)? mhpmcounter_q[656] : 
                (N350)? mhpmcounter_q[592] : 
                (N352)? mhpmcounter_q[528] : 
                (N354)? mhpmcounter_q[464] : 
                (N356)? mhpmcounter_q[400] : 
                (N358)? mhpmcounter_q[336] : 
                (N360)? mhpmcounter_q[272] : 
                (N362)? mhpmcounter_q[208] : 
                (N364)? mhpmcounter_q[144] : 
                (N366)? mhpmcounter_q[80] : 
                (N368)? mhpmcounter_q[16] : 1'b0;
  assign N254 = (N337)? mhpmcounter_q[1999] : 
                (N339)? mhpmcounter_q[1935] : 
                (N341)? mhpmcounter_q[1871] : 
                (N343)? mhpmcounter_q[1807] : 
                (N345)? mhpmcounter_q[1743] : 
                (N347)? mhpmcounter_q[1679] : 
                (N349)? mhpmcounter_q[1615] : 
                (N351)? mhpmcounter_q[1551] : 
                (N353)? mhpmcounter_q[1487] : 
                (N355)? mhpmcounter_q[1423] : 
                (N357)? mhpmcounter_q[1359] : 
                (N359)? mhpmcounter_q[1295] : 
                (N361)? mhpmcounter_q[1231] : 
                (N363)? mhpmcounter_q[1167] : 
                (N365)? mhpmcounter_q[1103] : 
                (N367)? mhpmcounter_q[1039] : 
                (N338)? mhpmcounter_q[975] : 
                (N340)? mhpmcounter_q[911] : 
                (N342)? mhpmcounter_q[847] : 
                (N344)? mhpmcounter_q[783] : 
                (N346)? mhpmcounter_q[719] : 
                (N348)? mhpmcounter_q[655] : 
                (N350)? mhpmcounter_q[591] : 
                (N352)? mhpmcounter_q[527] : 
                (N354)? mhpmcounter_q[463] : 
                (N356)? mhpmcounter_q[399] : 
                (N358)? mhpmcounter_q[335] : 
                (N360)? mhpmcounter_q[271] : 
                (N362)? mhpmcounter_q[207] : 
                (N364)? mhpmcounter_q[143] : 
                (N366)? mhpmcounter_q[79] : 
                (N368)? mhpmcounter_q[15] : 1'b0;
  assign N255 = (N337)? mhpmcounter_q[1998] : 
                (N339)? mhpmcounter_q[1934] : 
                (N341)? mhpmcounter_q[1870] : 
                (N343)? mhpmcounter_q[1806] : 
                (N345)? mhpmcounter_q[1742] : 
                (N347)? mhpmcounter_q[1678] : 
                (N349)? mhpmcounter_q[1614] : 
                (N351)? mhpmcounter_q[1550] : 
                (N353)? mhpmcounter_q[1486] : 
                (N355)? mhpmcounter_q[1422] : 
                (N357)? mhpmcounter_q[1358] : 
                (N359)? mhpmcounter_q[1294] : 
                (N361)? mhpmcounter_q[1230] : 
                (N363)? mhpmcounter_q[1166] : 
                (N365)? mhpmcounter_q[1102] : 
                (N367)? mhpmcounter_q[1038] : 
                (N338)? mhpmcounter_q[974] : 
                (N340)? mhpmcounter_q[910] : 
                (N342)? mhpmcounter_q[846] : 
                (N344)? mhpmcounter_q[782] : 
                (N346)? mhpmcounter_q[718] : 
                (N348)? mhpmcounter_q[654] : 
                (N350)? mhpmcounter_q[590] : 
                (N352)? mhpmcounter_q[526] : 
                (N354)? mhpmcounter_q[462] : 
                (N356)? mhpmcounter_q[398] : 
                (N358)? mhpmcounter_q[334] : 
                (N360)? mhpmcounter_q[270] : 
                (N362)? mhpmcounter_q[206] : 
                (N364)? mhpmcounter_q[142] : 
                (N366)? mhpmcounter_q[78] : 
                (N368)? mhpmcounter_q[14] : 1'b0;
  assign N256 = (N337)? mhpmcounter_q[1997] : 
                (N339)? mhpmcounter_q[1933] : 
                (N341)? mhpmcounter_q[1869] : 
                (N343)? mhpmcounter_q[1805] : 
                (N345)? mhpmcounter_q[1741] : 
                (N347)? mhpmcounter_q[1677] : 
                (N349)? mhpmcounter_q[1613] : 
                (N351)? mhpmcounter_q[1549] : 
                (N353)? mhpmcounter_q[1485] : 
                (N355)? mhpmcounter_q[1421] : 
                (N357)? mhpmcounter_q[1357] : 
                (N359)? mhpmcounter_q[1293] : 
                (N361)? mhpmcounter_q[1229] : 
                (N363)? mhpmcounter_q[1165] : 
                (N365)? mhpmcounter_q[1101] : 
                (N367)? mhpmcounter_q[1037] : 
                (N338)? mhpmcounter_q[973] : 
                (N340)? mhpmcounter_q[909] : 
                (N342)? mhpmcounter_q[845] : 
                (N344)? mhpmcounter_q[781] : 
                (N346)? mhpmcounter_q[717] : 
                (N348)? mhpmcounter_q[653] : 
                (N350)? mhpmcounter_q[589] : 
                (N352)? mhpmcounter_q[525] : 
                (N354)? mhpmcounter_q[461] : 
                (N356)? mhpmcounter_q[397] : 
                (N358)? mhpmcounter_q[333] : 
                (N360)? mhpmcounter_q[269] : 
                (N362)? mhpmcounter_q[205] : 
                (N364)? mhpmcounter_q[141] : 
                (N366)? mhpmcounter_q[77] : 
                (N368)? mhpmcounter_q[13] : 1'b0;
  assign N257 = (N337)? mhpmcounter_q[1996] : 
                (N339)? mhpmcounter_q[1932] : 
                (N341)? mhpmcounter_q[1868] : 
                (N343)? mhpmcounter_q[1804] : 
                (N345)? mhpmcounter_q[1740] : 
                (N347)? mhpmcounter_q[1676] : 
                (N349)? mhpmcounter_q[1612] : 
                (N351)? mhpmcounter_q[1548] : 
                (N353)? mhpmcounter_q[1484] : 
                (N355)? mhpmcounter_q[1420] : 
                (N357)? mhpmcounter_q[1356] : 
                (N359)? mhpmcounter_q[1292] : 
                (N361)? mhpmcounter_q[1228] : 
                (N363)? mhpmcounter_q[1164] : 
                (N365)? mhpmcounter_q[1100] : 
                (N367)? mhpmcounter_q[1036] : 
                (N338)? mhpmcounter_q[972] : 
                (N340)? mhpmcounter_q[908] : 
                (N342)? mhpmcounter_q[844] : 
                (N344)? mhpmcounter_q[780] : 
                (N346)? mhpmcounter_q[716] : 
                (N348)? mhpmcounter_q[652] : 
                (N350)? mhpmcounter_q[588] : 
                (N352)? mhpmcounter_q[524] : 
                (N354)? mhpmcounter_q[460] : 
                (N356)? mhpmcounter_q[396] : 
                (N358)? mhpmcounter_q[332] : 
                (N360)? mhpmcounter_q[268] : 
                (N362)? mhpmcounter_q[204] : 
                (N364)? mhpmcounter_q[140] : 
                (N366)? mhpmcounter_q[76] : 
                (N368)? mhpmcounter_q[12] : 1'b0;
  assign N258 = (N337)? mhpmcounter_q[1995] : 
                (N339)? mhpmcounter_q[1931] : 
                (N341)? mhpmcounter_q[1867] : 
                (N343)? mhpmcounter_q[1803] : 
                (N345)? mhpmcounter_q[1739] : 
                (N347)? mhpmcounter_q[1675] : 
                (N349)? mhpmcounter_q[1611] : 
                (N351)? mhpmcounter_q[1547] : 
                (N353)? mhpmcounter_q[1483] : 
                (N355)? mhpmcounter_q[1419] : 
                (N357)? mhpmcounter_q[1355] : 
                (N359)? mhpmcounter_q[1291] : 
                (N361)? mhpmcounter_q[1227] : 
                (N363)? mhpmcounter_q[1163] : 
                (N365)? mhpmcounter_q[1099] : 
                (N367)? mhpmcounter_q[1035] : 
                (N338)? mhpmcounter_q[971] : 
                (N340)? mhpmcounter_q[907] : 
                (N342)? mhpmcounter_q[843] : 
                (N344)? mhpmcounter_q[779] : 
                (N346)? mhpmcounter_q[715] : 
                (N348)? mhpmcounter_q[651] : 
                (N350)? mhpmcounter_q[587] : 
                (N352)? mhpmcounter_q[523] : 
                (N354)? mhpmcounter_q[459] : 
                (N356)? mhpmcounter_q[395] : 
                (N358)? mhpmcounter_q[331] : 
                (N360)? mhpmcounter_q[267] : 
                (N362)? mhpmcounter_q[203] : 
                (N364)? mhpmcounter_q[139] : 
                (N366)? mhpmcounter_q[75] : 
                (N368)? mhpmcounter_q[11] : 1'b0;
  assign N259 = (N337)? mhpmcounter_q[1994] : 
                (N339)? mhpmcounter_q[1930] : 
                (N341)? mhpmcounter_q[1866] : 
                (N343)? mhpmcounter_q[1802] : 
                (N345)? mhpmcounter_q[1738] : 
                (N347)? mhpmcounter_q[1674] : 
                (N349)? mhpmcounter_q[1610] : 
                (N351)? mhpmcounter_q[1546] : 
                (N353)? mhpmcounter_q[1482] : 
                (N355)? mhpmcounter_q[1418] : 
                (N357)? mhpmcounter_q[1354] : 
                (N359)? mhpmcounter_q[1290] : 
                (N361)? mhpmcounter_q[1226] : 
                (N363)? mhpmcounter_q[1162] : 
                (N365)? mhpmcounter_q[1098] : 
                (N367)? mhpmcounter_q[1034] : 
                (N338)? mhpmcounter_q[970] : 
                (N340)? mhpmcounter_q[906] : 
                (N342)? mhpmcounter_q[842] : 
                (N344)? mhpmcounter_q[778] : 
                (N346)? mhpmcounter_q[714] : 
                (N348)? mhpmcounter_q[650] : 
                (N350)? mhpmcounter_q[586] : 
                (N352)? mhpmcounter_q[522] : 
                (N354)? mhpmcounter_q[458] : 
                (N356)? mhpmcounter_q[394] : 
                (N358)? mhpmcounter_q[330] : 
                (N360)? mhpmcounter_q[266] : 
                (N362)? mhpmcounter_q[202] : 
                (N364)? mhpmcounter_q[138] : 
                (N366)? mhpmcounter_q[74] : 
                (N368)? mhpmcounter_q[10] : 1'b0;
  assign N260 = (N337)? mhpmcounter_q[1993] : 
                (N339)? mhpmcounter_q[1929] : 
                (N341)? mhpmcounter_q[1865] : 
                (N343)? mhpmcounter_q[1801] : 
                (N345)? mhpmcounter_q[1737] : 
                (N347)? mhpmcounter_q[1673] : 
                (N349)? mhpmcounter_q[1609] : 
                (N351)? mhpmcounter_q[1545] : 
                (N353)? mhpmcounter_q[1481] : 
                (N355)? mhpmcounter_q[1417] : 
                (N357)? mhpmcounter_q[1353] : 
                (N359)? mhpmcounter_q[1289] : 
                (N361)? mhpmcounter_q[1225] : 
                (N363)? mhpmcounter_q[1161] : 
                (N365)? mhpmcounter_q[1097] : 
                (N367)? mhpmcounter_q[1033] : 
                (N338)? mhpmcounter_q[969] : 
                (N340)? mhpmcounter_q[905] : 
                (N342)? mhpmcounter_q[841] : 
                (N344)? mhpmcounter_q[777] : 
                (N346)? mhpmcounter_q[713] : 
                (N348)? mhpmcounter_q[649] : 
                (N350)? mhpmcounter_q[585] : 
                (N352)? mhpmcounter_q[521] : 
                (N354)? mhpmcounter_q[457] : 
                (N356)? mhpmcounter_q[393] : 
                (N358)? mhpmcounter_q[329] : 
                (N360)? mhpmcounter_q[265] : 
                (N362)? mhpmcounter_q[201] : 
                (N364)? mhpmcounter_q[137] : 
                (N366)? mhpmcounter_q[73] : 
                (N368)? mhpmcounter_q[9] : 1'b0;
  assign N261 = (N337)? mhpmcounter_q[1992] : 
                (N339)? mhpmcounter_q[1928] : 
                (N341)? mhpmcounter_q[1864] : 
                (N343)? mhpmcounter_q[1800] : 
                (N345)? mhpmcounter_q[1736] : 
                (N347)? mhpmcounter_q[1672] : 
                (N349)? mhpmcounter_q[1608] : 
                (N351)? mhpmcounter_q[1544] : 
                (N353)? mhpmcounter_q[1480] : 
                (N355)? mhpmcounter_q[1416] : 
                (N357)? mhpmcounter_q[1352] : 
                (N359)? mhpmcounter_q[1288] : 
                (N361)? mhpmcounter_q[1224] : 
                (N363)? mhpmcounter_q[1160] : 
                (N365)? mhpmcounter_q[1096] : 
                (N367)? mhpmcounter_q[1032] : 
                (N338)? mhpmcounter_q[968] : 
                (N340)? mhpmcounter_q[904] : 
                (N342)? mhpmcounter_q[840] : 
                (N344)? mhpmcounter_q[776] : 
                (N346)? mhpmcounter_q[712] : 
                (N348)? mhpmcounter_q[648] : 
                (N350)? mhpmcounter_q[584] : 
                (N352)? mhpmcounter_q[520] : 
                (N354)? mhpmcounter_q[456] : 
                (N356)? mhpmcounter_q[392] : 
                (N358)? mhpmcounter_q[328] : 
                (N360)? mhpmcounter_q[264] : 
                (N362)? mhpmcounter_q[200] : 
                (N364)? mhpmcounter_q[136] : 
                (N366)? mhpmcounter_q[72] : 
                (N368)? mhpmcounter_q[8] : 1'b0;
  assign N262 = (N337)? mhpmcounter_q[1991] : 
                (N339)? mhpmcounter_q[1927] : 
                (N341)? mhpmcounter_q[1863] : 
                (N343)? mhpmcounter_q[1799] : 
                (N345)? mhpmcounter_q[1735] : 
                (N347)? mhpmcounter_q[1671] : 
                (N349)? mhpmcounter_q[1607] : 
                (N351)? mhpmcounter_q[1543] : 
                (N353)? mhpmcounter_q[1479] : 
                (N355)? mhpmcounter_q[1415] : 
                (N357)? mhpmcounter_q[1351] : 
                (N359)? mhpmcounter_q[1287] : 
                (N361)? mhpmcounter_q[1223] : 
                (N363)? mhpmcounter_q[1159] : 
                (N365)? mhpmcounter_q[1095] : 
                (N367)? mhpmcounter_q[1031] : 
                (N338)? mhpmcounter_q[967] : 
                (N340)? mhpmcounter_q[903] : 
                (N342)? mhpmcounter_q[839] : 
                (N344)? mhpmcounter_q[775] : 
                (N346)? mhpmcounter_q[711] : 
                (N348)? mhpmcounter_q[647] : 
                (N350)? mhpmcounter_q[583] : 
                (N352)? mhpmcounter_q[519] : 
                (N354)? mhpmcounter_q[455] : 
                (N356)? mhpmcounter_q[391] : 
                (N358)? mhpmcounter_q[327] : 
                (N360)? mhpmcounter_q[263] : 
                (N362)? mhpmcounter_q[199] : 
                (N364)? mhpmcounter_q[135] : 
                (N366)? mhpmcounter_q[71] : 
                (N368)? mhpmcounter_q[7] : 1'b0;
  assign N263 = (N337)? mhpmcounter_q[1990] : 
                (N339)? mhpmcounter_q[1926] : 
                (N341)? mhpmcounter_q[1862] : 
                (N343)? mhpmcounter_q[1798] : 
                (N345)? mhpmcounter_q[1734] : 
                (N347)? mhpmcounter_q[1670] : 
                (N349)? mhpmcounter_q[1606] : 
                (N351)? mhpmcounter_q[1542] : 
                (N353)? mhpmcounter_q[1478] : 
                (N355)? mhpmcounter_q[1414] : 
                (N357)? mhpmcounter_q[1350] : 
                (N359)? mhpmcounter_q[1286] : 
                (N361)? mhpmcounter_q[1222] : 
                (N363)? mhpmcounter_q[1158] : 
                (N365)? mhpmcounter_q[1094] : 
                (N367)? mhpmcounter_q[1030] : 
                (N338)? mhpmcounter_q[966] : 
                (N340)? mhpmcounter_q[902] : 
                (N342)? mhpmcounter_q[838] : 
                (N344)? mhpmcounter_q[774] : 
                (N346)? mhpmcounter_q[710] : 
                (N348)? mhpmcounter_q[646] : 
                (N350)? mhpmcounter_q[582] : 
                (N352)? mhpmcounter_q[518] : 
                (N354)? mhpmcounter_q[454] : 
                (N356)? mhpmcounter_q[390] : 
                (N358)? mhpmcounter_q[326] : 
                (N360)? mhpmcounter_q[262] : 
                (N362)? mhpmcounter_q[198] : 
                (N364)? mhpmcounter_q[134] : 
                (N366)? mhpmcounter_q[70] : 
                (N368)? mhpmcounter_q[6] : 1'b0;
  assign N264 = (N337)? mhpmcounter_q[1989] : 
                (N339)? mhpmcounter_q[1925] : 
                (N341)? mhpmcounter_q[1861] : 
                (N343)? mhpmcounter_q[1797] : 
                (N345)? mhpmcounter_q[1733] : 
                (N347)? mhpmcounter_q[1669] : 
                (N349)? mhpmcounter_q[1605] : 
                (N351)? mhpmcounter_q[1541] : 
                (N353)? mhpmcounter_q[1477] : 
                (N355)? mhpmcounter_q[1413] : 
                (N357)? mhpmcounter_q[1349] : 
                (N359)? mhpmcounter_q[1285] : 
                (N361)? mhpmcounter_q[1221] : 
                (N363)? mhpmcounter_q[1157] : 
                (N365)? mhpmcounter_q[1093] : 
                (N367)? mhpmcounter_q[1029] : 
                (N338)? mhpmcounter_q[965] : 
                (N340)? mhpmcounter_q[901] : 
                (N342)? mhpmcounter_q[837] : 
                (N344)? mhpmcounter_q[773] : 
                (N346)? mhpmcounter_q[709] : 
                (N348)? mhpmcounter_q[645] : 
                (N350)? mhpmcounter_q[581] : 
                (N352)? mhpmcounter_q[517] : 
                (N354)? mhpmcounter_q[453] : 
                (N356)? mhpmcounter_q[389] : 
                (N358)? mhpmcounter_q[325] : 
                (N360)? mhpmcounter_q[261] : 
                (N362)? mhpmcounter_q[197] : 
                (N364)? mhpmcounter_q[133] : 
                (N366)? mhpmcounter_q[69] : 
                (N368)? mhpmcounter_q[5] : 1'b0;
  assign N265 = (N337)? mhpmcounter_q[1988] : 
                (N339)? mhpmcounter_q[1924] : 
                (N341)? mhpmcounter_q[1860] : 
                (N343)? mhpmcounter_q[1796] : 
                (N345)? mhpmcounter_q[1732] : 
                (N347)? mhpmcounter_q[1668] : 
                (N349)? mhpmcounter_q[1604] : 
                (N351)? mhpmcounter_q[1540] : 
                (N353)? mhpmcounter_q[1476] : 
                (N355)? mhpmcounter_q[1412] : 
                (N357)? mhpmcounter_q[1348] : 
                (N359)? mhpmcounter_q[1284] : 
                (N361)? mhpmcounter_q[1220] : 
                (N363)? mhpmcounter_q[1156] : 
                (N365)? mhpmcounter_q[1092] : 
                (N367)? mhpmcounter_q[1028] : 
                (N338)? mhpmcounter_q[964] : 
                (N340)? mhpmcounter_q[900] : 
                (N342)? mhpmcounter_q[836] : 
                (N344)? mhpmcounter_q[772] : 
                (N346)? mhpmcounter_q[708] : 
                (N348)? mhpmcounter_q[644] : 
                (N350)? mhpmcounter_q[580] : 
                (N352)? mhpmcounter_q[516] : 
                (N354)? mhpmcounter_q[452] : 
                (N356)? mhpmcounter_q[388] : 
                (N358)? mhpmcounter_q[324] : 
                (N360)? mhpmcounter_q[260] : 
                (N362)? mhpmcounter_q[196] : 
                (N364)? mhpmcounter_q[132] : 
                (N366)? mhpmcounter_q[68] : 
                (N368)? mhpmcounter_q[4] : 1'b0;
  assign N266 = (N337)? mhpmcounter_q[1987] : 
                (N339)? mhpmcounter_q[1923] : 
                (N341)? mhpmcounter_q[1859] : 
                (N343)? mhpmcounter_q[1795] : 
                (N345)? mhpmcounter_q[1731] : 
                (N347)? mhpmcounter_q[1667] : 
                (N349)? mhpmcounter_q[1603] : 
                (N351)? mhpmcounter_q[1539] : 
                (N353)? mhpmcounter_q[1475] : 
                (N355)? mhpmcounter_q[1411] : 
                (N357)? mhpmcounter_q[1347] : 
                (N359)? mhpmcounter_q[1283] : 
                (N361)? mhpmcounter_q[1219] : 
                (N363)? mhpmcounter_q[1155] : 
                (N365)? mhpmcounter_q[1091] : 
                (N367)? mhpmcounter_q[1027] : 
                (N338)? mhpmcounter_q[963] : 
                (N340)? mhpmcounter_q[899] : 
                (N342)? mhpmcounter_q[835] : 
                (N344)? mhpmcounter_q[771] : 
                (N346)? mhpmcounter_q[707] : 
                (N348)? mhpmcounter_q[643] : 
                (N350)? mhpmcounter_q[579] : 
                (N352)? mhpmcounter_q[515] : 
                (N354)? mhpmcounter_q[451] : 
                (N356)? mhpmcounter_q[387] : 
                (N358)? mhpmcounter_q[323] : 
                (N360)? mhpmcounter_q[259] : 
                (N362)? mhpmcounter_q[195] : 
                (N364)? mhpmcounter_q[131] : 
                (N366)? mhpmcounter_q[67] : 
                (N368)? mhpmcounter_q[3] : 1'b0;
  assign N267 = (N337)? mhpmcounter_q[1986] : 
                (N339)? mhpmcounter_q[1922] : 
                (N341)? mhpmcounter_q[1858] : 
                (N343)? mhpmcounter_q[1794] : 
                (N345)? mhpmcounter_q[1730] : 
                (N347)? mhpmcounter_q[1666] : 
                (N349)? mhpmcounter_q[1602] : 
                (N351)? mhpmcounter_q[1538] : 
                (N353)? mhpmcounter_q[1474] : 
                (N355)? mhpmcounter_q[1410] : 
                (N357)? mhpmcounter_q[1346] : 
                (N359)? mhpmcounter_q[1282] : 
                (N361)? mhpmcounter_q[1218] : 
                (N363)? mhpmcounter_q[1154] : 
                (N365)? mhpmcounter_q[1090] : 
                (N367)? mhpmcounter_q[1026] : 
                (N338)? mhpmcounter_q[962] : 
                (N340)? mhpmcounter_q[898] : 
                (N342)? mhpmcounter_q[834] : 
                (N344)? mhpmcounter_q[770] : 
                (N346)? mhpmcounter_q[706] : 
                (N348)? mhpmcounter_q[642] : 
                (N350)? mhpmcounter_q[578] : 
                (N352)? mhpmcounter_q[514] : 
                (N354)? mhpmcounter_q[450] : 
                (N356)? mhpmcounter_q[386] : 
                (N358)? mhpmcounter_q[322] : 
                (N360)? mhpmcounter_q[258] : 
                (N362)? mhpmcounter_q[194] : 
                (N364)? mhpmcounter_q[130] : 
                (N366)? mhpmcounter_q[66] : 
                (N368)? mhpmcounter_q[2] : 1'b0;
  assign N268 = (N337)? mhpmcounter_q[1985] : 
                (N339)? mhpmcounter_q[1921] : 
                (N341)? mhpmcounter_q[1857] : 
                (N343)? mhpmcounter_q[1793] : 
                (N345)? mhpmcounter_q[1729] : 
                (N347)? mhpmcounter_q[1665] : 
                (N349)? mhpmcounter_q[1601] : 
                (N351)? mhpmcounter_q[1537] : 
                (N353)? mhpmcounter_q[1473] : 
                (N355)? mhpmcounter_q[1409] : 
                (N357)? mhpmcounter_q[1345] : 
                (N359)? mhpmcounter_q[1281] : 
                (N361)? mhpmcounter_q[1217] : 
                (N363)? mhpmcounter_q[1153] : 
                (N365)? mhpmcounter_q[1089] : 
                (N367)? mhpmcounter_q[1025] : 
                (N338)? mhpmcounter_q[961] : 
                (N340)? mhpmcounter_q[897] : 
                (N342)? mhpmcounter_q[833] : 
                (N344)? mhpmcounter_q[769] : 
                (N346)? mhpmcounter_q[705] : 
                (N348)? mhpmcounter_q[641] : 
                (N350)? mhpmcounter_q[577] : 
                (N352)? mhpmcounter_q[513] : 
                (N354)? mhpmcounter_q[449] : 
                (N356)? mhpmcounter_q[385] : 
                (N358)? mhpmcounter_q[321] : 
                (N360)? mhpmcounter_q[257] : 
                (N362)? mhpmcounter_q[193] : 
                (N364)? mhpmcounter_q[129] : 
                (N366)? mhpmcounter_q[65] : 
                (N368)? mhpmcounter_q[1] : 1'b0;
  assign N269 = (N337)? mhpmcounter_q[1984] : 
                (N339)? mhpmcounter_q[1920] : 
                (N341)? mhpmcounter_q[1856] : 
                (N343)? mhpmcounter_q[1792] : 
                (N345)? mhpmcounter_q[1728] : 
                (N347)? mhpmcounter_q[1664] : 
                (N349)? mhpmcounter_q[1600] : 
                (N351)? mhpmcounter_q[1536] : 
                (N353)? mhpmcounter_q[1472] : 
                (N355)? mhpmcounter_q[1408] : 
                (N357)? mhpmcounter_q[1344] : 
                (N359)? mhpmcounter_q[1280] : 
                (N361)? mhpmcounter_q[1216] : 
                (N363)? mhpmcounter_q[1152] : 
                (N365)? mhpmcounter_q[1088] : 
                (N367)? mhpmcounter_q[1024] : 
                (N338)? mhpmcounter_q[960] : 
                (N340)? mhpmcounter_q[896] : 
                (N342)? mhpmcounter_q[832] : 
                (N344)? mhpmcounter_q[768] : 
                (N346)? mhpmcounter_q[704] : 
                (N348)? mhpmcounter_q[640] : 
                (N350)? mhpmcounter_q[576] : 
                (N352)? mhpmcounter_q[512] : 
                (N354)? mhpmcounter_q[448] : 
                (N356)? mhpmcounter_q[384] : 
                (N358)? mhpmcounter_q[320] : 
                (N360)? mhpmcounter_q[256] : 
                (N362)? mhpmcounter_q[192] : 
                (N364)? mhpmcounter_q[128] : 
                (N366)? mhpmcounter_q[64] : 
                (N368)? mhpmcounter_q[0] : 1'b0;
  assign N270 = N10635 | N430;
  assign N271 = csr_addr_i[5] | N431;
  assign N272 = N270 | N460;
  assign N273 = N454 | N271;
  assign N274 = N280 | N450;
  assign N275 = N272 | N273;
  assign N276 = N275 | N274;
  assign N278 = N407 | N425;
  assign N280 = csr_addr_i[3] | N10658;
  assign N281 = N280 | N424;
  assign N282 = N407 | N281;
  assign N369 = (N337)? 1'b0 : 
                (N339)? 1'b0 : 
                (N341)? 1'b1 : 
                (N343)? 1'b0 : 
                (N345)? 1'b0 : 
                (N347)? 1'b0 : 
                (N349)? 1'b0 : 
                (N351)? 1'b0 : 
                (N353)? 1'b0 : 
                (N355)? 1'b0 : 
                (N357)? 1'b0 : 
                (N359)? 1'b0 : 
                (N361)? 1'b0 : 
                (N363)? 1'b0 : 
                (N365)? 1'b0 : 
                (N367)? 1'b0 : 
                (N338)? 1'b0 : 
                (N340)? 1'b0 : 
                (N342)? 1'b0 : 
                (N344)? 1'b0 : 
                (N346)? 1'b0 : 
                (N348)? 1'b0 : 
                (N350)? 1'b0 : 
                (N352)? 1'b0 : 
                (N354)? 1'b0 : 
                (N356)? 1'b0 : 
                (N358)? 1'b0 : 
                (N360)? 1'b0 : 
                (N362)? 1'b0 : 
                (N364)? 1'b0 : 
                (N366)? 1'b0 : 
                (N368)? 1'b0 : 1'b0;
  assign N370 = (N337)? 1'b1 : 
                (N339)? 1'b0 : 
                (N341)? 1'b0 : 
                (N343)? 1'b0 : 
                (N345)? 1'b0 : 
                (N347)? 1'b0 : 
                (N349)? 1'b0 : 
                (N351)? 1'b0 : 
                (N353)? 1'b0 : 
                (N355)? 1'b0 : 
                (N357)? 1'b0 : 
                (N359)? 1'b0 : 
                (N361)? 1'b0 : 
                (N363)? 1'b0 : 
                (N365)? 1'b0 : 
                (N367)? 1'b0 : 
                (N338)? 1'b0 : 
                (N340)? 1'b0 : 
                (N342)? 1'b0 : 
                (N344)? 1'b0 : 
                (N346)? 1'b0 : 
                (N348)? 1'b0 : 
                (N350)? 1'b0 : 
                (N352)? 1'b0 : 
                (N354)? 1'b0 : 
                (N356)? 1'b0 : 
                (N358)? 1'b0 : 
                (N360)? 1'b0 : 
                (N362)? 1'b0 : 
                (N364)? 1'b0 : 
                (N366)? 1'b0 : 
                (N368)? 1'b0 : 1'b0;
  assign N407 = N443 | N455;
  assign N408 = N407 | N451;
  assign N410 = N419 | N451;
  assign N412 = N419 | N425;
  assign N414 = N419 | N467;
  assign N417 = csr_addr_i[7] | N416;
  assign N418 = N417 | N462;
  assign N419 = N443 | N418;
  assign N420 = N419 | N437;
  assign N422 = N438 | N451;
  assign N424 = csr_addr_i[1] | N10623;
  assign N425 = N463 | N424;
  assign N426 = N438 | N425;
  assign N428 = N438 | N467;
  assign N432 = csr_addr_i[11] | N430;
  assign N433 = N10646 | N431;
  assign N434 = N10626 | N10623;
  assign N435 = N432 | N460;
  assign N436 = N461 | N433;
  assign N437 = N463 | N434;
  assign N438 = N435 | N436;
  assign N439 = N438 | N437;
  assign N441 = csr_addr_i[11] | csr_addr_i[10];
  assign N442 = N10646 | csr_addr_i[4];
  assign N443 = N441 | N460;
  assign N444 = N454 | N442;
  assign N445 = N443 | N444;
  assign N446 = N445 | N451;
  assign N448 = N456 | N451;
  assign N450 = csr_addr_i[1] | csr_addr_i[0];
  assign N451 = N463 | N450;
  assign N452 = N468 | N451;
  assign N454 = csr_addr_i[7] | csr_addr_i[6];
  assign N455 = N454 | N462;
  assign N456 = N465 | N455;
  assign N457 = N456 | N467;
  assign N459 = N10635 | csr_addr_i[10];
  assign N460 = N10636 | N10637;
  assign N461 = N10638 | csr_addr_i[6];
  assign N462 = csr_addr_i[5] | csr_addr_i[4];
  assign N463 = csr_addr_i[3] | csr_addr_i[2];
  assign N464 = N10626 | csr_addr_i[0];
  assign N465 = N459 | N460;
  assign N466 = N461 | N462;
  assign N467 = N463 | N464;
  assign N468 = N465 | N466;
  assign N469 = N468 | N467;
  assign dcsr_d[2] = N956;
  assign dcsr_d[3] = N957;
  assign dcsr_d[4] = N958;
  assign dcsr_d[5] = N959;
  assign dcsr_d[9] = N963;
  assign dcsr_d[10] = N964;
  assign dcsr_d[11] = N965;
  assign dcsr_d[12] = N966;
  assign dcsr_d[13] = N967;
  assign dcsr_d[14] = N968;
  assign dcsr_d[15] = N969;
  assign dcsr_d[16] = N970;
  assign dcsr_d[17] = N971;
  assign dcsr_d[18] = N972;
  assign dcsr_d[19] = N973;
  assign dcsr_d[20] = N974;
  assign dcsr_d[21] = N975;
  assign dcsr_d[22] = N976;
  assign dcsr_d[23] = N977;
  assign dcsr_d[24] = N978;
  assign dcsr_d[25] = N979;
  assign dcsr_d[26] = N980;
  assign dcsr_d[27] = N981;
  assign dcsr_d[28] = N982;
  assign dcsr_d[29] = N983;
  assign dcsr_d[30] = N984;
  assign dcsr_d[31] = N985;
  assign N1166 = csr_op_i[1] | N1172;
  assign N1168 = N1171 | csr_op_i[0];
  assign N1170 = csr_op_i[1] & csr_op_i[0];
  assign N1173 = N1171 & N1172;

  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[31] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[31] <= dscratch1_d[31];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[30] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[30] <= dscratch1_d[30];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[29] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[29] <= dscratch1_d[29];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[28] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[28] <= dscratch1_d[28];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[27] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[27] <= dscratch1_d[27];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[26] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[26] <= dscratch1_d[26];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[25] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[25] <= dscratch1_d[25];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[24] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[24] <= dscratch1_d[24];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[23] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[23] <= dscratch1_d[23];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[22] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[22] <= dscratch1_d[22];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[21] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[21] <= dscratch1_d[21];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[20] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[20] <= dscratch1_d[20];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[19] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[19] <= dscratch1_d[19];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[18] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[18] <= dscratch1_d[18];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[17] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[17] <= dscratch1_d[17];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[16] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[16] <= dscratch1_d[16];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[15] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[15] <= dscratch1_d[15];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[14] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[14] <= dscratch1_d[14];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[13] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[13] <= dscratch1_d[13];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[12] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[12] <= dscratch1_d[12];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[11] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[11] <= dscratch1_d[11];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[10] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[10] <= dscratch1_d[10];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[9] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[9] <= dscratch1_d[9];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[8] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[8] <= dscratch1_d[8];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[7] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[7] <= dscratch1_d[7];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[6] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[6] <= dscratch1_d[6];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[5] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[5] <= dscratch1_d[5];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[4] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[4] <= dscratch1_d[4];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[3] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[3] <= dscratch1_d[3];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[2] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[2] <= dscratch1_d[2];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[1] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[1] <= dscratch1_d[1];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch1_q[0] <= 1'b0;
    end else if(N10596) begin
      dscratch1_q[0] <= dscratch1_d[0];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      m_irq_enable_o <= 1'b0;
    end else if(1'b1) begin
      m_irq_enable_o <= mstatus_d_mie_;
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mstatus_q_mpie_ <= 1'b0;
    end else if(1'b1) begin
      mstatus_q_mpie_ <= mstatus_d_mpie_;
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mstatus_q_mpp__1_ <= 1'b1;
    end else if(1'b1) begin
      mstatus_q_mpp__1_ <= 1'b1;
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mstatus_q_mpp__0_ <= 1'b1;
    end else if(1'b1) begin
      mstatus_q_mpp__0_ <= 1'b1;
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[31] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[31] <= mscratch_d[31];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[30] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[30] <= mscratch_d[30];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[29] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[29] <= mscratch_d[29];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[28] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[28] <= mscratch_d[28];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[27] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[27] <= mscratch_d[27];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[26] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[26] <= mscratch_d[26];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[25] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[25] <= mscratch_d[25];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[24] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[24] <= mscratch_d[24];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[23] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[23] <= mscratch_d[23];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[22] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[22] <= mscratch_d[22];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[21] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[21] <= mscratch_d[21];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[20] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[20] <= mscratch_d[20];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[19] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[19] <= mscratch_d[19];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[18] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[18] <= mscratch_d[18];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[17] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[17] <= mscratch_d[17];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[16] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[16] <= mscratch_d[16];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[15] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[15] <= mscratch_d[15];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[14] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[14] <= mscratch_d[14];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[13] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[13] <= mscratch_d[13];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[12] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[12] <= mscratch_d[12];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[11] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[11] <= mscratch_d[11];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[10] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[10] <= mscratch_d[10];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[9] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[9] <= mscratch_d[9];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[8] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[8] <= mscratch_d[8];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[7] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[7] <= mscratch_d[7];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[6] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[6] <= mscratch_d[6];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[5] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[5] <= mscratch_d[5];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[4] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[4] <= mscratch_d[4];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[3] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[3] <= mscratch_d[3];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[2] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[2] <= mscratch_d[2];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[1] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[1] <= mscratch_d[1];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mscratch_q[0] <= 1'b0;
    end else if(N10609) begin
      mscratch_q[0] <= mscratch_d[0];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[31] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[31] <= mepc_d[31];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[30] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[30] <= mepc_d[30];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[29] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[29] <= mepc_d[29];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[28] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[28] <= mepc_d[28];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[27] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[27] <= mepc_d[27];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[26] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[26] <= mepc_d[26];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[25] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[25] <= mepc_d[25];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[24] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[24] <= mepc_d[24];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[23] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[23] <= mepc_d[23];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[22] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[22] <= mepc_d[22];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[21] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[21] <= mepc_d[21];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[20] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[20] <= mepc_d[20];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[19] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[19] <= mepc_d[19];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[18] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[18] <= mepc_d[18];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[17] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[17] <= mepc_d[17];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[16] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[16] <= mepc_d[16];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[15] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[15] <= mepc_d[15];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[14] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[14] <= mepc_d[14];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[13] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[13] <= mepc_d[13];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[12] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[12] <= mepc_d[12];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[11] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[11] <= mepc_d[11];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[10] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[10] <= mepc_d[10];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[9] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[9] <= mepc_d[9];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[8] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[8] <= mepc_d[8];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[7] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[7] <= mepc_d[7];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[6] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[6] <= mepc_d[6];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[5] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[5] <= mepc_d[5];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[4] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[4] <= mepc_d[4];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[3] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[3] <= mepc_d[3];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[2] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[2] <= mepc_d[2];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[1] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[1] <= mepc_d[1];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_mepc_o[0] <= 1'b0;
    end else if(1'b1) begin
      csr_mepc_o[0] <= mepc_d[0];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcause_q[5] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[5] <= mcause_d[5];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcause_q[4] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[4] <= mcause_d[4];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcause_q[3] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[3] <= mcause_d[3];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcause_q[2] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[2] <= mcause_d[2];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcause_q[1] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[1] <= mcause_d[1];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcause_q[0] <= 1'b0;
    end else if(1'b1) begin
      mcause_q[0] <= mcause_d[0];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[31] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[31] <= mtval_d[31];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[30] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[30] <= mtval_d[30];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[29] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[29] <= mtval_d[29];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[28] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[28] <= mtval_d[28];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[27] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[27] <= mtval_d[27];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[26] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[26] <= mtval_d[26];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[25] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[25] <= mtval_d[25];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[24] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[24] <= mtval_d[24];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[23] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[23] <= mtval_d[23];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[22] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[22] <= mtval_d[22];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[21] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[21] <= mtval_d[21];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[20] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[20] <= mtval_d[20];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[19] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[19] <= mtval_d[19];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[18] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[18] <= mtval_d[18];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[17] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[17] <= mtval_d[17];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[16] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[16] <= mtval_d[16];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[15] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[15] <= mtval_d[15];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[14] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[14] <= mtval_d[14];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[13] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[13] <= mtval_d[13];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[12] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[12] <= mtval_d[12];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[11] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[11] <= mtval_d[11];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[10] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[10] <= mtval_d[10];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[9] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[9] <= mtval_d[9];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[8] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[8] <= mtval_d[8];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[7] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[7] <= mtval_d[7];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[6] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[6] <= mtval_d[6];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[5] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[5] <= mtval_d[5];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[4] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[4] <= mtval_d[4];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[3] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[3] <= mtval_d[3];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[2] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[2] <= mtval_d[2];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[1] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[1] <= mtval_d[1];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mtval_q[0] <= 1'b0;
    end else if(1'b1) begin
      mtval_q[0] <= mtval_d[0];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_xdebugver__3_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_xdebugver__3_ <= dcsr_d[31];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_xdebugver__2_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_xdebugver__2_ <= dcsr_d[30];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_xdebugver__1_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_xdebugver__1_ <= dcsr_d[29];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_xdebugver__0_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_xdebugver__0_ <= dcsr_d[28];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_zero2__11_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero2__11_ <= dcsr_d[27];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_zero2__10_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero2__10_ <= dcsr_d[26];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_zero2__9_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero2__9_ <= dcsr_d[25];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_zero2__8_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero2__8_ <= dcsr_d[24];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_zero2__7_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero2__7_ <= dcsr_d[23];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_zero2__6_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero2__6_ <= dcsr_d[22];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_zero2__5_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero2__5_ <= dcsr_d[21];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_zero2__4_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero2__4_ <= dcsr_d[20];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_zero2__3_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero2__3_ <= dcsr_d[19];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_zero2__2_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero2__2_ <= dcsr_d[18];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_zero2__1_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero2__1_ <= dcsr_d[17];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_zero2__0_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero2__0_ <= dcsr_d[16];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      debug_ebreakm_o <= 1'b0;
    end else if(1'b1) begin
      debug_ebreakm_o <= dcsr_d[15];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_zero1_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero1_ <= dcsr_d[14];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_ebreaks_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_ebreaks_ <= dcsr_d[13];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_ebreaku_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_ebreaku_ <= dcsr_d[12];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_stepie_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_stepie_ <= dcsr_d[11];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_stopcount_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_stopcount_ <= dcsr_d[10];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_stoptime_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_stoptime_ <= dcsr_d[9];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_cause__2_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_cause__2_ <= dcsr_d[8];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_cause__1_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_cause__1_ <= dcsr_d[7];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_cause__0_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_cause__0_ <= dcsr_d[6];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_zero0_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_zero0_ <= dcsr_d[5];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_mprven_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_mprven_ <= dcsr_d[4];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_nmip_ <= 1'b0;
    end else if(1'b1) begin
      dcsr_q_nmip_ <= dcsr_d[3];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      debug_single_step_o <= 1'b0;
    end else if(1'b1) begin
      debug_single_step_o <= dcsr_d[2];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_prv__1_ <= 1'b1;
    end else if(1'b1) begin
      dcsr_q_prv__1_ <= dcsr_d[1];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dcsr_q_prv__0_ <= 1'b1;
    end else if(1'b1) begin
      dcsr_q_prv__0_ <= dcsr_d[0];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[31] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[31] <= depc_d[31];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[30] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[30] <= depc_d[30];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[29] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[29] <= depc_d[29];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[28] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[28] <= depc_d[28];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[27] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[27] <= depc_d[27];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[26] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[26] <= depc_d[26];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[25] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[25] <= depc_d[25];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[24] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[24] <= depc_d[24];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[23] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[23] <= depc_d[23];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[22] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[22] <= depc_d[22];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[21] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[21] <= depc_d[21];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[20] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[20] <= depc_d[20];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[19] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[19] <= depc_d[19];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[18] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[18] <= depc_d[18];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[17] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[17] <= depc_d[17];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[16] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[16] <= depc_d[16];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[15] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[15] <= depc_d[15];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[14] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[14] <= depc_d[14];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[13] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[13] <= depc_d[13];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[12] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[12] <= depc_d[12];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[11] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[11] <= depc_d[11];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[10] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[10] <= depc_d[10];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[9] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[9] <= depc_d[9];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[8] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[8] <= depc_d[8];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[7] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[7] <= depc_d[7];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[6] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[6] <= depc_d[6];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[5] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[5] <= depc_d[5];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[4] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[4] <= depc_d[4];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[3] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[3] <= depc_d[3];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[2] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[2] <= depc_d[2];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[1] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[1] <= depc_d[1];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      csr_depc_o[0] <= 1'b0;
    end else if(1'b1) begin
      csr_depc_o[0] <= depc_d[0];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[31] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[31] <= dscratch0_d[31];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[30] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[30] <= dscratch0_d[30];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[29] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[29] <= dscratch0_d[29];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[28] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[28] <= dscratch0_d[28];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[27] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[27] <= dscratch0_d[27];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[26] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[26] <= dscratch0_d[26];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[25] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[25] <= dscratch0_d[25];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[24] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[24] <= dscratch0_d[24];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[23] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[23] <= dscratch0_d[23];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[22] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[22] <= dscratch0_d[22];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[21] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[21] <= dscratch0_d[21];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[20] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[20] <= dscratch0_d[20];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[19] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[19] <= dscratch0_d[19];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[18] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[18] <= dscratch0_d[18];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[17] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[17] <= dscratch0_d[17];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[16] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[16] <= dscratch0_d[16];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[15] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[15] <= dscratch0_d[15];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[14] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[14] <= dscratch0_d[14];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[13] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[13] <= dscratch0_d[13];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[12] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[12] <= dscratch0_d[12];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[11] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[11] <= dscratch0_d[11];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[10] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[10] <= dscratch0_d[10];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[9] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[9] <= dscratch0_d[9];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[8] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[8] <= dscratch0_d[8];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[7] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[7] <= dscratch0_d[7];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[6] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[6] <= dscratch0_d[6];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[5] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[5] <= dscratch0_d[5];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[4] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[4] <= dscratch0_d[4];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[3] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[3] <= dscratch0_d[3];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[2] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[2] <= dscratch0_d[2];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[1] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[1] <= dscratch0_d[1];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      dscratch0_q[0] <= 1'b0;
    end else if(N10616) begin
      dscratch0_q[0] <= dscratch0_d[0];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[31] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[31] <= mcountinhibit_d[31];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[30] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[30] <= mcountinhibit_d[30];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[29] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[29] <= mcountinhibit_d[29];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[28] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[28] <= mcountinhibit_d[28];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[27] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[27] <= mcountinhibit_d[27];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[26] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[26] <= mcountinhibit_d[26];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[25] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[25] <= mcountinhibit_d[25];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[24] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[24] <= mcountinhibit_d[24];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[23] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[23] <= mcountinhibit_d[23];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[22] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[22] <= mcountinhibit_d[22];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[21] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[21] <= mcountinhibit_d[21];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[20] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[20] <= mcountinhibit_d[20];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[19] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[19] <= mcountinhibit_d[19];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[18] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[18] <= mcountinhibit_d[18];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[17] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[17] <= mcountinhibit_d[17];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[16] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[16] <= mcountinhibit_d[16];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[15] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[15] <= mcountinhibit_d[15];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[14] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[14] <= mcountinhibit_d[14];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[13] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[13] <= mcountinhibit_d[13];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[12] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[12] <= mcountinhibit_d[12];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[11] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[11] <= mcountinhibit_d[11];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[10] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[10] <= mcountinhibit_d[10];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[9] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[9] <= mcountinhibit_d[9];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[8] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[8] <= mcountinhibit_d[8];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[7] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[7] <= mcountinhibit_d[7];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[6] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[6] <= mcountinhibit_d[6];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[5] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[5] <= mcountinhibit_d[5];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[4] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[4] <= mcountinhibit_d[4];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[3] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[3] <= mcountinhibit_d[3];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[2] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[2] <= mcountinhibit_d[2];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[1] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[1] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mcountinhibit_q[0] <= 1'b0;
    end else if(1'b1) begin
      mcountinhibit_q[0] <= mcountinhibit_d_0;
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2047] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2047] <= mhpmcounter_d[2047];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2046] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2046] <= mhpmcounter_d[2046];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2045] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2045] <= mhpmcounter_d[2045];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2044] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2044] <= mhpmcounter_d[2044];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2043] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2043] <= mhpmcounter_d[2043];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2042] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2042] <= mhpmcounter_d[2042];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2041] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2041] <= mhpmcounter_d[2041];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2040] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2040] <= mhpmcounter_d[2040];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2039] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2039] <= mhpmcounter_d[2039];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2038] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2038] <= mhpmcounter_d[2038];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2037] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2037] <= mhpmcounter_d[2037];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2036] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2036] <= mhpmcounter_d[2036];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2035] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2035] <= mhpmcounter_d[2035];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2034] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2034] <= mhpmcounter_d[2034];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2033] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2033] <= mhpmcounter_d[2033];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2032] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2032] <= mhpmcounter_d[2032];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2031] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2031] <= mhpmcounter_d[2031];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2030] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2030] <= mhpmcounter_d[2030];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2029] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2029] <= mhpmcounter_d[2029];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2028] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2028] <= mhpmcounter_d[2028];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2027] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2027] <= mhpmcounter_d[2027];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2026] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2026] <= mhpmcounter_d[2026];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2025] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2025] <= mhpmcounter_d[2025];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2024] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2024] <= mhpmcounter_d[2024];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2023] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2023] <= mhpmcounter_d[2023];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2022] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2022] <= mhpmcounter_d[2022];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2021] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2021] <= mhpmcounter_d[2021];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2020] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2020] <= mhpmcounter_d[2020];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2019] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2019] <= mhpmcounter_d[2019];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2018] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2018] <= mhpmcounter_d[2018];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2017] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2017] <= mhpmcounter_d[2017];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2016] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2016] <= mhpmcounter_d[2016];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2015] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2015] <= mhpmcounter_d[2015];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2014] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2014] <= mhpmcounter_d[2014];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2013] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2013] <= mhpmcounter_d[2013];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2012] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2012] <= mhpmcounter_d[2012];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2011] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2011] <= mhpmcounter_d[2011];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2010] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2010] <= mhpmcounter_d[2010];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2009] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2009] <= mhpmcounter_d[2009];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2008] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2008] <= mhpmcounter_d[2008];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2007] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2007] <= mhpmcounter_d[2007];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2006] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2006] <= mhpmcounter_d[2006];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2005] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2005] <= mhpmcounter_d[2005];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2004] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2004] <= mhpmcounter_d[2004];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2003] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2003] <= mhpmcounter_d[2003];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2002] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2002] <= mhpmcounter_d[2002];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2001] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2001] <= mhpmcounter_d[2001];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2000] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2000] <= mhpmcounter_d[2000];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1999] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1999] <= mhpmcounter_d[1999];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1998] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1998] <= mhpmcounter_d[1998];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1997] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1997] <= mhpmcounter_d[1997];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1996] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1996] <= mhpmcounter_d[1996];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1995] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1995] <= mhpmcounter_d[1995];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1994] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1994] <= mhpmcounter_d[1994];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1993] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1993] <= mhpmcounter_d[1993];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1992] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1992] <= mhpmcounter_d[1992];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1991] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1991] <= mhpmcounter_d[1991];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1990] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1990] <= mhpmcounter_d[1990];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1989] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1989] <= mhpmcounter_d[1989];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1988] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1988] <= mhpmcounter_d[1988];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1987] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1987] <= mhpmcounter_d[1987];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1986] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1986] <= mhpmcounter_d[1986];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1985] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1985] <= mhpmcounter_d[1985];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1984] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1984] <= mhpmcounter_d[1984];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1983] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1983] <= mhpmcounter_d[1983];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1982] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1982] <= mhpmcounter_d[1982];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1981] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1981] <= mhpmcounter_d[1981];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1980] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1980] <= mhpmcounter_d[1980];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1979] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1979] <= mhpmcounter_d[1979];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1978] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1978] <= mhpmcounter_d[1978];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1977] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1977] <= mhpmcounter_d[1977];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1976] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1976] <= mhpmcounter_d[1976];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1975] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1975] <= mhpmcounter_d[1975];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1974] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1974] <= mhpmcounter_d[1974];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1973] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1973] <= mhpmcounter_d[1973];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1972] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1972] <= mhpmcounter_d[1972];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1971] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1971] <= mhpmcounter_d[1971];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1970] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1970] <= mhpmcounter_d[1970];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1969] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1969] <= mhpmcounter_d[1969];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1968] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1968] <= mhpmcounter_d[1968];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1967] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1967] <= mhpmcounter_d[1967];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1966] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1966] <= mhpmcounter_d[1966];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1965] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1965] <= mhpmcounter_d[1965];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1964] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1964] <= mhpmcounter_d[1964];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1963] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1963] <= mhpmcounter_d[1963];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1962] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1962] <= mhpmcounter_d[1962];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1961] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1961] <= mhpmcounter_d[1961];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1960] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1960] <= mhpmcounter_d[1960];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1959] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1959] <= mhpmcounter_d[1959];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1958] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1958] <= mhpmcounter_d[1958];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1957] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1957] <= mhpmcounter_d[1957];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1956] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1956] <= mhpmcounter_d[1956];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1955] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1955] <= mhpmcounter_d[1955];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1954] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1954] <= mhpmcounter_d[1954];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1953] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1953] <= mhpmcounter_d[1953];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1952] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1952] <= mhpmcounter_d[1952];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1951] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1951] <= mhpmcounter_d[1951];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1950] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1950] <= mhpmcounter_d[1950];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1949] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1949] <= mhpmcounter_d[1949];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1948] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1948] <= mhpmcounter_d[1948];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1947] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1947] <= mhpmcounter_d[1947];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1946] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1946] <= mhpmcounter_d[1946];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1945] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1945] <= mhpmcounter_d[1945];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1944] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1944] <= mhpmcounter_d[1944];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1943] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1943] <= mhpmcounter_d[1943];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1942] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1942] <= mhpmcounter_d[1942];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1941] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1941] <= mhpmcounter_d[1941];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1940] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1940] <= mhpmcounter_d[1940];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1939] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1939] <= mhpmcounter_d[1939];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1938] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1938] <= mhpmcounter_d[1938];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1937] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1937] <= mhpmcounter_d[1937];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1936] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1936] <= mhpmcounter_d[1936];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1935] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1935] <= mhpmcounter_d[1935];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1934] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1934] <= mhpmcounter_d[1934];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1933] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1933] <= mhpmcounter_d[1933];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1932] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1932] <= mhpmcounter_d[1932];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1931] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1931] <= mhpmcounter_d[1931];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1930] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1930] <= mhpmcounter_d[1930];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1929] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1929] <= mhpmcounter_d[1929];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1928] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1928] <= mhpmcounter_d[1928];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1927] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1927] <= mhpmcounter_d[1927];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1926] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1926] <= mhpmcounter_d[1926];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1925] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1925] <= mhpmcounter_d[1925];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1924] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1924] <= mhpmcounter_d[1924];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1923] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1923] <= mhpmcounter_d[1923];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1922] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1922] <= mhpmcounter_d[1922];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1921] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1921] <= mhpmcounter_d[1921];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1920] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1920] <= mhpmcounter_d[1920];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1919] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1919] <= mhpmcounter_d[1919];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1918] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1918] <= mhpmcounter_d[1918];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1917] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1917] <= mhpmcounter_d[1917];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1916] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1916] <= mhpmcounter_d[1916];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1915] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1915] <= mhpmcounter_d[1915];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1914] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1914] <= mhpmcounter_d[1914];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1913] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1913] <= mhpmcounter_d[1913];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1912] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1912] <= mhpmcounter_d[1912];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1911] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1911] <= mhpmcounter_d[1911];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1910] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1910] <= mhpmcounter_d[1910];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1909] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1909] <= mhpmcounter_d[1909];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1908] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1908] <= mhpmcounter_d[1908];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1907] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1907] <= mhpmcounter_d[1907];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1906] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1906] <= mhpmcounter_d[1906];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1905] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1905] <= mhpmcounter_d[1905];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1904] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1904] <= mhpmcounter_d[1904];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1903] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1903] <= mhpmcounter_d[1903];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1902] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1902] <= mhpmcounter_d[1902];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1901] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1901] <= mhpmcounter_d[1901];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1900] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1900] <= mhpmcounter_d[1900];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1899] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1899] <= mhpmcounter_d[1899];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1898] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1898] <= mhpmcounter_d[1898];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1897] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1897] <= mhpmcounter_d[1897];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1896] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1896] <= mhpmcounter_d[1896];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1895] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1895] <= mhpmcounter_d[1895];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1894] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1894] <= mhpmcounter_d[1894];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1893] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1893] <= mhpmcounter_d[1893];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1892] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1892] <= mhpmcounter_d[1892];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1891] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1891] <= mhpmcounter_d[1891];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1890] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1890] <= mhpmcounter_d[1890];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1889] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1889] <= mhpmcounter_d[1889];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1888] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1888] <= mhpmcounter_d[1888];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1887] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1887] <= mhpmcounter_d[1887];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1886] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1886] <= mhpmcounter_d[1886];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1885] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1885] <= mhpmcounter_d[1885];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1884] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1884] <= mhpmcounter_d[1884];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1883] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1883] <= mhpmcounter_d[1883];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1882] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1882] <= mhpmcounter_d[1882];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1881] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1881] <= mhpmcounter_d[1881];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1880] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1880] <= mhpmcounter_d[1880];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1879] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1879] <= mhpmcounter_d[1879];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1878] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1878] <= mhpmcounter_d[1878];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1877] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1877] <= mhpmcounter_d[1877];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1876] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1876] <= mhpmcounter_d[1876];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1875] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1875] <= mhpmcounter_d[1875];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1874] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1874] <= mhpmcounter_d[1874];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1873] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1873] <= mhpmcounter_d[1873];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1872] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1872] <= mhpmcounter_d[1872];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1871] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1871] <= mhpmcounter_d[1871];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1870] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1870] <= mhpmcounter_d[1870];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1869] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1869] <= mhpmcounter_d[1869];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1868] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1868] <= mhpmcounter_d[1868];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1867] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1867] <= mhpmcounter_d[1867];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1866] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1866] <= mhpmcounter_d[1866];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1865] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1865] <= mhpmcounter_d[1865];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1864] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1864] <= mhpmcounter_d[1864];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1863] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1863] <= mhpmcounter_d[1863];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1862] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1862] <= mhpmcounter_d[1862];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1861] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1861] <= mhpmcounter_d[1861];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1860] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1860] <= mhpmcounter_d[1860];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1859] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1859] <= mhpmcounter_d[1859];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1858] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1858] <= mhpmcounter_d[1858];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1857] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1857] <= mhpmcounter_d[1857];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1856] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1856] <= mhpmcounter_d[1856];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1855] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1855] <= mhpmcounter_d[1855];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1854] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1854] <= mhpmcounter_d[1854];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1853] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1853] <= mhpmcounter_d[1853];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1852] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1852] <= mhpmcounter_d[1852];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1851] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1851] <= mhpmcounter_d[1851];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1850] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1850] <= mhpmcounter_d[1850];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1849] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1849] <= mhpmcounter_d[1849];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1848] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1848] <= mhpmcounter_d[1848];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1847] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1847] <= mhpmcounter_d[1847];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1846] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1846] <= mhpmcounter_d[1846];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1845] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1845] <= mhpmcounter_d[1845];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1844] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1844] <= mhpmcounter_d[1844];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1843] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1843] <= mhpmcounter_d[1843];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1842] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1842] <= mhpmcounter_d[1842];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1841] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1841] <= mhpmcounter_d[1841];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1840] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1840] <= mhpmcounter_d[1840];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1839] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1839] <= mhpmcounter_d[1839];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1838] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1838] <= mhpmcounter_d[1838];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1837] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1837] <= mhpmcounter_d[1837];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1836] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1836] <= mhpmcounter_d[1836];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1835] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1835] <= mhpmcounter_d[1835];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1834] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1834] <= mhpmcounter_d[1834];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1833] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1833] <= mhpmcounter_d[1833];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1832] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1832] <= mhpmcounter_d[1832];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1831] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1831] <= mhpmcounter_d[1831];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1830] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1830] <= mhpmcounter_d[1830];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1829] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1829] <= mhpmcounter_d[1829];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1828] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1828] <= mhpmcounter_d[1828];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1827] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1827] <= mhpmcounter_d[1827];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1826] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1826] <= mhpmcounter_d[1826];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1825] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1825] <= mhpmcounter_d[1825];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1824] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1824] <= mhpmcounter_d[1824];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1823] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1823] <= mhpmcounter_d[1823];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1822] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1822] <= mhpmcounter_d[1822];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1821] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1821] <= mhpmcounter_d[1821];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1820] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1820] <= mhpmcounter_d[1820];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1819] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1819] <= mhpmcounter_d[1819];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1818] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1818] <= mhpmcounter_d[1818];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1817] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1817] <= mhpmcounter_d[1817];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1816] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1816] <= mhpmcounter_d[1816];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1815] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1815] <= mhpmcounter_d[1815];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1814] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1814] <= mhpmcounter_d[1814];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1813] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1813] <= mhpmcounter_d[1813];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1812] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1812] <= mhpmcounter_d[1812];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1811] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1811] <= mhpmcounter_d[1811];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1810] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1810] <= mhpmcounter_d[1810];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1809] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1809] <= mhpmcounter_d[1809];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1808] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1808] <= mhpmcounter_d[1808];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1807] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1807] <= mhpmcounter_d[1807];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1806] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1806] <= mhpmcounter_d[1806];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1805] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1805] <= mhpmcounter_d[1805];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1804] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1804] <= mhpmcounter_d[1804];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1803] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1803] <= mhpmcounter_d[1803];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1802] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1802] <= mhpmcounter_d[1802];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1801] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1801] <= mhpmcounter_d[1801];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1800] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1800] <= mhpmcounter_d[1800];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1799] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1799] <= mhpmcounter_d[1799];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1798] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1798] <= mhpmcounter_d[1798];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1797] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1797] <= mhpmcounter_d[1797];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1796] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1796] <= mhpmcounter_d[1796];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1795] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1795] <= mhpmcounter_d[1795];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1794] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1794] <= mhpmcounter_d[1794];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1793] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1793] <= mhpmcounter_d[1793];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1792] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1792] <= mhpmcounter_d[1792];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1791] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1791] <= mhpmcounter_d[1791];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1790] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1790] <= mhpmcounter_d[1790];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1789] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1789] <= mhpmcounter_d[1789];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1788] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1788] <= mhpmcounter_d[1788];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1787] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1787] <= mhpmcounter_d[1787];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1786] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1786] <= mhpmcounter_d[1786];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1785] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1785] <= mhpmcounter_d[1785];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1784] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1784] <= mhpmcounter_d[1784];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1783] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1783] <= mhpmcounter_d[1783];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1782] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1782] <= mhpmcounter_d[1782];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1781] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1781] <= mhpmcounter_d[1781];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1780] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1780] <= mhpmcounter_d[1780];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1779] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1779] <= mhpmcounter_d[1779];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1778] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1778] <= mhpmcounter_d[1778];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1777] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1777] <= mhpmcounter_d[1777];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1776] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1776] <= mhpmcounter_d[1776];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1775] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1775] <= mhpmcounter_d[1775];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1774] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1774] <= mhpmcounter_d[1774];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1773] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1773] <= mhpmcounter_d[1773];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1772] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1772] <= mhpmcounter_d[1772];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1771] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1771] <= mhpmcounter_d[1771];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1770] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1770] <= mhpmcounter_d[1770];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1769] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1769] <= mhpmcounter_d[1769];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1768] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1768] <= mhpmcounter_d[1768];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1767] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1767] <= mhpmcounter_d[1767];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1766] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1766] <= mhpmcounter_d[1766];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1765] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1765] <= mhpmcounter_d[1765];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1764] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1764] <= mhpmcounter_d[1764];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1763] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1763] <= mhpmcounter_d[1763];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1762] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1762] <= mhpmcounter_d[1762];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1761] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1761] <= mhpmcounter_d[1761];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1760] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1760] <= mhpmcounter_d[1760];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1759] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1759] <= mhpmcounter_d[1759];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1758] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1758] <= mhpmcounter_d[1758];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1757] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1757] <= mhpmcounter_d[1757];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1756] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1756] <= mhpmcounter_d[1756];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1755] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1755] <= mhpmcounter_d[1755];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1754] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1754] <= mhpmcounter_d[1754];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1753] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1753] <= mhpmcounter_d[1753];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1752] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1752] <= mhpmcounter_d[1752];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1751] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1751] <= mhpmcounter_d[1751];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1750] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1750] <= mhpmcounter_d[1750];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1749] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1749] <= mhpmcounter_d[1749];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1748] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1748] <= mhpmcounter_d[1748];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1747] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1747] <= mhpmcounter_d[1747];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1746] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1746] <= mhpmcounter_d[1746];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1745] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1745] <= mhpmcounter_d[1745];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1744] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1744] <= mhpmcounter_d[1744];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1743] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1743] <= mhpmcounter_d[1743];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1742] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1742] <= mhpmcounter_d[1742];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1741] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1741] <= mhpmcounter_d[1741];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1740] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1740] <= mhpmcounter_d[1740];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1739] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1739] <= mhpmcounter_d[1739];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1738] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1738] <= mhpmcounter_d[1738];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1737] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1737] <= mhpmcounter_d[1737];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1736] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1736] <= mhpmcounter_d[1736];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1735] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1735] <= mhpmcounter_d[1735];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1734] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1734] <= mhpmcounter_d[1734];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1733] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1733] <= mhpmcounter_d[1733];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1732] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1732] <= mhpmcounter_d[1732];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1731] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1731] <= mhpmcounter_d[1731];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1730] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1730] <= mhpmcounter_d[1730];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1729] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1729] <= mhpmcounter_d[1729];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1728] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1728] <= mhpmcounter_d[1728];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1727] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1727] <= mhpmcounter_d[1727];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1726] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1726] <= mhpmcounter_d[1726];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1725] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1725] <= mhpmcounter_d[1725];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1724] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1724] <= mhpmcounter_d[1724];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1723] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1723] <= mhpmcounter_d[1723];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1722] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1722] <= mhpmcounter_d[1722];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1721] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1721] <= mhpmcounter_d[1721];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1720] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1720] <= mhpmcounter_d[1720];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1719] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1719] <= mhpmcounter_d[1719];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1718] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1718] <= mhpmcounter_d[1718];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1717] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1717] <= mhpmcounter_d[1717];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1716] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1716] <= mhpmcounter_d[1716];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1715] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1715] <= mhpmcounter_d[1715];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1714] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1714] <= mhpmcounter_d[1714];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1713] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1713] <= mhpmcounter_d[1713];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1712] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1712] <= mhpmcounter_d[1712];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1711] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1711] <= mhpmcounter_d[1711];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1710] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1710] <= mhpmcounter_d[1710];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1709] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1709] <= mhpmcounter_d[1709];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1708] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1708] <= mhpmcounter_d[1708];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1707] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1707] <= mhpmcounter_d[1707];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1706] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1706] <= mhpmcounter_d[1706];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1705] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1705] <= mhpmcounter_d[1705];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1704] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1704] <= mhpmcounter_d[1704];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1703] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1703] <= mhpmcounter_d[1703];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1702] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1702] <= mhpmcounter_d[1702];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1701] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1701] <= mhpmcounter_d[1701];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1700] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1700] <= mhpmcounter_d[1700];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1699] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1699] <= mhpmcounter_d[1699];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1698] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1698] <= mhpmcounter_d[1698];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1697] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1697] <= mhpmcounter_d[1697];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1696] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1696] <= mhpmcounter_d[1696];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1695] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1695] <= mhpmcounter_d[1695];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1694] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1694] <= mhpmcounter_d[1694];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1693] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1693] <= mhpmcounter_d[1693];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1692] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1692] <= mhpmcounter_d[1692];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1691] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1691] <= mhpmcounter_d[1691];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1690] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1690] <= mhpmcounter_d[1690];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1689] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1689] <= mhpmcounter_d[1689];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1688] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1688] <= mhpmcounter_d[1688];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1687] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1687] <= mhpmcounter_d[1687];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1686] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1686] <= mhpmcounter_d[1686];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1685] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1685] <= mhpmcounter_d[1685];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1684] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1684] <= mhpmcounter_d[1684];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1683] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1683] <= mhpmcounter_d[1683];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1682] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1682] <= mhpmcounter_d[1682];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1681] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1681] <= mhpmcounter_d[1681];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1680] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1680] <= mhpmcounter_d[1680];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1679] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1679] <= mhpmcounter_d[1679];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1678] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1678] <= mhpmcounter_d[1678];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1677] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1677] <= mhpmcounter_d[1677];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1676] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1676] <= mhpmcounter_d[1676];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1675] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1675] <= mhpmcounter_d[1675];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1674] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1674] <= mhpmcounter_d[1674];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1673] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1673] <= mhpmcounter_d[1673];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1672] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1672] <= mhpmcounter_d[1672];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1671] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1671] <= mhpmcounter_d[1671];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1670] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1670] <= mhpmcounter_d[1670];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1669] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1669] <= mhpmcounter_d[1669];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1668] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1668] <= mhpmcounter_d[1668];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1667] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1667] <= mhpmcounter_d[1667];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1666] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1666] <= mhpmcounter_d[1666];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1665] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1665] <= mhpmcounter_d[1665];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1664] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1664] <= mhpmcounter_d[1664];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1663] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1663] <= mhpmcounter_d[1663];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1662] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1662] <= mhpmcounter_d[1662];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1661] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1661] <= mhpmcounter_d[1661];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1660] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1660] <= mhpmcounter_d[1660];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1659] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1659] <= mhpmcounter_d[1659];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1658] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1658] <= mhpmcounter_d[1658];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1657] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1657] <= mhpmcounter_d[1657];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1656] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1656] <= mhpmcounter_d[1656];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1655] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1655] <= mhpmcounter_d[1655];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1654] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1654] <= mhpmcounter_d[1654];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1653] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1653] <= mhpmcounter_d[1653];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1652] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1652] <= mhpmcounter_d[1652];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1651] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1651] <= mhpmcounter_d[1651];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1650] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1650] <= mhpmcounter_d[1650];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1649] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1649] <= mhpmcounter_d[1649];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1648] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1648] <= mhpmcounter_d[1648];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1647] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1647] <= mhpmcounter_d[1647];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1646] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1646] <= mhpmcounter_d[1646];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1645] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1645] <= mhpmcounter_d[1645];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1644] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1644] <= mhpmcounter_d[1644];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1643] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1643] <= mhpmcounter_d[1643];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1642] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1642] <= mhpmcounter_d[1642];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1641] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1641] <= mhpmcounter_d[1641];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1640] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1640] <= mhpmcounter_d[1640];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1639] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1639] <= mhpmcounter_d[1639];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1638] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1638] <= mhpmcounter_d[1638];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1637] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1637] <= mhpmcounter_d[1637];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1636] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1636] <= mhpmcounter_d[1636];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1635] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1635] <= mhpmcounter_d[1635];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1634] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1634] <= mhpmcounter_d[1634];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1633] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1633] <= mhpmcounter_d[1633];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1632] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1632] <= mhpmcounter_d[1632];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1631] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1631] <= mhpmcounter_d[1631];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1630] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1630] <= mhpmcounter_d[1630];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1629] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1629] <= mhpmcounter_d[1629];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1628] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1628] <= mhpmcounter_d[1628];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1627] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1627] <= mhpmcounter_d[1627];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1626] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1626] <= mhpmcounter_d[1626];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1625] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1625] <= mhpmcounter_d[1625];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1624] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1624] <= mhpmcounter_d[1624];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1623] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1623] <= mhpmcounter_d[1623];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1622] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1622] <= mhpmcounter_d[1622];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1621] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1621] <= mhpmcounter_d[1621];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1620] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1620] <= mhpmcounter_d[1620];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1619] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1619] <= mhpmcounter_d[1619];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1618] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1618] <= mhpmcounter_d[1618];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1617] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1617] <= mhpmcounter_d[1617];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1616] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1616] <= mhpmcounter_d[1616];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1615] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1615] <= mhpmcounter_d[1615];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1614] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1614] <= mhpmcounter_d[1614];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1613] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1613] <= mhpmcounter_d[1613];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1612] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1612] <= mhpmcounter_d[1612];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1611] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1611] <= mhpmcounter_d[1611];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1610] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1610] <= mhpmcounter_d[1610];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1609] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1609] <= mhpmcounter_d[1609];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1608] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1608] <= mhpmcounter_d[1608];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1607] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1607] <= mhpmcounter_d[1607];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1606] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1606] <= mhpmcounter_d[1606];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1605] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1605] <= mhpmcounter_d[1605];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1604] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1604] <= mhpmcounter_d[1604];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1603] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1603] <= mhpmcounter_d[1603];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1602] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1602] <= mhpmcounter_d[1602];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1601] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1601] <= mhpmcounter_d[1601];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1600] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1600] <= mhpmcounter_d[1600];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1599] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1599] <= mhpmcounter_d[1599];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1598] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1598] <= mhpmcounter_d[1598];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1597] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1597] <= mhpmcounter_d[1597];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1596] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1596] <= mhpmcounter_d[1596];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1595] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1595] <= mhpmcounter_d[1595];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1594] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1594] <= mhpmcounter_d[1594];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1593] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1593] <= mhpmcounter_d[1593];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1592] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1592] <= mhpmcounter_d[1592];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1591] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1591] <= mhpmcounter_d[1591];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1590] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1590] <= mhpmcounter_d[1590];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1589] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1589] <= mhpmcounter_d[1589];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1588] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1588] <= mhpmcounter_d[1588];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1587] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1587] <= mhpmcounter_d[1587];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1586] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1586] <= mhpmcounter_d[1586];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1585] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1585] <= mhpmcounter_d[1585];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1584] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1584] <= mhpmcounter_d[1584];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1583] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1583] <= mhpmcounter_d[1583];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1582] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1582] <= mhpmcounter_d[1582];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1581] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1581] <= mhpmcounter_d[1581];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1580] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1580] <= mhpmcounter_d[1580];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1579] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1579] <= mhpmcounter_d[1579];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1578] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1578] <= mhpmcounter_d[1578];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1577] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1577] <= mhpmcounter_d[1577];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1576] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1576] <= mhpmcounter_d[1576];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1575] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1575] <= mhpmcounter_d[1575];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1574] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1574] <= mhpmcounter_d[1574];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1573] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1573] <= mhpmcounter_d[1573];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1572] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1572] <= mhpmcounter_d[1572];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1571] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1571] <= mhpmcounter_d[1571];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1570] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1570] <= mhpmcounter_d[1570];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1569] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1569] <= mhpmcounter_d[1569];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1568] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1568] <= mhpmcounter_d[1568];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1567] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1567] <= mhpmcounter_d[1567];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1566] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1566] <= mhpmcounter_d[1566];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1565] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1565] <= mhpmcounter_d[1565];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1564] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1564] <= mhpmcounter_d[1564];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1563] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1563] <= mhpmcounter_d[1563];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1562] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1562] <= mhpmcounter_d[1562];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1561] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1561] <= mhpmcounter_d[1561];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1560] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1560] <= mhpmcounter_d[1560];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1559] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1559] <= mhpmcounter_d[1559];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1558] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1558] <= mhpmcounter_d[1558];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1557] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1557] <= mhpmcounter_d[1557];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1556] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1556] <= mhpmcounter_d[1556];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1555] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1555] <= mhpmcounter_d[1555];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1554] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1554] <= mhpmcounter_d[1554];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1553] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1553] <= mhpmcounter_d[1553];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1552] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1552] <= mhpmcounter_d[1552];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1551] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1551] <= mhpmcounter_d[1551];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1550] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1550] <= mhpmcounter_d[1550];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1549] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1549] <= mhpmcounter_d[1549];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1548] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1548] <= mhpmcounter_d[1548];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1547] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1547] <= mhpmcounter_d[1547];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1546] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1546] <= mhpmcounter_d[1546];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1545] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1545] <= mhpmcounter_d[1545];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1544] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1544] <= mhpmcounter_d[1544];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1543] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1543] <= mhpmcounter_d[1543];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1542] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1542] <= mhpmcounter_d[1542];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1541] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1541] <= mhpmcounter_d[1541];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1540] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1540] <= mhpmcounter_d[1540];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1539] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1539] <= mhpmcounter_d[1539];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1538] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1538] <= mhpmcounter_d[1538];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1537] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1537] <= mhpmcounter_d[1537];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1536] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1536] <= mhpmcounter_d[1536];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1535] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1535] <= mhpmcounter_d[1535];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1534] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1534] <= mhpmcounter_d[1534];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1533] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1533] <= mhpmcounter_d[1533];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1532] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1532] <= mhpmcounter_d[1532];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1531] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1531] <= mhpmcounter_d[1531];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1530] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1530] <= mhpmcounter_d[1530];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1529] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1529] <= mhpmcounter_d[1529];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1528] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1528] <= mhpmcounter_d[1528];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1527] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1527] <= mhpmcounter_d[1527];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1526] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1526] <= mhpmcounter_d[1526];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1525] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1525] <= mhpmcounter_d[1525];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1524] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1524] <= mhpmcounter_d[1524];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1523] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1523] <= mhpmcounter_d[1523];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1522] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1522] <= mhpmcounter_d[1522];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1521] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1521] <= mhpmcounter_d[1521];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1520] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1520] <= mhpmcounter_d[1520];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1519] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1519] <= mhpmcounter_d[1519];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1518] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1518] <= mhpmcounter_d[1518];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1517] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1517] <= mhpmcounter_d[1517];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1516] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1516] <= mhpmcounter_d[1516];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1515] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1515] <= mhpmcounter_d[1515];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1514] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1514] <= mhpmcounter_d[1514];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1513] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1513] <= mhpmcounter_d[1513];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1512] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1512] <= mhpmcounter_d[1512];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1511] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1511] <= mhpmcounter_d[1511];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1510] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1510] <= mhpmcounter_d[1510];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1509] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1509] <= mhpmcounter_d[1509];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1508] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1508] <= mhpmcounter_d[1508];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1507] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1507] <= mhpmcounter_d[1507];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1506] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1506] <= mhpmcounter_d[1506];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1505] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1505] <= mhpmcounter_d[1505];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1504] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1504] <= mhpmcounter_d[1504];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1503] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1503] <= mhpmcounter_d[1503];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1502] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1502] <= mhpmcounter_d[1502];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1501] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1501] <= mhpmcounter_d[1501];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1500] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1500] <= mhpmcounter_d[1500];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1499] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1499] <= mhpmcounter_d[1499];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1498] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1498] <= mhpmcounter_d[1498];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1497] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1497] <= mhpmcounter_d[1497];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1496] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1496] <= mhpmcounter_d[1496];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1495] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1495] <= mhpmcounter_d[1495];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1494] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1494] <= mhpmcounter_d[1494];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1493] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1493] <= mhpmcounter_d[1493];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1492] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1492] <= mhpmcounter_d[1492];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1491] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1491] <= mhpmcounter_d[1491];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1490] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1490] <= mhpmcounter_d[1490];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1489] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1489] <= mhpmcounter_d[1489];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1488] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1488] <= mhpmcounter_d[1488];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1487] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1487] <= mhpmcounter_d[1487];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1486] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1486] <= mhpmcounter_d[1486];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1485] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1485] <= mhpmcounter_d[1485];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1484] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1484] <= mhpmcounter_d[1484];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1483] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1483] <= mhpmcounter_d[1483];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1482] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1482] <= mhpmcounter_d[1482];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1481] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1481] <= mhpmcounter_d[1481];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1480] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1480] <= mhpmcounter_d[1480];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1479] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1479] <= mhpmcounter_d[1479];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1478] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1478] <= mhpmcounter_d[1478];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1477] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1477] <= mhpmcounter_d[1477];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1476] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1476] <= mhpmcounter_d[1476];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1475] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1475] <= mhpmcounter_d[1475];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1474] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1474] <= mhpmcounter_d[1474];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1473] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1473] <= mhpmcounter_d[1473];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1472] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1472] <= mhpmcounter_d[1472];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1471] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1471] <= mhpmcounter_d[1471];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1470] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1470] <= mhpmcounter_d[1470];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1469] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1469] <= mhpmcounter_d[1469];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1468] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1468] <= mhpmcounter_d[1468];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1467] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1467] <= mhpmcounter_d[1467];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1466] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1466] <= mhpmcounter_d[1466];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1465] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1465] <= mhpmcounter_d[1465];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1464] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1464] <= mhpmcounter_d[1464];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1463] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1463] <= mhpmcounter_d[1463];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1462] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1462] <= mhpmcounter_d[1462];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1461] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1461] <= mhpmcounter_d[1461];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1460] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1460] <= mhpmcounter_d[1460];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1459] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1459] <= mhpmcounter_d[1459];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1458] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1458] <= mhpmcounter_d[1458];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1457] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1457] <= mhpmcounter_d[1457];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1456] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1456] <= mhpmcounter_d[1456];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1455] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1455] <= mhpmcounter_d[1455];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1454] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1454] <= mhpmcounter_d[1454];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1453] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1453] <= mhpmcounter_d[1453];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1452] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1452] <= mhpmcounter_d[1452];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1451] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1451] <= mhpmcounter_d[1451];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1450] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1450] <= mhpmcounter_d[1450];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1449] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1449] <= mhpmcounter_d[1449];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1448] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1448] <= mhpmcounter_d[1448];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1447] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1447] <= mhpmcounter_d[1447];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1446] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1446] <= mhpmcounter_d[1446];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1445] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1445] <= mhpmcounter_d[1445];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1444] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1444] <= mhpmcounter_d[1444];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1443] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1443] <= mhpmcounter_d[1443];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1442] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1442] <= mhpmcounter_d[1442];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1441] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1441] <= mhpmcounter_d[1441];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1440] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1440] <= mhpmcounter_d[1440];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1439] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1439] <= mhpmcounter_d[1439];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1438] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1438] <= mhpmcounter_d[1438];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1437] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1437] <= mhpmcounter_d[1437];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1436] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1436] <= mhpmcounter_d[1436];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1435] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1435] <= mhpmcounter_d[1435];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1434] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1434] <= mhpmcounter_d[1434];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1433] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1433] <= mhpmcounter_d[1433];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1432] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1432] <= mhpmcounter_d[1432];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1431] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1431] <= mhpmcounter_d[1431];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1430] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1430] <= mhpmcounter_d[1430];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1429] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1429] <= mhpmcounter_d[1429];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1428] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1428] <= mhpmcounter_d[1428];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1427] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1427] <= mhpmcounter_d[1427];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1426] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1426] <= mhpmcounter_d[1426];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1425] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1425] <= mhpmcounter_d[1425];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1424] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1424] <= mhpmcounter_d[1424];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1423] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1423] <= mhpmcounter_d[1423];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1422] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1422] <= mhpmcounter_d[1422];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1421] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1421] <= mhpmcounter_d[1421];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1420] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1420] <= mhpmcounter_d[1420];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1419] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1419] <= mhpmcounter_d[1419];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1418] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1418] <= mhpmcounter_d[1418];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1417] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1417] <= mhpmcounter_d[1417];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1416] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1416] <= mhpmcounter_d[1416];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1415] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1415] <= mhpmcounter_d[1415];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1414] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1414] <= mhpmcounter_d[1414];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1413] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1413] <= mhpmcounter_d[1413];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1412] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1412] <= mhpmcounter_d[1412];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1411] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1411] <= mhpmcounter_d[1411];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1410] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1410] <= mhpmcounter_d[1410];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1409] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1409] <= mhpmcounter_d[1409];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1408] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1408] <= mhpmcounter_d[1408];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1407] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1407] <= mhpmcounter_d[1407];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1406] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1406] <= mhpmcounter_d[1406];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1405] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1405] <= mhpmcounter_d[1405];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1404] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1404] <= mhpmcounter_d[1404];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1403] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1403] <= mhpmcounter_d[1403];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1402] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1402] <= mhpmcounter_d[1402];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1401] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1401] <= mhpmcounter_d[1401];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1400] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1400] <= mhpmcounter_d[1400];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1399] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1399] <= mhpmcounter_d[1399];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1398] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1398] <= mhpmcounter_d[1398];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1397] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1397] <= mhpmcounter_d[1397];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1396] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1396] <= mhpmcounter_d[1396];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1395] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1395] <= mhpmcounter_d[1395];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1394] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1394] <= mhpmcounter_d[1394];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1393] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1393] <= mhpmcounter_d[1393];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1392] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1392] <= mhpmcounter_d[1392];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1391] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1391] <= mhpmcounter_d[1391];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1390] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1390] <= mhpmcounter_d[1390];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1389] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1389] <= mhpmcounter_d[1389];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1388] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1388] <= mhpmcounter_d[1388];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1387] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1387] <= mhpmcounter_d[1387];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1386] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1386] <= mhpmcounter_d[1386];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1385] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1385] <= mhpmcounter_d[1385];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1384] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1384] <= mhpmcounter_d[1384];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1383] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1383] <= mhpmcounter_d[1383];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1382] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1382] <= mhpmcounter_d[1382];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1381] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1381] <= mhpmcounter_d[1381];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1380] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1380] <= mhpmcounter_d[1380];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1379] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1379] <= mhpmcounter_d[1379];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1378] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1378] <= mhpmcounter_d[1378];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1377] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1377] <= mhpmcounter_d[1377];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1376] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1376] <= mhpmcounter_d[1376];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1375] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1375] <= mhpmcounter_d[1375];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1374] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1374] <= mhpmcounter_d[1374];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1373] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1373] <= mhpmcounter_d[1373];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1372] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1372] <= mhpmcounter_d[1372];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1371] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1371] <= mhpmcounter_d[1371];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1370] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1370] <= mhpmcounter_d[1370];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1369] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1369] <= mhpmcounter_d[1369];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1368] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1368] <= mhpmcounter_d[1368];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1367] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1367] <= mhpmcounter_d[1367];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1366] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1366] <= mhpmcounter_d[1366];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1365] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1365] <= mhpmcounter_d[1365];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1364] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1364] <= mhpmcounter_d[1364];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1363] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1363] <= mhpmcounter_d[1363];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1362] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1362] <= mhpmcounter_d[1362];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1361] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1361] <= mhpmcounter_d[1361];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1360] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1360] <= mhpmcounter_d[1360];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1359] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1359] <= mhpmcounter_d[1359];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1358] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1358] <= mhpmcounter_d[1358];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1357] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1357] <= mhpmcounter_d[1357];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1356] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1356] <= mhpmcounter_d[1356];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1355] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1355] <= mhpmcounter_d[1355];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1354] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1354] <= mhpmcounter_d[1354];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1353] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1353] <= mhpmcounter_d[1353];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1352] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1352] <= mhpmcounter_d[1352];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1351] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1351] <= mhpmcounter_d[1351];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1350] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1350] <= mhpmcounter_d[1350];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1349] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1349] <= mhpmcounter_d[1349];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1348] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1348] <= mhpmcounter_d[1348];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1347] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1347] <= mhpmcounter_d[1347];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1346] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1346] <= mhpmcounter_d[1346];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1345] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1345] <= mhpmcounter_d[1345];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1344] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1344] <= mhpmcounter_d[1344];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1343] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1343] <= mhpmcounter_d[1343];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1342] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1342] <= mhpmcounter_d[1342];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1341] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1341] <= mhpmcounter_d[1341];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1340] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1340] <= mhpmcounter_d[1340];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1339] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1339] <= mhpmcounter_d[1339];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1338] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1338] <= mhpmcounter_d[1338];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1337] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1337] <= mhpmcounter_d[1337];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1336] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1336] <= mhpmcounter_d[1336];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1335] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1335] <= mhpmcounter_d[1335];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1334] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1334] <= mhpmcounter_d[1334];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1333] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1333] <= mhpmcounter_d[1333];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1332] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1332] <= mhpmcounter_d[1332];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1331] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1331] <= mhpmcounter_d[1331];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1330] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1330] <= mhpmcounter_d[1330];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1329] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1329] <= mhpmcounter_d[1329];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1328] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1328] <= mhpmcounter_d[1328];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1327] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1327] <= mhpmcounter_d[1327];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1326] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1326] <= mhpmcounter_d[1326];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1325] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1325] <= mhpmcounter_d[1325];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1324] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1324] <= mhpmcounter_d[1324];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1323] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1323] <= mhpmcounter_d[1323];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1322] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1322] <= mhpmcounter_d[1322];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1321] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1321] <= mhpmcounter_d[1321];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1320] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1320] <= mhpmcounter_d[1320];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1319] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1319] <= mhpmcounter_d[1319];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1318] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1318] <= mhpmcounter_d[1318];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1317] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1317] <= mhpmcounter_d[1317];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1316] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1316] <= mhpmcounter_d[1316];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1315] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1315] <= mhpmcounter_d[1315];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1314] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1314] <= mhpmcounter_d[1314];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1313] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1313] <= mhpmcounter_d[1313];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1312] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1312] <= mhpmcounter_d[1312];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1311] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1311] <= mhpmcounter_d[1311];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1310] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1310] <= mhpmcounter_d[1310];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1309] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1309] <= mhpmcounter_d[1309];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1308] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1308] <= mhpmcounter_d[1308];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1307] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1307] <= mhpmcounter_d[1307];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1306] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1306] <= mhpmcounter_d[1306];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1305] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1305] <= mhpmcounter_d[1305];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1304] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1304] <= mhpmcounter_d[1304];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1303] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1303] <= mhpmcounter_d[1303];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1302] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1302] <= mhpmcounter_d[1302];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1301] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1301] <= mhpmcounter_d[1301];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1300] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1300] <= mhpmcounter_d[1300];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1299] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1299] <= mhpmcounter_d[1299];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1298] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1298] <= mhpmcounter_d[1298];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1297] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1297] <= mhpmcounter_d[1297];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1296] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1296] <= mhpmcounter_d[1296];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1295] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1295] <= mhpmcounter_d[1295];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1294] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1294] <= mhpmcounter_d[1294];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1293] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1293] <= mhpmcounter_d[1293];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1292] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1292] <= mhpmcounter_d[1292];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1291] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1291] <= mhpmcounter_d[1291];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1290] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1290] <= mhpmcounter_d[1290];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1289] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1289] <= mhpmcounter_d[1289];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1288] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1288] <= mhpmcounter_d[1288];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1287] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1287] <= mhpmcounter_d[1287];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1286] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1286] <= mhpmcounter_d[1286];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1285] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1285] <= mhpmcounter_d[1285];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1284] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1284] <= mhpmcounter_d[1284];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1283] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1283] <= mhpmcounter_d[1283];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1282] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1282] <= mhpmcounter_d[1282];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1281] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1281] <= mhpmcounter_d[1281];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1280] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1280] <= mhpmcounter_d[1280];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1279] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1279] <= mhpmcounter_d[1279];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1278] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1278] <= mhpmcounter_d[1278];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1277] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1277] <= mhpmcounter_d[1277];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1276] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1276] <= mhpmcounter_d[1276];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1275] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1275] <= mhpmcounter_d[1275];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1274] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1274] <= mhpmcounter_d[1274];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1273] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1273] <= mhpmcounter_d[1273];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1272] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1272] <= mhpmcounter_d[1272];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1271] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1271] <= mhpmcounter_d[1271];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1270] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1270] <= mhpmcounter_d[1270];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1269] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1269] <= mhpmcounter_d[1269];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1268] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1268] <= mhpmcounter_d[1268];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1267] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1267] <= mhpmcounter_d[1267];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1266] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1266] <= mhpmcounter_d[1266];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1265] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1265] <= mhpmcounter_d[1265];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1264] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1264] <= mhpmcounter_d[1264];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1263] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1263] <= mhpmcounter_d[1263];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1262] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1262] <= mhpmcounter_d[1262];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1261] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1261] <= mhpmcounter_d[1261];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1260] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1260] <= mhpmcounter_d[1260];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1259] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1259] <= mhpmcounter_d[1259];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1258] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1258] <= mhpmcounter_d[1258];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1257] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1257] <= mhpmcounter_d[1257];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1256] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1256] <= mhpmcounter_d[1256];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1255] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1255] <= mhpmcounter_d[1255];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1254] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1254] <= mhpmcounter_d[1254];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1253] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1253] <= mhpmcounter_d[1253];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1252] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1252] <= mhpmcounter_d[1252];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1251] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1251] <= mhpmcounter_d[1251];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1250] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1250] <= mhpmcounter_d[1250];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1249] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1249] <= mhpmcounter_d[1249];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1248] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1248] <= mhpmcounter_d[1248];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1247] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1247] <= mhpmcounter_d[1247];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1246] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1246] <= mhpmcounter_d[1246];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1245] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1245] <= mhpmcounter_d[1245];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1244] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1244] <= mhpmcounter_d[1244];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1243] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1243] <= mhpmcounter_d[1243];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1242] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1242] <= mhpmcounter_d[1242];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1241] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1241] <= mhpmcounter_d[1241];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1240] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1240] <= mhpmcounter_d[1240];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1239] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1239] <= mhpmcounter_d[1239];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1238] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1238] <= mhpmcounter_d[1238];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1237] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1237] <= mhpmcounter_d[1237];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1236] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1236] <= mhpmcounter_d[1236];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1235] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1235] <= mhpmcounter_d[1235];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1234] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1234] <= mhpmcounter_d[1234];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1233] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1233] <= mhpmcounter_d[1233];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1232] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1232] <= mhpmcounter_d[1232];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1231] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1231] <= mhpmcounter_d[1231];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1230] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1230] <= mhpmcounter_d[1230];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1229] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1229] <= mhpmcounter_d[1229];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1228] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1228] <= mhpmcounter_d[1228];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1227] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1227] <= mhpmcounter_d[1227];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1226] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1226] <= mhpmcounter_d[1226];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1225] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1225] <= mhpmcounter_d[1225];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1224] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1224] <= mhpmcounter_d[1224];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1223] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1223] <= mhpmcounter_d[1223];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1222] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1222] <= mhpmcounter_d[1222];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1221] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1221] <= mhpmcounter_d[1221];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1220] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1220] <= mhpmcounter_d[1220];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1219] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1219] <= mhpmcounter_d[1219];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1218] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1218] <= mhpmcounter_d[1218];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1217] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1217] <= mhpmcounter_d[1217];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1216] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1216] <= mhpmcounter_d[1216];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1215] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1215] <= mhpmcounter_d[1215];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1214] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1214] <= mhpmcounter_d[1214];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1213] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1213] <= mhpmcounter_d[1213];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1212] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1212] <= mhpmcounter_d[1212];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1211] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1211] <= mhpmcounter_d[1211];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1210] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1210] <= mhpmcounter_d[1210];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1209] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1209] <= mhpmcounter_d[1209];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1208] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1208] <= mhpmcounter_d[1208];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1207] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1207] <= mhpmcounter_d[1207];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1206] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1206] <= mhpmcounter_d[1206];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1205] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1205] <= mhpmcounter_d[1205];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1204] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1204] <= mhpmcounter_d[1204];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1203] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1203] <= mhpmcounter_d[1203];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1202] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1202] <= mhpmcounter_d[1202];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1201] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1201] <= mhpmcounter_d[1201];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1200] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1200] <= mhpmcounter_d[1200];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1199] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1199] <= mhpmcounter_d[1199];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1198] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1198] <= mhpmcounter_d[1198];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1197] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1197] <= mhpmcounter_d[1197];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1196] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1196] <= mhpmcounter_d[1196];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1195] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1195] <= mhpmcounter_d[1195];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1194] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1194] <= mhpmcounter_d[1194];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1193] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1193] <= mhpmcounter_d[1193];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1192] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1192] <= mhpmcounter_d[1192];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1191] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1191] <= mhpmcounter_d[1191];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1190] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1190] <= mhpmcounter_d[1190];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1189] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1189] <= mhpmcounter_d[1189];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1188] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1188] <= mhpmcounter_d[1188];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1187] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1187] <= mhpmcounter_d[1187];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1186] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1186] <= mhpmcounter_d[1186];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1185] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1185] <= mhpmcounter_d[1185];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1184] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1184] <= mhpmcounter_d[1184];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1183] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1183] <= mhpmcounter_d[1183];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1182] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1182] <= mhpmcounter_d[1182];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1181] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1181] <= mhpmcounter_d[1181];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1180] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1180] <= mhpmcounter_d[1180];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1179] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1179] <= mhpmcounter_d[1179];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1178] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1178] <= mhpmcounter_d[1178];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1177] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1177] <= mhpmcounter_d[1177];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1176] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1176] <= mhpmcounter_d[1176];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1175] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1175] <= mhpmcounter_d[1175];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1174] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1174] <= mhpmcounter_d[1174];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1173] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1173] <= mhpmcounter_d[1173];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1172] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1172] <= mhpmcounter_d[1172];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1171] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1171] <= mhpmcounter_d[1171];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1170] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1170] <= mhpmcounter_d[1170];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1169] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1169] <= mhpmcounter_d[1169];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1168] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1168] <= mhpmcounter_d[1168];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1167] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1167] <= mhpmcounter_d[1167];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1166] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1166] <= mhpmcounter_d[1166];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1165] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1165] <= mhpmcounter_d[1165];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1164] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1164] <= mhpmcounter_d[1164];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1163] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1163] <= mhpmcounter_d[1163];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1162] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1162] <= mhpmcounter_d[1162];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1161] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1161] <= mhpmcounter_d[1161];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1160] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1160] <= mhpmcounter_d[1160];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1159] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1159] <= mhpmcounter_d[1159];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1158] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1158] <= mhpmcounter_d[1158];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1157] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1157] <= mhpmcounter_d[1157];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1156] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1156] <= mhpmcounter_d[1156];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1155] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1155] <= mhpmcounter_d[1155];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1154] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1154] <= mhpmcounter_d[1154];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1153] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1153] <= mhpmcounter_d[1153];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1152] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1152] <= mhpmcounter_d[1152];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1151] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1151] <= mhpmcounter_d[1151];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1150] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1150] <= mhpmcounter_d[1150];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1149] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1149] <= mhpmcounter_d[1149];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1148] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1148] <= mhpmcounter_d[1148];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1147] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1147] <= mhpmcounter_d[1147];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1146] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1146] <= mhpmcounter_d[1146];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1145] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1145] <= mhpmcounter_d[1145];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1144] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1144] <= mhpmcounter_d[1144];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1143] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1143] <= mhpmcounter_d[1143];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1142] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1142] <= mhpmcounter_d[1142];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1141] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1141] <= mhpmcounter_d[1141];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1140] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1140] <= mhpmcounter_d[1140];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1139] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1139] <= mhpmcounter_d[1139];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1138] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1138] <= mhpmcounter_d[1138];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1137] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1137] <= mhpmcounter_d[1137];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1136] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1136] <= mhpmcounter_d[1136];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1135] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1135] <= mhpmcounter_d[1135];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1134] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1134] <= mhpmcounter_d[1134];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1133] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1133] <= mhpmcounter_d[1133];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1132] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1132] <= mhpmcounter_d[1132];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1131] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1131] <= mhpmcounter_d[1131];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1130] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1130] <= mhpmcounter_d[1130];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1129] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1129] <= mhpmcounter_d[1129];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1128] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1128] <= mhpmcounter_d[1128];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1127] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1127] <= mhpmcounter_d[1127];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1126] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1126] <= mhpmcounter_d[1126];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1125] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1125] <= mhpmcounter_d[1125];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1124] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1124] <= mhpmcounter_d[1124];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1123] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1123] <= mhpmcounter_d[1123];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1122] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1122] <= mhpmcounter_d[1122];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1121] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1121] <= mhpmcounter_d[1121];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1120] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1120] <= mhpmcounter_d[1120];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1119] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1119] <= mhpmcounter_d[1119];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1118] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1118] <= mhpmcounter_d[1118];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1117] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1117] <= mhpmcounter_d[1117];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1116] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1116] <= mhpmcounter_d[1116];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1115] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1115] <= mhpmcounter_d[1115];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1114] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1114] <= mhpmcounter_d[1114];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1113] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1113] <= mhpmcounter_d[1113];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1112] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1112] <= mhpmcounter_d[1112];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1111] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1111] <= mhpmcounter_d[1111];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1110] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1110] <= mhpmcounter_d[1110];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1109] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1109] <= mhpmcounter_d[1109];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1108] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1108] <= mhpmcounter_d[1108];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1107] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1107] <= mhpmcounter_d[1107];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1106] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1106] <= mhpmcounter_d[1106];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1105] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1105] <= mhpmcounter_d[1105];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1104] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1104] <= mhpmcounter_d[1104];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1103] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1103] <= mhpmcounter_d[1103];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1102] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1102] <= mhpmcounter_d[1102];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1101] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1101] <= mhpmcounter_d[1101];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1100] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1100] <= mhpmcounter_d[1100];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1099] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1099] <= mhpmcounter_d[1099];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1098] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1098] <= mhpmcounter_d[1098];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1097] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1097] <= mhpmcounter_d[1097];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1096] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1096] <= mhpmcounter_d[1096];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1095] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1095] <= mhpmcounter_d[1095];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1094] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1094] <= mhpmcounter_d[1094];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1093] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1093] <= mhpmcounter_d[1093];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1092] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1092] <= mhpmcounter_d[1092];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1091] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1091] <= mhpmcounter_d[1091];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1090] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1090] <= mhpmcounter_d[1090];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1089] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1089] <= mhpmcounter_d[1089];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1088] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1088] <= mhpmcounter_d[1088];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1087] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1087] <= mhpmcounter_d[1087];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1086] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1086] <= mhpmcounter_d[1086];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1085] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1085] <= mhpmcounter_d[1085];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1084] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1084] <= mhpmcounter_d[1084];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1083] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1083] <= mhpmcounter_d[1083];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1082] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1082] <= mhpmcounter_d[1082];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1081] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1081] <= mhpmcounter_d[1081];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1080] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1080] <= mhpmcounter_d[1080];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1079] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1079] <= mhpmcounter_d[1079];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1078] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1078] <= mhpmcounter_d[1078];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1077] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1077] <= mhpmcounter_d[1077];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1076] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1076] <= mhpmcounter_d[1076];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1075] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1075] <= mhpmcounter_d[1075];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1074] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1074] <= mhpmcounter_d[1074];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1073] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1073] <= mhpmcounter_d[1073];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1072] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1072] <= mhpmcounter_d[1072];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1071] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1071] <= mhpmcounter_d[1071];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1070] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1070] <= mhpmcounter_d[1070];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1069] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1069] <= mhpmcounter_d[1069];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1068] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1068] <= mhpmcounter_d[1068];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1067] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1067] <= mhpmcounter_d[1067];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1066] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1066] <= mhpmcounter_d[1066];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1065] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1065] <= mhpmcounter_d[1065];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1064] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1064] <= mhpmcounter_d[1064];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1063] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1063] <= mhpmcounter_d[1063];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1062] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1062] <= mhpmcounter_d[1062];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1061] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1061] <= mhpmcounter_d[1061];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1060] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1060] <= mhpmcounter_d[1060];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1059] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1059] <= mhpmcounter_d[1059];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1058] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1058] <= mhpmcounter_d[1058];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1057] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1057] <= mhpmcounter_d[1057];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1056] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1056] <= mhpmcounter_d[1056];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1055] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1055] <= mhpmcounter_d[1055];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1054] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1054] <= mhpmcounter_d[1054];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1053] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1053] <= mhpmcounter_d[1053];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1052] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1052] <= mhpmcounter_d[1052];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1051] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1051] <= mhpmcounter_d[1051];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1050] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1050] <= mhpmcounter_d[1050];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1049] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1049] <= mhpmcounter_d[1049];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1048] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1048] <= mhpmcounter_d[1048];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1047] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1047] <= mhpmcounter_d[1047];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1046] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1046] <= mhpmcounter_d[1046];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1045] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1045] <= mhpmcounter_d[1045];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1044] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1044] <= mhpmcounter_d[1044];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1043] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1043] <= mhpmcounter_d[1043];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1042] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1042] <= mhpmcounter_d[1042];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1041] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1041] <= mhpmcounter_d[1041];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1040] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1040] <= mhpmcounter_d[1040];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1039] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1039] <= mhpmcounter_d[1039];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1038] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1038] <= mhpmcounter_d[1038];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1037] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1037] <= mhpmcounter_d[1037];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1036] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1036] <= mhpmcounter_d[1036];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1035] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1035] <= mhpmcounter_d[1035];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1034] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1034] <= mhpmcounter_d[1034];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1033] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1033] <= mhpmcounter_d[1033];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1032] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1032] <= mhpmcounter_d[1032];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1031] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1031] <= mhpmcounter_d[1031];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1030] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1030] <= mhpmcounter_d[1030];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1029] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1029] <= mhpmcounter_d[1029];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1028] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1028] <= mhpmcounter_d[1028];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1027] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1027] <= mhpmcounter_d[1027];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1026] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1026] <= mhpmcounter_d[1026];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1025] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1025] <= mhpmcounter_d[1025];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1024] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1024] <= mhpmcounter_d[1024];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1023] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1023] <= mhpmcounter_d[1023];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1022] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1022] <= mhpmcounter_d[1022];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1021] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1021] <= mhpmcounter_d[1021];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1020] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1020] <= mhpmcounter_d[1020];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1019] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1019] <= mhpmcounter_d[1019];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1018] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1018] <= mhpmcounter_d[1018];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1017] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1017] <= mhpmcounter_d[1017];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1016] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1016] <= mhpmcounter_d[1016];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1015] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1015] <= mhpmcounter_d[1015];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1014] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1014] <= mhpmcounter_d[1014];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1013] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1013] <= mhpmcounter_d[1013];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1012] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1012] <= mhpmcounter_d[1012];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1011] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1011] <= mhpmcounter_d[1011];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1010] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1010] <= mhpmcounter_d[1010];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1009] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1009] <= mhpmcounter_d[1009];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1008] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1008] <= mhpmcounter_d[1008];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1007] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1007] <= mhpmcounter_d[1007];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1006] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1006] <= mhpmcounter_d[1006];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1005] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1005] <= mhpmcounter_d[1005];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1004] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1004] <= mhpmcounter_d[1004];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1003] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1003] <= mhpmcounter_d[1003];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1002] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1002] <= mhpmcounter_d[1002];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1001] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1001] <= mhpmcounter_d[1001];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1000] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1000] <= mhpmcounter_d[1000];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[999] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[999] <= mhpmcounter_d[999];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[998] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[998] <= mhpmcounter_d[998];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[997] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[997] <= mhpmcounter_d[997];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[996] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[996] <= mhpmcounter_d[996];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[995] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[995] <= mhpmcounter_d[995];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[994] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[994] <= mhpmcounter_d[994];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[993] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[993] <= mhpmcounter_d[993];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[992] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[992] <= mhpmcounter_d[992];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[991] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[991] <= mhpmcounter_d[991];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[990] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[990] <= mhpmcounter_d[990];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[989] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[989] <= mhpmcounter_d[989];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[988] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[988] <= mhpmcounter_d[988];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[987] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[987] <= mhpmcounter_d[987];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[986] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[986] <= mhpmcounter_d[986];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[985] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[985] <= mhpmcounter_d[985];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[984] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[984] <= mhpmcounter_d[984];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[983] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[983] <= mhpmcounter_d[983];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[982] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[982] <= mhpmcounter_d[982];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[981] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[981] <= mhpmcounter_d[981];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[980] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[980] <= mhpmcounter_d[980];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[979] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[979] <= mhpmcounter_d[979];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[978] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[978] <= mhpmcounter_d[978];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[977] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[977] <= mhpmcounter_d[977];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[976] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[976] <= mhpmcounter_d[976];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[975] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[975] <= mhpmcounter_d[975];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[974] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[974] <= mhpmcounter_d[974];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[973] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[973] <= mhpmcounter_d[973];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[972] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[972] <= mhpmcounter_d[972];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[971] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[971] <= mhpmcounter_d[971];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[970] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[970] <= mhpmcounter_d[970];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[969] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[969] <= mhpmcounter_d[969];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[968] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[968] <= mhpmcounter_d[968];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[967] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[967] <= mhpmcounter_d[967];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[966] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[966] <= mhpmcounter_d[966];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[965] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[965] <= mhpmcounter_d[965];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[964] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[964] <= mhpmcounter_d[964];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[963] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[963] <= mhpmcounter_d[963];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[962] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[962] <= mhpmcounter_d[962];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[961] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[961] <= mhpmcounter_d[961];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[960] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[960] <= mhpmcounter_d[960];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[959] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[959] <= mhpmcounter_d[959];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[958] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[958] <= mhpmcounter_d[958];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[957] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[957] <= mhpmcounter_d[957];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[956] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[956] <= mhpmcounter_d[956];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[955] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[955] <= mhpmcounter_d[955];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[954] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[954] <= mhpmcounter_d[954];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[953] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[953] <= mhpmcounter_d[953];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[952] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[952] <= mhpmcounter_d[952];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[951] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[951] <= mhpmcounter_d[951];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[950] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[950] <= mhpmcounter_d[950];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[949] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[949] <= mhpmcounter_d[949];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[948] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[948] <= mhpmcounter_d[948];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[947] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[947] <= mhpmcounter_d[947];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[946] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[946] <= mhpmcounter_d[946];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[945] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[945] <= mhpmcounter_d[945];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[944] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[944] <= mhpmcounter_d[944];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[943] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[943] <= mhpmcounter_d[943];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[942] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[942] <= mhpmcounter_d[942];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[941] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[941] <= mhpmcounter_d[941];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[940] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[940] <= mhpmcounter_d[940];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[939] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[939] <= mhpmcounter_d[939];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[938] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[938] <= mhpmcounter_d[938];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[937] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[937] <= mhpmcounter_d[937];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[936] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[936] <= mhpmcounter_d[936];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[935] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[935] <= mhpmcounter_d[935];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[934] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[934] <= mhpmcounter_d[934];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[933] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[933] <= mhpmcounter_d[933];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[932] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[932] <= mhpmcounter_d[932];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[931] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[931] <= mhpmcounter_d[931];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[930] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[930] <= mhpmcounter_d[930];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[929] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[929] <= mhpmcounter_d[929];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[928] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[928] <= mhpmcounter_d[928];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[927] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[927] <= mhpmcounter_d[927];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[926] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[926] <= mhpmcounter_d[926];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[925] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[925] <= mhpmcounter_d[925];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[924] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[924] <= mhpmcounter_d[924];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[923] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[923] <= mhpmcounter_d[923];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[922] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[922] <= mhpmcounter_d[922];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[921] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[921] <= mhpmcounter_d[921];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[920] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[920] <= mhpmcounter_d[920];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[919] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[919] <= mhpmcounter_d[919];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[918] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[918] <= mhpmcounter_d[918];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[917] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[917] <= mhpmcounter_d[917];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[916] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[916] <= mhpmcounter_d[916];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[915] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[915] <= mhpmcounter_d[915];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[914] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[914] <= mhpmcounter_d[914];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[913] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[913] <= mhpmcounter_d[913];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[912] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[912] <= mhpmcounter_d[912];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[911] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[911] <= mhpmcounter_d[911];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[910] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[910] <= mhpmcounter_d[910];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[909] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[909] <= mhpmcounter_d[909];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[908] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[908] <= mhpmcounter_d[908];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[907] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[907] <= mhpmcounter_d[907];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[906] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[906] <= mhpmcounter_d[906];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[905] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[905] <= mhpmcounter_d[905];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[904] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[904] <= mhpmcounter_d[904];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[903] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[903] <= mhpmcounter_d[903];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[902] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[902] <= mhpmcounter_d[902];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[901] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[901] <= mhpmcounter_d[901];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[900] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[900] <= mhpmcounter_d[900];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[899] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[899] <= mhpmcounter_d[899];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[898] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[898] <= mhpmcounter_d[898];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[897] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[897] <= mhpmcounter_d[897];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[896] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[896] <= mhpmcounter_d[896];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[895] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[895] <= mhpmcounter_d[895];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[894] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[894] <= mhpmcounter_d[894];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[893] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[893] <= mhpmcounter_d[893];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[892] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[892] <= mhpmcounter_d[892];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[891] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[891] <= mhpmcounter_d[891];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[890] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[890] <= mhpmcounter_d[890];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[889] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[889] <= mhpmcounter_d[889];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[888] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[888] <= mhpmcounter_d[888];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[887] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[887] <= mhpmcounter_d[887];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[886] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[886] <= mhpmcounter_d[886];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[885] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[885] <= mhpmcounter_d[885];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[884] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[884] <= mhpmcounter_d[884];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[883] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[883] <= mhpmcounter_d[883];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[882] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[882] <= mhpmcounter_d[882];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[881] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[881] <= mhpmcounter_d[881];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[880] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[880] <= mhpmcounter_d[880];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[879] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[879] <= mhpmcounter_d[879];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[878] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[878] <= mhpmcounter_d[878];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[877] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[877] <= mhpmcounter_d[877];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[876] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[876] <= mhpmcounter_d[876];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[875] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[875] <= mhpmcounter_d[875];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[874] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[874] <= mhpmcounter_d[874];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[873] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[873] <= mhpmcounter_d[873];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[872] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[872] <= mhpmcounter_d[872];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[871] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[871] <= mhpmcounter_d[871];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[870] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[870] <= mhpmcounter_d[870];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[869] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[869] <= mhpmcounter_d[869];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[868] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[868] <= mhpmcounter_d[868];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[867] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[867] <= mhpmcounter_d[867];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[866] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[866] <= mhpmcounter_d[866];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[865] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[865] <= mhpmcounter_d[865];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[864] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[864] <= mhpmcounter_d[864];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[863] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[863] <= mhpmcounter_d[863];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[862] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[862] <= mhpmcounter_d[862];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[861] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[861] <= mhpmcounter_d[861];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[860] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[860] <= mhpmcounter_d[860];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[859] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[859] <= mhpmcounter_d[859];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[858] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[858] <= mhpmcounter_d[858];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[857] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[857] <= mhpmcounter_d[857];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[856] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[856] <= mhpmcounter_d[856];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[855] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[855] <= mhpmcounter_d[855];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[854] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[854] <= mhpmcounter_d[854];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[853] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[853] <= mhpmcounter_d[853];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[852] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[852] <= mhpmcounter_d[852];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[851] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[851] <= mhpmcounter_d[851];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[850] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[850] <= mhpmcounter_d[850];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[849] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[849] <= mhpmcounter_d[849];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[848] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[848] <= mhpmcounter_d[848];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[847] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[847] <= mhpmcounter_d[847];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[846] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[846] <= mhpmcounter_d[846];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[845] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[845] <= mhpmcounter_d[845];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[844] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[844] <= mhpmcounter_d[844];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[843] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[843] <= mhpmcounter_d[843];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[842] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[842] <= mhpmcounter_d[842];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[841] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[841] <= mhpmcounter_d[841];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[840] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[840] <= mhpmcounter_d[840];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[839] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[839] <= mhpmcounter_d[839];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[838] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[838] <= mhpmcounter_d[838];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[837] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[837] <= mhpmcounter_d[837];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[836] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[836] <= mhpmcounter_d[836];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[835] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[835] <= mhpmcounter_d[835];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[834] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[834] <= mhpmcounter_d[834];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[833] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[833] <= mhpmcounter_d[833];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[832] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[832] <= mhpmcounter_d[832];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[831] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[831] <= mhpmcounter_d[831];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[830] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[830] <= mhpmcounter_d[830];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[829] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[829] <= mhpmcounter_d[829];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[828] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[828] <= mhpmcounter_d[828];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[827] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[827] <= mhpmcounter_d[827];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[826] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[826] <= mhpmcounter_d[826];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[825] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[825] <= mhpmcounter_d[825];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[824] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[824] <= mhpmcounter_d[824];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[823] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[823] <= mhpmcounter_d[823];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[822] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[822] <= mhpmcounter_d[822];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[821] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[821] <= mhpmcounter_d[821];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[820] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[820] <= mhpmcounter_d[820];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[819] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[819] <= mhpmcounter_d[819];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[818] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[818] <= mhpmcounter_d[818];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[817] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[817] <= mhpmcounter_d[817];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[816] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[816] <= mhpmcounter_d[816];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[815] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[815] <= mhpmcounter_d[815];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[814] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[814] <= mhpmcounter_d[814];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[813] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[813] <= mhpmcounter_d[813];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[812] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[812] <= mhpmcounter_d[812];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[811] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[811] <= mhpmcounter_d[811];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[810] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[810] <= mhpmcounter_d[810];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[809] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[809] <= mhpmcounter_d[809];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[808] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[808] <= mhpmcounter_d[808];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[807] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[807] <= mhpmcounter_d[807];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[806] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[806] <= mhpmcounter_d[806];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[805] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[805] <= mhpmcounter_d[805];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[804] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[804] <= mhpmcounter_d[804];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[803] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[803] <= mhpmcounter_d[803];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[802] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[802] <= mhpmcounter_d[802];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[801] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[801] <= mhpmcounter_d[801];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[800] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[800] <= mhpmcounter_d[800];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[799] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[799] <= mhpmcounter_d[799];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[798] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[798] <= mhpmcounter_d[798];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[797] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[797] <= mhpmcounter_d[797];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[796] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[796] <= mhpmcounter_d[796];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[795] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[795] <= mhpmcounter_d[795];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[794] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[794] <= mhpmcounter_d[794];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[793] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[793] <= mhpmcounter_d[793];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[792] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[792] <= mhpmcounter_d[792];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[791] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[791] <= mhpmcounter_d[791];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[790] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[790] <= mhpmcounter_d[790];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[789] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[789] <= mhpmcounter_d[789];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[788] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[788] <= mhpmcounter_d[788];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[787] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[787] <= mhpmcounter_d[787];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[786] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[786] <= mhpmcounter_d[786];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[785] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[785] <= mhpmcounter_d[785];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[784] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[784] <= mhpmcounter_d[784];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[783] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[783] <= mhpmcounter_d[783];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[782] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[782] <= mhpmcounter_d[782];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[781] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[781] <= mhpmcounter_d[781];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[780] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[780] <= mhpmcounter_d[780];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[779] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[779] <= mhpmcounter_d[779];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[778] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[778] <= mhpmcounter_d[778];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[777] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[777] <= mhpmcounter_d[777];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[776] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[776] <= mhpmcounter_d[776];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[775] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[775] <= mhpmcounter_d[775];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[774] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[774] <= mhpmcounter_d[774];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[773] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[773] <= mhpmcounter_d[773];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[772] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[772] <= mhpmcounter_d[772];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[771] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[771] <= mhpmcounter_d[771];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[770] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[770] <= mhpmcounter_d[770];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[769] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[769] <= mhpmcounter_d[769];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[768] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[768] <= mhpmcounter_d[768];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[767] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[767] <= mhpmcounter_d[767];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[766] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[766] <= mhpmcounter_d[766];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[765] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[765] <= mhpmcounter_d[765];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[764] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[764] <= mhpmcounter_d[764];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[763] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[763] <= mhpmcounter_d[763];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[762] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[762] <= mhpmcounter_d[762];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[761] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[761] <= mhpmcounter_d[761];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[760] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[760] <= mhpmcounter_d[760];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[759] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[759] <= mhpmcounter_d[759];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[758] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[758] <= mhpmcounter_d[758];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[757] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[757] <= mhpmcounter_d[757];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[756] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[756] <= mhpmcounter_d[756];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[755] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[755] <= mhpmcounter_d[755];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[754] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[754] <= mhpmcounter_d[754];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[753] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[753] <= mhpmcounter_d[753];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[752] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[752] <= mhpmcounter_d[752];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[751] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[751] <= mhpmcounter_d[751];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[750] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[750] <= mhpmcounter_d[750];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[749] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[749] <= mhpmcounter_d[749];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[748] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[748] <= mhpmcounter_d[748];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[747] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[747] <= mhpmcounter_d[747];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[746] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[746] <= mhpmcounter_d[746];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[745] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[745] <= mhpmcounter_d[745];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[744] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[744] <= mhpmcounter_d[744];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[743] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[743] <= mhpmcounter_d[743];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[742] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[742] <= mhpmcounter_d[742];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[741] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[741] <= mhpmcounter_d[741];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[740] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[740] <= mhpmcounter_d[740];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[739] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[739] <= mhpmcounter_d[739];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[738] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[738] <= mhpmcounter_d[738];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[737] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[737] <= mhpmcounter_d[737];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[736] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[736] <= mhpmcounter_d[736];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[735] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[735] <= mhpmcounter_d[735];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[734] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[734] <= mhpmcounter_d[734];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[733] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[733] <= mhpmcounter_d[733];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[732] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[732] <= mhpmcounter_d[732];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[731] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[731] <= mhpmcounter_d[731];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[730] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[730] <= mhpmcounter_d[730];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[729] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[729] <= mhpmcounter_d[729];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[728] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[728] <= mhpmcounter_d[728];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[727] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[727] <= mhpmcounter_d[727];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[726] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[726] <= mhpmcounter_d[726];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[725] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[725] <= mhpmcounter_d[725];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[724] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[724] <= mhpmcounter_d[724];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[723] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[723] <= mhpmcounter_d[723];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[722] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[722] <= mhpmcounter_d[722];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[721] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[721] <= mhpmcounter_d[721];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[720] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[720] <= mhpmcounter_d[720];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[719] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[719] <= mhpmcounter_d[719];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[718] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[718] <= mhpmcounter_d[718];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[717] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[717] <= mhpmcounter_d[717];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[716] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[716] <= mhpmcounter_d[716];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[715] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[715] <= mhpmcounter_d[715];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[714] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[714] <= mhpmcounter_d[714];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[713] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[713] <= mhpmcounter_d[713];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[712] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[712] <= mhpmcounter_d[712];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[711] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[711] <= mhpmcounter_d[711];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[710] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[710] <= mhpmcounter_d[710];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[709] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[709] <= mhpmcounter_d[709];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[708] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[708] <= mhpmcounter_d[708];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[707] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[707] <= mhpmcounter_d[707];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[706] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[706] <= mhpmcounter_d[706];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[705] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[705] <= mhpmcounter_d[705];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[704] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[704] <= mhpmcounter_d[704];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[703] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[703] <= mhpmcounter_d[703];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[702] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[702] <= mhpmcounter_d[702];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[701] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[701] <= mhpmcounter_d[701];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[700] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[700] <= mhpmcounter_d[700];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[699] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[699] <= mhpmcounter_d[699];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[698] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[698] <= mhpmcounter_d[698];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[697] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[697] <= mhpmcounter_d[697];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[696] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[696] <= mhpmcounter_d[696];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[695] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[695] <= mhpmcounter_d[695];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[694] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[694] <= mhpmcounter_d[694];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[693] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[693] <= mhpmcounter_d[693];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[692] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[692] <= mhpmcounter_d[692];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[691] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[691] <= mhpmcounter_d[691];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[690] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[690] <= mhpmcounter_d[690];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[689] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[689] <= mhpmcounter_d[689];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[688] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[688] <= mhpmcounter_d[688];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[687] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[687] <= mhpmcounter_d[687];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[686] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[686] <= mhpmcounter_d[686];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[685] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[685] <= mhpmcounter_d[685];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[684] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[684] <= mhpmcounter_d[684];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[683] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[683] <= mhpmcounter_d[683];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[682] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[682] <= mhpmcounter_d[682];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[681] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[681] <= mhpmcounter_d[681];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[680] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[680] <= mhpmcounter_d[680];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[679] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[679] <= mhpmcounter_d[679];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[678] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[678] <= mhpmcounter_d[678];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[677] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[677] <= mhpmcounter_d[677];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[676] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[676] <= mhpmcounter_d[676];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[675] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[675] <= mhpmcounter_d[675];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[674] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[674] <= mhpmcounter_d[674];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[673] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[673] <= mhpmcounter_d[673];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[672] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[672] <= mhpmcounter_d[672];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[671] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[671] <= mhpmcounter_d[671];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[670] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[670] <= mhpmcounter_d[670];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[669] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[669] <= mhpmcounter_d[669];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[668] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[668] <= mhpmcounter_d[668];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[667] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[667] <= mhpmcounter_d[667];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[666] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[666] <= mhpmcounter_d[666];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[665] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[665] <= mhpmcounter_d[665];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[664] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[664] <= mhpmcounter_d[664];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[663] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[663] <= mhpmcounter_d[663];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[662] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[662] <= mhpmcounter_d[662];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[661] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[661] <= mhpmcounter_d[661];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[660] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[660] <= mhpmcounter_d[660];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[659] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[659] <= mhpmcounter_d[659];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[658] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[658] <= mhpmcounter_d[658];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[657] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[657] <= mhpmcounter_d[657];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[656] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[656] <= mhpmcounter_d[656];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[655] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[655] <= mhpmcounter_d[655];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[654] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[654] <= mhpmcounter_d[654];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[653] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[653] <= mhpmcounter_d[653];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[652] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[652] <= mhpmcounter_d[652];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[651] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[651] <= mhpmcounter_d[651];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[650] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[650] <= mhpmcounter_d[650];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[649] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[649] <= mhpmcounter_d[649];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[648] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[648] <= mhpmcounter_d[648];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[647] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[647] <= mhpmcounter_d[647];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[646] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[646] <= mhpmcounter_d[646];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[645] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[645] <= mhpmcounter_d[645];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[644] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[644] <= mhpmcounter_d[644];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[643] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[643] <= mhpmcounter_d[643];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[642] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[642] <= mhpmcounter_d[642];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[641] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[641] <= mhpmcounter_d[641];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[640] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[640] <= mhpmcounter_d[640];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[639] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[639] <= mhpmcounter_d[639];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[638] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[638] <= mhpmcounter_d[638];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[637] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[637] <= mhpmcounter_d[637];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[636] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[636] <= mhpmcounter_d[636];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[635] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[635] <= mhpmcounter_d[635];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[634] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[634] <= mhpmcounter_d[634];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[633] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[633] <= mhpmcounter_d[633];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[632] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[632] <= mhpmcounter_d[632];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[631] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[631] <= mhpmcounter_d[631];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[630] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[630] <= mhpmcounter_d[630];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[629] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[629] <= mhpmcounter_d[629];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[628] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[628] <= mhpmcounter_d[628];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[627] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[627] <= mhpmcounter_d[627];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[626] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[626] <= mhpmcounter_d[626];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[625] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[625] <= mhpmcounter_d[625];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[624] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[624] <= mhpmcounter_d[624];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[623] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[623] <= mhpmcounter_d[623];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[622] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[622] <= mhpmcounter_d[622];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[621] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[621] <= mhpmcounter_d[621];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[620] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[620] <= mhpmcounter_d[620];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[619] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[619] <= mhpmcounter_d[619];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[618] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[618] <= mhpmcounter_d[618];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[617] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[617] <= mhpmcounter_d[617];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[616] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[616] <= mhpmcounter_d[616];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[615] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[615] <= mhpmcounter_d[615];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[614] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[614] <= mhpmcounter_d[614];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[613] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[613] <= mhpmcounter_d[613];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[612] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[612] <= mhpmcounter_d[612];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[611] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[611] <= mhpmcounter_d[611];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[610] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[610] <= mhpmcounter_d[610];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[609] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[609] <= mhpmcounter_d[609];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[608] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[608] <= mhpmcounter_d[608];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[607] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[607] <= mhpmcounter_d[607];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[606] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[606] <= mhpmcounter_d[606];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[605] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[605] <= mhpmcounter_d[605];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[604] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[604] <= mhpmcounter_d[604];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[603] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[603] <= mhpmcounter_d[603];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[602] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[602] <= mhpmcounter_d[602];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[601] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[601] <= mhpmcounter_d[601];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[600] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[600] <= mhpmcounter_d[600];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[599] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[599] <= mhpmcounter_d[599];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[598] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[598] <= mhpmcounter_d[598];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[597] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[597] <= mhpmcounter_d[597];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[596] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[596] <= mhpmcounter_d[596];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[595] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[595] <= mhpmcounter_d[595];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[594] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[594] <= mhpmcounter_d[594];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[593] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[593] <= mhpmcounter_d[593];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[592] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[592] <= mhpmcounter_d[592];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[591] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[591] <= mhpmcounter_d[591];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[590] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[590] <= mhpmcounter_d[590];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[589] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[589] <= mhpmcounter_d[589];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[588] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[588] <= mhpmcounter_d[588];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[587] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[587] <= mhpmcounter_d[587];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[586] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[586] <= mhpmcounter_d[586];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[585] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[585] <= mhpmcounter_d[585];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[584] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[584] <= mhpmcounter_d[584];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[583] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[583] <= mhpmcounter_d[583];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[582] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[582] <= mhpmcounter_d[582];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[581] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[581] <= mhpmcounter_d[581];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[580] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[580] <= mhpmcounter_d[580];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[579] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[579] <= mhpmcounter_d[579];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[578] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[578] <= mhpmcounter_d[578];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[577] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[577] <= mhpmcounter_d[577];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[576] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[576] <= mhpmcounter_d[576];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[575] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[575] <= mhpmcounter_d[575];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[574] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[574] <= mhpmcounter_d[574];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[573] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[573] <= mhpmcounter_d[573];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[572] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[572] <= mhpmcounter_d[572];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[571] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[571] <= mhpmcounter_d[571];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[570] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[570] <= mhpmcounter_d[570];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[569] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[569] <= mhpmcounter_d[569];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[568] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[568] <= mhpmcounter_d[568];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[567] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[567] <= mhpmcounter_d[567];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[566] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[566] <= mhpmcounter_d[566];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[565] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[565] <= mhpmcounter_d[565];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[564] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[564] <= mhpmcounter_d[564];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[563] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[563] <= mhpmcounter_d[563];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[562] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[562] <= mhpmcounter_d[562];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[561] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[561] <= mhpmcounter_d[561];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[560] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[560] <= mhpmcounter_d[560];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[559] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[559] <= mhpmcounter_d[559];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[558] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[558] <= mhpmcounter_d[558];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[557] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[557] <= mhpmcounter_d[557];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[556] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[556] <= mhpmcounter_d[556];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[555] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[555] <= mhpmcounter_d[555];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[554] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[554] <= mhpmcounter_d[554];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[553] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[553] <= mhpmcounter_d[553];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[552] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[552] <= mhpmcounter_d[552];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[551] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[551] <= mhpmcounter_d[551];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[550] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[550] <= mhpmcounter_d[550];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[549] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[549] <= mhpmcounter_d[549];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[548] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[548] <= mhpmcounter_d[548];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[547] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[547] <= mhpmcounter_d[547];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[546] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[546] <= mhpmcounter_d[546];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[545] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[545] <= mhpmcounter_d[545];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[544] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[544] <= mhpmcounter_d[544];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[543] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[543] <= mhpmcounter_d[543];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[542] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[542] <= mhpmcounter_d[542];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[541] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[541] <= mhpmcounter_d[541];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[540] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[540] <= mhpmcounter_d[540];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[539] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[539] <= mhpmcounter_d[539];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[538] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[538] <= mhpmcounter_d[538];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[537] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[537] <= mhpmcounter_d[537];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[536] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[536] <= mhpmcounter_d[536];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[535] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[535] <= mhpmcounter_d[535];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[534] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[534] <= mhpmcounter_d[534];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[533] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[533] <= mhpmcounter_d[533];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[532] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[532] <= mhpmcounter_d[532];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[531] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[531] <= mhpmcounter_d[531];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[530] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[530] <= mhpmcounter_d[530];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[529] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[529] <= mhpmcounter_d[529];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[528] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[528] <= mhpmcounter_d[528];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[527] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[527] <= mhpmcounter_d[527];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[526] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[526] <= mhpmcounter_d[526];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[525] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[525] <= mhpmcounter_d[525];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[524] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[524] <= mhpmcounter_d[524];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[523] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[523] <= mhpmcounter_d[523];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[522] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[522] <= mhpmcounter_d[522];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[521] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[521] <= mhpmcounter_d[521];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[520] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[520] <= mhpmcounter_d[520];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[519] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[519] <= mhpmcounter_d[519];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[518] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[518] <= mhpmcounter_d[518];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[517] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[517] <= mhpmcounter_d[517];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[516] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[516] <= mhpmcounter_d[516];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[515] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[515] <= mhpmcounter_d[515];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[514] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[514] <= mhpmcounter_d[514];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[513] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[513] <= mhpmcounter_d[513];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[512] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[512] <= mhpmcounter_d[512];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[511] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[511] <= mhpmcounter_d[511];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[510] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[510] <= mhpmcounter_d[510];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[509] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[509] <= mhpmcounter_d[509];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[508] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[508] <= mhpmcounter_d[508];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[507] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[507] <= mhpmcounter_d[507];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[506] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[506] <= mhpmcounter_d[506];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[505] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[505] <= mhpmcounter_d[505];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[504] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[504] <= mhpmcounter_d[504];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[503] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[503] <= mhpmcounter_d[503];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[502] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[502] <= mhpmcounter_d[502];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[501] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[501] <= mhpmcounter_d[501];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[500] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[500] <= mhpmcounter_d[500];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[499] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[499] <= mhpmcounter_d[499];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[498] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[498] <= mhpmcounter_d[498];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[497] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[497] <= mhpmcounter_d[497];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[496] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[496] <= mhpmcounter_d[496];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[495] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[495] <= mhpmcounter_d[495];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[494] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[494] <= mhpmcounter_d[494];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[493] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[493] <= mhpmcounter_d[493];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[492] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[492] <= mhpmcounter_d[492];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[491] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[491] <= mhpmcounter_d[491];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[490] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[490] <= mhpmcounter_d[490];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[489] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[489] <= mhpmcounter_d[489];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[488] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[488] <= mhpmcounter_d[488];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[487] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[487] <= mhpmcounter_d[487];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[486] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[486] <= mhpmcounter_d[486];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[485] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[485] <= mhpmcounter_d[485];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[484] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[484] <= mhpmcounter_d[484];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[483] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[483] <= mhpmcounter_d[483];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[482] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[482] <= mhpmcounter_d[482];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[481] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[481] <= mhpmcounter_d[481];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[480] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[480] <= mhpmcounter_d[480];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[479] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[479] <= mhpmcounter_d[479];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[478] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[478] <= mhpmcounter_d[478];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[477] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[477] <= mhpmcounter_d[477];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[476] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[476] <= mhpmcounter_d[476];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[475] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[475] <= mhpmcounter_d[475];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[474] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[474] <= mhpmcounter_d[474];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[473] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[473] <= mhpmcounter_d[473];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[472] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[472] <= mhpmcounter_d[472];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[471] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[471] <= mhpmcounter_d[471];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[470] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[470] <= mhpmcounter_d[470];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[469] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[469] <= mhpmcounter_d[469];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[468] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[468] <= mhpmcounter_d[468];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[467] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[467] <= mhpmcounter_d[467];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[466] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[466] <= mhpmcounter_d[466];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[465] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[465] <= mhpmcounter_d[465];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[464] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[464] <= mhpmcounter_d[464];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[463] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[463] <= mhpmcounter_d[463];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[462] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[462] <= mhpmcounter_d[462];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[461] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[461] <= mhpmcounter_d[461];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[460] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[460] <= mhpmcounter_d[460];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[459] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[459] <= mhpmcounter_d[459];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[458] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[458] <= mhpmcounter_d[458];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[457] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[457] <= mhpmcounter_d[457];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[456] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[456] <= mhpmcounter_d[456];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[455] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[455] <= mhpmcounter_d[455];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[454] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[454] <= mhpmcounter_d[454];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[453] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[453] <= mhpmcounter_d[453];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[452] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[452] <= mhpmcounter_d[452];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[451] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[451] <= mhpmcounter_d[451];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[450] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[450] <= mhpmcounter_d[450];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[449] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[449] <= mhpmcounter_d[449];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[448] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[448] <= mhpmcounter_d[448];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[447] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[447] <= mhpmcounter_d[447];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[446] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[446] <= mhpmcounter_d[446];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[445] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[445] <= mhpmcounter_d[445];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[444] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[444] <= mhpmcounter_d[444];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[443] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[443] <= mhpmcounter_d[443];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[442] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[442] <= mhpmcounter_d[442];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[441] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[441] <= mhpmcounter_d[441];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[440] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[440] <= mhpmcounter_d[440];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[439] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[439] <= mhpmcounter_d[439];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[438] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[438] <= mhpmcounter_d[438];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[437] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[437] <= mhpmcounter_d[437];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[436] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[436] <= mhpmcounter_d[436];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[435] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[435] <= mhpmcounter_d[435];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[434] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[434] <= mhpmcounter_d[434];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[433] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[433] <= mhpmcounter_d[433];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[432] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[432] <= mhpmcounter_d[432];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[431] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[431] <= mhpmcounter_d[431];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[430] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[430] <= mhpmcounter_d[430];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[429] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[429] <= mhpmcounter_d[429];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[428] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[428] <= mhpmcounter_d[428];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[427] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[427] <= mhpmcounter_d[427];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[426] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[426] <= mhpmcounter_d[426];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[425] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[425] <= mhpmcounter_d[425];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[424] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[424] <= mhpmcounter_d[424];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[423] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[423] <= mhpmcounter_d[423];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[422] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[422] <= mhpmcounter_d[422];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[421] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[421] <= mhpmcounter_d[421];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[420] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[420] <= mhpmcounter_d[420];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[419] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[419] <= mhpmcounter_d[419];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[418] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[418] <= mhpmcounter_d[418];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[417] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[417] <= mhpmcounter_d[417];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[416] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[416] <= mhpmcounter_d[416];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[415] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[415] <= mhpmcounter_d[415];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[414] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[414] <= mhpmcounter_d[414];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[413] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[413] <= mhpmcounter_d[413];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[412] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[412] <= mhpmcounter_d[412];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[411] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[411] <= mhpmcounter_d[411];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[410] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[410] <= mhpmcounter_d[410];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[409] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[409] <= mhpmcounter_d[409];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[408] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[408] <= mhpmcounter_d[408];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[407] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[407] <= mhpmcounter_d[407];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[406] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[406] <= mhpmcounter_d[406];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[405] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[405] <= mhpmcounter_d[405];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[404] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[404] <= mhpmcounter_d[404];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[403] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[403] <= mhpmcounter_d[403];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[402] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[402] <= mhpmcounter_d[402];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[401] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[401] <= mhpmcounter_d[401];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[400] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[400] <= mhpmcounter_d[400];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[399] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[399] <= mhpmcounter_d[399];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[398] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[398] <= mhpmcounter_d[398];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[397] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[397] <= mhpmcounter_d[397];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[396] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[396] <= mhpmcounter_d[396];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[395] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[395] <= mhpmcounter_d[395];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[394] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[394] <= mhpmcounter_d[394];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[393] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[393] <= mhpmcounter_d[393];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[392] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[392] <= mhpmcounter_d[392];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[391] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[391] <= mhpmcounter_d[391];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[390] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[390] <= mhpmcounter_d[390];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[389] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[389] <= mhpmcounter_d[389];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[388] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[388] <= mhpmcounter_d[388];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[387] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[387] <= mhpmcounter_d[387];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[386] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[386] <= mhpmcounter_d[386];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[385] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[385] <= mhpmcounter_d[385];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[384] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[384] <= mhpmcounter_d[384];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[383] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[383] <= mhpmcounter_d[383];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[382] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[382] <= mhpmcounter_d[382];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[381] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[381] <= mhpmcounter_d[381];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[380] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[380] <= mhpmcounter_d[380];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[379] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[379] <= mhpmcounter_d[379];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[378] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[378] <= mhpmcounter_d[378];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[377] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[377] <= mhpmcounter_d[377];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[376] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[376] <= mhpmcounter_d[376];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[375] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[375] <= mhpmcounter_d[375];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[374] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[374] <= mhpmcounter_d[374];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[373] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[373] <= mhpmcounter_d[373];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[372] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[372] <= mhpmcounter_d[372];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[371] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[371] <= mhpmcounter_d[371];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[370] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[370] <= mhpmcounter_d[370];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[369] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[369] <= mhpmcounter_d[369];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[368] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[368] <= mhpmcounter_d[368];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[367] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[367] <= mhpmcounter_d[367];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[366] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[366] <= mhpmcounter_d[366];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[365] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[365] <= mhpmcounter_d[365];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[364] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[364] <= mhpmcounter_d[364];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[363] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[363] <= mhpmcounter_d[363];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[362] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[362] <= mhpmcounter_d[362];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[361] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[361] <= mhpmcounter_d[361];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[360] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[360] <= mhpmcounter_d[360];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[359] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[359] <= mhpmcounter_d[359];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[358] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[358] <= mhpmcounter_d[358];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[357] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[357] <= mhpmcounter_d[357];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[356] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[356] <= mhpmcounter_d[356];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[355] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[355] <= mhpmcounter_d[355];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[354] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[354] <= mhpmcounter_d[354];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[353] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[353] <= mhpmcounter_d[353];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[352] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[352] <= mhpmcounter_d[352];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[351] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[351] <= mhpmcounter_d[351];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[350] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[350] <= mhpmcounter_d[350];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[349] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[349] <= mhpmcounter_d[349];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[348] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[348] <= mhpmcounter_d[348];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[347] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[347] <= mhpmcounter_d[347];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[346] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[346] <= mhpmcounter_d[346];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[345] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[345] <= mhpmcounter_d[345];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[344] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[344] <= mhpmcounter_d[344];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[343] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[343] <= mhpmcounter_d[343];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[342] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[342] <= mhpmcounter_d[342];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[341] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[341] <= mhpmcounter_d[341];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[340] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[340] <= mhpmcounter_d[340];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[339] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[339] <= mhpmcounter_d[339];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[338] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[338] <= mhpmcounter_d[338];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[337] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[337] <= mhpmcounter_d[337];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[336] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[336] <= mhpmcounter_d[336];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[335] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[335] <= mhpmcounter_d[335];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[334] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[334] <= mhpmcounter_d[334];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[333] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[333] <= mhpmcounter_d[333];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[332] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[332] <= mhpmcounter_d[332];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[331] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[331] <= mhpmcounter_d[331];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[330] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[330] <= mhpmcounter_d[330];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[329] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[329] <= mhpmcounter_d[329];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[328] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[328] <= mhpmcounter_d[328];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[327] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[327] <= mhpmcounter_d[327];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[326] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[326] <= mhpmcounter_d[326];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[325] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[325] <= mhpmcounter_d[325];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[324] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[324] <= mhpmcounter_d[324];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[323] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[323] <= mhpmcounter_d[323];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[322] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[322] <= mhpmcounter_d[322];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[321] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[321] <= mhpmcounter_d[321];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[320] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[320] <= mhpmcounter_d[320];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[319] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[319] <= mhpmcounter_d[319];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[318] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[318] <= mhpmcounter_d[318];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[317] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[317] <= mhpmcounter_d[317];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[316] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[316] <= mhpmcounter_d[316];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[315] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[315] <= mhpmcounter_d[315];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[314] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[314] <= mhpmcounter_d[314];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[313] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[313] <= mhpmcounter_d[313];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[312] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[312] <= mhpmcounter_d[312];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[311] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[311] <= mhpmcounter_d[311];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[310] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[310] <= mhpmcounter_d[310];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[309] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[309] <= mhpmcounter_d[309];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[308] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[308] <= mhpmcounter_d[308];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[307] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[307] <= mhpmcounter_d[307];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[306] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[306] <= mhpmcounter_d[306];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[305] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[305] <= mhpmcounter_d[305];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[304] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[304] <= mhpmcounter_d[304];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[303] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[303] <= mhpmcounter_d[303];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[302] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[302] <= mhpmcounter_d[302];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[301] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[301] <= mhpmcounter_d[301];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[300] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[300] <= mhpmcounter_d[300];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[299] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[299] <= mhpmcounter_d[299];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[298] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[298] <= mhpmcounter_d[298];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[297] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[297] <= mhpmcounter_d[297];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[296] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[296] <= mhpmcounter_d[296];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[295] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[295] <= mhpmcounter_d[295];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[294] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[294] <= mhpmcounter_d[294];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[293] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[293] <= mhpmcounter_d[293];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[292] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[292] <= mhpmcounter_d[292];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[291] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[291] <= mhpmcounter_d[291];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[290] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[290] <= mhpmcounter_d[290];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[289] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[289] <= mhpmcounter_d[289];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[288] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[288] <= mhpmcounter_d[288];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[287] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[287] <= mhpmcounter_d[287];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[286] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[286] <= mhpmcounter_d[286];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[285] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[285] <= mhpmcounter_d[285];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[284] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[284] <= mhpmcounter_d[284];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[283] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[283] <= mhpmcounter_d[283];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[282] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[282] <= mhpmcounter_d[282];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[281] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[281] <= mhpmcounter_d[281];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[280] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[280] <= mhpmcounter_d[280];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[279] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[279] <= mhpmcounter_d[279];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[278] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[278] <= mhpmcounter_d[278];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[277] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[277] <= mhpmcounter_d[277];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[276] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[276] <= mhpmcounter_d[276];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[275] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[275] <= mhpmcounter_d[275];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[274] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[274] <= mhpmcounter_d[274];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[273] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[273] <= mhpmcounter_d[273];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[272] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[272] <= mhpmcounter_d[272];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[271] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[271] <= mhpmcounter_d[271];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[270] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[270] <= mhpmcounter_d[270];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[269] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[269] <= mhpmcounter_d[269];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[268] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[268] <= mhpmcounter_d[268];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[267] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[267] <= mhpmcounter_d[267];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[266] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[266] <= mhpmcounter_d[266];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[265] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[265] <= mhpmcounter_d[265];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[264] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[264] <= mhpmcounter_d[264];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[263] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[263] <= mhpmcounter_d[263];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[262] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[262] <= mhpmcounter_d[262];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[261] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[261] <= mhpmcounter_d[261];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[260] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[260] <= mhpmcounter_d[260];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[259] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[259] <= mhpmcounter_d[259];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[258] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[258] <= mhpmcounter_d[258];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[257] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[257] <= mhpmcounter_d[257];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[256] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[256] <= mhpmcounter_d[256];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[255] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[255] <= mhpmcounter_d[255];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[254] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[254] <= mhpmcounter_d[254];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[253] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[253] <= mhpmcounter_d[253];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[252] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[252] <= mhpmcounter_d[252];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[251] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[251] <= mhpmcounter_d[251];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[250] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[250] <= mhpmcounter_d[250];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[249] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[249] <= mhpmcounter_d[249];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[248] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[248] <= mhpmcounter_d[248];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[247] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[247] <= mhpmcounter_d[247];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[246] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[246] <= mhpmcounter_d[246];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[245] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[245] <= mhpmcounter_d[245];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[244] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[244] <= mhpmcounter_d[244];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[243] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[243] <= mhpmcounter_d[243];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[242] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[242] <= mhpmcounter_d[242];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[241] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[241] <= mhpmcounter_d[241];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[240] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[240] <= mhpmcounter_d[240];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[239] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[239] <= mhpmcounter_d[239];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[238] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[238] <= mhpmcounter_d[238];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[237] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[237] <= mhpmcounter_d[237];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[236] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[236] <= mhpmcounter_d[236];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[235] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[235] <= mhpmcounter_d[235];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[234] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[234] <= mhpmcounter_d[234];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[233] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[233] <= mhpmcounter_d[233];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[232] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[232] <= mhpmcounter_d[232];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[231] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[231] <= mhpmcounter_d[231];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[230] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[230] <= mhpmcounter_d[230];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[229] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[229] <= mhpmcounter_d[229];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[228] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[228] <= mhpmcounter_d[228];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[227] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[227] <= mhpmcounter_d[227];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[226] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[226] <= mhpmcounter_d[226];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[225] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[225] <= mhpmcounter_d[225];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[224] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[224] <= mhpmcounter_d[224];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[223] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[223] <= mhpmcounter_d[223];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[222] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[222] <= mhpmcounter_d[222];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[221] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[221] <= mhpmcounter_d[221];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[220] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[220] <= mhpmcounter_d[220];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[219] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[219] <= mhpmcounter_d[219];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[218] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[218] <= mhpmcounter_d[218];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[217] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[217] <= mhpmcounter_d[217];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[216] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[216] <= mhpmcounter_d[216];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[215] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[215] <= mhpmcounter_d[215];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[214] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[214] <= mhpmcounter_d[214];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[213] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[213] <= mhpmcounter_d[213];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[212] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[212] <= mhpmcounter_d[212];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[211] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[211] <= mhpmcounter_d[211];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[210] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[210] <= mhpmcounter_d[210];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[209] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[209] <= mhpmcounter_d[209];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[208] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[208] <= mhpmcounter_d[208];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[207] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[207] <= mhpmcounter_d[207];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[206] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[206] <= mhpmcounter_d[206];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[205] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[205] <= mhpmcounter_d[205];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[204] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[204] <= mhpmcounter_d[204];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[203] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[203] <= mhpmcounter_d[203];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[202] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[202] <= mhpmcounter_d[202];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[201] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[201] <= mhpmcounter_d[201];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[200] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[200] <= mhpmcounter_d[200];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[199] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[199] <= mhpmcounter_d[199];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[198] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[198] <= mhpmcounter_d[198];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[197] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[197] <= mhpmcounter_d[197];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[196] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[196] <= mhpmcounter_d[196];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[195] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[195] <= mhpmcounter_d[195];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[194] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[194] <= mhpmcounter_d[194];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[193] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[193] <= mhpmcounter_d[193];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[192] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[192] <= mhpmcounter_d[192];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[191] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[191] <= mhpmcounter_d[191];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[190] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[190] <= mhpmcounter_d[190];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[189] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[189] <= mhpmcounter_d[189];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[188] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[188] <= mhpmcounter_d[188];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[187] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[187] <= mhpmcounter_d[187];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[186] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[186] <= mhpmcounter_d[186];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[185] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[185] <= mhpmcounter_d[185];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[184] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[184] <= mhpmcounter_d[184];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[183] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[183] <= mhpmcounter_d[183];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[182] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[182] <= mhpmcounter_d[182];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[181] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[181] <= mhpmcounter_d[181];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[180] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[180] <= mhpmcounter_d[180];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[179] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[179] <= mhpmcounter_d[179];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[178] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[178] <= mhpmcounter_d[178];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[177] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[177] <= mhpmcounter_d[177];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[176] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[176] <= mhpmcounter_d[176];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[175] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[175] <= mhpmcounter_d[175];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[174] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[174] <= mhpmcounter_d[174];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[173] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[173] <= mhpmcounter_d[173];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[172] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[172] <= mhpmcounter_d[172];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[171] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[171] <= mhpmcounter_d[171];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[170] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[170] <= mhpmcounter_d[170];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[169] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[169] <= mhpmcounter_d[169];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[168] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[168] <= mhpmcounter_d[168];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[167] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[167] <= mhpmcounter_d[167];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[166] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[166] <= mhpmcounter_d[166];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[165] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[165] <= mhpmcounter_d[165];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[164] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[164] <= mhpmcounter_d[164];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[163] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[163] <= mhpmcounter_d[163];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[162] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[162] <= mhpmcounter_d[162];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[161] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[161] <= mhpmcounter_d[161];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[160] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[160] <= mhpmcounter_d[160];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[159] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[159] <= mhpmcounter_d[159];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[158] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[158] <= mhpmcounter_d[158];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[157] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[157] <= mhpmcounter_d[157];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[156] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[156] <= mhpmcounter_d[156];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[155] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[155] <= mhpmcounter_d[155];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[154] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[154] <= mhpmcounter_d[154];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[153] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[153] <= mhpmcounter_d[153];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[152] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[152] <= mhpmcounter_d[152];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[151] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[151] <= mhpmcounter_d[151];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[150] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[150] <= mhpmcounter_d[150];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[149] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[149] <= mhpmcounter_d[149];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[148] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[148] <= mhpmcounter_d[148];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[147] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[147] <= mhpmcounter_d[147];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[146] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[146] <= mhpmcounter_d[146];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[145] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[145] <= mhpmcounter_d[145];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[144] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[144] <= mhpmcounter_d[144];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[143] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[143] <= mhpmcounter_d[143];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[142] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[142] <= mhpmcounter_d[142];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[141] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[141] <= mhpmcounter_d[141];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[140] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[140] <= mhpmcounter_d[140];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[139] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[139] <= mhpmcounter_d[139];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[138] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[138] <= mhpmcounter_d[138];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[137] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[137] <= mhpmcounter_d[137];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[136] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[136] <= mhpmcounter_d[136];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[135] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[135] <= mhpmcounter_d[135];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[134] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[134] <= mhpmcounter_d[134];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[133] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[133] <= mhpmcounter_d[133];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[132] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[132] <= mhpmcounter_d[132];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[131] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[131] <= mhpmcounter_d[131];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[130] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[130] <= mhpmcounter_d[130];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[129] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[129] <= mhpmcounter_d[129];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[128] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[128] <= mhpmcounter_d[128];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[127] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[127] <= mhpmcounter_d[127];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[126] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[126] <= mhpmcounter_d[126];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[125] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[125] <= mhpmcounter_d[125];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[124] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[124] <= mhpmcounter_d[124];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[123] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[123] <= mhpmcounter_d[123];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[122] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[122] <= mhpmcounter_d[122];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[121] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[121] <= mhpmcounter_d[121];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[120] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[120] <= mhpmcounter_d[120];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[119] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[119] <= mhpmcounter_d[119];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[118] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[118] <= mhpmcounter_d[118];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[117] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[117] <= mhpmcounter_d[117];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[116] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[116] <= mhpmcounter_d[116];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[115] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[115] <= mhpmcounter_d[115];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[114] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[114] <= mhpmcounter_d[114];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[113] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[113] <= mhpmcounter_d[113];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[112] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[112] <= mhpmcounter_d[112];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[111] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[111] <= mhpmcounter_d[111];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[110] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[110] <= mhpmcounter_d[110];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[109] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[109] <= mhpmcounter_d[109];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[108] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[108] <= mhpmcounter_d[108];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[107] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[107] <= mhpmcounter_d[107];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[106] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[106] <= mhpmcounter_d[106];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[105] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[105] <= mhpmcounter_d[105];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[104] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[104] <= mhpmcounter_d[104];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[103] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[103] <= mhpmcounter_d[103];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[102] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[102] <= mhpmcounter_d[102];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[101] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[101] <= mhpmcounter_d[101];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[100] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[100] <= mhpmcounter_d[100];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[99] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[99] <= mhpmcounter_d[99];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[98] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[98] <= mhpmcounter_d[98];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[97] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[97] <= mhpmcounter_d[97];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[96] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[96] <= mhpmcounter_d[96];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[95] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[95] <= mhpmcounter_d[95];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[94] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[94] <= mhpmcounter_d[94];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[93] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[93] <= mhpmcounter_d[93];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[92] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[92] <= mhpmcounter_d[92];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[91] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[91] <= mhpmcounter_d[91];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[90] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[90] <= mhpmcounter_d[90];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[89] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[89] <= mhpmcounter_d[89];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[88] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[88] <= mhpmcounter_d[88];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[87] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[87] <= mhpmcounter_d[87];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[86] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[86] <= mhpmcounter_d[86];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[85] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[85] <= mhpmcounter_d[85];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[84] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[84] <= mhpmcounter_d[84];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[83] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[83] <= mhpmcounter_d[83];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[82] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[82] <= mhpmcounter_d[82];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[81] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[81] <= mhpmcounter_d[81];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[80] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[80] <= mhpmcounter_d[80];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[79] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[79] <= mhpmcounter_d[79];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[78] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[78] <= mhpmcounter_d[78];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[77] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[77] <= mhpmcounter_d[77];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[76] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[76] <= mhpmcounter_d[76];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[75] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[75] <= mhpmcounter_d[75];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[74] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[74] <= mhpmcounter_d[74];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[73] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[73] <= mhpmcounter_d[73];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[72] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[72] <= mhpmcounter_d[72];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[71] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[71] <= mhpmcounter_d[71];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[70] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[70] <= mhpmcounter_d[70];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[69] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[69] <= mhpmcounter_d[69];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[68] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[68] <= mhpmcounter_d[68];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[67] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[67] <= mhpmcounter_d[67];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[66] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[66] <= mhpmcounter_d[66];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[65] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[65] <= mhpmcounter_d[65];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[64] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[64] <= mhpmcounter_d[64];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[63] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[63] <= mhpmcounter_d[63];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[62] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[62] <= mhpmcounter_d[62];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[61] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[61] <= mhpmcounter_d[61];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[60] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[60] <= mhpmcounter_d[60];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[59] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[59] <= mhpmcounter_d[59];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[58] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[58] <= mhpmcounter_d[58];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[57] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[57] <= mhpmcounter_d[57];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[56] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[56] <= mhpmcounter_d[56];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[55] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[55] <= mhpmcounter_d[55];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[54] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[54] <= mhpmcounter_d[54];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[53] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[53] <= mhpmcounter_d[53];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[52] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[52] <= mhpmcounter_d[52];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[51] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[51] <= mhpmcounter_d[51];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[50] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[50] <= mhpmcounter_d[50];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[49] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[49] <= mhpmcounter_d[49];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[48] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[48] <= mhpmcounter_d[48];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[47] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[47] <= mhpmcounter_d[47];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[46] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[46] <= mhpmcounter_d[46];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[45] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[45] <= mhpmcounter_d[45];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[44] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[44] <= mhpmcounter_d[44];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[43] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[43] <= mhpmcounter_d[43];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[42] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[42] <= mhpmcounter_d[42];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[41] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[41] <= mhpmcounter_d[41];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[40] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[40] <= mhpmcounter_d[40];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[39] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[39] <= mhpmcounter_d[39];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[38] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[38] <= mhpmcounter_d[38];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[37] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[37] <= mhpmcounter_d[37];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[36] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[36] <= mhpmcounter_d[36];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[35] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[35] <= mhpmcounter_d[35];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[34] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[34] <= mhpmcounter_d[34];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[33] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[33] <= mhpmcounter_d[33];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[32] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[32] <= mhpmcounter_d[32];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[31] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[31] <= mhpmcounter_d[31];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[30] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[30] <= mhpmcounter_d[30];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[29] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[29] <= mhpmcounter_d[29];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[28] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[28] <= mhpmcounter_d[28];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[27] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[27] <= mhpmcounter_d[27];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[26] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[26] <= mhpmcounter_d[26];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[25] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[25] <= mhpmcounter_d[25];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[24] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[24] <= mhpmcounter_d[24];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[23] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[23] <= mhpmcounter_d[23];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[22] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[22] <= mhpmcounter_d[22];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[21] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[21] <= mhpmcounter_d[21];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[20] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[20] <= mhpmcounter_d[20];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[19] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[19] <= mhpmcounter_d[19];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[18] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[18] <= mhpmcounter_d[18];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[17] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[17] <= mhpmcounter_d[17];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[16] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[16] <= mhpmcounter_d[16];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[15] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[15] <= mhpmcounter_d[15];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[14] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[14] <= mhpmcounter_d[14];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[13] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[13] <= mhpmcounter_d[13];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[12] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[12] <= mhpmcounter_d[12];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[11] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[11] <= mhpmcounter_d[11];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[10] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[10] <= mhpmcounter_d[10];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[9] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[9] <= mhpmcounter_d[9];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[8] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[8] <= mhpmcounter_d[8];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[7] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[7] <= mhpmcounter_d[7];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[6] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[6] <= mhpmcounter_d[6];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[5] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[5] <= mhpmcounter_d[5];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[4] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[4] <= mhpmcounter_d[4];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[3] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[3] <= mhpmcounter_d[3];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[2] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[2] <= mhpmcounter_d[2];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[1] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[1] <= mhpmcounter_d[1];
    end 
  end


  always @(posedge clk_i or posedge N1238) begin
    if(N1238) begin
      mhpmcounter_q[0] <= 1'b0;
    end else if(1'b1) begin
      mhpmcounter_q[0] <= mhpmcounter_d[0];
    end 
  end

  assign N10617 = csr_addr_i[10] & csr_addr_i[11];
  assign N10618 = csr_addr_i[3] | csr_addr_i[4];
  assign N10619 = csr_addr_i[2] | N10618;
  assign N10620 = csr_addr_i[1] | N10619;
  assign N10621 = csr_addr_i[0] | N10620;
  assign N10622 = ~N10621;
  assign N10623 = ~csr_addr_i[0];
  assign N10624 = N10623 | N10620;
  assign N10625 = ~N10624;
  assign N10626 = ~csr_addr_i[1];
  assign N10627 = N10626 | N10619;
  assign N10628 = csr_addr_i[0] | N10627;
  assign N10629 = ~N10628;
  assign N10630 = ~csr_wdata_int[0];
  assign N10631 = csr_addr_i[7] | N10641;
  assign N10632 = csr_addr_i[6] | N10631;
  assign N10633 = csr_addr_i[5] | N10632;
  assign N10634 = ~N10633;
  assign N10635 = ~csr_addr_i[11];
  assign N10636 = ~csr_addr_i[9];
  assign N10637 = ~csr_addr_i[8];
  assign N10638 = ~csr_addr_i[7];
  assign N10639 = csr_addr_i[10] | N10635;
  assign N10640 = N10636 | N10639;
  assign N10641 = N10637 | N10640;
  assign N10642 = N10638 | N10641;
  assign N10643 = csr_addr_i[6] | N10642;
  assign N10644 = csr_addr_i[5] | N10643;
  assign N10645 = ~N10644;
  assign N10646 = ~csr_addr_i[5];
  assign N10647 = csr_addr_i[10] | csr_addr_i[11];
  assign N10648 = N10636 | N10647;
  assign N10649 = N10637 | N10648;
  assign N10650 = csr_addr_i[7] | N10649;
  assign N10651 = csr_addr_i[6] | N10650;
  assign N10652 = N10646 | N10651;
  assign N10653 = ~N10652;
  assign { N10357, N10356, N10355, N10354, N10353, N10352, N10351, N10350, N10349, N10348, N10347, N10346, N10345, N10344, N10343, N10342, N10341, N10340, N10339, N10338, N10337, N10336, N10335, N10334, N10333, N10332, N10331, N10330, N10329, N10328, N10327, N10326, N10325, N10324, N10323, N10322, N10321, N10320, N10319, N10318, N10317, N10316, N10315, N10314, N10313, N10312, N10311, N10310, N10309, N10308, N10307, N10306, N10305, N10304, N10303, N10302, N10301, N10300, N10299, N10298, N10297, N10296, N10295, N10294 } = mhpmcounter_q[63:0] + 1'b1;
  assign { N10065, N10064, N10063, N10062, N10061, N10060, N10059, N10058, N10057, N10056, N10055, N10054, N10053, N10052, N10051, N10050, N10049, N10048, N10047, N10046, N10045, N10044, N10043, N10042, N10041, N10040, N10039, N10038, N10037, N10036, N10035, N10034, N10033, N10032, N10031, N10030, N10029, N10028, N10027, N10026, N10025, N10024, N10023, N10022, N10021, N10020, N10019, N10018, N10017, N10016, N10015, N10014, N10013, N10012, N10011, N10010, N10009, N10008, N10007, N10006, N10005, N10004, N10003, N10002 } = mhpmcounter_q[127:64] + 1'b1;
  assign { N9773, N9772, N9771, N9770, N9769, N9768, N9767, N9766, N9765, N9764, N9763, N9762, N9761, N9760, N9759, N9758, N9757, N9756, N9755, N9754, N9753, N9752, N9751, N9750, N9749, N9748, N9747, N9746, N9745, N9744, N9743, N9742, N9741, N9740, N9739, N9738, N9737, N9736, N9735, N9734, N9733, N9732, N9731, N9730, N9729, N9728, N9727, N9726, N9725, N9724, N9723, N9722, N9721, N9720, N9719, N9718, N9717, N9716, N9715, N9714, N9713, N9712, N9711, N9710 } = mhpmcounter_q[191:128] + 1'b1;
  assign { N9481, N9480, N9479, N9478, N9477, N9476, N9475, N9474, N9473, N9472, N9471, N9470, N9469, N9468, N9467, N9466, N9465, N9464, N9463, N9462, N9461, N9460, N9459, N9458, N9457, N9456, N9455, N9454, N9453, N9452, N9451, N9450, N9449, N9448, N9447, N9446, N9445, N9444, N9443, N9442, N9441, N9440, N9439, N9438, N9437, N9436, N9435, N9434, N9433, N9432, N9431, N9430, N9429, N9428, N9427, N9426, N9425, N9424, N9423, N9422, N9421, N9420, N9419, N9418 } = mhpmcounter_q[255:192] + 1'b1;
  assign { N9189, N9188, N9187, N9186, N9185, N9184, N9183, N9182, N9181, N9180, N9179, N9178, N9177, N9176, N9175, N9174, N9173, N9172, N9171, N9170, N9169, N9168, N9167, N9166, N9165, N9164, N9163, N9162, N9161, N9160, N9159, N9158, N9157, N9156, N9155, N9154, N9153, N9152, N9151, N9150, N9149, N9148, N9147, N9146, N9145, N9144, N9143, N9142, N9141, N9140, N9139, N9138, N9137, N9136, N9135, N9134, N9133, N9132, N9131, N9130, N9129, N9128, N9127, N9126 } = mhpmcounter_q[319:256] + 1'b1;
  assign { N8897, N8896, N8895, N8894, N8893, N8892, N8891, N8890, N8889, N8888, N8887, N8886, N8885, N8884, N8883, N8882, N8881, N8880, N8879, N8878, N8877, N8876, N8875, N8874, N8873, N8872, N8871, N8870, N8869, N8868, N8867, N8866, N8865, N8864, N8863, N8862, N8861, N8860, N8859, N8858, N8857, N8856, N8855, N8854, N8853, N8852, N8851, N8850, N8849, N8848, N8847, N8846, N8845, N8844, N8843, N8842, N8841, N8840, N8839, N8838, N8837, N8836, N8835, N8834 } = mhpmcounter_q[383:320] + 1'b1;
  assign { N8605, N8604, N8603, N8602, N8601, N8600, N8599, N8598, N8597, N8596, N8595, N8594, N8593, N8592, N8591, N8590, N8589, N8588, N8587, N8586, N8585, N8584, N8583, N8582, N8581, N8580, N8579, N8578, N8577, N8576, N8575, N8574, N8573, N8572, N8571, N8570, N8569, N8568, N8567, N8566, N8565, N8564, N8563, N8562, N8561, N8560, N8559, N8558, N8557, N8556, N8555, N8554, N8553, N8552, N8551, N8550, N8549, N8548, N8547, N8546, N8545, N8544, N8543, N8542 } = mhpmcounter_q[447:384] + 1'b1;
  assign { N8313, N8312, N8311, N8310, N8309, N8308, N8307, N8306, N8305, N8304, N8303, N8302, N8301, N8300, N8299, N8298, N8297, N8296, N8295, N8294, N8293, N8292, N8291, N8290, N8289, N8288, N8287, N8286, N8285, N8284, N8283, N8282, N8281, N8280, N8279, N8278, N8277, N8276, N8275, N8274, N8273, N8272, N8271, N8270, N8269, N8268, N8267, N8266, N8265, N8264, N8263, N8262, N8261, N8260, N8259, N8258, N8257, N8256, N8255, N8254, N8253, N8252, N8251, N8250 } = mhpmcounter_q[511:448] + 1'b1;
  assign { N8021, N8020, N8019, N8018, N8017, N8016, N8015, N8014, N8013, N8012, N8011, N8010, N8009, N8008, N8007, N8006, N8005, N8004, N8003, N8002, N8001, N8000, N7999, N7998, N7997, N7996, N7995, N7994, N7993, N7992, N7991, N7990, N7989, N7988, N7987, N7986, N7985, N7984, N7983, N7982, N7981, N7980, N7979, N7978, N7977, N7976, N7975, N7974, N7973, N7972, N7971, N7970, N7969, N7968, N7967, N7966, N7965, N7964, N7963, N7962, N7961, N7960, N7959, N7958 } = mhpmcounter_q[575:512] + 1'b1;
  assign { N7729, N7728, N7727, N7726, N7725, N7724, N7723, N7722, N7721, N7720, N7719, N7718, N7717, N7716, N7715, N7714, N7713, N7712, N7711, N7710, N7709, N7708, N7707, N7706, N7705, N7704, N7703, N7702, N7701, N7700, N7699, N7698, N7697, N7696, N7695, N7694, N7693, N7692, N7691, N7690, N7689, N7688, N7687, N7686, N7685, N7684, N7683, N7682, N7681, N7680, N7679, N7678, N7677, N7676, N7675, N7674, N7673, N7672, N7671, N7670, N7669, N7668, N7667, N7666 } = mhpmcounter_q[639:576] + 1'b1;
  assign { N7437, N7436, N7435, N7434, N7433, N7432, N7431, N7430, N7429, N7428, N7427, N7426, N7425, N7424, N7423, N7422, N7421, N7420, N7419, N7418, N7417, N7416, N7415, N7414, N7413, N7412, N7411, N7410, N7409, N7408, N7407, N7406, N7405, N7404, N7403, N7402, N7401, N7400, N7399, N7398, N7397, N7396, N7395, N7394, N7393, N7392, N7391, N7390, N7389, N7388, N7387, N7386, N7385, N7384, N7383, N7382, N7381, N7380, N7379, N7378, N7377, N7376, N7375, N7374 } = mhpmcounter_q[703:640] + 1'b1;
  assign { N7145, N7144, N7143, N7142, N7141, N7140, N7139, N7138, N7137, N7136, N7135, N7134, N7133, N7132, N7131, N7130, N7129, N7128, N7127, N7126, N7125, N7124, N7123, N7122, N7121, N7120, N7119, N7118, N7117, N7116, N7115, N7114, N7113, N7112, N7111, N7110, N7109, N7108, N7107, N7106, N7105, N7104, N7103, N7102, N7101, N7100, N7099, N7098, N7097, N7096, N7095, N7094, N7093, N7092, N7091, N7090, N7089, N7088, N7087, N7086, N7085, N7084, N7083, N7082 } = mhpmcounter_q[767:704] + 1'b1;
  assign { N6853, N6852, N6851, N6850, N6849, N6848, N6847, N6846, N6845, N6844, N6843, N6842, N6841, N6840, N6839, N6838, N6837, N6836, N6835, N6834, N6833, N6832, N6831, N6830, N6829, N6828, N6827, N6826, N6825, N6824, N6823, N6822, N6821, N6820, N6819, N6818, N6817, N6816, N6815, N6814, N6813, N6812, N6811, N6810, N6809, N6808, N6807, N6806, N6805, N6804, N6803, N6802, N6801, N6800, N6799, N6798, N6797, N6796, N6795, N6794, N6793, N6792, N6791, N6790 } = mhpmcounter_q[831:768] + 1'b1;
  assign { N6561, N6560, N6559, N6558, N6557, N6556, N6555, N6554, N6553, N6552, N6551, N6550, N6549, N6548, N6547, N6546, N6545, N6544, N6543, N6542, N6541, N6540, N6539, N6538, N6537, N6536, N6535, N6534, N6533, N6532, N6531, N6530, N6529, N6528, N6527, N6526, N6525, N6524, N6523, N6522, N6521, N6520, N6519, N6518, N6517, N6516, N6515, N6514, N6513, N6512, N6511, N6510, N6509, N6508, N6507, N6506, N6505, N6504, N6503, N6502, N6501, N6500, N6499, N6498 } = mhpmcounter_q[895:832] + 1'b1;
  assign { N6269, N6268, N6267, N6266, N6265, N6264, N6263, N6262, N6261, N6260, N6259, N6258, N6257, N6256, N6255, N6254, N6253, N6252, N6251, N6250, N6249, N6248, N6247, N6246, N6245, N6244, N6243, N6242, N6241, N6240, N6239, N6238, N6237, N6236, N6235, N6234, N6233, N6232, N6231, N6230, N6229, N6228, N6227, N6226, N6225, N6224, N6223, N6222, N6221, N6220, N6219, N6218, N6217, N6216, N6215, N6214, N6213, N6212, N6211, N6210, N6209, N6208, N6207, N6206 } = mhpmcounter_q[959:896] + 1'b1;
  assign { N5977, N5976, N5975, N5974, N5973, N5972, N5971, N5970, N5969, N5968, N5967, N5966, N5965, N5964, N5963, N5962, N5961, N5960, N5959, N5958, N5957, N5956, N5955, N5954, N5953, N5952, N5951, N5950, N5949, N5948, N5947, N5946, N5945, N5944, N5943, N5942, N5941, N5940, N5939, N5938, N5937, N5936, N5935, N5934, N5933, N5932, N5931, N5930, N5929, N5928, N5927, N5926, N5925, N5924, N5923, N5922, N5921, N5920, N5919, N5918, N5917, N5916, N5915, N5914 } = mhpmcounter_q[1023:960] + 1'b1;
  assign { N5685, N5684, N5683, N5682, N5681, N5680, N5679, N5678, N5677, N5676, N5675, N5674, N5673, N5672, N5671, N5670, N5669, N5668, N5667, N5666, N5665, N5664, N5663, N5662, N5661, N5660, N5659, N5658, N5657, N5656, N5655, N5654, N5653, N5652, N5651, N5650, N5649, N5648, N5647, N5646, N5645, N5644, N5643, N5642, N5641, N5640, N5639, N5638, N5637, N5636, N5635, N5634, N5633, N5632, N5631, N5630, N5629, N5628, N5627, N5626, N5625, N5624, N5623, N5622 } = mhpmcounter_q[1087:1024] + 1'b1;
  assign { N5393, N5392, N5391, N5390, N5389, N5388, N5387, N5386, N5385, N5384, N5383, N5382, N5381, N5380, N5379, N5378, N5377, N5376, N5375, N5374, N5373, N5372, N5371, N5370, N5369, N5368, N5367, N5366, N5365, N5364, N5363, N5362, N5361, N5360, N5359, N5358, N5357, N5356, N5355, N5354, N5353, N5352, N5351, N5350, N5349, N5348, N5347, N5346, N5345, N5344, N5343, N5342, N5341, N5340, N5339, N5338, N5337, N5336, N5335, N5334, N5333, N5332, N5331, N5330 } = mhpmcounter_q[1151:1088] + 1'b1;
  assign { N5101, N5100, N5099, N5098, N5097, N5096, N5095, N5094, N5093, N5092, N5091, N5090, N5089, N5088, N5087, N5086, N5085, N5084, N5083, N5082, N5081, N5080, N5079, N5078, N5077, N5076, N5075, N5074, N5073, N5072, N5071, N5070, N5069, N5068, N5067, N5066, N5065, N5064, N5063, N5062, N5061, N5060, N5059, N5058, N5057, N5056, N5055, N5054, N5053, N5052, N5051, N5050, N5049, N5048, N5047, N5046, N5045, N5044, N5043, N5042, N5041, N5040, N5039, N5038 } = mhpmcounter_q[1215:1152] + 1'b1;
  assign { N4809, N4808, N4807, N4806, N4805, N4804, N4803, N4802, N4801, N4800, N4799, N4798, N4797, N4796, N4795, N4794, N4793, N4792, N4791, N4790, N4789, N4788, N4787, N4786, N4785, N4784, N4783, N4782, N4781, N4780, N4779, N4778, N4777, N4776, N4775, N4774, N4773, N4772, N4771, N4770, N4769, N4768, N4767, N4766, N4765, N4764, N4763, N4762, N4761, N4760, N4759, N4758, N4757, N4756, N4755, N4754, N4753, N4752, N4751, N4750, N4749, N4748, N4747, N4746 } = mhpmcounter_q[1279:1216] + 1'b1;
  assign { N4517, N4516, N4515, N4514, N4513, N4512, N4511, N4510, N4509, N4508, N4507, N4506, N4505, N4504, N4503, N4502, N4501, N4500, N4499, N4498, N4497, N4496, N4495, N4494, N4493, N4492, N4491, N4490, N4489, N4488, N4487, N4486, N4485, N4484, N4483, N4482, N4481, N4480, N4479, N4478, N4477, N4476, N4475, N4474, N4473, N4472, N4471, N4470, N4469, N4468, N4467, N4466, N4465, N4464, N4463, N4462, N4461, N4460, N4459, N4458, N4457, N4456, N4455, N4454 } = mhpmcounter_q[1343:1280] + 1'b1;
  assign { N4225, N4224, N4223, N4222, N4221, N4220, N4219, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4211, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4203, N4202, N4201, N4200, N4199, N4198, N4197, N4196, N4195, N4194, N4193, N4192, N4191, N4190, N4189, N4188, N4187, N4186, N4185, N4184, N4183, N4182, N4181, N4180, N4179, N4178, N4177, N4176, N4175, N4174, N4173, N4172, N4171, N4170, N4169, N4168, N4167, N4166, N4165, N4164, N4163, N4162 } = mhpmcounter_q[1407:1344] + 1'b1;
  assign { N3933, N3932, N3931, N3930, N3929, N3928, N3927, N3926, N3925, N3924, N3923, N3922, N3921, N3920, N3919, N3918, N3917, N3916, N3915, N3914, N3913, N3912, N3911, N3910, N3909, N3908, N3907, N3906, N3905, N3904, N3903, N3902, N3901, N3900, N3899, N3898, N3897, N3896, N3895, N3894, N3893, N3892, N3891, N3890, N3889, N3888, N3887, N3886, N3885, N3884, N3883, N3882, N3881, N3880, N3879, N3878, N3877, N3876, N3875, N3874, N3873, N3872, N3871, N3870 } = mhpmcounter_q[1471:1408] + 1'b1;
  assign { N3641, N3640, N3639, N3638, N3637, N3636, N3635, N3634, N3633, N3632, N3631, N3630, N3629, N3628, N3627, N3626, N3625, N3624, N3623, N3622, N3621, N3620, N3619, N3618, N3617, N3616, N3615, N3614, N3613, N3612, N3611, N3610, N3609, N3608, N3607, N3606, N3605, N3604, N3603, N3602, N3601, N3600, N3599, N3598, N3597, N3596, N3595, N3594, N3593, N3592, N3591, N3590, N3589, N3588, N3587, N3586, N3585, N3584, N3583, N3582, N3581, N3580, N3579, N3578 } = mhpmcounter_q[1535:1472] + 1'b1;
  assign { N3349, N3348, N3347, N3346, N3345, N3344, N3343, N3342, N3341, N3340, N3339, N3338, N3337, N3336, N3335, N3334, N3333, N3332, N3331, N3330, N3329, N3328, N3327, N3326, N3325, N3324, N3323, N3322, N3321, N3320, N3319, N3318, N3317, N3316, N3315, N3314, N3313, N3312, N3311, N3310, N3309, N3308, N3307, N3306, N3305, N3304, N3303, N3302, N3301, N3300, N3299, N3298, N3297, N3296, N3295, N3294, N3293, N3292, N3291, N3290, N3289, N3288, N3287, N3286 } = mhpmcounter_q[1599:1536] + 1'b1;
  assign { N3057, N3056, N3055, N3054, N3053, N3052, N3051, N3050, N3049, N3048, N3047, N3046, N3045, N3044, N3043, N3042, N3041, N3040, N3039, N3038, N3037, N3036, N3035, N3034, N3033, N3032, N3031, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N3023, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N3015, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N3007, N3006, N3005, N3004, N3003, N3002, N3001, N3000, N2999, N2998, N2997, N2996, N2995, N2994 } = mhpmcounter_q[1663:1600] + 1'b1;
  assign { N2765, N2764, N2763, N2762, N2761, N2760, N2759, N2758, N2757, N2756, N2755, N2754, N2753, N2752, N2751, N2750, N2749, N2748, N2747, N2746, N2745, N2744, N2743, N2742, N2741, N2740, N2739, N2738, N2737, N2736, N2735, N2734, N2733, N2732, N2731, N2730, N2729, N2728, N2727, N2726, N2725, N2724, N2723, N2722, N2721, N2720, N2719, N2718, N2717, N2716, N2715, N2714, N2713, N2712, N2711, N2710, N2709, N2708, N2707, N2706, N2705, N2704, N2703, N2702 } = mhpmcounter_q[1727:1664] + 1'b1;
  assign { N2473, N2472, N2471, N2470, N2469, N2468, N2467, N2466, N2465, N2464, N2463, N2462, N2461, N2460, N2459, N2458, N2457, N2456, N2455, N2454, N2453, N2452, N2451, N2450, N2449, N2448, N2447, N2446, N2445, N2444, N2443, N2442, N2441, N2440, N2439, N2438, N2437, N2436, N2435, N2434, N2433, N2432, N2431, N2430, N2429, N2428, N2427, N2426, N2425, N2424, N2423, N2422, N2421, N2420, N2419, N2418, N2417, N2416, N2415, N2414, N2413, N2412, N2411, N2410 } = mhpmcounter_q[1791:1728] + 1'b1;
  assign { N2181, N2180, N2179, N2178, N2177, N2176, N2175, N2174, N2173, N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, N2158, N2157, N2156, N2155, N2154, N2153, N2152, N2151, N2150, N2149, N2148, N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140, N2139, N2138, N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, N2123, N2122, N2121, N2120, N2119, N2118 } = mhpmcounter_q[1855:1792] + 1'b1;
  assign { N1889, N1888, N1887, N1886, N1885, N1884, N1883, N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862, N1861, N1860, N1859, N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835, N1834, N1833, N1832, N1831, N1830, N1829, N1828, N1827, N1826 } = mhpmcounter_q[1919:1856] + 1'b1;
  assign { N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534 } = mhpmcounter_q[1983:1920] + 1'b1;
  assign { N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242 } = mhpmcounter_q[2047:1984] + 1'b1;
  assign N10654 = csr_addr_i[3] & csr_addr_i[4];
  assign N10655 = N0 & csr_addr_i[4];
  assign N0 = ~csr_addr_i[3];
  assign N10656 = csr_addr_i[3] & N1;
  assign N1 = ~csr_addr_i[4];
  assign N10657 = N2 & N3;
  assign N2 = ~csr_addr_i[3];
  assign N3 = ~csr_addr_i[4];
  assign N10658 = ~csr_addr_i[2];
  assign N10659 = csr_addr_i[0] & csr_addr_i[1];
  assign N10660 = N4 & csr_addr_i[1];
  assign N4 = ~csr_addr_i[0];
  assign N10661 = csr_addr_i[0] & N5;
  assign N5 = ~csr_addr_i[1];
  assign N10662 = N6 & N7;
  assign N6 = ~csr_addr_i[0];
  assign N7 = ~csr_addr_i[1];
  assign N10663 = csr_addr_i[2] & N10659;
  assign N10664 = csr_addr_i[2] & N10660;
  assign N10665 = csr_addr_i[2] & N10661;
  assign N10666 = csr_addr_i[2] & N10662;
  assign N10667 = N10658 & N10659;
  assign N10668 = N10658 & N10660;
  assign N10669 = N10658 & N10661;
  assign N10670 = N10658 & N10662;
  assign N753 = N10654 & N10663;
  assign N752 = N10654 & N10664;
  assign N751 = N10654 & N10665;
  assign N750 = N10654 & N10666;
  assign N749 = N10654 & N10667;
  assign N748 = N10654 & N10668;
  assign N747 = N10654 & N10669;
  assign N746 = N10654 & N10670;
  assign N745 = N10655 & N10663;
  assign N744 = N10655 & N10664;
  assign N743 = N10655 & N10665;
  assign N742 = N10655 & N10666;
  assign N741 = N10655 & N10667;
  assign N740 = N10655 & N10668;
  assign N739 = N10655 & N10669;
  assign N738 = N10655 & N10670;
  assign N737 = N10656 & N10663;
  assign N736 = N10656 & N10664;
  assign N735 = N10656 & N10665;
  assign N734 = N10656 & N10666;
  assign N733 = N10656 & N10667;
  assign N732 = N10656 & N10668;
  assign N731 = N10656 & N10669;
  assign N730 = N10656 & N10670;
  assign N729 = N10657 & N10663;
  assign N728 = N10657 & N10664;
  assign N727 = N10657 & N10665;
  assign N726 = N10657 & N10666;
  assign N725 = N10657 & N10667;
  assign N724 = N10657 & N10668;
  assign N723 = N10657 & N10669;
  assign N722 = N10657 & N10670;
  assign N373 = (N8)? csr_access_i : 
                (N372)? 1'b0 : 1'b0;
  assign N8 = N371;
  assign { N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374 } = (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N369, 1'b0, N370 } : 
                                                                                                                                                                                                              (N10)? { N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269 } : 
                                                                                                                                                                                                              (N11)? { N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237 } : 
                                                                                                                                                                                                              (N303)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N9 = N10653;
  assign N10 = N10634;
  assign N11 = N10645;
  assign N406 = (N9)? N373 : 
                (N10)? N373 : 
                (N11)? N373 : 
                (N303)? csr_access_i : 1'b0;
  assign csr_rdata_o = (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, cluster_id_i, 1'b0, core_id_i } : 
                       (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mstatus_q_mpp__1_, mstatus_q_mpp__0_, 1'b0, 1'b0, 1'b0, mstatus_q_mpie_, 1'b0, 1'b0, 1'b0, m_irq_enable_o, 1'b0, 1'b0, 1'b0 } : 
                       (N14)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                       (N15)? mscratch_q : 
                       (N16)? csr_mtvec_i : 
                       (N17)? csr_mepc_o : 
                       (N18)? { mcause_q[5:5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mcause_q[4:0] } : 
                       (N19)? mtval_q : 
                       (N20)? { dcsr_q_xdebugver__3_, dcsr_q_xdebugver__2_, dcsr_q_xdebugver__1_, dcsr_q_xdebugver__0_, dcsr_q_zero2__11_, dcsr_q_zero2__10_, dcsr_q_zero2__9_, dcsr_q_zero2__8_, dcsr_q_zero2__7_, dcsr_q_zero2__6_, dcsr_q_zero2__5_, dcsr_q_zero2__4_, dcsr_q_zero2__3_, dcsr_q_zero2__2_, dcsr_q_zero2__1_, dcsr_q_zero2__0_, debug_ebreakm_o, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__2_, dcsr_q_cause__1_, dcsr_q_cause__0_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, debug_single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                       (N21)? csr_depc_o : 
                       (N22)? dscratch0_q : 
                       (N23)? dscratch1_q : 
                       (N24)? mcountinhibit : 
                       (N25)? mhpmcounter_q[2015:1984] : 
                       (N26)? mhpmcounter_q[2047:2016] : 
                       (N27)? mhpmcounter_q[1887:1856] : 
                       (N28)? mhpmcounter_q[1919:1888] : 
                       (N300)? { N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374 } : 1'b0;
  assign N12 = N277;
  assign N13 = N409;
  assign N14 = N279;
  assign N15 = N411;
  assign N16 = N283;
  assign N17 = N413;
  assign N18 = N415;
  assign N19 = N421;
  assign N20 = N423;
  assign N21 = N427;
  assign N22 = N429;
  assign N23 = N440;
  assign N24 = N447;
  assign N25 = N449;
  assign N26 = N453;
  assign N27 = N458;
  assign N28 = N470;
  assign illegal_csr = (N12)? 1'b0 : 
                       (N13)? 1'b0 : 
                       (N14)? 1'b0 : 
                       (N15)? 1'b0 : 
                       (N16)? 1'b0 : 
                       (N17)? 1'b0 : 
                       (N18)? 1'b0 : 
                       (N19)? 1'b0 : 
                       (N20)? 1'b0 : 
                       (N21)? 1'b0 : 
                       (N22)? 1'b0 : 
                       (N23)? 1'b0 : 
                       (N24)? 1'b0 : 
                       (N25)? 1'b0 : 
                       (N26)? 1'b0 : 
                       (N27)? 1'b0 : 
                       (N28)? 1'b0 : 
                       (N300)? N406 : 1'b0;
  assign { N487, N486 } = (N29)? { csr_wdata_int[3:3], csr_wdata_int[7:7] } : 
                          (N30)? { m_irq_enable_o, mstatus_q_mpie_ } : 1'b0;
  assign N29 = csr_we_int;
  assign N30 = N485;
  assign { N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488 } = (N29)? csr_wdata_int : 
                                                                                                                                                                                                              (N30)? mscratch_q : 1'b0;
  assign { N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520 } = (N29)? { csr_wdata_int[31:1], 1'b0 } : 
                                                                                                                                                                                                              (N30)? csr_mepc_o : 1'b0;
  assign { N557, N556, N555, N554, N553, N552 } = (N29)? { csr_wdata_int[31:31], csr_wdata_int[4:0] } : 
                                                  (N30)? mcause_q : 1'b0;
  assign { N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558 } = (N29)? csr_wdata_int : 
                                                                                                                                                                                                              (N30)? mtval_q : 1'b0;
  assign { N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590 } = (N29)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, csr_wdata_int[15:15], 1'b0, csr_wdata_int[13:11], 1'b0, 1'b0, csr_wdata_int[8:6], 1'b0, 1'b0, 1'b0, csr_wdata_int[2:2], 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N30)? { dcsr_q_xdebugver__3_, dcsr_q_xdebugver__2_, dcsr_q_xdebugver__1_, dcsr_q_xdebugver__0_, dcsr_q_zero2__11_, dcsr_q_zero2__10_, dcsr_q_zero2__9_, dcsr_q_zero2__8_, dcsr_q_zero2__7_, dcsr_q_zero2__6_, dcsr_q_zero2__5_, dcsr_q_zero2__4_, dcsr_q_zero2__3_, dcsr_q_zero2__2_, dcsr_q_zero2__1_, dcsr_q_zero2__0_, debug_ebreakm_o, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__2_, dcsr_q_cause__1_, dcsr_q_cause__0_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, debug_single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 1'b0;
  assign { N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624 } = (N31)? csr_wdata_int : 
                                                                                                                                                                                                              (N623)? csr_depc_o : 1'b0;
  assign N31 = N622;
  assign { N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656 } = (N29)? csr_wdata_int : 
                                                                                                                                                                                                              (N30)? dscratch0_q : 1'b0;
  assign { N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688 } = (N29)? csr_wdata_int : 
                                                                                                                                                                                                              (N30)? dscratch1_q : 1'b0;
  assign { N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754 } = (N10)? { N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722 } : 
                                                                                                                                                                                                              (N32)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                              (N33)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N32 = N10633;
  assign N33 = 1'b0;
  assign { N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786 } = (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                              (N11)? { N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722 } : 
                                                                                                                                                                                                              (N721)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818 } = (N29)? { N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786 } : 
                                                                                                                                                                                                              (N30)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850 } = (N29)? { N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754 } : 
                                                                                                                                                                                                              (N30)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N883, N882 } = (N13)? { N487, N486 } : 
                          (N15)? { m_irq_enable_o, mstatus_q_mpie_ } : 
                          (N17)? { m_irq_enable_o, mstatus_q_mpie_ } : 
                          (N18)? { m_irq_enable_o, mstatus_q_mpie_ } : 
                          (N19)? { m_irq_enable_o, mstatus_q_mpie_ } : 
                          (N20)? { m_irq_enable_o, mstatus_q_mpie_ } : 
                          (N21)? { m_irq_enable_o, mstatus_q_mpie_ } : 
                          (N22)? { m_irq_enable_o, mstatus_q_mpie_ } : 
                          (N23)? { m_irq_enable_o, mstatus_q_mpie_ } : 
                          (N24)? { m_irq_enable_o, mstatus_q_mpie_ } : 
                          (N25)? { m_irq_enable_o, mstatus_q_mpie_ } : 
                          (N26)? { m_irq_enable_o, mstatus_q_mpie_ } : 
                          (N27)? { m_irq_enable_o, mstatus_q_mpie_ } : 
                          (N28)? { m_irq_enable_o, mstatus_q_mpie_ } : 
                          (N484)? { m_irq_enable_o, mstatus_q_mpie_ } : 1'b0;
  assign mscratch_d = (N15)? { N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488 } : 
                      (N484)? mscratch_q : 1'b0;
  assign { N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884 } = (N13)? csr_mepc_o : 
                                                                                                                                                                                                              (N15)? csr_mepc_o : 
                                                                                                                                                                                                              (N17)? { N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520 } : 
                                                                                                                                                                                                              (N18)? csr_mepc_o : 
                                                                                                                                                                                                              (N19)? csr_mepc_o : 
                                                                                                                                                                                                              (N20)? csr_mepc_o : 
                                                                                                                                                                                                              (N21)? csr_mepc_o : 
                                                                                                                                                                                                              (N22)? csr_mepc_o : 
                                                                                                                                                                                                              (N23)? csr_mepc_o : 
                                                                                                                                                                                                              (N24)? csr_mepc_o : 
                                                                                                                                                                                                              (N25)? csr_mepc_o : 
                                                                                                                                                                                                              (N26)? csr_mepc_o : 
                                                                                                                                                                                                              (N27)? csr_mepc_o : 
                                                                                                                                                                                                              (N28)? csr_mepc_o : 
                                                                                                                                                                                                              (N484)? csr_mepc_o : 1'b0;
  assign { N921, N920, N919, N918, N917, N916 } = (N13)? mcause_q : 
                                                  (N15)? mcause_q : 
                                                  (N17)? mcause_q : 
                                                  (N18)? { N557, N556, N555, N554, N553, N552 } : 
                                                  (N19)? mcause_q : 
                                                  (N20)? mcause_q : 
                                                  (N21)? mcause_q : 
                                                  (N22)? mcause_q : 
                                                  (N23)? mcause_q : 
                                                  (N24)? mcause_q : 
                                                  (N25)? mcause_q : 
                                                  (N26)? mcause_q : 
                                                  (N27)? mcause_q : 
                                                  (N28)? mcause_q : 
                                                  (N484)? mcause_q : 1'b0;
  assign { N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922 } = (N13)? mtval_q : 
                                                                                                                                                                                                              (N15)? mtval_q : 
                                                                                                                                                                                                              (N17)? mtval_q : 
                                                                                                                                                                                                              (N18)? mtval_q : 
                                                                                                                                                                                                              (N19)? { N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558 } : 
                                                                                                                                                                                                              (N20)? mtval_q : 
                                                                                                                                                                                                              (N21)? mtval_q : 
                                                                                                                                                                                                              (N22)? mtval_q : 
                                                                                                                                                                                                              (N23)? mtval_q : 
                                                                                                                                                                                                              (N24)? mtval_q : 
                                                                                                                                                                                                              (N25)? mtval_q : 
                                                                                                                                                                                                              (N26)? mtval_q : 
                                                                                                                                                                                                              (N27)? mtval_q : 
                                                                                                                                                                                                              (N28)? mtval_q : 
                                                                                                                                                                                                              (N484)? mtval_q : 1'b0;
  assign { N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954 } = (N13)? { dcsr_q_xdebugver__3_, dcsr_q_xdebugver__2_, dcsr_q_xdebugver__1_, dcsr_q_xdebugver__0_, dcsr_q_zero2__11_, dcsr_q_zero2__10_, dcsr_q_zero2__9_, dcsr_q_zero2__8_, dcsr_q_zero2__7_, dcsr_q_zero2__6_, dcsr_q_zero2__5_, dcsr_q_zero2__4_, dcsr_q_zero2__3_, dcsr_q_zero2__2_, dcsr_q_zero2__1_, dcsr_q_zero2__0_, debug_ebreakm_o, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__2_, dcsr_q_cause__1_, dcsr_q_cause__0_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, debug_single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                              (N15)? { dcsr_q_xdebugver__3_, dcsr_q_xdebugver__2_, dcsr_q_xdebugver__1_, dcsr_q_xdebugver__0_, dcsr_q_zero2__11_, dcsr_q_zero2__10_, dcsr_q_zero2__9_, dcsr_q_zero2__8_, dcsr_q_zero2__7_, dcsr_q_zero2__6_, dcsr_q_zero2__5_, dcsr_q_zero2__4_, dcsr_q_zero2__3_, dcsr_q_zero2__2_, dcsr_q_zero2__1_, dcsr_q_zero2__0_, debug_ebreakm_o, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__2_, dcsr_q_cause__1_, dcsr_q_cause__0_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, debug_single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                              (N17)? { dcsr_q_xdebugver__3_, dcsr_q_xdebugver__2_, dcsr_q_xdebugver__1_, dcsr_q_xdebugver__0_, dcsr_q_zero2__11_, dcsr_q_zero2__10_, dcsr_q_zero2__9_, dcsr_q_zero2__8_, dcsr_q_zero2__7_, dcsr_q_zero2__6_, dcsr_q_zero2__5_, dcsr_q_zero2__4_, dcsr_q_zero2__3_, dcsr_q_zero2__2_, dcsr_q_zero2__1_, dcsr_q_zero2__0_, debug_ebreakm_o, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__2_, dcsr_q_cause__1_, dcsr_q_cause__0_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, debug_single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                              (N18)? { dcsr_q_xdebugver__3_, dcsr_q_xdebugver__2_, dcsr_q_xdebugver__1_, dcsr_q_xdebugver__0_, dcsr_q_zero2__11_, dcsr_q_zero2__10_, dcsr_q_zero2__9_, dcsr_q_zero2__8_, dcsr_q_zero2__7_, dcsr_q_zero2__6_, dcsr_q_zero2__5_, dcsr_q_zero2__4_, dcsr_q_zero2__3_, dcsr_q_zero2__2_, dcsr_q_zero2__1_, dcsr_q_zero2__0_, debug_ebreakm_o, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__2_, dcsr_q_cause__1_, dcsr_q_cause__0_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, debug_single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                              (N19)? { dcsr_q_xdebugver__3_, dcsr_q_xdebugver__2_, dcsr_q_xdebugver__1_, dcsr_q_xdebugver__0_, dcsr_q_zero2__11_, dcsr_q_zero2__10_, dcsr_q_zero2__9_, dcsr_q_zero2__8_, dcsr_q_zero2__7_, dcsr_q_zero2__6_, dcsr_q_zero2__5_, dcsr_q_zero2__4_, dcsr_q_zero2__3_, dcsr_q_zero2__2_, dcsr_q_zero2__1_, dcsr_q_zero2__0_, debug_ebreakm_o, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__2_, dcsr_q_cause__1_, dcsr_q_cause__0_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, debug_single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                              (N20)? { N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590 } : 
                                                                                                                                                                                                              (N21)? { dcsr_q_xdebugver__3_, dcsr_q_xdebugver__2_, dcsr_q_xdebugver__1_, dcsr_q_xdebugver__0_, dcsr_q_zero2__11_, dcsr_q_zero2__10_, dcsr_q_zero2__9_, dcsr_q_zero2__8_, dcsr_q_zero2__7_, dcsr_q_zero2__6_, dcsr_q_zero2__5_, dcsr_q_zero2__4_, dcsr_q_zero2__3_, dcsr_q_zero2__2_, dcsr_q_zero2__1_, dcsr_q_zero2__0_, debug_ebreakm_o, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__2_, dcsr_q_cause__1_, dcsr_q_cause__0_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, debug_single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                              (N22)? { dcsr_q_xdebugver__3_, dcsr_q_xdebugver__2_, dcsr_q_xdebugver__1_, dcsr_q_xdebugver__0_, dcsr_q_zero2__11_, dcsr_q_zero2__10_, dcsr_q_zero2__9_, dcsr_q_zero2__8_, dcsr_q_zero2__7_, dcsr_q_zero2__6_, dcsr_q_zero2__5_, dcsr_q_zero2__4_, dcsr_q_zero2__3_, dcsr_q_zero2__2_, dcsr_q_zero2__1_, dcsr_q_zero2__0_, debug_ebreakm_o, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__2_, dcsr_q_cause__1_, dcsr_q_cause__0_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, debug_single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                              (N23)? { dcsr_q_xdebugver__3_, dcsr_q_xdebugver__2_, dcsr_q_xdebugver__1_, dcsr_q_xdebugver__0_, dcsr_q_zero2__11_, dcsr_q_zero2__10_, dcsr_q_zero2__9_, dcsr_q_zero2__8_, dcsr_q_zero2__7_, dcsr_q_zero2__6_, dcsr_q_zero2__5_, dcsr_q_zero2__4_, dcsr_q_zero2__3_, dcsr_q_zero2__2_, dcsr_q_zero2__1_, dcsr_q_zero2__0_, debug_ebreakm_o, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__2_, dcsr_q_cause__1_, dcsr_q_cause__0_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, debug_single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                              (N24)? { dcsr_q_xdebugver__3_, dcsr_q_xdebugver__2_, dcsr_q_xdebugver__1_, dcsr_q_xdebugver__0_, dcsr_q_zero2__11_, dcsr_q_zero2__10_, dcsr_q_zero2__9_, dcsr_q_zero2__8_, dcsr_q_zero2__7_, dcsr_q_zero2__6_, dcsr_q_zero2__5_, dcsr_q_zero2__4_, dcsr_q_zero2__3_, dcsr_q_zero2__2_, dcsr_q_zero2__1_, dcsr_q_zero2__0_, debug_ebreakm_o, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__2_, dcsr_q_cause__1_, dcsr_q_cause__0_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, debug_single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                              (N25)? { dcsr_q_xdebugver__3_, dcsr_q_xdebugver__2_, dcsr_q_xdebugver__1_, dcsr_q_xdebugver__0_, dcsr_q_zero2__11_, dcsr_q_zero2__10_, dcsr_q_zero2__9_, dcsr_q_zero2__8_, dcsr_q_zero2__7_, dcsr_q_zero2__6_, dcsr_q_zero2__5_, dcsr_q_zero2__4_, dcsr_q_zero2__3_, dcsr_q_zero2__2_, dcsr_q_zero2__1_, dcsr_q_zero2__0_, debug_ebreakm_o, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__2_, dcsr_q_cause__1_, dcsr_q_cause__0_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, debug_single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                              (N26)? { dcsr_q_xdebugver__3_, dcsr_q_xdebugver__2_, dcsr_q_xdebugver__1_, dcsr_q_xdebugver__0_, dcsr_q_zero2__11_, dcsr_q_zero2__10_, dcsr_q_zero2__9_, dcsr_q_zero2__8_, dcsr_q_zero2__7_, dcsr_q_zero2__6_, dcsr_q_zero2__5_, dcsr_q_zero2__4_, dcsr_q_zero2__3_, dcsr_q_zero2__2_, dcsr_q_zero2__1_, dcsr_q_zero2__0_, debug_ebreakm_o, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__2_, dcsr_q_cause__1_, dcsr_q_cause__0_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, debug_single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                              (N27)? { dcsr_q_xdebugver__3_, dcsr_q_xdebugver__2_, dcsr_q_xdebugver__1_, dcsr_q_xdebugver__0_, dcsr_q_zero2__11_, dcsr_q_zero2__10_, dcsr_q_zero2__9_, dcsr_q_zero2__8_, dcsr_q_zero2__7_, dcsr_q_zero2__6_, dcsr_q_zero2__5_, dcsr_q_zero2__4_, dcsr_q_zero2__3_, dcsr_q_zero2__2_, dcsr_q_zero2__1_, dcsr_q_zero2__0_, debug_ebreakm_o, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__2_, dcsr_q_cause__1_, dcsr_q_cause__0_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, debug_single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                              (N28)? { dcsr_q_xdebugver__3_, dcsr_q_xdebugver__2_, dcsr_q_xdebugver__1_, dcsr_q_xdebugver__0_, dcsr_q_zero2__11_, dcsr_q_zero2__10_, dcsr_q_zero2__9_, dcsr_q_zero2__8_, dcsr_q_zero2__7_, dcsr_q_zero2__6_, dcsr_q_zero2__5_, dcsr_q_zero2__4_, dcsr_q_zero2__3_, dcsr_q_zero2__2_, dcsr_q_zero2__1_, dcsr_q_zero2__0_, debug_ebreakm_o, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__2_, dcsr_q_cause__1_, dcsr_q_cause__0_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, debug_single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 
                                                                                                                                                                                                              (N484)? { dcsr_q_xdebugver__3_, dcsr_q_xdebugver__2_, dcsr_q_xdebugver__1_, dcsr_q_xdebugver__0_, dcsr_q_zero2__11_, dcsr_q_zero2__10_, dcsr_q_zero2__9_, dcsr_q_zero2__8_, dcsr_q_zero2__7_, dcsr_q_zero2__6_, dcsr_q_zero2__5_, dcsr_q_zero2__4_, dcsr_q_zero2__3_, dcsr_q_zero2__2_, dcsr_q_zero2__1_, dcsr_q_zero2__0_, debug_ebreakm_o, dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_ebreaku_, dcsr_q_stepie_, dcsr_q_stopcount_, dcsr_q_stoptime_, dcsr_q_cause__2_, dcsr_q_cause__1_, dcsr_q_cause__0_, dcsr_q_zero0_, dcsr_q_mprven_, dcsr_q_nmip_, debug_single_step_o, dcsr_q_prv__1_, dcsr_q_prv__0_ } : 1'b0;
  assign { N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986 } = (N13)? csr_depc_o : 
                                                                                                                                                                                                                                (N15)? csr_depc_o : 
                                                                                                                                                                                                                                (N17)? csr_depc_o : 
                                                                                                                                                                                                                                (N18)? csr_depc_o : 
                                                                                                                                                                                                                                (N19)? csr_depc_o : 
                                                                                                                                                                                                                                (N20)? csr_depc_o : 
                                                                                                                                                                                                                                (N21)? { N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624 } : 
                                                                                                                                                                                                                                (N22)? csr_depc_o : 
                                                                                                                                                                                                                                (N23)? csr_depc_o : 
                                                                                                                                                                                                                                (N24)? csr_depc_o : 
                                                                                                                                                                                                                                (N25)? csr_depc_o : 
                                                                                                                                                                                                                                (N26)? csr_depc_o : 
                                                                                                                                                                                                                                (N27)? csr_depc_o : 
                                                                                                                                                                                                                                (N28)? csr_depc_o : 
                                                                                                                                                                                                                                (N484)? csr_depc_o : 1'b0;
  assign dscratch0_d = (N22)? { N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656 } : 
                       (N484)? dscratch0_q : 1'b0;
  assign dscratch1_d = (N23)? { N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688 } : 
                       (N484)? dscratch1_q : 1'b0;
  assign mcountinhibit_we = (N13)? 1'b0 : 
                            (N15)? 1'b0 : 
                            (N17)? 1'b0 : 
                            (N18)? 1'b0 : 
                            (N19)? 1'b0 : 
                            (N20)? 1'b0 : 
                            (N21)? 1'b0 : 
                            (N22)? 1'b0 : 
                            (N23)? 1'b0 : 
                            (N24)? csr_we_int : 
                            (N25)? 1'b0 : 
                            (N26)? 1'b0 : 
                            (N27)? 1'b0 : 
                            (N28)? 1'b0 : 
                            (N484)? 1'b0 : 1'b0;
  assign { mhpmcounter_we[2:2], mhpmcounter_we[0:0] } = (N13)? { 1'b0, 1'b0 } : 
                                                        (N15)? { 1'b0, 1'b0 } : 
                                                        (N17)? { 1'b0, 1'b0 } : 
                                                        (N18)? { 1'b0, 1'b0 } : 
                                                        (N19)? { 1'b0, 1'b0 } : 
                                                        (N20)? { 1'b0, 1'b0 } : 
                                                        (N21)? { 1'b0, 1'b0 } : 
                                                        (N22)? { 1'b0, 1'b0 } : 
                                                        (N23)? { 1'b0, 1'b0 } : 
                                                        (N24)? { 1'b0, 1'b0 } : 
                                                        (N25)? { 1'b0, csr_we_int } : 
                                                        (N26)? { 1'b0, 1'b0 } : 
                                                        (N27)? { csr_we_int, 1'b0 } : 
                                                        (N28)? { 1'b0, 1'b0 } : 
                                                        (N484)? { N852, N850 } : 1'b0;
  assign { mhpmcounter_we[31:3], mhpmcounter_we[1:1] } = (N484)? { N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N851 } : 
                                                         (N1018)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { mhpmcounterh_we[2:2], mhpmcounterh_we[0:0] } = (N13)? { 1'b0, 1'b0 } : 
                                                          (N15)? { 1'b0, 1'b0 } : 
                                                          (N17)? { 1'b0, 1'b0 } : 
                                                          (N18)? { 1'b0, 1'b0 } : 
                                                          (N19)? { 1'b0, 1'b0 } : 
                                                          (N20)? { 1'b0, 1'b0 } : 
                                                          (N21)? { 1'b0, 1'b0 } : 
                                                          (N22)? { 1'b0, 1'b0 } : 
                                                          (N23)? { 1'b0, 1'b0 } : 
                                                          (N24)? { 1'b0, 1'b0 } : 
                                                          (N25)? { 1'b0, 1'b0 } : 
                                                          (N26)? { 1'b0, csr_we_int } : 
                                                          (N27)? { 1'b0, 1'b0 } : 
                                                          (N28)? { csr_we_int, 1'b0 } : 
                                                          (N484)? { N820, N818 } : 1'b0;
  assign { mhpmcounterh_we[31:3], mhpmcounterh_we[1:1] } = (N484)? { N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N819 } : 
                                                           (N1018)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023 } = (N34)? pc_if_i : 
                                                                                                                                                                                                                                              (N1022)? pc_id_i : 
                                                                                                                                                                                                                                              (N33)? pc_id_i : 1'b0;
  assign N34 = csr_save_if_i;
  assign { N1060, N1059, N1058, N1057, N1056 } = (N35)? { debug_cause_i, 1'b1, 1'b1 } : 
                                                 (N36)? { N962, N961, N960, N955, N954 } : 1'b0;
  assign N35 = debug_csr_save_i;
  assign N36 = N1055;
  assign { N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061 } = (N35)? { N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023 } : 
                                                                                                                                                                                                                                              (N36)? { N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986 } : 1'b0;
  assign { N1094, N1093 } = (N35)? { N883, N882 } : 
                            (N36)? { 1'b0, m_irq_enable_o } : 1'b0;
  assign { N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095 } = (N35)? { N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884 } : 
                                                                                                                                                                                                                                              (N36)? { N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023 } : 1'b0;
  assign { N1132, N1131, N1130, N1129, N1128, N1127 } = (N35)? { N921, N920, N919, N918, N917, N916 } : 
                                                        (N36)? csr_mcause_i : 1'b0;
  assign { N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133 } = (N35)? { N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922 } : 
                                                                                                                                                                                                                                              (N36)? csr_mtval_i : 1'b0;
  assign mcause_d = (N37)? { N1132, N1131, N1130, N1129, N1128, N1127 } : 
                    (N1165)? { N921, N920, N919, N918, N917, N916 } : 
                    (N33)? { N921, N920, N919, N918, N917, N916 } : 
                    (N33)? { N921, N920, N919, N918, N917, N916 } : 1'b0;
  assign N37 = csr_save_cause_i;
  assign mtval_d = (N37)? { N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133 } : 
                   (N1165)? { N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922 } : 
                   (N33)? { N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922 } : 
                   (N33)? { N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922 } : 1'b0;
  assign { dcsr_d[8:6], dcsr_d[1:0] } = (N37)? { N1060, N1059, N1058, N1057, N1056 } : 
                                        (N1165)? { N962, N961, N960, N955, N954 } : 
                                        (N33)? { N962, N961, N960, N955, N954 } : 
                                        (N33)? { N962, N961, N960, N955, N954 } : 1'b0;
  assign depc_d = (N37)? { N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061 } : 
                  (N1165)? { N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986 } : 
                  (N33)? { N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986 } : 
                  (N33)? { N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986 } : 1'b0;
  assign { mstatus_d_mie_, mstatus_d_mpie_ } = (N37)? { N1094, N1093 } : 
                                               (N38)? { mstatus_q_mpie_, 1'b1 } : 
                                               (N39)? { mstatus_q_mpie_, 1'b1 } : 
                                               (N1021)? { N883, N882 } : 1'b0;
  assign N38 = csr_restore_mret_i;
  assign N39 = csr_restore_dret_i;
  assign mepc_d = (N37)? { N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095 } : 
                  (N1165)? { N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884 } : 
                  (N33)? { N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884 } : 
                  (N33)? { N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884 } : 1'b0;
  assign csr_wdata_int = (N40)? csr_wdata_i : 
                         (N41)? { N1174, N1175, N1176, N1177, N1178, N1179, N1180, N1181, N1182, N1183, N1184, N1185, N1186, N1187, N1188, N1189, N1190, N1191, N1192, N1193, N1194, N1195, N1196, N1197, N1198, N1199, N1200, N1201, N1202, N1203, N1204, N1205 } : 
                         (N42)? { N1206, N1207, N1208, N1209, N1210, N1211, N1212, N1213, N1214, N1215, N1216, N1217, N1218, N1219, N1220, N1221, N1222, N1223, N1224, N1225, N1226, N1227, N1228, N1229, N1230, N1231, N1232, N1233, N1234, N1235, N1236, N1237 } : 
                         (N43)? csr_wdata_i : 1'b0;
  assign N40 = N1167;
  assign N41 = N1169;
  assign N42 = N1170;
  assign N43 = N1173;
  assign csr_wreq = (N40)? 1'b1 : 
                    (N41)? 1'b1 : 
                    (N42)? 1'b1 : 
                    (N43)? 1'b0 : 1'b0;
  assign { mcountinhibit_d, mcountinhibit_d_0 } = (N44)? { csr_wdata_int[31:2], csr_wdata_int[0:0] } : 
                                                  (N45)? { mcountinhibit_q[31:2], mcountinhibit_q[0:0] } : 1'b0;
  assign N44 = mcountinhibit_we;
  assign N45 = N1239;
  assign { N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370 } = (N46)? { N1306, N1307, N1308, N1309, N1310, N1311, N1312, N1313, N1314, N1315, N1316, N1317, N1318, N1319, N1320, N1321, N1322, N1323, N1324, N1325, N1326, N1327, N1328, N1329, N1330, N1331, N1332, N1333, N1334, N1335, N1336, N1337, N1338, N1339, N1340, N1341, N1342, N1343, N1344, N1345, N1346, N1347, N1348, N1349, N1350, N1351, N1352, N1353, N1354, N1355, N1356, N1357, N1358, N1359, N1360, N1361, N1362, N1363, N1364, N1365, N1366, N1367, N1368, N1369 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1241)? mhpmcounter_q[2047:1984] : 1'b0;
  assign N46 = N1240;
  assign { N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500 } = (N47)? { N1468, N1469, N1470, N1471, N1472, N1473, N1474, N1475, N1476, N1477, N1478, N1479, N1480, N1481, N1482, N1483, N1484, N1485, N1486, N1487, N1488, N1489, N1490, N1491, N1492, N1493, N1494, N1495, N1496, N1497, N1498, N1499 } : 
                                                                                                                                                                                                                                              (N48)? { N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402 } : 1'b0;
  assign N47 = mhpmcounterh_we[0];
  assign N48 = N1467;
  assign mhpmcounter_d[2047:1984] = (N49)? { N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1435, N1436, N1437, N1438, N1439, N1440, N1441, N1442, N1443, N1444, N1445, N1446, N1447, N1448, N1449, N1450, N1451, N1452, N1453, N1454, N1455, N1456, N1457, N1458, N1459, N1460, N1461, N1462, N1463, N1464, N1465, N1466 } : 
                                    (N50)? { N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370 } : 1'b0;
  assign N49 = mhpmcounter_we[0];
  assign N50 = N1434;
  assign { N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694, N1693, N1692, N1691, N1690, N1689, N1688, N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662 } = (N51)? { N1598, N1599, N1600, N1601, N1602, N1603, N1604, N1605, N1606, N1607, N1608, N1609, N1610, N1611, N1612, N1613, N1614, N1615, N1616, N1617, N1618, N1619, N1620, N1621, N1622, N1623, N1624, N1625, N1626, N1627, N1628, N1629, N1630, N1631, N1632, N1633, N1634, N1635, N1636, N1637, N1638, N1639, N1640, N1641, N1642, N1643, N1644, N1645, N1646, N1647, N1648, N1649, N1650, N1651, N1652, N1653, N1654, N1655, N1656, N1657, N1658, N1659, N1660, N1661 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1533)? mhpmcounter_q[1983:1920] : 1'b0;
  assign N51 = N1532;
  assign { N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792 } = (N52)? { N1760, N1761, N1762, N1763, N1764, N1765, N1766, N1767, N1768, N1769, N1770, N1771, N1772, N1773, N1774, N1775, N1776, N1777, N1778, N1779, N1780, N1781, N1782, N1783, N1784, N1785, N1786, N1787, N1788, N1789, N1790, N1791 } : 
                                                                                                                                                                                                                                              (N53)? { N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694 } : 1'b0;
  assign N52 = mhpmcounterh_we[1];
  assign N53 = N1759;
  assign mhpmcounter_d[1983:1920] = (N54)? { N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694, N1727, N1728, N1729, N1730, N1731, N1732, N1733, N1734, N1735, N1736, N1737, N1738, N1739, N1740, N1741, N1742, N1743, N1744, N1745, N1746, N1747, N1748, N1749, N1750, N1751, N1752, N1753, N1754, N1755, N1756, N1757, N1758 } : 
                                    (N55)? { N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1693, N1692, N1691, N1690, N1689, N1688, N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662 } : 1'b0;
  assign N54 = mhpmcounter_we[1];
  assign N55 = N1726;
  assign { N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, N2008, N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954 } = (N56)? { N1890, N1891, N1892, N1893, N1894, N1895, N1896, N1897, N1898, N1899, N1900, N1901, N1902, N1903, N1904, N1905, N1906, N1907, N1908, N1909, N1910, N1911, N1912, N1913, N1914, N1915, N1916, N1917, N1918, N1919, N1920, N1921, N1922, N1923, N1924, N1925, N1926, N1927, N1928, N1929, N1930, N1931, N1932, N1933, N1934, N1935, N1936, N1937, N1938, N1939, N1940, N1941, N1942, N1943, N1944, N1945, N1946, N1947, N1948, N1949, N1950, N1951, N1952, N1953 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1825)? mhpmcounter_q[1919:1856] : 1'b0;
  assign N56 = N1824;
  assign { N2115, N2114, N2113, N2112, N2111, N2110, N2109, N2108, N2107, N2106, N2105, N2104, N2103, N2102, N2101, N2100, N2099, N2098, N2097, N2096, N2095, N2094, N2093, N2092, N2091, N2090, N2089, N2088, N2087, N2086, N2085, N2084 } = (N57)? { N2052, N2053, N2054, N2055, N2056, N2057, N2058, N2059, N2060, N2061, N2062, N2063, N2064, N2065, N2066, N2067, N2068, N2069, N2070, N2071, N2072, N2073, N2074, N2075, N2076, N2077, N2078, N2079, N2080, N2081, N2082, N2083 } : 
                                                                                                                                                                                                                                              (N58)? { N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, N2008, N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986 } : 1'b0;
  assign N57 = mhpmcounterh_we[2];
  assign N58 = N2051;
  assign mhpmcounter_d[1919:1856] = (N59)? { N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, N2008, N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986, N2019, N2020, N2021, N2022, N2023, N2024, N2025, N2026, N2027, N2028, N2029, N2030, N2031, N2032, N2033, N2034, N2035, N2036, N2037, N2038, N2039, N2040, N2041, N2042, N2043, N2044, N2045, N2046, N2047, N2048, N2049, N2050 } : 
                                    (N60)? { N2115, N2114, N2113, N2112, N2111, N2110, N2109, N2108, N2107, N2106, N2105, N2104, N2103, N2102, N2101, N2100, N2099, N2098, N2097, N2096, N2095, N2094, N2093, N2092, N2091, N2090, N2089, N2088, N2087, N2086, N2085, N2084, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954 } : 1'b0;
  assign N59 = mhpmcounter_we[2];
  assign N60 = N2018;
  assign { N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277, N2276, N2275, N2274, N2273, N2272, N2271, N2270, N2269, N2268, N2267, N2266, N2265, N2264, N2263, N2262, N2261, N2260, N2259, N2258, N2257, N2256, N2255, N2254, N2253, N2252, N2251, N2250, N2249, N2248, N2247, N2246 } = (N61)? { N2182, N2183, N2184, N2185, N2186, N2187, N2188, N2189, N2190, N2191, N2192, N2193, N2194, N2195, N2196, N2197, N2198, N2199, N2200, N2201, N2202, N2203, N2204, N2205, N2206, N2207, N2208, N2209, N2210, N2211, N2212, N2213, N2214, N2215, N2216, N2217, N2218, N2219, N2220, N2221, N2222, N2223, N2224, N2225, N2226, N2227, N2228, N2229, N2230, N2231, N2232, N2233, N2234, N2235, N2236, N2237, N2238, N2239, N2240, N2241, N2242, N2243, N2244, N2245 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2117)? mhpmcounter_q[1855:1792] : 1'b0;
  assign N61 = N2116;
  assign { N2407, N2406, N2405, N2404, N2403, N2402, N2401, N2400, N2399, N2398, N2397, N2396, N2395, N2394, N2393, N2392, N2391, N2390, N2389, N2388, N2387, N2386, N2385, N2384, N2383, N2382, N2381, N2380, N2379, N2378, N2377, N2376 } = (N62)? { N2344, N2345, N2346, N2347, N2348, N2349, N2350, N2351, N2352, N2353, N2354, N2355, N2356, N2357, N2358, N2359, N2360, N2361, N2362, N2363, N2364, N2365, N2366, N2367, N2368, N2369, N2370, N2371, N2372, N2373, N2374, N2375 } : 
                                                                                                                                                                                                                                              (N63)? { N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278 } : 1'b0;
  assign N62 = mhpmcounterh_we[3];
  assign N63 = N2343;
  assign mhpmcounter_d[1855:1792] = (N64)? { N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2311, N2312, N2313, N2314, N2315, N2316, N2317, N2318, N2319, N2320, N2321, N2322, N2323, N2324, N2325, N2326, N2327, N2328, N2329, N2330, N2331, N2332, N2333, N2334, N2335, N2336, N2337, N2338, N2339, N2340, N2341, N2342 } : 
                                    (N65)? { N2407, N2406, N2405, N2404, N2403, N2402, N2401, N2400, N2399, N2398, N2397, N2396, N2395, N2394, N2393, N2392, N2391, N2390, N2389, N2388, N2387, N2386, N2385, N2384, N2383, N2382, N2381, N2380, N2379, N2378, N2377, N2376, N2277, N2276, N2275, N2274, N2273, N2272, N2271, N2270, N2269, N2268, N2267, N2266, N2265, N2264, N2263, N2262, N2261, N2260, N2259, N2258, N2257, N2256, N2255, N2254, N2253, N2252, N2251, N2250, N2249, N2248, N2247, N2246 } : 1'b0;
  assign N64 = mhpmcounter_we[3];
  assign N65 = N2310;
  assign { N2601, N2600, N2599, N2598, N2597, N2596, N2595, N2594, N2593, N2592, N2591, N2590, N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579, N2578, N2577, N2576, N2575, N2574, N2573, N2572, N2571, N2570, N2569, N2568, N2567, N2566, N2565, N2564, N2563, N2562, N2561, N2560, N2559, N2558, N2557, N2556, N2555, N2554, N2553, N2552, N2551, N2550, N2549, N2548, N2547, N2546, N2545, N2544, N2543, N2542, N2541, N2540, N2539, N2538 } = (N66)? { N2474, N2475, N2476, N2477, N2478, N2479, N2480, N2481, N2482, N2483, N2484, N2485, N2486, N2487, N2488, N2489, N2490, N2491, N2492, N2493, N2494, N2495, N2496, N2497, N2498, N2499, N2500, N2501, N2502, N2503, N2504, N2505, N2506, N2507, N2508, N2509, N2510, N2511, N2512, N2513, N2514, N2515, N2516, N2517, N2518, N2519, N2520, N2521, N2522, N2523, N2524, N2525, N2526, N2527, N2528, N2529, N2530, N2531, N2532, N2533, N2534, N2535, N2536, N2537 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2409)? mhpmcounter_q[1791:1728] : 1'b0;
  assign N66 = N2408;
  assign { N2699, N2698, N2697, N2696, N2695, N2694, N2693, N2692, N2691, N2690, N2689, N2688, N2687, N2686, N2685, N2684, N2683, N2682, N2681, N2680, N2679, N2678, N2677, N2676, N2675, N2674, N2673, N2672, N2671, N2670, N2669, N2668 } = (N67)? { N2636, N2637, N2638, N2639, N2640, N2641, N2642, N2643, N2644, N2645, N2646, N2647, N2648, N2649, N2650, N2651, N2652, N2653, N2654, N2655, N2656, N2657, N2658, N2659, N2660, N2661, N2662, N2663, N2664, N2665, N2666, N2667 } : 
                                                                                                                                                                                                                                              (N68)? { N2601, N2600, N2599, N2598, N2597, N2596, N2595, N2594, N2593, N2592, N2591, N2590, N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579, N2578, N2577, N2576, N2575, N2574, N2573, N2572, N2571, N2570 } : 1'b0;
  assign N67 = mhpmcounterh_we[4];
  assign N68 = N2635;
  assign mhpmcounter_d[1791:1728] = (N69)? { N2601, N2600, N2599, N2598, N2597, N2596, N2595, N2594, N2593, N2592, N2591, N2590, N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579, N2578, N2577, N2576, N2575, N2574, N2573, N2572, N2571, N2570, N2603, N2604, N2605, N2606, N2607, N2608, N2609, N2610, N2611, N2612, N2613, N2614, N2615, N2616, N2617, N2618, N2619, N2620, N2621, N2622, N2623, N2624, N2625, N2626, N2627, N2628, N2629, N2630, N2631, N2632, N2633, N2634 } : 
                                    (N70)? { N2699, N2698, N2697, N2696, N2695, N2694, N2693, N2692, N2691, N2690, N2689, N2688, N2687, N2686, N2685, N2684, N2683, N2682, N2681, N2680, N2679, N2678, N2677, N2676, N2675, N2674, N2673, N2672, N2671, N2670, N2669, N2668, N2569, N2568, N2567, N2566, N2565, N2564, N2563, N2562, N2561, N2560, N2559, N2558, N2557, N2556, N2555, N2554, N2553, N2552, N2551, N2550, N2549, N2548, N2547, N2546, N2545, N2544, N2543, N2542, N2541, N2540, N2539, N2538 } : 1'b0;
  assign N69 = mhpmcounter_we[4];
  assign N70 = N2602;
  assign { N2893, N2892, N2891, N2890, N2889, N2888, N2887, N2886, N2885, N2884, N2883, N2882, N2881, N2880, N2879, N2878, N2877, N2876, N2875, N2874, N2873, N2872, N2871, N2870, N2869, N2868, N2867, N2866, N2865, N2864, N2863, N2862, N2861, N2860, N2859, N2858, N2857, N2856, N2855, N2854, N2853, N2852, N2851, N2850, N2849, N2848, N2847, N2846, N2845, N2844, N2843, N2842, N2841, N2840, N2839, N2838, N2837, N2836, N2835, N2834, N2833, N2832, N2831, N2830 } = (N71)? { N2766, N2767, N2768, N2769, N2770, N2771, N2772, N2773, N2774, N2775, N2776, N2777, N2778, N2779, N2780, N2781, N2782, N2783, N2784, N2785, N2786, N2787, N2788, N2789, N2790, N2791, N2792, N2793, N2794, N2795, N2796, N2797, N2798, N2799, N2800, N2801, N2802, N2803, N2804, N2805, N2806, N2807, N2808, N2809, N2810, N2811, N2812, N2813, N2814, N2815, N2816, N2817, N2818, N2819, N2820, N2821, N2822, N2823, N2824, N2825, N2826, N2827, N2828, N2829 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2701)? mhpmcounter_q[1727:1664] : 1'b0;
  assign N71 = N2700;
  assign { N2991, N2990, N2989, N2988, N2987, N2986, N2985, N2984, N2983, N2982, N2981, N2980, N2979, N2978, N2977, N2976, N2975, N2974, N2973, N2972, N2971, N2970, N2969, N2968, N2967, N2966, N2965, N2964, N2963, N2962, N2961, N2960 } = (N72)? { N2928, N2929, N2930, N2931, N2932, N2933, N2934, N2935, N2936, N2937, N2938, N2939, N2940, N2941, N2942, N2943, N2944, N2945, N2946, N2947, N2948, N2949, N2950, N2951, N2952, N2953, N2954, N2955, N2956, N2957, N2958, N2959 } : 
                                                                                                                                                                                                                                              (N73)? { N2893, N2892, N2891, N2890, N2889, N2888, N2887, N2886, N2885, N2884, N2883, N2882, N2881, N2880, N2879, N2878, N2877, N2876, N2875, N2874, N2873, N2872, N2871, N2870, N2869, N2868, N2867, N2866, N2865, N2864, N2863, N2862 } : 1'b0;
  assign N72 = mhpmcounterh_we[5];
  assign N73 = N2927;
  assign mhpmcounter_d[1727:1664] = (N74)? { N2893, N2892, N2891, N2890, N2889, N2888, N2887, N2886, N2885, N2884, N2883, N2882, N2881, N2880, N2879, N2878, N2877, N2876, N2875, N2874, N2873, N2872, N2871, N2870, N2869, N2868, N2867, N2866, N2865, N2864, N2863, N2862, N2895, N2896, N2897, N2898, N2899, N2900, N2901, N2902, N2903, N2904, N2905, N2906, N2907, N2908, N2909, N2910, N2911, N2912, N2913, N2914, N2915, N2916, N2917, N2918, N2919, N2920, N2921, N2922, N2923, N2924, N2925, N2926 } : 
                                    (N75)? { N2991, N2990, N2989, N2988, N2987, N2986, N2985, N2984, N2983, N2982, N2981, N2980, N2979, N2978, N2977, N2976, N2975, N2974, N2973, N2972, N2971, N2970, N2969, N2968, N2967, N2966, N2965, N2964, N2963, N2962, N2961, N2960, N2861, N2860, N2859, N2858, N2857, N2856, N2855, N2854, N2853, N2852, N2851, N2850, N2849, N2848, N2847, N2846, N2845, N2844, N2843, N2842, N2841, N2840, N2839, N2838, N2837, N2836, N2835, N2834, N2833, N2832, N2831, N2830 } : 1'b0;
  assign N74 = mhpmcounter_we[5];
  assign N75 = N2894;
  assign { N3185, N3184, N3183, N3182, N3181, N3180, N3179, N3178, N3177, N3176, N3175, N3174, N3173, N3172, N3171, N3170, N3169, N3168, N3167, N3166, N3165, N3164, N3163, N3162, N3161, N3160, N3159, N3158, N3157, N3156, N3155, N3154, N3153, N3152, N3151, N3150, N3149, N3148, N3147, N3146, N3145, N3144, N3143, N3142, N3141, N3140, N3139, N3138, N3137, N3136, N3135, N3134, N3133, N3132, N3131, N3130, N3129, N3128, N3127, N3126, N3125, N3124, N3123, N3122 } = (N76)? { N3058, N3059, N3060, N3061, N3062, N3063, N3064, N3065, N3066, N3067, N3068, N3069, N3070, N3071, N3072, N3073, N3074, N3075, N3076, N3077, N3078, N3079, N3080, N3081, N3082, N3083, N3084, N3085, N3086, N3087, N3088, N3089, N3090, N3091, N3092, N3093, N3094, N3095, N3096, N3097, N3098, N3099, N3100, N3101, N3102, N3103, N3104, N3105, N3106, N3107, N3108, N3109, N3110, N3111, N3112, N3113, N3114, N3115, N3116, N3117, N3118, N3119, N3120, N3121 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2993)? mhpmcounter_q[1663:1600] : 1'b0;
  assign N76 = N2992;
  assign { N3283, N3282, N3281, N3280, N3279, N3278, N3277, N3276, N3275, N3274, N3273, N3272, N3271, N3270, N3269, N3268, N3267, N3266, N3265, N3264, N3263, N3262, N3261, N3260, N3259, N3258, N3257, N3256, N3255, N3254, N3253, N3252 } = (N77)? { N3220, N3221, N3222, N3223, N3224, N3225, N3226, N3227, N3228, N3229, N3230, N3231, N3232, N3233, N3234, N3235, N3236, N3237, N3238, N3239, N3240, N3241, N3242, N3243, N3244, N3245, N3246, N3247, N3248, N3249, N3250, N3251 } : 
                                                                                                                                                                                                                                              (N78)? { N3185, N3184, N3183, N3182, N3181, N3180, N3179, N3178, N3177, N3176, N3175, N3174, N3173, N3172, N3171, N3170, N3169, N3168, N3167, N3166, N3165, N3164, N3163, N3162, N3161, N3160, N3159, N3158, N3157, N3156, N3155, N3154 } : 1'b0;
  assign N77 = mhpmcounterh_we[6];
  assign N78 = N3219;
  assign mhpmcounter_d[1663:1600] = (N79)? { N3185, N3184, N3183, N3182, N3181, N3180, N3179, N3178, N3177, N3176, N3175, N3174, N3173, N3172, N3171, N3170, N3169, N3168, N3167, N3166, N3165, N3164, N3163, N3162, N3161, N3160, N3159, N3158, N3157, N3156, N3155, N3154, N3187, N3188, N3189, N3190, N3191, N3192, N3193, N3194, N3195, N3196, N3197, N3198, N3199, N3200, N3201, N3202, N3203, N3204, N3205, N3206, N3207, N3208, N3209, N3210, N3211, N3212, N3213, N3214, N3215, N3216, N3217, N3218 } : 
                                    (N80)? { N3283, N3282, N3281, N3280, N3279, N3278, N3277, N3276, N3275, N3274, N3273, N3272, N3271, N3270, N3269, N3268, N3267, N3266, N3265, N3264, N3263, N3262, N3261, N3260, N3259, N3258, N3257, N3256, N3255, N3254, N3253, N3252, N3153, N3152, N3151, N3150, N3149, N3148, N3147, N3146, N3145, N3144, N3143, N3142, N3141, N3140, N3139, N3138, N3137, N3136, N3135, N3134, N3133, N3132, N3131, N3130, N3129, N3128, N3127, N3126, N3125, N3124, N3123, N3122 } : 1'b0;
  assign N79 = mhpmcounter_we[6];
  assign N80 = N3186;
  assign { N3477, N3476, N3475, N3474, N3473, N3472, N3471, N3470, N3469, N3468, N3467, N3466, N3465, N3464, N3463, N3462, N3461, N3460, N3459, N3458, N3457, N3456, N3455, N3454, N3453, N3452, N3451, N3450, N3449, N3448, N3447, N3446, N3445, N3444, N3443, N3442, N3441, N3440, N3439, N3438, N3437, N3436, N3435, N3434, N3433, N3432, N3431, N3430, N3429, N3428, N3427, N3426, N3425, N3424, N3423, N3422, N3421, N3420, N3419, N3418, N3417, N3416, N3415, N3414 } = (N81)? { N3350, N3351, N3352, N3353, N3354, N3355, N3356, N3357, N3358, N3359, N3360, N3361, N3362, N3363, N3364, N3365, N3366, N3367, N3368, N3369, N3370, N3371, N3372, N3373, N3374, N3375, N3376, N3377, N3378, N3379, N3380, N3381, N3382, N3383, N3384, N3385, N3386, N3387, N3388, N3389, N3390, N3391, N3392, N3393, N3394, N3395, N3396, N3397, N3398, N3399, N3400, N3401, N3402, N3403, N3404, N3405, N3406, N3407, N3408, N3409, N3410, N3411, N3412, N3413 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3285)? mhpmcounter_q[1599:1536] : 1'b0;
  assign N81 = N3284;
  assign { N3575, N3574, N3573, N3572, N3571, N3570, N3569, N3568, N3567, N3566, N3565, N3564, N3563, N3562, N3561, N3560, N3559, N3558, N3557, N3556, N3555, N3554, N3553, N3552, N3551, N3550, N3549, N3548, N3547, N3546, N3545, N3544 } = (N82)? { N3512, N3513, N3514, N3515, N3516, N3517, N3518, N3519, N3520, N3521, N3522, N3523, N3524, N3525, N3526, N3527, N3528, N3529, N3530, N3531, N3532, N3533, N3534, N3535, N3536, N3537, N3538, N3539, N3540, N3541, N3542, N3543 } : 
                                                                                                                                                                                                                                              (N83)? { N3477, N3476, N3475, N3474, N3473, N3472, N3471, N3470, N3469, N3468, N3467, N3466, N3465, N3464, N3463, N3462, N3461, N3460, N3459, N3458, N3457, N3456, N3455, N3454, N3453, N3452, N3451, N3450, N3449, N3448, N3447, N3446 } : 1'b0;
  assign N82 = mhpmcounterh_we[7];
  assign N83 = N3511;
  assign mhpmcounter_d[1599:1536] = (N84)? { N3477, N3476, N3475, N3474, N3473, N3472, N3471, N3470, N3469, N3468, N3467, N3466, N3465, N3464, N3463, N3462, N3461, N3460, N3459, N3458, N3457, N3456, N3455, N3454, N3453, N3452, N3451, N3450, N3449, N3448, N3447, N3446, N3479, N3480, N3481, N3482, N3483, N3484, N3485, N3486, N3487, N3488, N3489, N3490, N3491, N3492, N3493, N3494, N3495, N3496, N3497, N3498, N3499, N3500, N3501, N3502, N3503, N3504, N3505, N3506, N3507, N3508, N3509, N3510 } : 
                                    (N85)? { N3575, N3574, N3573, N3572, N3571, N3570, N3569, N3568, N3567, N3566, N3565, N3564, N3563, N3562, N3561, N3560, N3559, N3558, N3557, N3556, N3555, N3554, N3553, N3552, N3551, N3550, N3549, N3548, N3547, N3546, N3545, N3544, N3445, N3444, N3443, N3442, N3441, N3440, N3439, N3438, N3437, N3436, N3435, N3434, N3433, N3432, N3431, N3430, N3429, N3428, N3427, N3426, N3425, N3424, N3423, N3422, N3421, N3420, N3419, N3418, N3417, N3416, N3415, N3414 } : 1'b0;
  assign N84 = mhpmcounter_we[7];
  assign N85 = N3478;
  assign { N3769, N3768, N3767, N3766, N3765, N3764, N3763, N3762, N3761, N3760, N3759, N3758, N3757, N3756, N3755, N3754, N3753, N3752, N3751, N3750, N3749, N3748, N3747, N3746, N3745, N3744, N3743, N3742, N3741, N3740, N3739, N3738, N3737, N3736, N3735, N3734, N3733, N3732, N3731, N3730, N3729, N3728, N3727, N3726, N3725, N3724, N3723, N3722, N3721, N3720, N3719, N3718, N3717, N3716, N3715, N3714, N3713, N3712, N3711, N3710, N3709, N3708, N3707, N3706 } = (N86)? { N3642, N3643, N3644, N3645, N3646, N3647, N3648, N3649, N3650, N3651, N3652, N3653, N3654, N3655, N3656, N3657, N3658, N3659, N3660, N3661, N3662, N3663, N3664, N3665, N3666, N3667, N3668, N3669, N3670, N3671, N3672, N3673, N3674, N3675, N3676, N3677, N3678, N3679, N3680, N3681, N3682, N3683, N3684, N3685, N3686, N3687, N3688, N3689, N3690, N3691, N3692, N3693, N3694, N3695, N3696, N3697, N3698, N3699, N3700, N3701, N3702, N3703, N3704, N3705 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3577)? mhpmcounter_q[1535:1472] : 1'b0;
  assign N86 = N3576;
  assign { N3867, N3866, N3865, N3864, N3863, N3862, N3861, N3860, N3859, N3858, N3857, N3856, N3855, N3854, N3853, N3852, N3851, N3850, N3849, N3848, N3847, N3846, N3845, N3844, N3843, N3842, N3841, N3840, N3839, N3838, N3837, N3836 } = (N87)? { N3804, N3805, N3806, N3807, N3808, N3809, N3810, N3811, N3812, N3813, N3814, N3815, N3816, N3817, N3818, N3819, N3820, N3821, N3822, N3823, N3824, N3825, N3826, N3827, N3828, N3829, N3830, N3831, N3832, N3833, N3834, N3835 } : 
                                                                                                                                                                                                                                              (N88)? { N3769, N3768, N3767, N3766, N3765, N3764, N3763, N3762, N3761, N3760, N3759, N3758, N3757, N3756, N3755, N3754, N3753, N3752, N3751, N3750, N3749, N3748, N3747, N3746, N3745, N3744, N3743, N3742, N3741, N3740, N3739, N3738 } : 1'b0;
  assign N87 = mhpmcounterh_we[8];
  assign N88 = N3803;
  assign mhpmcounter_d[1535:1472] = (N89)? { N3769, N3768, N3767, N3766, N3765, N3764, N3763, N3762, N3761, N3760, N3759, N3758, N3757, N3756, N3755, N3754, N3753, N3752, N3751, N3750, N3749, N3748, N3747, N3746, N3745, N3744, N3743, N3742, N3741, N3740, N3739, N3738, N3771, N3772, N3773, N3774, N3775, N3776, N3777, N3778, N3779, N3780, N3781, N3782, N3783, N3784, N3785, N3786, N3787, N3788, N3789, N3790, N3791, N3792, N3793, N3794, N3795, N3796, N3797, N3798, N3799, N3800, N3801, N3802 } : 
                                    (N90)? { N3867, N3866, N3865, N3864, N3863, N3862, N3861, N3860, N3859, N3858, N3857, N3856, N3855, N3854, N3853, N3852, N3851, N3850, N3849, N3848, N3847, N3846, N3845, N3844, N3843, N3842, N3841, N3840, N3839, N3838, N3837, N3836, N3737, N3736, N3735, N3734, N3733, N3732, N3731, N3730, N3729, N3728, N3727, N3726, N3725, N3724, N3723, N3722, N3721, N3720, N3719, N3718, N3717, N3716, N3715, N3714, N3713, N3712, N3711, N3710, N3709, N3708, N3707, N3706 } : 1'b0;
  assign N89 = mhpmcounter_we[8];
  assign N90 = N3770;
  assign { N4061, N4060, N4059, N4058, N4057, N4056, N4055, N4054, N4053, N4052, N4051, N4050, N4049, N4048, N4047, N4046, N4045, N4044, N4043, N4042, N4041, N4040, N4039, N4038, N4037, N4036, N4035, N4034, N4033, N4032, N4031, N4030, N4029, N4028, N4027, N4026, N4025, N4024, N4023, N4022, N4021, N4020, N4019, N4018, N4017, N4016, N4015, N4014, N4013, N4012, N4011, N4010, N4009, N4008, N4007, N4006, N4005, N4004, N4003, N4002, N4001, N4000, N3999, N3998 } = (N91)? { N3934, N3935, N3936, N3937, N3938, N3939, N3940, N3941, N3942, N3943, N3944, N3945, N3946, N3947, N3948, N3949, N3950, N3951, N3952, N3953, N3954, N3955, N3956, N3957, N3958, N3959, N3960, N3961, N3962, N3963, N3964, N3965, N3966, N3967, N3968, N3969, N3970, N3971, N3972, N3973, N3974, N3975, N3976, N3977, N3978, N3979, N3980, N3981, N3982, N3983, N3984, N3985, N3986, N3987, N3988, N3989, N3990, N3991, N3992, N3993, N3994, N3995, N3996, N3997 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3869)? mhpmcounter_q[1471:1408] : 1'b0;
  assign N91 = N3868;
  assign { N4159, N4158, N4157, N4156, N4155, N4154, N4153, N4152, N4151, N4150, N4149, N4148, N4147, N4146, N4145, N4144, N4143, N4142, N4141, N4140, N4139, N4138, N4137, N4136, N4135, N4134, N4133, N4132, N4131, N4130, N4129, N4128 } = (N92)? { N4096, N4097, N4098, N4099, N4100, N4101, N4102, N4103, N4104, N4105, N4106, N4107, N4108, N4109, N4110, N4111, N4112, N4113, N4114, N4115, N4116, N4117, N4118, N4119, N4120, N4121, N4122, N4123, N4124, N4125, N4126, N4127 } : 
                                                                                                                                                                                                                                              (N93)? { N4061, N4060, N4059, N4058, N4057, N4056, N4055, N4054, N4053, N4052, N4051, N4050, N4049, N4048, N4047, N4046, N4045, N4044, N4043, N4042, N4041, N4040, N4039, N4038, N4037, N4036, N4035, N4034, N4033, N4032, N4031, N4030 } : 1'b0;
  assign N92 = mhpmcounterh_we[9];
  assign N93 = N4095;
  assign mhpmcounter_d[1471:1408] = (N94)? { N4061, N4060, N4059, N4058, N4057, N4056, N4055, N4054, N4053, N4052, N4051, N4050, N4049, N4048, N4047, N4046, N4045, N4044, N4043, N4042, N4041, N4040, N4039, N4038, N4037, N4036, N4035, N4034, N4033, N4032, N4031, N4030, N4063, N4064, N4065, N4066, N4067, N4068, N4069, N4070, N4071, N4072, N4073, N4074, N4075, N4076, N4077, N4078, N4079, N4080, N4081, N4082, N4083, N4084, N4085, N4086, N4087, N4088, N4089, N4090, N4091, N4092, N4093, N4094 } : 
                                    (N95)? { N4159, N4158, N4157, N4156, N4155, N4154, N4153, N4152, N4151, N4150, N4149, N4148, N4147, N4146, N4145, N4144, N4143, N4142, N4141, N4140, N4139, N4138, N4137, N4136, N4135, N4134, N4133, N4132, N4131, N4130, N4129, N4128, N4029, N4028, N4027, N4026, N4025, N4024, N4023, N4022, N4021, N4020, N4019, N4018, N4017, N4016, N4015, N4014, N4013, N4012, N4011, N4010, N4009, N4008, N4007, N4006, N4005, N4004, N4003, N4002, N4001, N4000, N3999, N3998 } : 1'b0;
  assign N94 = mhpmcounter_we[9];
  assign N95 = N4062;
  assign { N4353, N4352, N4351, N4350, N4349, N4348, N4347, N4346, N4345, N4344, N4343, N4342, N4341, N4340, N4339, N4338, N4337, N4336, N4335, N4334, N4333, N4332, N4331, N4330, N4329, N4328, N4327, N4326, N4325, N4324, N4323, N4322, N4321, N4320, N4319, N4318, N4317, N4316, N4315, N4314, N4313, N4312, N4311, N4310, N4309, N4308, N4307, N4306, N4305, N4304, N4303, N4302, N4301, N4300, N4299, N4298, N4297, N4296, N4295, N4294, N4293, N4292, N4291, N4290 } = (N96)? { N4226, N4227, N4228, N4229, N4230, N4231, N4232, N4233, N4234, N4235, N4236, N4237, N4238, N4239, N4240, N4241, N4242, N4243, N4244, N4245, N4246, N4247, N4248, N4249, N4250, N4251, N4252, N4253, N4254, N4255, N4256, N4257, N4258, N4259, N4260, N4261, N4262, N4263, N4264, N4265, N4266, N4267, N4268, N4269, N4270, N4271, N4272, N4273, N4274, N4275, N4276, N4277, N4278, N4279, N4280, N4281, N4282, N4283, N4284, N4285, N4286, N4287, N4288, N4289 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4161)? mhpmcounter_q[1407:1344] : 1'b0;
  assign N96 = N4160;
  assign { N4451, N4450, N4449, N4448, N4447, N4446, N4445, N4444, N4443, N4442, N4441, N4440, N4439, N4438, N4437, N4436, N4435, N4434, N4433, N4432, N4431, N4430, N4429, N4428, N4427, N4426, N4425, N4424, N4423, N4422, N4421, N4420 } = (N97)? { N4388, N4389, N4390, N4391, N4392, N4393, N4394, N4395, N4396, N4397, N4398, N4399, N4400, N4401, N4402, N4403, N4404, N4405, N4406, N4407, N4408, N4409, N4410, N4411, N4412, N4413, N4414, N4415, N4416, N4417, N4418, N4419 } : 
                                                                                                                                                                                                                                              (N98)? { N4353, N4352, N4351, N4350, N4349, N4348, N4347, N4346, N4345, N4344, N4343, N4342, N4341, N4340, N4339, N4338, N4337, N4336, N4335, N4334, N4333, N4332, N4331, N4330, N4329, N4328, N4327, N4326, N4325, N4324, N4323, N4322 } : 1'b0;
  assign N97 = mhpmcounterh_we[10];
  assign N98 = N4387;
  assign mhpmcounter_d[1407:1344] = (N99)? { N4353, N4352, N4351, N4350, N4349, N4348, N4347, N4346, N4345, N4344, N4343, N4342, N4341, N4340, N4339, N4338, N4337, N4336, N4335, N4334, N4333, N4332, N4331, N4330, N4329, N4328, N4327, N4326, N4325, N4324, N4323, N4322, N4355, N4356, N4357, N4358, N4359, N4360, N4361, N4362, N4363, N4364, N4365, N4366, N4367, N4368, N4369, N4370, N4371, N4372, N4373, N4374, N4375, N4376, N4377, N4378, N4379, N4380, N4381, N4382, N4383, N4384, N4385, N4386 } : 
                                    (N100)? { N4451, N4450, N4449, N4448, N4447, N4446, N4445, N4444, N4443, N4442, N4441, N4440, N4439, N4438, N4437, N4436, N4435, N4434, N4433, N4432, N4431, N4430, N4429, N4428, N4427, N4426, N4425, N4424, N4423, N4422, N4421, N4420, N4321, N4320, N4319, N4318, N4317, N4316, N4315, N4314, N4313, N4312, N4311, N4310, N4309, N4308, N4307, N4306, N4305, N4304, N4303, N4302, N4301, N4300, N4299, N4298, N4297, N4296, N4295, N4294, N4293, N4292, N4291, N4290 } : 1'b0;
  assign N99 = mhpmcounter_we[10];
  assign N100 = N4354;
  assign { N4645, N4644, N4643, N4642, N4641, N4640, N4639, N4638, N4637, N4636, N4635, N4634, N4633, N4632, N4631, N4630, N4629, N4628, N4627, N4626, N4625, N4624, N4623, N4622, N4621, N4620, N4619, N4618, N4617, N4616, N4615, N4614, N4613, N4612, N4611, N4610, N4609, N4608, N4607, N4606, N4605, N4604, N4603, N4602, N4601, N4600, N4599, N4598, N4597, N4596, N4595, N4594, N4593, N4592, N4591, N4590, N4589, N4588, N4587, N4586, N4585, N4584, N4583, N4582 } = (N101)? { N4518, N4519, N4520, N4521, N4522, N4523, N4524, N4525, N4526, N4527, N4528, N4529, N4530, N4531, N4532, N4533, N4534, N4535, N4536, N4537, N4538, N4539, N4540, N4541, N4542, N4543, N4544, N4545, N4546, N4547, N4548, N4549, N4550, N4551, N4552, N4553, N4554, N4555, N4556, N4557, N4558, N4559, N4560, N4561, N4562, N4563, N4564, N4565, N4566, N4567, N4568, N4569, N4570, N4571, N4572, N4573, N4574, N4575, N4576, N4577, N4578, N4579, N4580, N4581 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4453)? mhpmcounter_q[1343:1280] : 1'b0;
  assign N101 = N4452;
  assign { N4743, N4742, N4741, N4740, N4739, N4738, N4737, N4736, N4735, N4734, N4733, N4732, N4731, N4730, N4729, N4728, N4727, N4726, N4725, N4724, N4723, N4722, N4721, N4720, N4719, N4718, N4717, N4716, N4715, N4714, N4713, N4712 } = (N102)? { N4680, N4681, N4682, N4683, N4684, N4685, N4686, N4687, N4688, N4689, N4690, N4691, N4692, N4693, N4694, N4695, N4696, N4697, N4698, N4699, N4700, N4701, N4702, N4703, N4704, N4705, N4706, N4707, N4708, N4709, N4710, N4711 } : 
                                                                                                                                                                                                                                              (N103)? { N4645, N4644, N4643, N4642, N4641, N4640, N4639, N4638, N4637, N4636, N4635, N4634, N4633, N4632, N4631, N4630, N4629, N4628, N4627, N4626, N4625, N4624, N4623, N4622, N4621, N4620, N4619, N4618, N4617, N4616, N4615, N4614 } : 1'b0;
  assign N102 = mhpmcounterh_we[11];
  assign N103 = N4679;
  assign mhpmcounter_d[1343:1280] = (N104)? { N4645, N4644, N4643, N4642, N4641, N4640, N4639, N4638, N4637, N4636, N4635, N4634, N4633, N4632, N4631, N4630, N4629, N4628, N4627, N4626, N4625, N4624, N4623, N4622, N4621, N4620, N4619, N4618, N4617, N4616, N4615, N4614, N4647, N4648, N4649, N4650, N4651, N4652, N4653, N4654, N4655, N4656, N4657, N4658, N4659, N4660, N4661, N4662, N4663, N4664, N4665, N4666, N4667, N4668, N4669, N4670, N4671, N4672, N4673, N4674, N4675, N4676, N4677, N4678 } : 
                                    (N105)? { N4743, N4742, N4741, N4740, N4739, N4738, N4737, N4736, N4735, N4734, N4733, N4732, N4731, N4730, N4729, N4728, N4727, N4726, N4725, N4724, N4723, N4722, N4721, N4720, N4719, N4718, N4717, N4716, N4715, N4714, N4713, N4712, N4613, N4612, N4611, N4610, N4609, N4608, N4607, N4606, N4605, N4604, N4603, N4602, N4601, N4600, N4599, N4598, N4597, N4596, N4595, N4594, N4593, N4592, N4591, N4590, N4589, N4588, N4587, N4586, N4585, N4584, N4583, N4582 } : 1'b0;
  assign N104 = mhpmcounter_we[11];
  assign N105 = N4646;
  assign { N4937, N4936, N4935, N4934, N4933, N4932, N4931, N4930, N4929, N4928, N4927, N4926, N4925, N4924, N4923, N4922, N4921, N4920, N4919, N4918, N4917, N4916, N4915, N4914, N4913, N4912, N4911, N4910, N4909, N4908, N4907, N4906, N4905, N4904, N4903, N4902, N4901, N4900, N4899, N4898, N4897, N4896, N4895, N4894, N4893, N4892, N4891, N4890, N4889, N4888, N4887, N4886, N4885, N4884, N4883, N4882, N4881, N4880, N4879, N4878, N4877, N4876, N4875, N4874 } = (N106)? { N4810, N4811, N4812, N4813, N4814, N4815, N4816, N4817, N4818, N4819, N4820, N4821, N4822, N4823, N4824, N4825, N4826, N4827, N4828, N4829, N4830, N4831, N4832, N4833, N4834, N4835, N4836, N4837, N4838, N4839, N4840, N4841, N4842, N4843, N4844, N4845, N4846, N4847, N4848, N4849, N4850, N4851, N4852, N4853, N4854, N4855, N4856, N4857, N4858, N4859, N4860, N4861, N4862, N4863, N4864, N4865, N4866, N4867, N4868, N4869, N4870, N4871, N4872, N4873 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4745)? mhpmcounter_q[1279:1216] : 1'b0;
  assign N106 = N4744;
  assign { N5035, N5034, N5033, N5032, N5031, N5030, N5029, N5028, N5027, N5026, N5025, N5024, N5023, N5022, N5021, N5020, N5019, N5018, N5017, N5016, N5015, N5014, N5013, N5012, N5011, N5010, N5009, N5008, N5007, N5006, N5005, N5004 } = (N107)? { N4972, N4973, N4974, N4975, N4976, N4977, N4978, N4979, N4980, N4981, N4982, N4983, N4984, N4985, N4986, N4987, N4988, N4989, N4990, N4991, N4992, N4993, N4994, N4995, N4996, N4997, N4998, N4999, N5000, N5001, N5002, N5003 } : 
                                                                                                                                                                                                                                              (N108)? { N4937, N4936, N4935, N4934, N4933, N4932, N4931, N4930, N4929, N4928, N4927, N4926, N4925, N4924, N4923, N4922, N4921, N4920, N4919, N4918, N4917, N4916, N4915, N4914, N4913, N4912, N4911, N4910, N4909, N4908, N4907, N4906 } : 1'b0;
  assign N107 = mhpmcounterh_we[12];
  assign N108 = N4971;
  assign mhpmcounter_d[1279:1216] = (N109)? { N4937, N4936, N4935, N4934, N4933, N4932, N4931, N4930, N4929, N4928, N4927, N4926, N4925, N4924, N4923, N4922, N4921, N4920, N4919, N4918, N4917, N4916, N4915, N4914, N4913, N4912, N4911, N4910, N4909, N4908, N4907, N4906, N4939, N4940, N4941, N4942, N4943, N4944, N4945, N4946, N4947, N4948, N4949, N4950, N4951, N4952, N4953, N4954, N4955, N4956, N4957, N4958, N4959, N4960, N4961, N4962, N4963, N4964, N4965, N4966, N4967, N4968, N4969, N4970 } : 
                                    (N110)? { N5035, N5034, N5033, N5032, N5031, N5030, N5029, N5028, N5027, N5026, N5025, N5024, N5023, N5022, N5021, N5020, N5019, N5018, N5017, N5016, N5015, N5014, N5013, N5012, N5011, N5010, N5009, N5008, N5007, N5006, N5005, N5004, N4905, N4904, N4903, N4902, N4901, N4900, N4899, N4898, N4897, N4896, N4895, N4894, N4893, N4892, N4891, N4890, N4889, N4888, N4887, N4886, N4885, N4884, N4883, N4882, N4881, N4880, N4879, N4878, N4877, N4876, N4875, N4874 } : 1'b0;
  assign N109 = mhpmcounter_we[12];
  assign N110 = N4938;
  assign { N5229, N5228, N5227, N5226, N5225, N5224, N5223, N5222, N5221, N5220, N5219, N5218, N5217, N5216, N5215, N5214, N5213, N5212, N5211, N5210, N5209, N5208, N5207, N5206, N5205, N5204, N5203, N5202, N5201, N5200, N5199, N5198, N5197, N5196, N5195, N5194, N5193, N5192, N5191, N5190, N5189, N5188, N5187, N5186, N5185, N5184, N5183, N5182, N5181, N5180, N5179, N5178, N5177, N5176, N5175, N5174, N5173, N5172, N5171, N5170, N5169, N5168, N5167, N5166 } = (N111)? { N5102, N5103, N5104, N5105, N5106, N5107, N5108, N5109, N5110, N5111, N5112, N5113, N5114, N5115, N5116, N5117, N5118, N5119, N5120, N5121, N5122, N5123, N5124, N5125, N5126, N5127, N5128, N5129, N5130, N5131, N5132, N5133, N5134, N5135, N5136, N5137, N5138, N5139, N5140, N5141, N5142, N5143, N5144, N5145, N5146, N5147, N5148, N5149, N5150, N5151, N5152, N5153, N5154, N5155, N5156, N5157, N5158, N5159, N5160, N5161, N5162, N5163, N5164, N5165 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5037)? mhpmcounter_q[1215:1152] : 1'b0;
  assign N111 = N5036;
  assign { N5327, N5326, N5325, N5324, N5323, N5322, N5321, N5320, N5319, N5318, N5317, N5316, N5315, N5314, N5313, N5312, N5311, N5310, N5309, N5308, N5307, N5306, N5305, N5304, N5303, N5302, N5301, N5300, N5299, N5298, N5297, N5296 } = (N112)? { N5264, N5265, N5266, N5267, N5268, N5269, N5270, N5271, N5272, N5273, N5274, N5275, N5276, N5277, N5278, N5279, N5280, N5281, N5282, N5283, N5284, N5285, N5286, N5287, N5288, N5289, N5290, N5291, N5292, N5293, N5294, N5295 } : 
                                                                                                                                                                                                                                              (N113)? { N5229, N5228, N5227, N5226, N5225, N5224, N5223, N5222, N5221, N5220, N5219, N5218, N5217, N5216, N5215, N5214, N5213, N5212, N5211, N5210, N5209, N5208, N5207, N5206, N5205, N5204, N5203, N5202, N5201, N5200, N5199, N5198 } : 1'b0;
  assign N112 = mhpmcounterh_we[13];
  assign N113 = N5263;
  assign mhpmcounter_d[1215:1152] = (N114)? { N5229, N5228, N5227, N5226, N5225, N5224, N5223, N5222, N5221, N5220, N5219, N5218, N5217, N5216, N5215, N5214, N5213, N5212, N5211, N5210, N5209, N5208, N5207, N5206, N5205, N5204, N5203, N5202, N5201, N5200, N5199, N5198, N5231, N5232, N5233, N5234, N5235, N5236, N5237, N5238, N5239, N5240, N5241, N5242, N5243, N5244, N5245, N5246, N5247, N5248, N5249, N5250, N5251, N5252, N5253, N5254, N5255, N5256, N5257, N5258, N5259, N5260, N5261, N5262 } : 
                                    (N115)? { N5327, N5326, N5325, N5324, N5323, N5322, N5321, N5320, N5319, N5318, N5317, N5316, N5315, N5314, N5313, N5312, N5311, N5310, N5309, N5308, N5307, N5306, N5305, N5304, N5303, N5302, N5301, N5300, N5299, N5298, N5297, N5296, N5197, N5196, N5195, N5194, N5193, N5192, N5191, N5190, N5189, N5188, N5187, N5186, N5185, N5184, N5183, N5182, N5181, N5180, N5179, N5178, N5177, N5176, N5175, N5174, N5173, N5172, N5171, N5170, N5169, N5168, N5167, N5166 } : 1'b0;
  assign N114 = mhpmcounter_we[13];
  assign N115 = N5230;
  assign { N5521, N5520, N5519, N5518, N5517, N5516, N5515, N5514, N5513, N5512, N5511, N5510, N5509, N5508, N5507, N5506, N5505, N5504, N5503, N5502, N5501, N5500, N5499, N5498, N5497, N5496, N5495, N5494, N5493, N5492, N5491, N5490, N5489, N5488, N5487, N5486, N5485, N5484, N5483, N5482, N5481, N5480, N5479, N5478, N5477, N5476, N5475, N5474, N5473, N5472, N5471, N5470, N5469, N5468, N5467, N5466, N5465, N5464, N5463, N5462, N5461, N5460, N5459, N5458 } = (N116)? { N5394, N5395, N5396, N5397, N5398, N5399, N5400, N5401, N5402, N5403, N5404, N5405, N5406, N5407, N5408, N5409, N5410, N5411, N5412, N5413, N5414, N5415, N5416, N5417, N5418, N5419, N5420, N5421, N5422, N5423, N5424, N5425, N5426, N5427, N5428, N5429, N5430, N5431, N5432, N5433, N5434, N5435, N5436, N5437, N5438, N5439, N5440, N5441, N5442, N5443, N5444, N5445, N5446, N5447, N5448, N5449, N5450, N5451, N5452, N5453, N5454, N5455, N5456, N5457 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5329)? mhpmcounter_q[1151:1088] : 1'b0;
  assign N116 = N5328;
  assign { N5619, N5618, N5617, N5616, N5615, N5614, N5613, N5612, N5611, N5610, N5609, N5608, N5607, N5606, N5605, N5604, N5603, N5602, N5601, N5600, N5599, N5598, N5597, N5596, N5595, N5594, N5593, N5592, N5591, N5590, N5589, N5588 } = (N117)? { N5556, N5557, N5558, N5559, N5560, N5561, N5562, N5563, N5564, N5565, N5566, N5567, N5568, N5569, N5570, N5571, N5572, N5573, N5574, N5575, N5576, N5577, N5578, N5579, N5580, N5581, N5582, N5583, N5584, N5585, N5586, N5587 } : 
                                                                                                                                                                                                                                              (N118)? { N5521, N5520, N5519, N5518, N5517, N5516, N5515, N5514, N5513, N5512, N5511, N5510, N5509, N5508, N5507, N5506, N5505, N5504, N5503, N5502, N5501, N5500, N5499, N5498, N5497, N5496, N5495, N5494, N5493, N5492, N5491, N5490 } : 1'b0;
  assign N117 = mhpmcounterh_we[14];
  assign N118 = N5555;
  assign mhpmcounter_d[1151:1088] = (N119)? { N5521, N5520, N5519, N5518, N5517, N5516, N5515, N5514, N5513, N5512, N5511, N5510, N5509, N5508, N5507, N5506, N5505, N5504, N5503, N5502, N5501, N5500, N5499, N5498, N5497, N5496, N5495, N5494, N5493, N5492, N5491, N5490, N5523, N5524, N5525, N5526, N5527, N5528, N5529, N5530, N5531, N5532, N5533, N5534, N5535, N5536, N5537, N5538, N5539, N5540, N5541, N5542, N5543, N5544, N5545, N5546, N5547, N5548, N5549, N5550, N5551, N5552, N5553, N5554 } : 
                                    (N120)? { N5619, N5618, N5617, N5616, N5615, N5614, N5613, N5612, N5611, N5610, N5609, N5608, N5607, N5606, N5605, N5604, N5603, N5602, N5601, N5600, N5599, N5598, N5597, N5596, N5595, N5594, N5593, N5592, N5591, N5590, N5589, N5588, N5489, N5488, N5487, N5486, N5485, N5484, N5483, N5482, N5481, N5480, N5479, N5478, N5477, N5476, N5475, N5474, N5473, N5472, N5471, N5470, N5469, N5468, N5467, N5466, N5465, N5464, N5463, N5462, N5461, N5460, N5459, N5458 } : 1'b0;
  assign N119 = mhpmcounter_we[14];
  assign N120 = N5522;
  assign { N5813, N5812, N5811, N5810, N5809, N5808, N5807, N5806, N5805, N5804, N5803, N5802, N5801, N5800, N5799, N5798, N5797, N5796, N5795, N5794, N5793, N5792, N5791, N5790, N5789, N5788, N5787, N5786, N5785, N5784, N5783, N5782, N5781, N5780, N5779, N5778, N5777, N5776, N5775, N5774, N5773, N5772, N5771, N5770, N5769, N5768, N5767, N5766, N5765, N5764, N5763, N5762, N5761, N5760, N5759, N5758, N5757, N5756, N5755, N5754, N5753, N5752, N5751, N5750 } = (N121)? { N5686, N5687, N5688, N5689, N5690, N5691, N5692, N5693, N5694, N5695, N5696, N5697, N5698, N5699, N5700, N5701, N5702, N5703, N5704, N5705, N5706, N5707, N5708, N5709, N5710, N5711, N5712, N5713, N5714, N5715, N5716, N5717, N5718, N5719, N5720, N5721, N5722, N5723, N5724, N5725, N5726, N5727, N5728, N5729, N5730, N5731, N5732, N5733, N5734, N5735, N5736, N5737, N5738, N5739, N5740, N5741, N5742, N5743, N5744, N5745, N5746, N5747, N5748, N5749 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5621)? mhpmcounter_q[1087:1024] : 1'b0;
  assign N121 = N5620;
  assign { N5911, N5910, N5909, N5908, N5907, N5906, N5905, N5904, N5903, N5902, N5901, N5900, N5899, N5898, N5897, N5896, N5895, N5894, N5893, N5892, N5891, N5890, N5889, N5888, N5887, N5886, N5885, N5884, N5883, N5882, N5881, N5880 } = (N122)? { N5848, N5849, N5850, N5851, N5852, N5853, N5854, N5855, N5856, N5857, N5858, N5859, N5860, N5861, N5862, N5863, N5864, N5865, N5866, N5867, N5868, N5869, N5870, N5871, N5872, N5873, N5874, N5875, N5876, N5877, N5878, N5879 } : 
                                                                                                                                                                                                                                              (N123)? { N5813, N5812, N5811, N5810, N5809, N5808, N5807, N5806, N5805, N5804, N5803, N5802, N5801, N5800, N5799, N5798, N5797, N5796, N5795, N5794, N5793, N5792, N5791, N5790, N5789, N5788, N5787, N5786, N5785, N5784, N5783, N5782 } : 1'b0;
  assign N122 = mhpmcounterh_we[15];
  assign N123 = N5847;
  assign mhpmcounter_d[1087:1024] = (N124)? { N5813, N5812, N5811, N5810, N5809, N5808, N5807, N5806, N5805, N5804, N5803, N5802, N5801, N5800, N5799, N5798, N5797, N5796, N5795, N5794, N5793, N5792, N5791, N5790, N5789, N5788, N5787, N5786, N5785, N5784, N5783, N5782, N5815, N5816, N5817, N5818, N5819, N5820, N5821, N5822, N5823, N5824, N5825, N5826, N5827, N5828, N5829, N5830, N5831, N5832, N5833, N5834, N5835, N5836, N5837, N5838, N5839, N5840, N5841, N5842, N5843, N5844, N5845, N5846 } : 
                                    (N125)? { N5911, N5910, N5909, N5908, N5907, N5906, N5905, N5904, N5903, N5902, N5901, N5900, N5899, N5898, N5897, N5896, N5895, N5894, N5893, N5892, N5891, N5890, N5889, N5888, N5887, N5886, N5885, N5884, N5883, N5882, N5881, N5880, N5781, N5780, N5779, N5778, N5777, N5776, N5775, N5774, N5773, N5772, N5771, N5770, N5769, N5768, N5767, N5766, N5765, N5764, N5763, N5762, N5761, N5760, N5759, N5758, N5757, N5756, N5755, N5754, N5753, N5752, N5751, N5750 } : 1'b0;
  assign N124 = mhpmcounter_we[15];
  assign N125 = N5814;
  assign { N6105, N6104, N6103, N6102, N6101, N6100, N6099, N6098, N6097, N6096, N6095, N6094, N6093, N6092, N6091, N6090, N6089, N6088, N6087, N6086, N6085, N6084, N6083, N6082, N6081, N6080, N6079, N6078, N6077, N6076, N6075, N6074, N6073, N6072, N6071, N6070, N6069, N6068, N6067, N6066, N6065, N6064, N6063, N6062, N6061, N6060, N6059, N6058, N6057, N6056, N6055, N6054, N6053, N6052, N6051, N6050, N6049, N6048, N6047, N6046, N6045, N6044, N6043, N6042 } = (N126)? { N5978, N5979, N5980, N5981, N5982, N5983, N5984, N5985, N5986, N5987, N5988, N5989, N5990, N5991, N5992, N5993, N5994, N5995, N5996, N5997, N5998, N5999, N6000, N6001, N6002, N6003, N6004, N6005, N6006, N6007, N6008, N6009, N6010, N6011, N6012, N6013, N6014, N6015, N6016, N6017, N6018, N6019, N6020, N6021, N6022, N6023, N6024, N6025, N6026, N6027, N6028, N6029, N6030, N6031, N6032, N6033, N6034, N6035, N6036, N6037, N6038, N6039, N6040, N6041 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5913)? mhpmcounter_q[1023:960] : 1'b0;
  assign N126 = N5912;
  assign { N6203, N6202, N6201, N6200, N6199, N6198, N6197, N6196, N6195, N6194, N6193, N6192, N6191, N6190, N6189, N6188, N6187, N6186, N6185, N6184, N6183, N6182, N6181, N6180, N6179, N6178, N6177, N6176, N6175, N6174, N6173, N6172 } = (N127)? { N6140, N6141, N6142, N6143, N6144, N6145, N6146, N6147, N6148, N6149, N6150, N6151, N6152, N6153, N6154, N6155, N6156, N6157, N6158, N6159, N6160, N6161, N6162, N6163, N6164, N6165, N6166, N6167, N6168, N6169, N6170, N6171 } : 
                                                                                                                                                                                                                                              (N128)? { N6105, N6104, N6103, N6102, N6101, N6100, N6099, N6098, N6097, N6096, N6095, N6094, N6093, N6092, N6091, N6090, N6089, N6088, N6087, N6086, N6085, N6084, N6083, N6082, N6081, N6080, N6079, N6078, N6077, N6076, N6075, N6074 } : 1'b0;
  assign N127 = mhpmcounterh_we[16];
  assign N128 = N6139;
  assign mhpmcounter_d[1023:960] = (N129)? { N6105, N6104, N6103, N6102, N6101, N6100, N6099, N6098, N6097, N6096, N6095, N6094, N6093, N6092, N6091, N6090, N6089, N6088, N6087, N6086, N6085, N6084, N6083, N6082, N6081, N6080, N6079, N6078, N6077, N6076, N6075, N6074, N6107, N6108, N6109, N6110, N6111, N6112, N6113, N6114, N6115, N6116, N6117, N6118, N6119, N6120, N6121, N6122, N6123, N6124, N6125, N6126, N6127, N6128, N6129, N6130, N6131, N6132, N6133, N6134, N6135, N6136, N6137, N6138 } : 
                                   (N130)? { N6203, N6202, N6201, N6200, N6199, N6198, N6197, N6196, N6195, N6194, N6193, N6192, N6191, N6190, N6189, N6188, N6187, N6186, N6185, N6184, N6183, N6182, N6181, N6180, N6179, N6178, N6177, N6176, N6175, N6174, N6173, N6172, N6073, N6072, N6071, N6070, N6069, N6068, N6067, N6066, N6065, N6064, N6063, N6062, N6061, N6060, N6059, N6058, N6057, N6056, N6055, N6054, N6053, N6052, N6051, N6050, N6049, N6048, N6047, N6046, N6045, N6044, N6043, N6042 } : 1'b0;
  assign N129 = mhpmcounter_we[16];
  assign N130 = N6106;
  assign { N6397, N6396, N6395, N6394, N6393, N6392, N6391, N6390, N6389, N6388, N6387, N6386, N6385, N6384, N6383, N6382, N6381, N6380, N6379, N6378, N6377, N6376, N6375, N6374, N6373, N6372, N6371, N6370, N6369, N6368, N6367, N6366, N6365, N6364, N6363, N6362, N6361, N6360, N6359, N6358, N6357, N6356, N6355, N6354, N6353, N6352, N6351, N6350, N6349, N6348, N6347, N6346, N6345, N6344, N6343, N6342, N6341, N6340, N6339, N6338, N6337, N6336, N6335, N6334 } = (N131)? { N6270, N6271, N6272, N6273, N6274, N6275, N6276, N6277, N6278, N6279, N6280, N6281, N6282, N6283, N6284, N6285, N6286, N6287, N6288, N6289, N6290, N6291, N6292, N6293, N6294, N6295, N6296, N6297, N6298, N6299, N6300, N6301, N6302, N6303, N6304, N6305, N6306, N6307, N6308, N6309, N6310, N6311, N6312, N6313, N6314, N6315, N6316, N6317, N6318, N6319, N6320, N6321, N6322, N6323, N6324, N6325, N6326, N6327, N6328, N6329, N6330, N6331, N6332, N6333 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6205)? mhpmcounter_q[959:896] : 1'b0;
  assign N131 = N6204;
  assign { N6495, N6494, N6493, N6492, N6491, N6490, N6489, N6488, N6487, N6486, N6485, N6484, N6483, N6482, N6481, N6480, N6479, N6478, N6477, N6476, N6475, N6474, N6473, N6472, N6471, N6470, N6469, N6468, N6467, N6466, N6465, N6464 } = (N132)? { N6432, N6433, N6434, N6435, N6436, N6437, N6438, N6439, N6440, N6441, N6442, N6443, N6444, N6445, N6446, N6447, N6448, N6449, N6450, N6451, N6452, N6453, N6454, N6455, N6456, N6457, N6458, N6459, N6460, N6461, N6462, N6463 } : 
                                                                                                                                                                                                                                              (N133)? { N6397, N6396, N6395, N6394, N6393, N6392, N6391, N6390, N6389, N6388, N6387, N6386, N6385, N6384, N6383, N6382, N6381, N6380, N6379, N6378, N6377, N6376, N6375, N6374, N6373, N6372, N6371, N6370, N6369, N6368, N6367, N6366 } : 1'b0;
  assign N132 = mhpmcounterh_we[17];
  assign N133 = N6431;
  assign mhpmcounter_d[959:896] = (N134)? { N6397, N6396, N6395, N6394, N6393, N6392, N6391, N6390, N6389, N6388, N6387, N6386, N6385, N6384, N6383, N6382, N6381, N6380, N6379, N6378, N6377, N6376, N6375, N6374, N6373, N6372, N6371, N6370, N6369, N6368, N6367, N6366, N6399, N6400, N6401, N6402, N6403, N6404, N6405, N6406, N6407, N6408, N6409, N6410, N6411, N6412, N6413, N6414, N6415, N6416, N6417, N6418, N6419, N6420, N6421, N6422, N6423, N6424, N6425, N6426, N6427, N6428, N6429, N6430 } : 
                                  (N135)? { N6495, N6494, N6493, N6492, N6491, N6490, N6489, N6488, N6487, N6486, N6485, N6484, N6483, N6482, N6481, N6480, N6479, N6478, N6477, N6476, N6475, N6474, N6473, N6472, N6471, N6470, N6469, N6468, N6467, N6466, N6465, N6464, N6365, N6364, N6363, N6362, N6361, N6360, N6359, N6358, N6357, N6356, N6355, N6354, N6353, N6352, N6351, N6350, N6349, N6348, N6347, N6346, N6345, N6344, N6343, N6342, N6341, N6340, N6339, N6338, N6337, N6336, N6335, N6334 } : 1'b0;
  assign N134 = mhpmcounter_we[17];
  assign N135 = N6398;
  assign { N6689, N6688, N6687, N6686, N6685, N6684, N6683, N6682, N6681, N6680, N6679, N6678, N6677, N6676, N6675, N6674, N6673, N6672, N6671, N6670, N6669, N6668, N6667, N6666, N6665, N6664, N6663, N6662, N6661, N6660, N6659, N6658, N6657, N6656, N6655, N6654, N6653, N6652, N6651, N6650, N6649, N6648, N6647, N6646, N6645, N6644, N6643, N6642, N6641, N6640, N6639, N6638, N6637, N6636, N6635, N6634, N6633, N6632, N6631, N6630, N6629, N6628, N6627, N6626 } = (N136)? { N6562, N6563, N6564, N6565, N6566, N6567, N6568, N6569, N6570, N6571, N6572, N6573, N6574, N6575, N6576, N6577, N6578, N6579, N6580, N6581, N6582, N6583, N6584, N6585, N6586, N6587, N6588, N6589, N6590, N6591, N6592, N6593, N6594, N6595, N6596, N6597, N6598, N6599, N6600, N6601, N6602, N6603, N6604, N6605, N6606, N6607, N6608, N6609, N6610, N6611, N6612, N6613, N6614, N6615, N6616, N6617, N6618, N6619, N6620, N6621, N6622, N6623, N6624, N6625 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6497)? mhpmcounter_q[895:832] : 1'b0;
  assign N136 = N6496;
  assign { N6787, N6786, N6785, N6784, N6783, N6782, N6781, N6780, N6779, N6778, N6777, N6776, N6775, N6774, N6773, N6772, N6771, N6770, N6769, N6768, N6767, N6766, N6765, N6764, N6763, N6762, N6761, N6760, N6759, N6758, N6757, N6756 } = (N137)? { N6724, N6725, N6726, N6727, N6728, N6729, N6730, N6731, N6732, N6733, N6734, N6735, N6736, N6737, N6738, N6739, N6740, N6741, N6742, N6743, N6744, N6745, N6746, N6747, N6748, N6749, N6750, N6751, N6752, N6753, N6754, N6755 } : 
                                                                                                                                                                                                                                              (N138)? { N6689, N6688, N6687, N6686, N6685, N6684, N6683, N6682, N6681, N6680, N6679, N6678, N6677, N6676, N6675, N6674, N6673, N6672, N6671, N6670, N6669, N6668, N6667, N6666, N6665, N6664, N6663, N6662, N6661, N6660, N6659, N6658 } : 1'b0;
  assign N137 = mhpmcounterh_we[18];
  assign N138 = N6723;
  assign mhpmcounter_d[895:832] = (N139)? { N6689, N6688, N6687, N6686, N6685, N6684, N6683, N6682, N6681, N6680, N6679, N6678, N6677, N6676, N6675, N6674, N6673, N6672, N6671, N6670, N6669, N6668, N6667, N6666, N6665, N6664, N6663, N6662, N6661, N6660, N6659, N6658, N6691, N6692, N6693, N6694, N6695, N6696, N6697, N6698, N6699, N6700, N6701, N6702, N6703, N6704, N6705, N6706, N6707, N6708, N6709, N6710, N6711, N6712, N6713, N6714, N6715, N6716, N6717, N6718, N6719, N6720, N6721, N6722 } : 
                                  (N140)? { N6787, N6786, N6785, N6784, N6783, N6782, N6781, N6780, N6779, N6778, N6777, N6776, N6775, N6774, N6773, N6772, N6771, N6770, N6769, N6768, N6767, N6766, N6765, N6764, N6763, N6762, N6761, N6760, N6759, N6758, N6757, N6756, N6657, N6656, N6655, N6654, N6653, N6652, N6651, N6650, N6649, N6648, N6647, N6646, N6645, N6644, N6643, N6642, N6641, N6640, N6639, N6638, N6637, N6636, N6635, N6634, N6633, N6632, N6631, N6630, N6629, N6628, N6627, N6626 } : 1'b0;
  assign N139 = mhpmcounter_we[18];
  assign N140 = N6690;
  assign { N6981, N6980, N6979, N6978, N6977, N6976, N6975, N6974, N6973, N6972, N6971, N6970, N6969, N6968, N6967, N6966, N6965, N6964, N6963, N6962, N6961, N6960, N6959, N6958, N6957, N6956, N6955, N6954, N6953, N6952, N6951, N6950, N6949, N6948, N6947, N6946, N6945, N6944, N6943, N6942, N6941, N6940, N6939, N6938, N6937, N6936, N6935, N6934, N6933, N6932, N6931, N6930, N6929, N6928, N6927, N6926, N6925, N6924, N6923, N6922, N6921, N6920, N6919, N6918 } = (N141)? { N6854, N6855, N6856, N6857, N6858, N6859, N6860, N6861, N6862, N6863, N6864, N6865, N6866, N6867, N6868, N6869, N6870, N6871, N6872, N6873, N6874, N6875, N6876, N6877, N6878, N6879, N6880, N6881, N6882, N6883, N6884, N6885, N6886, N6887, N6888, N6889, N6890, N6891, N6892, N6893, N6894, N6895, N6896, N6897, N6898, N6899, N6900, N6901, N6902, N6903, N6904, N6905, N6906, N6907, N6908, N6909, N6910, N6911, N6912, N6913, N6914, N6915, N6916, N6917 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6789)? mhpmcounter_q[831:768] : 1'b0;
  assign N141 = N6788;
  assign { N7079, N7078, N7077, N7076, N7075, N7074, N7073, N7072, N7071, N7070, N7069, N7068, N7067, N7066, N7065, N7064, N7063, N7062, N7061, N7060, N7059, N7058, N7057, N7056, N7055, N7054, N7053, N7052, N7051, N7050, N7049, N7048 } = (N142)? { N7016, N7017, N7018, N7019, N7020, N7021, N7022, N7023, N7024, N7025, N7026, N7027, N7028, N7029, N7030, N7031, N7032, N7033, N7034, N7035, N7036, N7037, N7038, N7039, N7040, N7041, N7042, N7043, N7044, N7045, N7046, N7047 } : 
                                                                                                                                                                                                                                              (N143)? { N6981, N6980, N6979, N6978, N6977, N6976, N6975, N6974, N6973, N6972, N6971, N6970, N6969, N6968, N6967, N6966, N6965, N6964, N6963, N6962, N6961, N6960, N6959, N6958, N6957, N6956, N6955, N6954, N6953, N6952, N6951, N6950 } : 1'b0;
  assign N142 = mhpmcounterh_we[19];
  assign N143 = N7015;
  assign mhpmcounter_d[831:768] = (N144)? { N6981, N6980, N6979, N6978, N6977, N6976, N6975, N6974, N6973, N6972, N6971, N6970, N6969, N6968, N6967, N6966, N6965, N6964, N6963, N6962, N6961, N6960, N6959, N6958, N6957, N6956, N6955, N6954, N6953, N6952, N6951, N6950, N6983, N6984, N6985, N6986, N6987, N6988, N6989, N6990, N6991, N6992, N6993, N6994, N6995, N6996, N6997, N6998, N6999, N7000, N7001, N7002, N7003, N7004, N7005, N7006, N7007, N7008, N7009, N7010, N7011, N7012, N7013, N7014 } : 
                                  (N145)? { N7079, N7078, N7077, N7076, N7075, N7074, N7073, N7072, N7071, N7070, N7069, N7068, N7067, N7066, N7065, N7064, N7063, N7062, N7061, N7060, N7059, N7058, N7057, N7056, N7055, N7054, N7053, N7052, N7051, N7050, N7049, N7048, N6949, N6948, N6947, N6946, N6945, N6944, N6943, N6942, N6941, N6940, N6939, N6938, N6937, N6936, N6935, N6934, N6933, N6932, N6931, N6930, N6929, N6928, N6927, N6926, N6925, N6924, N6923, N6922, N6921, N6920, N6919, N6918 } : 1'b0;
  assign N144 = mhpmcounter_we[19];
  assign N145 = N6982;
  assign { N7273, N7272, N7271, N7270, N7269, N7268, N7267, N7266, N7265, N7264, N7263, N7262, N7261, N7260, N7259, N7258, N7257, N7256, N7255, N7254, N7253, N7252, N7251, N7250, N7249, N7248, N7247, N7246, N7245, N7244, N7243, N7242, N7241, N7240, N7239, N7238, N7237, N7236, N7235, N7234, N7233, N7232, N7231, N7230, N7229, N7228, N7227, N7226, N7225, N7224, N7223, N7222, N7221, N7220, N7219, N7218, N7217, N7216, N7215, N7214, N7213, N7212, N7211, N7210 } = (N146)? { N7146, N7147, N7148, N7149, N7150, N7151, N7152, N7153, N7154, N7155, N7156, N7157, N7158, N7159, N7160, N7161, N7162, N7163, N7164, N7165, N7166, N7167, N7168, N7169, N7170, N7171, N7172, N7173, N7174, N7175, N7176, N7177, N7178, N7179, N7180, N7181, N7182, N7183, N7184, N7185, N7186, N7187, N7188, N7189, N7190, N7191, N7192, N7193, N7194, N7195, N7196, N7197, N7198, N7199, N7200, N7201, N7202, N7203, N7204, N7205, N7206, N7207, N7208, N7209 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N7081)? mhpmcounter_q[767:704] : 1'b0;
  assign N146 = N7080;
  assign { N7371, N7370, N7369, N7368, N7367, N7366, N7365, N7364, N7363, N7362, N7361, N7360, N7359, N7358, N7357, N7356, N7355, N7354, N7353, N7352, N7351, N7350, N7349, N7348, N7347, N7346, N7345, N7344, N7343, N7342, N7341, N7340 } = (N147)? { N7308, N7309, N7310, N7311, N7312, N7313, N7314, N7315, N7316, N7317, N7318, N7319, N7320, N7321, N7322, N7323, N7324, N7325, N7326, N7327, N7328, N7329, N7330, N7331, N7332, N7333, N7334, N7335, N7336, N7337, N7338, N7339 } : 
                                                                                                                                                                                                                                              (N148)? { N7273, N7272, N7271, N7270, N7269, N7268, N7267, N7266, N7265, N7264, N7263, N7262, N7261, N7260, N7259, N7258, N7257, N7256, N7255, N7254, N7253, N7252, N7251, N7250, N7249, N7248, N7247, N7246, N7245, N7244, N7243, N7242 } : 1'b0;
  assign N147 = mhpmcounterh_we[20];
  assign N148 = N7307;
  assign mhpmcounter_d[767:704] = (N149)? { N7273, N7272, N7271, N7270, N7269, N7268, N7267, N7266, N7265, N7264, N7263, N7262, N7261, N7260, N7259, N7258, N7257, N7256, N7255, N7254, N7253, N7252, N7251, N7250, N7249, N7248, N7247, N7246, N7245, N7244, N7243, N7242, N7275, N7276, N7277, N7278, N7279, N7280, N7281, N7282, N7283, N7284, N7285, N7286, N7287, N7288, N7289, N7290, N7291, N7292, N7293, N7294, N7295, N7296, N7297, N7298, N7299, N7300, N7301, N7302, N7303, N7304, N7305, N7306 } : 
                                  (N150)? { N7371, N7370, N7369, N7368, N7367, N7366, N7365, N7364, N7363, N7362, N7361, N7360, N7359, N7358, N7357, N7356, N7355, N7354, N7353, N7352, N7351, N7350, N7349, N7348, N7347, N7346, N7345, N7344, N7343, N7342, N7341, N7340, N7241, N7240, N7239, N7238, N7237, N7236, N7235, N7234, N7233, N7232, N7231, N7230, N7229, N7228, N7227, N7226, N7225, N7224, N7223, N7222, N7221, N7220, N7219, N7218, N7217, N7216, N7215, N7214, N7213, N7212, N7211, N7210 } : 1'b0;
  assign N149 = mhpmcounter_we[20];
  assign N150 = N7274;
  assign { N7565, N7564, N7563, N7562, N7561, N7560, N7559, N7558, N7557, N7556, N7555, N7554, N7553, N7552, N7551, N7550, N7549, N7548, N7547, N7546, N7545, N7544, N7543, N7542, N7541, N7540, N7539, N7538, N7537, N7536, N7535, N7534, N7533, N7532, N7531, N7530, N7529, N7528, N7527, N7526, N7525, N7524, N7523, N7522, N7521, N7520, N7519, N7518, N7517, N7516, N7515, N7514, N7513, N7512, N7511, N7510, N7509, N7508, N7507, N7506, N7505, N7504, N7503, N7502 } = (N151)? { N7438, N7439, N7440, N7441, N7442, N7443, N7444, N7445, N7446, N7447, N7448, N7449, N7450, N7451, N7452, N7453, N7454, N7455, N7456, N7457, N7458, N7459, N7460, N7461, N7462, N7463, N7464, N7465, N7466, N7467, N7468, N7469, N7470, N7471, N7472, N7473, N7474, N7475, N7476, N7477, N7478, N7479, N7480, N7481, N7482, N7483, N7484, N7485, N7486, N7487, N7488, N7489, N7490, N7491, N7492, N7493, N7494, N7495, N7496, N7497, N7498, N7499, N7500, N7501 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N7373)? mhpmcounter_q[703:640] : 1'b0;
  assign N151 = N7372;
  assign { N7663, N7662, N7661, N7660, N7659, N7658, N7657, N7656, N7655, N7654, N7653, N7652, N7651, N7650, N7649, N7648, N7647, N7646, N7645, N7644, N7643, N7642, N7641, N7640, N7639, N7638, N7637, N7636, N7635, N7634, N7633, N7632 } = (N152)? { N7600, N7601, N7602, N7603, N7604, N7605, N7606, N7607, N7608, N7609, N7610, N7611, N7612, N7613, N7614, N7615, N7616, N7617, N7618, N7619, N7620, N7621, N7622, N7623, N7624, N7625, N7626, N7627, N7628, N7629, N7630, N7631 } : 
                                                                                                                                                                                                                                              (N153)? { N7565, N7564, N7563, N7562, N7561, N7560, N7559, N7558, N7557, N7556, N7555, N7554, N7553, N7552, N7551, N7550, N7549, N7548, N7547, N7546, N7545, N7544, N7543, N7542, N7541, N7540, N7539, N7538, N7537, N7536, N7535, N7534 } : 1'b0;
  assign N152 = mhpmcounterh_we[21];
  assign N153 = N7599;
  assign mhpmcounter_d[703:640] = (N154)? { N7565, N7564, N7563, N7562, N7561, N7560, N7559, N7558, N7557, N7556, N7555, N7554, N7553, N7552, N7551, N7550, N7549, N7548, N7547, N7546, N7545, N7544, N7543, N7542, N7541, N7540, N7539, N7538, N7537, N7536, N7535, N7534, N7567, N7568, N7569, N7570, N7571, N7572, N7573, N7574, N7575, N7576, N7577, N7578, N7579, N7580, N7581, N7582, N7583, N7584, N7585, N7586, N7587, N7588, N7589, N7590, N7591, N7592, N7593, N7594, N7595, N7596, N7597, N7598 } : 
                                  (N155)? { N7663, N7662, N7661, N7660, N7659, N7658, N7657, N7656, N7655, N7654, N7653, N7652, N7651, N7650, N7649, N7648, N7647, N7646, N7645, N7644, N7643, N7642, N7641, N7640, N7639, N7638, N7637, N7636, N7635, N7634, N7633, N7632, N7533, N7532, N7531, N7530, N7529, N7528, N7527, N7526, N7525, N7524, N7523, N7522, N7521, N7520, N7519, N7518, N7517, N7516, N7515, N7514, N7513, N7512, N7511, N7510, N7509, N7508, N7507, N7506, N7505, N7504, N7503, N7502 } : 1'b0;
  assign N154 = mhpmcounter_we[21];
  assign N155 = N7566;
  assign { N7857, N7856, N7855, N7854, N7853, N7852, N7851, N7850, N7849, N7848, N7847, N7846, N7845, N7844, N7843, N7842, N7841, N7840, N7839, N7838, N7837, N7836, N7835, N7834, N7833, N7832, N7831, N7830, N7829, N7828, N7827, N7826, N7825, N7824, N7823, N7822, N7821, N7820, N7819, N7818, N7817, N7816, N7815, N7814, N7813, N7812, N7811, N7810, N7809, N7808, N7807, N7806, N7805, N7804, N7803, N7802, N7801, N7800, N7799, N7798, N7797, N7796, N7795, N7794 } = (N156)? { N7730, N7731, N7732, N7733, N7734, N7735, N7736, N7737, N7738, N7739, N7740, N7741, N7742, N7743, N7744, N7745, N7746, N7747, N7748, N7749, N7750, N7751, N7752, N7753, N7754, N7755, N7756, N7757, N7758, N7759, N7760, N7761, N7762, N7763, N7764, N7765, N7766, N7767, N7768, N7769, N7770, N7771, N7772, N7773, N7774, N7775, N7776, N7777, N7778, N7779, N7780, N7781, N7782, N7783, N7784, N7785, N7786, N7787, N7788, N7789, N7790, N7791, N7792, N7793 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N7665)? mhpmcounter_q[639:576] : 1'b0;
  assign N156 = N7664;
  assign { N7955, N7954, N7953, N7952, N7951, N7950, N7949, N7948, N7947, N7946, N7945, N7944, N7943, N7942, N7941, N7940, N7939, N7938, N7937, N7936, N7935, N7934, N7933, N7932, N7931, N7930, N7929, N7928, N7927, N7926, N7925, N7924 } = (N157)? { N7892, N7893, N7894, N7895, N7896, N7897, N7898, N7899, N7900, N7901, N7902, N7903, N7904, N7905, N7906, N7907, N7908, N7909, N7910, N7911, N7912, N7913, N7914, N7915, N7916, N7917, N7918, N7919, N7920, N7921, N7922, N7923 } : 
                                                                                                                                                                                                                                              (N158)? { N7857, N7856, N7855, N7854, N7853, N7852, N7851, N7850, N7849, N7848, N7847, N7846, N7845, N7844, N7843, N7842, N7841, N7840, N7839, N7838, N7837, N7836, N7835, N7834, N7833, N7832, N7831, N7830, N7829, N7828, N7827, N7826 } : 1'b0;
  assign N157 = mhpmcounterh_we[22];
  assign N158 = N7891;
  assign mhpmcounter_d[639:576] = (N159)? { N7857, N7856, N7855, N7854, N7853, N7852, N7851, N7850, N7849, N7848, N7847, N7846, N7845, N7844, N7843, N7842, N7841, N7840, N7839, N7838, N7837, N7836, N7835, N7834, N7833, N7832, N7831, N7830, N7829, N7828, N7827, N7826, N7859, N7860, N7861, N7862, N7863, N7864, N7865, N7866, N7867, N7868, N7869, N7870, N7871, N7872, N7873, N7874, N7875, N7876, N7877, N7878, N7879, N7880, N7881, N7882, N7883, N7884, N7885, N7886, N7887, N7888, N7889, N7890 } : 
                                  (N160)? { N7955, N7954, N7953, N7952, N7951, N7950, N7949, N7948, N7947, N7946, N7945, N7944, N7943, N7942, N7941, N7940, N7939, N7938, N7937, N7936, N7935, N7934, N7933, N7932, N7931, N7930, N7929, N7928, N7927, N7926, N7925, N7924, N7825, N7824, N7823, N7822, N7821, N7820, N7819, N7818, N7817, N7816, N7815, N7814, N7813, N7812, N7811, N7810, N7809, N7808, N7807, N7806, N7805, N7804, N7803, N7802, N7801, N7800, N7799, N7798, N7797, N7796, N7795, N7794 } : 1'b0;
  assign N159 = mhpmcounter_we[22];
  assign N160 = N7858;
  assign { N8149, N8148, N8147, N8146, N8145, N8144, N8143, N8142, N8141, N8140, N8139, N8138, N8137, N8136, N8135, N8134, N8133, N8132, N8131, N8130, N8129, N8128, N8127, N8126, N8125, N8124, N8123, N8122, N8121, N8120, N8119, N8118, N8117, N8116, N8115, N8114, N8113, N8112, N8111, N8110, N8109, N8108, N8107, N8106, N8105, N8104, N8103, N8102, N8101, N8100, N8099, N8098, N8097, N8096, N8095, N8094, N8093, N8092, N8091, N8090, N8089, N8088, N8087, N8086 } = (N161)? { N8022, N8023, N8024, N8025, N8026, N8027, N8028, N8029, N8030, N8031, N8032, N8033, N8034, N8035, N8036, N8037, N8038, N8039, N8040, N8041, N8042, N8043, N8044, N8045, N8046, N8047, N8048, N8049, N8050, N8051, N8052, N8053, N8054, N8055, N8056, N8057, N8058, N8059, N8060, N8061, N8062, N8063, N8064, N8065, N8066, N8067, N8068, N8069, N8070, N8071, N8072, N8073, N8074, N8075, N8076, N8077, N8078, N8079, N8080, N8081, N8082, N8083, N8084, N8085 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N7957)? mhpmcounter_q[575:512] : 1'b0;
  assign N161 = N7956;
  assign { N8247, N8246, N8245, N8244, N8243, N8242, N8241, N8240, N8239, N8238, N8237, N8236, N8235, N8234, N8233, N8232, N8231, N8230, N8229, N8228, N8227, N8226, N8225, N8224, N8223, N8222, N8221, N8220, N8219, N8218, N8217, N8216 } = (N162)? { N8184, N8185, N8186, N8187, N8188, N8189, N8190, N8191, N8192, N8193, N8194, N8195, N8196, N8197, N8198, N8199, N8200, N8201, N8202, N8203, N8204, N8205, N8206, N8207, N8208, N8209, N8210, N8211, N8212, N8213, N8214, N8215 } : 
                                                                                                                                                                                                                                              (N163)? { N8149, N8148, N8147, N8146, N8145, N8144, N8143, N8142, N8141, N8140, N8139, N8138, N8137, N8136, N8135, N8134, N8133, N8132, N8131, N8130, N8129, N8128, N8127, N8126, N8125, N8124, N8123, N8122, N8121, N8120, N8119, N8118 } : 1'b0;
  assign N162 = mhpmcounterh_we[23];
  assign N163 = N8183;
  assign mhpmcounter_d[575:512] = (N164)? { N8149, N8148, N8147, N8146, N8145, N8144, N8143, N8142, N8141, N8140, N8139, N8138, N8137, N8136, N8135, N8134, N8133, N8132, N8131, N8130, N8129, N8128, N8127, N8126, N8125, N8124, N8123, N8122, N8121, N8120, N8119, N8118, N8151, N8152, N8153, N8154, N8155, N8156, N8157, N8158, N8159, N8160, N8161, N8162, N8163, N8164, N8165, N8166, N8167, N8168, N8169, N8170, N8171, N8172, N8173, N8174, N8175, N8176, N8177, N8178, N8179, N8180, N8181, N8182 } : 
                                  (N165)? { N8247, N8246, N8245, N8244, N8243, N8242, N8241, N8240, N8239, N8238, N8237, N8236, N8235, N8234, N8233, N8232, N8231, N8230, N8229, N8228, N8227, N8226, N8225, N8224, N8223, N8222, N8221, N8220, N8219, N8218, N8217, N8216, N8117, N8116, N8115, N8114, N8113, N8112, N8111, N8110, N8109, N8108, N8107, N8106, N8105, N8104, N8103, N8102, N8101, N8100, N8099, N8098, N8097, N8096, N8095, N8094, N8093, N8092, N8091, N8090, N8089, N8088, N8087, N8086 } : 1'b0;
  assign N164 = mhpmcounter_we[23];
  assign N165 = N8150;
  assign { N8441, N8440, N8439, N8438, N8437, N8436, N8435, N8434, N8433, N8432, N8431, N8430, N8429, N8428, N8427, N8426, N8425, N8424, N8423, N8422, N8421, N8420, N8419, N8418, N8417, N8416, N8415, N8414, N8413, N8412, N8411, N8410, N8409, N8408, N8407, N8406, N8405, N8404, N8403, N8402, N8401, N8400, N8399, N8398, N8397, N8396, N8395, N8394, N8393, N8392, N8391, N8390, N8389, N8388, N8387, N8386, N8385, N8384, N8383, N8382, N8381, N8380, N8379, N8378 } = (N166)? { N8314, N8315, N8316, N8317, N8318, N8319, N8320, N8321, N8322, N8323, N8324, N8325, N8326, N8327, N8328, N8329, N8330, N8331, N8332, N8333, N8334, N8335, N8336, N8337, N8338, N8339, N8340, N8341, N8342, N8343, N8344, N8345, N8346, N8347, N8348, N8349, N8350, N8351, N8352, N8353, N8354, N8355, N8356, N8357, N8358, N8359, N8360, N8361, N8362, N8363, N8364, N8365, N8366, N8367, N8368, N8369, N8370, N8371, N8372, N8373, N8374, N8375, N8376, N8377 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N8249)? mhpmcounter_q[511:448] : 1'b0;
  assign N166 = N8248;
  assign { N8539, N8538, N8537, N8536, N8535, N8534, N8533, N8532, N8531, N8530, N8529, N8528, N8527, N8526, N8525, N8524, N8523, N8522, N8521, N8520, N8519, N8518, N8517, N8516, N8515, N8514, N8513, N8512, N8511, N8510, N8509, N8508 } = (N167)? { N8476, N8477, N8478, N8479, N8480, N8481, N8482, N8483, N8484, N8485, N8486, N8487, N8488, N8489, N8490, N8491, N8492, N8493, N8494, N8495, N8496, N8497, N8498, N8499, N8500, N8501, N8502, N8503, N8504, N8505, N8506, N8507 } : 
                                                                                                                                                                                                                                              (N168)? { N8441, N8440, N8439, N8438, N8437, N8436, N8435, N8434, N8433, N8432, N8431, N8430, N8429, N8428, N8427, N8426, N8425, N8424, N8423, N8422, N8421, N8420, N8419, N8418, N8417, N8416, N8415, N8414, N8413, N8412, N8411, N8410 } : 1'b0;
  assign N167 = mhpmcounterh_we[24];
  assign N168 = N8475;
  assign mhpmcounter_d[511:448] = (N169)? { N8441, N8440, N8439, N8438, N8437, N8436, N8435, N8434, N8433, N8432, N8431, N8430, N8429, N8428, N8427, N8426, N8425, N8424, N8423, N8422, N8421, N8420, N8419, N8418, N8417, N8416, N8415, N8414, N8413, N8412, N8411, N8410, N8443, N8444, N8445, N8446, N8447, N8448, N8449, N8450, N8451, N8452, N8453, N8454, N8455, N8456, N8457, N8458, N8459, N8460, N8461, N8462, N8463, N8464, N8465, N8466, N8467, N8468, N8469, N8470, N8471, N8472, N8473, N8474 } : 
                                  (N170)? { N8539, N8538, N8537, N8536, N8535, N8534, N8533, N8532, N8531, N8530, N8529, N8528, N8527, N8526, N8525, N8524, N8523, N8522, N8521, N8520, N8519, N8518, N8517, N8516, N8515, N8514, N8513, N8512, N8511, N8510, N8509, N8508, N8409, N8408, N8407, N8406, N8405, N8404, N8403, N8402, N8401, N8400, N8399, N8398, N8397, N8396, N8395, N8394, N8393, N8392, N8391, N8390, N8389, N8388, N8387, N8386, N8385, N8384, N8383, N8382, N8381, N8380, N8379, N8378 } : 1'b0;
  assign N169 = mhpmcounter_we[24];
  assign N170 = N8442;
  assign { N8733, N8732, N8731, N8730, N8729, N8728, N8727, N8726, N8725, N8724, N8723, N8722, N8721, N8720, N8719, N8718, N8717, N8716, N8715, N8714, N8713, N8712, N8711, N8710, N8709, N8708, N8707, N8706, N8705, N8704, N8703, N8702, N8701, N8700, N8699, N8698, N8697, N8696, N8695, N8694, N8693, N8692, N8691, N8690, N8689, N8688, N8687, N8686, N8685, N8684, N8683, N8682, N8681, N8680, N8679, N8678, N8677, N8676, N8675, N8674, N8673, N8672, N8671, N8670 } = (N171)? { N8606, N8607, N8608, N8609, N8610, N8611, N8612, N8613, N8614, N8615, N8616, N8617, N8618, N8619, N8620, N8621, N8622, N8623, N8624, N8625, N8626, N8627, N8628, N8629, N8630, N8631, N8632, N8633, N8634, N8635, N8636, N8637, N8638, N8639, N8640, N8641, N8642, N8643, N8644, N8645, N8646, N8647, N8648, N8649, N8650, N8651, N8652, N8653, N8654, N8655, N8656, N8657, N8658, N8659, N8660, N8661, N8662, N8663, N8664, N8665, N8666, N8667, N8668, N8669 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N8541)? mhpmcounter_q[447:384] : 1'b0;
  assign N171 = N8540;
  assign { N8831, N8830, N8829, N8828, N8827, N8826, N8825, N8824, N8823, N8822, N8821, N8820, N8819, N8818, N8817, N8816, N8815, N8814, N8813, N8812, N8811, N8810, N8809, N8808, N8807, N8806, N8805, N8804, N8803, N8802, N8801, N8800 } = (N172)? { N8768, N8769, N8770, N8771, N8772, N8773, N8774, N8775, N8776, N8777, N8778, N8779, N8780, N8781, N8782, N8783, N8784, N8785, N8786, N8787, N8788, N8789, N8790, N8791, N8792, N8793, N8794, N8795, N8796, N8797, N8798, N8799 } : 
                                                                                                                                                                                                                                              (N173)? { N8733, N8732, N8731, N8730, N8729, N8728, N8727, N8726, N8725, N8724, N8723, N8722, N8721, N8720, N8719, N8718, N8717, N8716, N8715, N8714, N8713, N8712, N8711, N8710, N8709, N8708, N8707, N8706, N8705, N8704, N8703, N8702 } : 1'b0;
  assign N172 = mhpmcounterh_we[25];
  assign N173 = N8767;
  assign mhpmcounter_d[447:384] = (N174)? { N8733, N8732, N8731, N8730, N8729, N8728, N8727, N8726, N8725, N8724, N8723, N8722, N8721, N8720, N8719, N8718, N8717, N8716, N8715, N8714, N8713, N8712, N8711, N8710, N8709, N8708, N8707, N8706, N8705, N8704, N8703, N8702, N8735, N8736, N8737, N8738, N8739, N8740, N8741, N8742, N8743, N8744, N8745, N8746, N8747, N8748, N8749, N8750, N8751, N8752, N8753, N8754, N8755, N8756, N8757, N8758, N8759, N8760, N8761, N8762, N8763, N8764, N8765, N8766 } : 
                                  (N175)? { N8831, N8830, N8829, N8828, N8827, N8826, N8825, N8824, N8823, N8822, N8821, N8820, N8819, N8818, N8817, N8816, N8815, N8814, N8813, N8812, N8811, N8810, N8809, N8808, N8807, N8806, N8805, N8804, N8803, N8802, N8801, N8800, N8701, N8700, N8699, N8698, N8697, N8696, N8695, N8694, N8693, N8692, N8691, N8690, N8689, N8688, N8687, N8686, N8685, N8684, N8683, N8682, N8681, N8680, N8679, N8678, N8677, N8676, N8675, N8674, N8673, N8672, N8671, N8670 } : 1'b0;
  assign N174 = mhpmcounter_we[25];
  assign N175 = N8734;
  assign { N9025, N9024, N9023, N9022, N9021, N9020, N9019, N9018, N9017, N9016, N9015, N9014, N9013, N9012, N9011, N9010, N9009, N9008, N9007, N9006, N9005, N9004, N9003, N9002, N9001, N9000, N8999, N8998, N8997, N8996, N8995, N8994, N8993, N8992, N8991, N8990, N8989, N8988, N8987, N8986, N8985, N8984, N8983, N8982, N8981, N8980, N8979, N8978, N8977, N8976, N8975, N8974, N8973, N8972, N8971, N8970, N8969, N8968, N8967, N8966, N8965, N8964, N8963, N8962 } = (N176)? { N8898, N8899, N8900, N8901, N8902, N8903, N8904, N8905, N8906, N8907, N8908, N8909, N8910, N8911, N8912, N8913, N8914, N8915, N8916, N8917, N8918, N8919, N8920, N8921, N8922, N8923, N8924, N8925, N8926, N8927, N8928, N8929, N8930, N8931, N8932, N8933, N8934, N8935, N8936, N8937, N8938, N8939, N8940, N8941, N8942, N8943, N8944, N8945, N8946, N8947, N8948, N8949, N8950, N8951, N8952, N8953, N8954, N8955, N8956, N8957, N8958, N8959, N8960, N8961 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N8833)? mhpmcounter_q[383:320] : 1'b0;
  assign N176 = N8832;
  assign { N9123, N9122, N9121, N9120, N9119, N9118, N9117, N9116, N9115, N9114, N9113, N9112, N9111, N9110, N9109, N9108, N9107, N9106, N9105, N9104, N9103, N9102, N9101, N9100, N9099, N9098, N9097, N9096, N9095, N9094, N9093, N9092 } = (N177)? { N9060, N9061, N9062, N9063, N9064, N9065, N9066, N9067, N9068, N9069, N9070, N9071, N9072, N9073, N9074, N9075, N9076, N9077, N9078, N9079, N9080, N9081, N9082, N9083, N9084, N9085, N9086, N9087, N9088, N9089, N9090, N9091 } : 
                                                                                                                                                                                                                                              (N178)? { N9025, N9024, N9023, N9022, N9021, N9020, N9019, N9018, N9017, N9016, N9015, N9014, N9013, N9012, N9011, N9010, N9009, N9008, N9007, N9006, N9005, N9004, N9003, N9002, N9001, N9000, N8999, N8998, N8997, N8996, N8995, N8994 } : 1'b0;
  assign N177 = mhpmcounterh_we[26];
  assign N178 = N9059;
  assign mhpmcounter_d[383:320] = (N179)? { N9025, N9024, N9023, N9022, N9021, N9020, N9019, N9018, N9017, N9016, N9015, N9014, N9013, N9012, N9011, N9010, N9009, N9008, N9007, N9006, N9005, N9004, N9003, N9002, N9001, N9000, N8999, N8998, N8997, N8996, N8995, N8994, N9027, N9028, N9029, N9030, N9031, N9032, N9033, N9034, N9035, N9036, N9037, N9038, N9039, N9040, N9041, N9042, N9043, N9044, N9045, N9046, N9047, N9048, N9049, N9050, N9051, N9052, N9053, N9054, N9055, N9056, N9057, N9058 } : 
                                  (N180)? { N9123, N9122, N9121, N9120, N9119, N9118, N9117, N9116, N9115, N9114, N9113, N9112, N9111, N9110, N9109, N9108, N9107, N9106, N9105, N9104, N9103, N9102, N9101, N9100, N9099, N9098, N9097, N9096, N9095, N9094, N9093, N9092, N8993, N8992, N8991, N8990, N8989, N8988, N8987, N8986, N8985, N8984, N8983, N8982, N8981, N8980, N8979, N8978, N8977, N8976, N8975, N8974, N8973, N8972, N8971, N8970, N8969, N8968, N8967, N8966, N8965, N8964, N8963, N8962 } : 1'b0;
  assign N179 = mhpmcounter_we[26];
  assign N180 = N9026;
  assign { N9317, N9316, N9315, N9314, N9313, N9312, N9311, N9310, N9309, N9308, N9307, N9306, N9305, N9304, N9303, N9302, N9301, N9300, N9299, N9298, N9297, N9296, N9295, N9294, N9293, N9292, N9291, N9290, N9289, N9288, N9287, N9286, N9285, N9284, N9283, N9282, N9281, N9280, N9279, N9278, N9277, N9276, N9275, N9274, N9273, N9272, N9271, N9270, N9269, N9268, N9267, N9266, N9265, N9264, N9263, N9262, N9261, N9260, N9259, N9258, N9257, N9256, N9255, N9254 } = (N181)? { N9190, N9191, N9192, N9193, N9194, N9195, N9196, N9197, N9198, N9199, N9200, N9201, N9202, N9203, N9204, N9205, N9206, N9207, N9208, N9209, N9210, N9211, N9212, N9213, N9214, N9215, N9216, N9217, N9218, N9219, N9220, N9221, N9222, N9223, N9224, N9225, N9226, N9227, N9228, N9229, N9230, N9231, N9232, N9233, N9234, N9235, N9236, N9237, N9238, N9239, N9240, N9241, N9242, N9243, N9244, N9245, N9246, N9247, N9248, N9249, N9250, N9251, N9252, N9253 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N9125)? mhpmcounter_q[319:256] : 1'b0;
  assign N181 = N9124;
  assign { N9415, N9414, N9413, N9412, N9411, N9410, N9409, N9408, N9407, N9406, N9405, N9404, N9403, N9402, N9401, N9400, N9399, N9398, N9397, N9396, N9395, N9394, N9393, N9392, N9391, N9390, N9389, N9388, N9387, N9386, N9385, N9384 } = (N182)? { N9352, N9353, N9354, N9355, N9356, N9357, N9358, N9359, N9360, N9361, N9362, N9363, N9364, N9365, N9366, N9367, N9368, N9369, N9370, N9371, N9372, N9373, N9374, N9375, N9376, N9377, N9378, N9379, N9380, N9381, N9382, N9383 } : 
                                                                                                                                                                                                                                              (N183)? { N9317, N9316, N9315, N9314, N9313, N9312, N9311, N9310, N9309, N9308, N9307, N9306, N9305, N9304, N9303, N9302, N9301, N9300, N9299, N9298, N9297, N9296, N9295, N9294, N9293, N9292, N9291, N9290, N9289, N9288, N9287, N9286 } : 1'b0;
  assign N182 = mhpmcounterh_we[27];
  assign N183 = N9351;
  assign mhpmcounter_d[319:256] = (N184)? { N9317, N9316, N9315, N9314, N9313, N9312, N9311, N9310, N9309, N9308, N9307, N9306, N9305, N9304, N9303, N9302, N9301, N9300, N9299, N9298, N9297, N9296, N9295, N9294, N9293, N9292, N9291, N9290, N9289, N9288, N9287, N9286, N9319, N9320, N9321, N9322, N9323, N9324, N9325, N9326, N9327, N9328, N9329, N9330, N9331, N9332, N9333, N9334, N9335, N9336, N9337, N9338, N9339, N9340, N9341, N9342, N9343, N9344, N9345, N9346, N9347, N9348, N9349, N9350 } : 
                                  (N185)? { N9415, N9414, N9413, N9412, N9411, N9410, N9409, N9408, N9407, N9406, N9405, N9404, N9403, N9402, N9401, N9400, N9399, N9398, N9397, N9396, N9395, N9394, N9393, N9392, N9391, N9390, N9389, N9388, N9387, N9386, N9385, N9384, N9285, N9284, N9283, N9282, N9281, N9280, N9279, N9278, N9277, N9276, N9275, N9274, N9273, N9272, N9271, N9270, N9269, N9268, N9267, N9266, N9265, N9264, N9263, N9262, N9261, N9260, N9259, N9258, N9257, N9256, N9255, N9254 } : 1'b0;
  assign N184 = mhpmcounter_we[27];
  assign N185 = N9318;
  assign { N9609, N9608, N9607, N9606, N9605, N9604, N9603, N9602, N9601, N9600, N9599, N9598, N9597, N9596, N9595, N9594, N9593, N9592, N9591, N9590, N9589, N9588, N9587, N9586, N9585, N9584, N9583, N9582, N9581, N9580, N9579, N9578, N9577, N9576, N9575, N9574, N9573, N9572, N9571, N9570, N9569, N9568, N9567, N9566, N9565, N9564, N9563, N9562, N9561, N9560, N9559, N9558, N9557, N9556, N9555, N9554, N9553, N9552, N9551, N9550, N9549, N9548, N9547, N9546 } = (N186)? { N9482, N9483, N9484, N9485, N9486, N9487, N9488, N9489, N9490, N9491, N9492, N9493, N9494, N9495, N9496, N9497, N9498, N9499, N9500, N9501, N9502, N9503, N9504, N9505, N9506, N9507, N9508, N9509, N9510, N9511, N9512, N9513, N9514, N9515, N9516, N9517, N9518, N9519, N9520, N9521, N9522, N9523, N9524, N9525, N9526, N9527, N9528, N9529, N9530, N9531, N9532, N9533, N9534, N9535, N9536, N9537, N9538, N9539, N9540, N9541, N9542, N9543, N9544, N9545 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N9417)? mhpmcounter_q[255:192] : 1'b0;
  assign N186 = N9416;
  assign { N9707, N9706, N9705, N9704, N9703, N9702, N9701, N9700, N9699, N9698, N9697, N9696, N9695, N9694, N9693, N9692, N9691, N9690, N9689, N9688, N9687, N9686, N9685, N9684, N9683, N9682, N9681, N9680, N9679, N9678, N9677, N9676 } = (N187)? { N9644, N9645, N9646, N9647, N9648, N9649, N9650, N9651, N9652, N9653, N9654, N9655, N9656, N9657, N9658, N9659, N9660, N9661, N9662, N9663, N9664, N9665, N9666, N9667, N9668, N9669, N9670, N9671, N9672, N9673, N9674, N9675 } : 
                                                                                                                                                                                                                                              (N188)? { N9609, N9608, N9607, N9606, N9605, N9604, N9603, N9602, N9601, N9600, N9599, N9598, N9597, N9596, N9595, N9594, N9593, N9592, N9591, N9590, N9589, N9588, N9587, N9586, N9585, N9584, N9583, N9582, N9581, N9580, N9579, N9578 } : 1'b0;
  assign N187 = mhpmcounterh_we[28];
  assign N188 = N9643;
  assign mhpmcounter_d[255:192] = (N189)? { N9609, N9608, N9607, N9606, N9605, N9604, N9603, N9602, N9601, N9600, N9599, N9598, N9597, N9596, N9595, N9594, N9593, N9592, N9591, N9590, N9589, N9588, N9587, N9586, N9585, N9584, N9583, N9582, N9581, N9580, N9579, N9578, N9611, N9612, N9613, N9614, N9615, N9616, N9617, N9618, N9619, N9620, N9621, N9622, N9623, N9624, N9625, N9626, N9627, N9628, N9629, N9630, N9631, N9632, N9633, N9634, N9635, N9636, N9637, N9638, N9639, N9640, N9641, N9642 } : 
                                  (N190)? { N9707, N9706, N9705, N9704, N9703, N9702, N9701, N9700, N9699, N9698, N9697, N9696, N9695, N9694, N9693, N9692, N9691, N9690, N9689, N9688, N9687, N9686, N9685, N9684, N9683, N9682, N9681, N9680, N9679, N9678, N9677, N9676, N9577, N9576, N9575, N9574, N9573, N9572, N9571, N9570, N9569, N9568, N9567, N9566, N9565, N9564, N9563, N9562, N9561, N9560, N9559, N9558, N9557, N9556, N9555, N9554, N9553, N9552, N9551, N9550, N9549, N9548, N9547, N9546 } : 1'b0;
  assign N189 = mhpmcounter_we[28];
  assign N190 = N9610;
  assign { N9901, N9900, N9899, N9898, N9897, N9896, N9895, N9894, N9893, N9892, N9891, N9890, N9889, N9888, N9887, N9886, N9885, N9884, N9883, N9882, N9881, N9880, N9879, N9878, N9877, N9876, N9875, N9874, N9873, N9872, N9871, N9870, N9869, N9868, N9867, N9866, N9865, N9864, N9863, N9862, N9861, N9860, N9859, N9858, N9857, N9856, N9855, N9854, N9853, N9852, N9851, N9850, N9849, N9848, N9847, N9846, N9845, N9844, N9843, N9842, N9841, N9840, N9839, N9838 } = (N191)? { N9774, N9775, N9776, N9777, N9778, N9779, N9780, N9781, N9782, N9783, N9784, N9785, N9786, N9787, N9788, N9789, N9790, N9791, N9792, N9793, N9794, N9795, N9796, N9797, N9798, N9799, N9800, N9801, N9802, N9803, N9804, N9805, N9806, N9807, N9808, N9809, N9810, N9811, N9812, N9813, N9814, N9815, N9816, N9817, N9818, N9819, N9820, N9821, N9822, N9823, N9824, N9825, N9826, N9827, N9828, N9829, N9830, N9831, N9832, N9833, N9834, N9835, N9836, N9837 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N9709)? mhpmcounter_q[191:128] : 1'b0;
  assign N191 = N9708;
  assign { N9999, N9998, N9997, N9996, N9995, N9994, N9993, N9992, N9991, N9990, N9989, N9988, N9987, N9986, N9985, N9984, N9983, N9982, N9981, N9980, N9979, N9978, N9977, N9976, N9975, N9974, N9973, N9972, N9971, N9970, N9969, N9968 } = (N192)? { N9936, N9937, N9938, N9939, N9940, N9941, N9942, N9943, N9944, N9945, N9946, N9947, N9948, N9949, N9950, N9951, N9952, N9953, N9954, N9955, N9956, N9957, N9958, N9959, N9960, N9961, N9962, N9963, N9964, N9965, N9966, N9967 } : 
                                                                                                                                                                                                                                              (N193)? { N9901, N9900, N9899, N9898, N9897, N9896, N9895, N9894, N9893, N9892, N9891, N9890, N9889, N9888, N9887, N9886, N9885, N9884, N9883, N9882, N9881, N9880, N9879, N9878, N9877, N9876, N9875, N9874, N9873, N9872, N9871, N9870 } : 1'b0;
  assign N192 = mhpmcounterh_we[29];
  assign N193 = N9935;
  assign mhpmcounter_d[191:128] = (N194)? { N9901, N9900, N9899, N9898, N9897, N9896, N9895, N9894, N9893, N9892, N9891, N9890, N9889, N9888, N9887, N9886, N9885, N9884, N9883, N9882, N9881, N9880, N9879, N9878, N9877, N9876, N9875, N9874, N9873, N9872, N9871, N9870, N9903, N9904, N9905, N9906, N9907, N9908, N9909, N9910, N9911, N9912, N9913, N9914, N9915, N9916, N9917, N9918, N9919, N9920, N9921, N9922, N9923, N9924, N9925, N9926, N9927, N9928, N9929, N9930, N9931, N9932, N9933, N9934 } : 
                                  (N195)? { N9999, N9998, N9997, N9996, N9995, N9994, N9993, N9992, N9991, N9990, N9989, N9988, N9987, N9986, N9985, N9984, N9983, N9982, N9981, N9980, N9979, N9978, N9977, N9976, N9975, N9974, N9973, N9972, N9971, N9970, N9969, N9968, N9869, N9868, N9867, N9866, N9865, N9864, N9863, N9862, N9861, N9860, N9859, N9858, N9857, N9856, N9855, N9854, N9853, N9852, N9851, N9850, N9849, N9848, N9847, N9846, N9845, N9844, N9843, N9842, N9841, N9840, N9839, N9838 } : 1'b0;
  assign N194 = mhpmcounter_we[29];
  assign N195 = N9902;
  assign { N10193, N10192, N10191, N10190, N10189, N10188, N10187, N10186, N10185, N10184, N10183, N10182, N10181, N10180, N10179, N10178, N10177, N10176, N10175, N10174, N10173, N10172, N10171, N10170, N10169, N10168, N10167, N10166, N10165, N10164, N10163, N10162, N10161, N10160, N10159, N10158, N10157, N10156, N10155, N10154, N10153, N10152, N10151, N10150, N10149, N10148, N10147, N10146, N10145, N10144, N10143, N10142, N10141, N10140, N10139, N10138, N10137, N10136, N10135, N10134, N10133, N10132, N10131, N10130 } = (N196)? { N10066, N10067, N10068, N10069, N10070, N10071, N10072, N10073, N10074, N10075, N10076, N10077, N10078, N10079, N10080, N10081, N10082, N10083, N10084, N10085, N10086, N10087, N10088, N10089, N10090, N10091, N10092, N10093, N10094, N10095, N10096, N10097, N10098, N10099, N10100, N10101, N10102, N10103, N10104, N10105, N10106, N10107, N10108, N10109, N10110, N10111, N10112, N10113, N10114, N10115, N10116, N10117, N10118, N10119, N10120, N10121, N10122, N10123, N10124, N10125, N10126, N10127, N10128, N10129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N10001)? mhpmcounter_q[127:64] : 1'b0;
  assign N196 = N10000;
  assign { N10291, N10290, N10289, N10288, N10287, N10286, N10285, N10284, N10283, N10282, N10281, N10280, N10279, N10278, N10277, N10276, N10275, N10274, N10273, N10272, N10271, N10270, N10269, N10268, N10267, N10266, N10265, N10264, N10263, N10262, N10261, N10260 } = (N197)? { N10228, N10229, N10230, N10231, N10232, N10233, N10234, N10235, N10236, N10237, N10238, N10239, N10240, N10241, N10242, N10243, N10244, N10245, N10246, N10247, N10248, N10249, N10250, N10251, N10252, N10253, N10254, N10255, N10256, N10257, N10258, N10259 } : 
                                                                                                                                                                                                                                                                              (N198)? { N10193, N10192, N10191, N10190, N10189, N10188, N10187, N10186, N10185, N10184, N10183, N10182, N10181, N10180, N10179, N10178, N10177, N10176, N10175, N10174, N10173, N10172, N10171, N10170, N10169, N10168, N10167, N10166, N10165, N10164, N10163, N10162 } : 1'b0;
  assign N197 = mhpmcounterh_we[30];
  assign N198 = N10227;
  assign mhpmcounter_d[127:64] = (N199)? { N10193, N10192, N10191, N10190, N10189, N10188, N10187, N10186, N10185, N10184, N10183, N10182, N10181, N10180, N10179, N10178, N10177, N10176, N10175, N10174, N10173, N10172, N10171, N10170, N10169, N10168, N10167, N10166, N10165, N10164, N10163, N10162, N10195, N10196, N10197, N10198, N10199, N10200, N10201, N10202, N10203, N10204, N10205, N10206, N10207, N10208, N10209, N10210, N10211, N10212, N10213, N10214, N10215, N10216, N10217, N10218, N10219, N10220, N10221, N10222, N10223, N10224, N10225, N10226 } : 
                                 (N200)? { N10291, N10290, N10289, N10288, N10287, N10286, N10285, N10284, N10283, N10282, N10281, N10280, N10279, N10278, N10277, N10276, N10275, N10274, N10273, N10272, N10271, N10270, N10269, N10268, N10267, N10266, N10265, N10264, N10263, N10262, N10261, N10260, N10161, N10160, N10159, N10158, N10157, N10156, N10155, N10154, N10153, N10152, N10151, N10150, N10149, N10148, N10147, N10146, N10145, N10144, N10143, N10142, N10141, N10140, N10139, N10138, N10137, N10136, N10135, N10134, N10133, N10132, N10131, N10130 } : 1'b0;
  assign N199 = mhpmcounter_we[30];
  assign N200 = N10194;
  assign { N10485, N10484, N10483, N10482, N10481, N10480, N10479, N10478, N10477, N10476, N10475, N10474, N10473, N10472, N10471, N10470, N10469, N10468, N10467, N10466, N10465, N10464, N10463, N10462, N10461, N10460, N10459, N10458, N10457, N10456, N10455, N10454, N10453, N10452, N10451, N10450, N10449, N10448, N10447, N10446, N10445, N10444, N10443, N10442, N10441, N10440, N10439, N10438, N10437, N10436, N10435, N10434, N10433, N10432, N10431, N10430, N10429, N10428, N10427, N10426, N10425, N10424, N10423, N10422 } = (N201)? { N10358, N10359, N10360, N10361, N10362, N10363, N10364, N10365, N10366, N10367, N10368, N10369, N10370, N10371, N10372, N10373, N10374, N10375, N10376, N10377, N10378, N10379, N10380, N10381, N10382, N10383, N10384, N10385, N10386, N10387, N10388, N10389, N10390, N10391, N10392, N10393, N10394, N10395, N10396, N10397, N10398, N10399, N10400, N10401, N10402, N10403, N10404, N10405, N10406, N10407, N10408, N10409, N10410, N10411, N10412, N10413, N10414, N10415, N10416, N10417, N10418, N10419, N10420, N10421 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N10293)? mhpmcounter_q[63:0] : 1'b0;
  assign N201 = N10292;
  assign { N10583, N10582, N10581, N10580, N10579, N10578, N10577, N10576, N10575, N10574, N10573, N10572, N10571, N10570, N10569, N10568, N10567, N10566, N10565, N10564, N10563, N10562, N10561, N10560, N10559, N10558, N10557, N10556, N10555, N10554, N10553, N10552 } = (N202)? { N10520, N10521, N10522, N10523, N10524, N10525, N10526, N10527, N10528, N10529, N10530, N10531, N10532, N10533, N10534, N10535, N10536, N10537, N10538, N10539, N10540, N10541, N10542, N10543, N10544, N10545, N10546, N10547, N10548, N10549, N10550, N10551 } : 
                                                                                                                                                                                                                                                                              (N203)? { N10485, N10484, N10483, N10482, N10481, N10480, N10479, N10478, N10477, N10476, N10475, N10474, N10473, N10472, N10471, N10470, N10469, N10468, N10467, N10466, N10465, N10464, N10463, N10462, N10461, N10460, N10459, N10458, N10457, N10456, N10455, N10454 } : 1'b0;
  assign N202 = mhpmcounterh_we[31];
  assign N203 = N10519;
  assign mhpmcounter_d[63:0] = (N204)? { N10485, N10484, N10483, N10482, N10481, N10480, N10479, N10478, N10477, N10476, N10475, N10474, N10473, N10472, N10471, N10470, N10469, N10468, N10467, N10466, N10465, N10464, N10463, N10462, N10461, N10460, N10459, N10458, N10457, N10456, N10455, N10454, N10487, N10488, N10489, N10490, N10491, N10492, N10493, N10494, N10495, N10496, N10497, N10498, N10499, N10500, N10501, N10502, N10503, N10504, N10505, N10506, N10507, N10508, N10509, N10510, N10511, N10512, N10513, N10514, N10515, N10516, N10517, N10518 } : 
                               (N205)? { N10583, N10582, N10581, N10580, N10579, N10578, N10577, N10576, N10575, N10574, N10573, N10572, N10571, N10570, N10569, N10568, N10567, N10566, N10565, N10564, N10563, N10562, N10561, N10560, N10559, N10558, N10557, N10556, N10555, N10554, N10553, N10552, N10453, N10452, N10451, N10450, N10449, N10448, N10447, N10446, N10445, N10444, N10443, N10442, N10441, N10440, N10439, N10438, N10437, N10436, N10435, N10434, N10433, N10432, N10431, N10430, N10429, N10428, N10427, N10426, N10425, N10424, N10423, N10422 } : 1'b0;
  assign N204 = mhpmcounter_we[31];
  assign N205 = N10486;
  assign illegal_csr_write = N10617 & csr_wreq;
  assign illegal_csr_insn_o = N10671 | 1'b0;
  assign N10671 = illegal_csr | illegal_csr_write;
  assign N277 = ~N276;
  assign N279 = ~N278;
  assign N283 = ~N282;
  assign N284 = N409 | N277;
  assign N285 = N279 | N284;
  assign N286 = N411 | N285;
  assign N287 = N283 | N286;
  assign N288 = N413 | N287;
  assign N289 = N415 | N288;
  assign N290 = N421 | N289;
  assign N291 = N423 | N290;
  assign N292 = N427 | N291;
  assign N293 = N429 | N292;
  assign N294 = N440 | N293;
  assign N295 = N447 | N294;
  assign N296 = N449 | N295;
  assign N297 = N453 | N296;
  assign N298 = N458 | N297;
  assign N299 = N470 | N298;
  assign N300 = ~N299;
  assign N301 = N10634 | N10653;
  assign N302 = N10645 | N301;
  assign N303 = ~N302;
  assign N304 = ~csr_addr_i[0];
  assign N305 = ~csr_addr_i[1];
  assign N306 = N304 & N305;
  assign N307 = N304 & csr_addr_i[1];
  assign N308 = csr_addr_i[0] & N305;
  assign N309 = csr_addr_i[0] & csr_addr_i[1];
  assign N310 = ~csr_addr_i[2];
  assign N311 = N306 & N310;
  assign N312 = N306 & csr_addr_i[2];
  assign N313 = N308 & N310;
  assign N314 = N308 & csr_addr_i[2];
  assign N315 = N307 & N310;
  assign N316 = N307 & csr_addr_i[2];
  assign N317 = N309 & N310;
  assign N318 = N309 & csr_addr_i[2];
  assign N319 = ~csr_addr_i[3];
  assign N320 = N311 & N319;
  assign N321 = N311 & csr_addr_i[3];
  assign N322 = N313 & N319;
  assign N323 = N313 & csr_addr_i[3];
  assign N324 = N315 & N319;
  assign N325 = N315 & csr_addr_i[3];
  assign N326 = N317 & N319;
  assign N327 = N317 & csr_addr_i[3];
  assign N328 = N312 & N319;
  assign N329 = N312 & csr_addr_i[3];
  assign N330 = N314 & N319;
  assign N331 = N314 & csr_addr_i[3];
  assign N332 = N316 & N319;
  assign N333 = N316 & csr_addr_i[3];
  assign N334 = N318 & N319;
  assign N335 = N318 & csr_addr_i[3];
  assign N336 = ~csr_addr_i[4];
  assign N337 = N320 & N336;
  assign N338 = N320 & csr_addr_i[4];
  assign N339 = N322 & N336;
  assign N340 = N322 & csr_addr_i[4];
  assign N341 = N324 & N336;
  assign N342 = N324 & csr_addr_i[4];
  assign N343 = N326 & N336;
  assign N344 = N326 & csr_addr_i[4];
  assign N345 = N328 & N336;
  assign N346 = N328 & csr_addr_i[4];
  assign N347 = N330 & N336;
  assign N348 = N330 & csr_addr_i[4];
  assign N349 = N332 & N336;
  assign N350 = N332 & csr_addr_i[4];
  assign N351 = N334 & N336;
  assign N352 = N334 & csr_addr_i[4];
  assign N353 = N321 & N336;
  assign N354 = N321 & csr_addr_i[4];
  assign N355 = N323 & N336;
  assign N356 = N323 & csr_addr_i[4];
  assign N357 = N325 & N336;
  assign N358 = N325 & csr_addr_i[4];
  assign N359 = N327 & N336;
  assign N360 = N327 & csr_addr_i[4];
  assign N361 = N329 & N336;
  assign N362 = N329 & csr_addr_i[4];
  assign N363 = N331 & N336;
  assign N364 = N331 & csr_addr_i[4];
  assign N365 = N333 & N336;
  assign N366 = N333 & csr_addr_i[4];
  assign N367 = N335 & N336;
  assign N368 = N335 & csr_addr_i[4];
  assign N371 = N10672 | N10629;
  assign N10672 = N10622 | N10625;
  assign N372 = ~N371;
  assign N409 = ~N408;
  assign N411 = ~N410;
  assign N413 = ~N412;
  assign N415 = ~N414;
  assign N416 = ~csr_addr_i[6];
  assign N421 = ~N420;
  assign N423 = ~N422;
  assign N427 = ~N426;
  assign N429 = ~N428;
  assign N430 = ~csr_addr_i[10];
  assign N431 = ~csr_addr_i[4];
  assign N440 = ~N439;
  assign N447 = ~N446;
  assign N449 = ~N448;
  assign N453 = ~N452;
  assign N458 = ~N457;
  assign N470 = ~N469;
  assign N471 = N411 | N409;
  assign N472 = N413 | N471;
  assign N473 = N415 | N472;
  assign N474 = N421 | N473;
  assign N475 = N423 | N474;
  assign N476 = N427 | N475;
  assign N477 = N429 | N476;
  assign N478 = N440 | N477;
  assign N479 = N447 | N478;
  assign N480 = N449 | N479;
  assign N481 = N453 | N480;
  assign N482 = N458 | N481;
  assign N483 = N470 | N482;
  assign N484 = ~N483;
  assign N485 = ~csr_we_int;
  assign N622 = csr_we_int & N10630;
  assign N623 = ~N622;
  assign N720 = N10645 | N10634;
  assign N721 = ~N720;
  assign N1018 = N483;
  assign N1019 = csr_restore_mret_i | csr_save_cause_i;
  assign N1020 = csr_restore_dret_i | N1019;
  assign N1021 = ~N1020;
  assign N1022 = ~csr_save_if_i;
  assign N1055 = ~debug_csr_save_i;
  assign N1165 = ~csr_save_cause_i;
  assign N1167 = ~N1166;
  assign N1169 = ~N1168;
  assign N1171 = ~csr_op_i[1];
  assign N1172 = ~csr_op_i[0];
  assign N1174 = csr_wdata_i[31] | csr_rdata_o[31];
  assign N1175 = csr_wdata_i[30] | csr_rdata_o[30];
  assign N1176 = csr_wdata_i[29] | csr_rdata_o[29];
  assign N1177 = csr_wdata_i[28] | csr_rdata_o[28];
  assign N1178 = csr_wdata_i[27] | csr_rdata_o[27];
  assign N1179 = csr_wdata_i[26] | csr_rdata_o[26];
  assign N1180 = csr_wdata_i[25] | csr_rdata_o[25];
  assign N1181 = csr_wdata_i[24] | csr_rdata_o[24];
  assign N1182 = csr_wdata_i[23] | csr_rdata_o[23];
  assign N1183 = csr_wdata_i[22] | csr_rdata_o[22];
  assign N1184 = csr_wdata_i[21] | csr_rdata_o[21];
  assign N1185 = csr_wdata_i[20] | csr_rdata_o[20];
  assign N1186 = csr_wdata_i[19] | csr_rdata_o[19];
  assign N1187 = csr_wdata_i[18] | csr_rdata_o[18];
  assign N1188 = csr_wdata_i[17] | csr_rdata_o[17];
  assign N1189 = csr_wdata_i[16] | csr_rdata_o[16];
  assign N1190 = csr_wdata_i[15] | csr_rdata_o[15];
  assign N1191 = csr_wdata_i[14] | csr_rdata_o[14];
  assign N1192 = csr_wdata_i[13] | csr_rdata_o[13];
  assign N1193 = csr_wdata_i[12] | csr_rdata_o[12];
  assign N1194 = csr_wdata_i[11] | csr_rdata_o[11];
  assign N1195 = csr_wdata_i[10] | csr_rdata_o[10];
  assign N1196 = csr_wdata_i[9] | csr_rdata_o[9];
  assign N1197 = csr_wdata_i[8] | csr_rdata_o[8];
  assign N1198 = csr_wdata_i[7] | csr_rdata_o[7];
  assign N1199 = csr_wdata_i[6] | csr_rdata_o[6];
  assign N1200 = csr_wdata_i[5] | csr_rdata_o[5];
  assign N1201 = csr_wdata_i[4] | csr_rdata_o[4];
  assign N1202 = csr_wdata_i[3] | csr_rdata_o[3];
  assign N1203 = csr_wdata_i[2] | csr_rdata_o[2];
  assign N1204 = csr_wdata_i[1] | csr_rdata_o[1];
  assign N1205 = csr_wdata_i[0] | csr_rdata_o[0];
  assign N1206 = N10673 & csr_rdata_o[31];
  assign N10673 = ~csr_wdata_i[31];
  assign N1207 = N10674 & csr_rdata_o[30];
  assign N10674 = ~csr_wdata_i[30];
  assign N1208 = N10675 & csr_rdata_o[29];
  assign N10675 = ~csr_wdata_i[29];
  assign N1209 = N10676 & csr_rdata_o[28];
  assign N10676 = ~csr_wdata_i[28];
  assign N1210 = N10677 & csr_rdata_o[27];
  assign N10677 = ~csr_wdata_i[27];
  assign N1211 = N10678 & csr_rdata_o[26];
  assign N10678 = ~csr_wdata_i[26];
  assign N1212 = N10679 & csr_rdata_o[25];
  assign N10679 = ~csr_wdata_i[25];
  assign N1213 = N10680 & csr_rdata_o[24];
  assign N10680 = ~csr_wdata_i[24];
  assign N1214 = N10681 & csr_rdata_o[23];
  assign N10681 = ~csr_wdata_i[23];
  assign N1215 = N10682 & csr_rdata_o[22];
  assign N10682 = ~csr_wdata_i[22];
  assign N1216 = N10683 & csr_rdata_o[21];
  assign N10683 = ~csr_wdata_i[21];
  assign N1217 = N10684 & csr_rdata_o[20];
  assign N10684 = ~csr_wdata_i[20];
  assign N1218 = N10685 & csr_rdata_o[19];
  assign N10685 = ~csr_wdata_i[19];
  assign N1219 = N10686 & csr_rdata_o[18];
  assign N10686 = ~csr_wdata_i[18];
  assign N1220 = N10687 & csr_rdata_o[17];
  assign N10687 = ~csr_wdata_i[17];
  assign N1221 = N10688 & csr_rdata_o[16];
  assign N10688 = ~csr_wdata_i[16];
  assign N1222 = N10689 & csr_rdata_o[15];
  assign N10689 = ~csr_wdata_i[15];
  assign N1223 = N10690 & csr_rdata_o[14];
  assign N10690 = ~csr_wdata_i[14];
  assign N1224 = N10691 & csr_rdata_o[13];
  assign N10691 = ~csr_wdata_i[13];
  assign N1225 = N10692 & csr_rdata_o[12];
  assign N10692 = ~csr_wdata_i[12];
  assign N1226 = N10693 & csr_rdata_o[11];
  assign N10693 = ~csr_wdata_i[11];
  assign N1227 = N10694 & csr_rdata_o[10];
  assign N10694 = ~csr_wdata_i[10];
  assign N1228 = N10695 & csr_rdata_o[9];
  assign N10695 = ~csr_wdata_i[9];
  assign N1229 = N10696 & csr_rdata_o[8];
  assign N10696 = ~csr_wdata_i[8];
  assign N1230 = N10697 & csr_rdata_o[7];
  assign N10697 = ~csr_wdata_i[7];
  assign N1231 = N10698 & csr_rdata_o[6];
  assign N10698 = ~csr_wdata_i[6];
  assign N1232 = N10699 & csr_rdata_o[5];
  assign N10699 = ~csr_wdata_i[5];
  assign N1233 = N10700 & csr_rdata_o[4];
  assign N10700 = ~csr_wdata_i[4];
  assign N1234 = N10701 & csr_rdata_o[3];
  assign N10701 = ~csr_wdata_i[3];
  assign N1235 = N10702 & csr_rdata_o[2];
  assign N10702 = ~csr_wdata_i[2];
  assign N1236 = N10703 & csr_rdata_o[1];
  assign N10703 = ~csr_wdata_i[1];
  assign N1237 = N10704 & csr_rdata_o[0];
  assign N10704 = ~csr_wdata_i[0];
  assign csr_we_int = csr_wreq & instr_new_id_i;
  assign N1238 = ~rst_ni;
  assign N1239 = ~mcountinhibit_we;
  assign mcountinhibit[31] = mcountinhibit_q[31] | 1'b1;
  assign mcountinhibit[30] = mcountinhibit_q[30] | 1'b1;
  assign mcountinhibit[29] = mcountinhibit_q[29] | 1'b1;
  assign mcountinhibit[28] = mcountinhibit_q[28] | 1'b1;
  assign mcountinhibit[27] = mcountinhibit_q[27] | 1'b1;
  assign mcountinhibit[26] = mcountinhibit_q[26] | 1'b1;
  assign mcountinhibit[25] = mcountinhibit_q[25] | 1'b1;
  assign mcountinhibit[24] = mcountinhibit_q[24] | 1'b1;
  assign mcountinhibit[23] = mcountinhibit_q[23] | 1'b1;
  assign mcountinhibit[22] = mcountinhibit_q[22] | 1'b1;
  assign mcountinhibit[21] = mcountinhibit_q[21] | 1'b1;
  assign mcountinhibit[20] = mcountinhibit_q[20] | 1'b1;
  assign mcountinhibit[19] = mcountinhibit_q[19] | 1'b1;
  assign mcountinhibit[18] = mcountinhibit_q[18] | 1'b1;
  assign mcountinhibit[17] = mcountinhibit_q[17] | 1'b1;
  assign mcountinhibit[16] = mcountinhibit_q[16] | 1'b1;
  assign mcountinhibit[15] = mcountinhibit_q[15] | 1'b1;
  assign mcountinhibit[14] = mcountinhibit_q[14] | 1'b1;
  assign mcountinhibit[13] = mcountinhibit_q[13] | 1'b1;
  assign mcountinhibit[12] = mcountinhibit_q[12] | 1'b1;
  assign mcountinhibit[11] = mcountinhibit_q[11] | 1'b1;
  assign mcountinhibit[10] = mcountinhibit_q[10] | 1'b1;
  assign mcountinhibit[9] = mcountinhibit_q[9] | 1'b1;
  assign mcountinhibit[8] = mcountinhibit_q[8] | 1'b1;
  assign mcountinhibit[7] = mcountinhibit_q[7] | 1'b1;
  assign mcountinhibit[6] = mcountinhibit_q[6] | 1'b1;
  assign mcountinhibit[5] = mcountinhibit_q[5] | 1'b1;
  assign mcountinhibit[4] = mcountinhibit_q[4] | 1'b1;
  assign mcountinhibit[3] = mcountinhibit_q[3] | 1'b1;
  assign mcountinhibit[2] = mcountinhibit_q[2] | 1'b0;
  assign mcountinhibit[1] = mcountinhibit_q[1] | 1'b0;
  assign mcountinhibit[0] = mcountinhibit_q[0] | 1'b0;
  assign N1240 = 1'b1 & N10705;
  assign N10705 = ~mcountinhibit[0];
  assign N1241 = ~N1240;
  assign N1306 = 1'b1 & N1305;
  assign N1307 = 1'b1 & N1304;
  assign N1308 = 1'b1 & N1303;
  assign N1309 = 1'b1 & N1302;
  assign N1310 = 1'b1 & N1301;
  assign N1311 = 1'b1 & N1300;
  assign N1312 = 1'b1 & N1299;
  assign N1313 = 1'b1 & N1298;
  assign N1314 = 1'b1 & N1297;
  assign N1315 = 1'b1 & N1296;
  assign N1316 = 1'b1 & N1295;
  assign N1317 = 1'b1 & N1294;
  assign N1318 = 1'b1 & N1293;
  assign N1319 = 1'b1 & N1292;
  assign N1320 = 1'b1 & N1291;
  assign N1321 = 1'b1 & N1290;
  assign N1322 = 1'b1 & N1289;
  assign N1323 = 1'b1 & N1288;
  assign N1324 = 1'b1 & N1287;
  assign N1325 = 1'b1 & N1286;
  assign N1326 = 1'b1 & N1285;
  assign N1327 = 1'b1 & N1284;
  assign N1328 = 1'b1 & N1283;
  assign N1329 = 1'b1 & N1282;
  assign N1330 = 1'b1 & N1281;
  assign N1331 = 1'b1 & N1280;
  assign N1332 = 1'b1 & N1279;
  assign N1333 = 1'b1 & N1278;
  assign N1334 = 1'b1 & N1277;
  assign N1335 = 1'b1 & N1276;
  assign N1336 = 1'b1 & N1275;
  assign N1337 = 1'b1 & N1274;
  assign N1338 = 1'b1 & N1273;
  assign N1339 = 1'b1 & N1272;
  assign N1340 = 1'b1 & N1271;
  assign N1341 = 1'b1 & N1270;
  assign N1342 = 1'b1 & N1269;
  assign N1343 = 1'b1 & N1268;
  assign N1344 = 1'b1 & N1267;
  assign N1345 = 1'b1 & N1266;
  assign N1346 = 1'b1 & N1265;
  assign N1347 = 1'b1 & N1264;
  assign N1348 = 1'b1 & N1263;
  assign N1349 = 1'b1 & N1262;
  assign N1350 = 1'b1 & N1261;
  assign N1351 = 1'b1 & N1260;
  assign N1352 = 1'b1 & N1259;
  assign N1353 = 1'b1 & N1258;
  assign N1354 = 1'b1 & N1257;
  assign N1355 = 1'b1 & N1256;
  assign N1356 = 1'b1 & N1255;
  assign N1357 = 1'b1 & N1254;
  assign N1358 = 1'b1 & N1253;
  assign N1359 = 1'b1 & N1252;
  assign N1360 = 1'b1 & N1251;
  assign N1361 = 1'b1 & N1250;
  assign N1362 = 1'b1 & N1249;
  assign N1363 = 1'b1 & N1248;
  assign N1364 = 1'b1 & N1247;
  assign N1365 = 1'b1 & N1246;
  assign N1366 = 1'b1 & N1245;
  assign N1367 = 1'b1 & N1244;
  assign N1368 = 1'b1 & N1243;
  assign N1369 = 1'b1 & N1242;
  assign N1434 = ~mhpmcounter_we[0];
  assign N1435 = 1'b1 & csr_wdata_int[31];
  assign N1436 = 1'b1 & csr_wdata_int[30];
  assign N1437 = 1'b1 & csr_wdata_int[29];
  assign N1438 = 1'b1 & csr_wdata_int[28];
  assign N1439 = 1'b1 & csr_wdata_int[27];
  assign N1440 = 1'b1 & csr_wdata_int[26];
  assign N1441 = 1'b1 & csr_wdata_int[25];
  assign N1442 = 1'b1 & csr_wdata_int[24];
  assign N1443 = 1'b1 & csr_wdata_int[23];
  assign N1444 = 1'b1 & csr_wdata_int[22];
  assign N1445 = 1'b1 & csr_wdata_int[21];
  assign N1446 = 1'b1 & csr_wdata_int[20];
  assign N1447 = 1'b1 & csr_wdata_int[19];
  assign N1448 = 1'b1 & csr_wdata_int[18];
  assign N1449 = 1'b1 & csr_wdata_int[17];
  assign N1450 = 1'b1 & csr_wdata_int[16];
  assign N1451 = 1'b1 & csr_wdata_int[15];
  assign N1452 = 1'b1 & csr_wdata_int[14];
  assign N1453 = 1'b1 & csr_wdata_int[13];
  assign N1454 = 1'b1 & csr_wdata_int[12];
  assign N1455 = 1'b1 & csr_wdata_int[11];
  assign N1456 = 1'b1 & csr_wdata_int[10];
  assign N1457 = 1'b1 & csr_wdata_int[9];
  assign N1458 = 1'b1 & csr_wdata_int[8];
  assign N1459 = 1'b1 & csr_wdata_int[7];
  assign N1460 = 1'b1 & csr_wdata_int[6];
  assign N1461 = 1'b1 & csr_wdata_int[5];
  assign N1462 = 1'b1 & csr_wdata_int[4];
  assign N1463 = 1'b1 & csr_wdata_int[3];
  assign N1464 = 1'b1 & csr_wdata_int[2];
  assign N1465 = 1'b1 & csr_wdata_int[1];
  assign N1466 = 1'b1 & csr_wdata_int[0];
  assign N1467 = ~mhpmcounterh_we[0];
  assign N1468 = 1'b1 & csr_wdata_int[31];
  assign N1469 = 1'b1 & csr_wdata_int[30];
  assign N1470 = 1'b1 & csr_wdata_int[29];
  assign N1471 = 1'b1 & csr_wdata_int[28];
  assign N1472 = 1'b1 & csr_wdata_int[27];
  assign N1473 = 1'b1 & csr_wdata_int[26];
  assign N1474 = 1'b1 & csr_wdata_int[25];
  assign N1475 = 1'b1 & csr_wdata_int[24];
  assign N1476 = 1'b1 & csr_wdata_int[23];
  assign N1477 = 1'b1 & csr_wdata_int[22];
  assign N1478 = 1'b1 & csr_wdata_int[21];
  assign N1479 = 1'b1 & csr_wdata_int[20];
  assign N1480 = 1'b1 & csr_wdata_int[19];
  assign N1481 = 1'b1 & csr_wdata_int[18];
  assign N1482 = 1'b1 & csr_wdata_int[17];
  assign N1483 = 1'b1 & csr_wdata_int[16];
  assign N1484 = 1'b1 & csr_wdata_int[15];
  assign N1485 = 1'b1 & csr_wdata_int[14];
  assign N1486 = 1'b1 & csr_wdata_int[13];
  assign N1487 = 1'b1 & csr_wdata_int[12];
  assign N1488 = 1'b1 & csr_wdata_int[11];
  assign N1489 = 1'b1 & csr_wdata_int[10];
  assign N1490 = 1'b1 & csr_wdata_int[9];
  assign N1491 = 1'b1 & csr_wdata_int[8];
  assign N1492 = 1'b1 & csr_wdata_int[7];
  assign N1493 = 1'b1 & csr_wdata_int[6];
  assign N1494 = 1'b1 & csr_wdata_int[5];
  assign N1495 = 1'b1 & csr_wdata_int[4];
  assign N1496 = 1'b1 & csr_wdata_int[3];
  assign N1497 = 1'b1 & csr_wdata_int[2];
  assign N1498 = 1'b1 & csr_wdata_int[1];
  assign N1499 = 1'b1 & csr_wdata_int[0];
  assign N1532 = 1'b0 & N10706;
  assign N10706 = ~mcountinhibit[1];
  assign N1533 = ~N1532;
  assign N1598 = 1'b1 & N1597;
  assign N1599 = 1'b1 & N1596;
  assign N1600 = 1'b1 & N1595;
  assign N1601 = 1'b1 & N1594;
  assign N1602 = 1'b1 & N1593;
  assign N1603 = 1'b1 & N1592;
  assign N1604 = 1'b1 & N1591;
  assign N1605 = 1'b1 & N1590;
  assign N1606 = 1'b1 & N1589;
  assign N1607 = 1'b1 & N1588;
  assign N1608 = 1'b1 & N1587;
  assign N1609 = 1'b1 & N1586;
  assign N1610 = 1'b1 & N1585;
  assign N1611 = 1'b1 & N1584;
  assign N1612 = 1'b1 & N1583;
  assign N1613 = 1'b1 & N1582;
  assign N1614 = 1'b1 & N1581;
  assign N1615 = 1'b1 & N1580;
  assign N1616 = 1'b1 & N1579;
  assign N1617 = 1'b1 & N1578;
  assign N1618 = 1'b1 & N1577;
  assign N1619 = 1'b1 & N1576;
  assign N1620 = 1'b1 & N1575;
  assign N1621 = 1'b1 & N1574;
  assign N1622 = 1'b1 & N1573;
  assign N1623 = 1'b1 & N1572;
  assign N1624 = 1'b1 & N1571;
  assign N1625 = 1'b1 & N1570;
  assign N1626 = 1'b1 & N1569;
  assign N1627 = 1'b1 & N1568;
  assign N1628 = 1'b1 & N1567;
  assign N1629 = 1'b1 & N1566;
  assign N1630 = 1'b1 & N1565;
  assign N1631 = 1'b1 & N1564;
  assign N1632 = 1'b1 & N1563;
  assign N1633 = 1'b1 & N1562;
  assign N1634 = 1'b1 & N1561;
  assign N1635 = 1'b1 & N1560;
  assign N1636 = 1'b1 & N1559;
  assign N1637 = 1'b1 & N1558;
  assign N1638 = 1'b1 & N1557;
  assign N1639 = 1'b1 & N1556;
  assign N1640 = 1'b1 & N1555;
  assign N1641 = 1'b1 & N1554;
  assign N1642 = 1'b1 & N1553;
  assign N1643 = 1'b1 & N1552;
  assign N1644 = 1'b1 & N1551;
  assign N1645 = 1'b1 & N1550;
  assign N1646 = 1'b1 & N1549;
  assign N1647 = 1'b1 & N1548;
  assign N1648 = 1'b1 & N1547;
  assign N1649 = 1'b1 & N1546;
  assign N1650 = 1'b1 & N1545;
  assign N1651 = 1'b1 & N1544;
  assign N1652 = 1'b1 & N1543;
  assign N1653 = 1'b1 & N1542;
  assign N1654 = 1'b1 & N1541;
  assign N1655 = 1'b1 & N1540;
  assign N1656 = 1'b1 & N1539;
  assign N1657 = 1'b1 & N1538;
  assign N1658 = 1'b1 & N1537;
  assign N1659 = 1'b1 & N1536;
  assign N1660 = 1'b1 & N1535;
  assign N1661 = 1'b1 & N1534;
  assign N1726 = ~mhpmcounter_we[1];
  assign N1727 = 1'b1 & csr_wdata_int[31];
  assign N1728 = 1'b1 & csr_wdata_int[30];
  assign N1729 = 1'b1 & csr_wdata_int[29];
  assign N1730 = 1'b1 & csr_wdata_int[28];
  assign N1731 = 1'b1 & csr_wdata_int[27];
  assign N1732 = 1'b1 & csr_wdata_int[26];
  assign N1733 = 1'b1 & csr_wdata_int[25];
  assign N1734 = 1'b1 & csr_wdata_int[24];
  assign N1735 = 1'b1 & csr_wdata_int[23];
  assign N1736 = 1'b1 & csr_wdata_int[22];
  assign N1737 = 1'b1 & csr_wdata_int[21];
  assign N1738 = 1'b1 & csr_wdata_int[20];
  assign N1739 = 1'b1 & csr_wdata_int[19];
  assign N1740 = 1'b1 & csr_wdata_int[18];
  assign N1741 = 1'b1 & csr_wdata_int[17];
  assign N1742 = 1'b1 & csr_wdata_int[16];
  assign N1743 = 1'b1 & csr_wdata_int[15];
  assign N1744 = 1'b1 & csr_wdata_int[14];
  assign N1745 = 1'b1 & csr_wdata_int[13];
  assign N1746 = 1'b1 & csr_wdata_int[12];
  assign N1747 = 1'b1 & csr_wdata_int[11];
  assign N1748 = 1'b1 & csr_wdata_int[10];
  assign N1749 = 1'b1 & csr_wdata_int[9];
  assign N1750 = 1'b1 & csr_wdata_int[8];
  assign N1751 = 1'b1 & csr_wdata_int[7];
  assign N1752 = 1'b1 & csr_wdata_int[6];
  assign N1753 = 1'b1 & csr_wdata_int[5];
  assign N1754 = 1'b1 & csr_wdata_int[4];
  assign N1755 = 1'b1 & csr_wdata_int[3];
  assign N1756 = 1'b1 & csr_wdata_int[2];
  assign N1757 = 1'b1 & csr_wdata_int[1];
  assign N1758 = 1'b1 & csr_wdata_int[0];
  assign N1759 = ~mhpmcounterh_we[1];
  assign N1760 = 1'b1 & csr_wdata_int[31];
  assign N1761 = 1'b1 & csr_wdata_int[30];
  assign N1762 = 1'b1 & csr_wdata_int[29];
  assign N1763 = 1'b1 & csr_wdata_int[28];
  assign N1764 = 1'b1 & csr_wdata_int[27];
  assign N1765 = 1'b1 & csr_wdata_int[26];
  assign N1766 = 1'b1 & csr_wdata_int[25];
  assign N1767 = 1'b1 & csr_wdata_int[24];
  assign N1768 = 1'b1 & csr_wdata_int[23];
  assign N1769 = 1'b1 & csr_wdata_int[22];
  assign N1770 = 1'b1 & csr_wdata_int[21];
  assign N1771 = 1'b1 & csr_wdata_int[20];
  assign N1772 = 1'b1 & csr_wdata_int[19];
  assign N1773 = 1'b1 & csr_wdata_int[18];
  assign N1774 = 1'b1 & csr_wdata_int[17];
  assign N1775 = 1'b1 & csr_wdata_int[16];
  assign N1776 = 1'b1 & csr_wdata_int[15];
  assign N1777 = 1'b1 & csr_wdata_int[14];
  assign N1778 = 1'b1 & csr_wdata_int[13];
  assign N1779 = 1'b1 & csr_wdata_int[12];
  assign N1780 = 1'b1 & csr_wdata_int[11];
  assign N1781 = 1'b1 & csr_wdata_int[10];
  assign N1782 = 1'b1 & csr_wdata_int[9];
  assign N1783 = 1'b1 & csr_wdata_int[8];
  assign N1784 = 1'b1 & csr_wdata_int[7];
  assign N1785 = 1'b1 & csr_wdata_int[6];
  assign N1786 = 1'b1 & csr_wdata_int[5];
  assign N1787 = 1'b1 & csr_wdata_int[4];
  assign N1788 = 1'b1 & csr_wdata_int[3];
  assign N1789 = 1'b1 & csr_wdata_int[2];
  assign N1790 = 1'b1 & csr_wdata_int[1];
  assign N1791 = 1'b1 & csr_wdata_int[0];
  assign N1824 = instr_ret_i & N10707;
  assign N10707 = ~mcountinhibit[2];
  assign N1825 = ~N1824;
  assign N1890 = 1'b1 & N1889;
  assign N1891 = 1'b1 & N1888;
  assign N1892 = 1'b1 & N1887;
  assign N1893 = 1'b1 & N1886;
  assign N1894 = 1'b1 & N1885;
  assign N1895 = 1'b1 & N1884;
  assign N1896 = 1'b1 & N1883;
  assign N1897 = 1'b1 & N1882;
  assign N1898 = 1'b1 & N1881;
  assign N1899 = 1'b1 & N1880;
  assign N1900 = 1'b1 & N1879;
  assign N1901 = 1'b1 & N1878;
  assign N1902 = 1'b1 & N1877;
  assign N1903 = 1'b1 & N1876;
  assign N1904 = 1'b1 & N1875;
  assign N1905 = 1'b1 & N1874;
  assign N1906 = 1'b1 & N1873;
  assign N1907 = 1'b1 & N1872;
  assign N1908 = 1'b1 & N1871;
  assign N1909 = 1'b1 & N1870;
  assign N1910 = 1'b1 & N1869;
  assign N1911 = 1'b1 & N1868;
  assign N1912 = 1'b1 & N1867;
  assign N1913 = 1'b1 & N1866;
  assign N1914 = 1'b1 & N1865;
  assign N1915 = 1'b1 & N1864;
  assign N1916 = 1'b1 & N1863;
  assign N1917 = 1'b1 & N1862;
  assign N1918 = 1'b1 & N1861;
  assign N1919 = 1'b1 & N1860;
  assign N1920 = 1'b1 & N1859;
  assign N1921 = 1'b1 & N1858;
  assign N1922 = 1'b1 & N1857;
  assign N1923 = 1'b1 & N1856;
  assign N1924 = 1'b1 & N1855;
  assign N1925 = 1'b1 & N1854;
  assign N1926 = 1'b1 & N1853;
  assign N1927 = 1'b1 & N1852;
  assign N1928 = 1'b1 & N1851;
  assign N1929 = 1'b1 & N1850;
  assign N1930 = 1'b1 & N1849;
  assign N1931 = 1'b1 & N1848;
  assign N1932 = 1'b1 & N1847;
  assign N1933 = 1'b1 & N1846;
  assign N1934 = 1'b1 & N1845;
  assign N1935 = 1'b1 & N1844;
  assign N1936 = 1'b1 & N1843;
  assign N1937 = 1'b1 & N1842;
  assign N1938 = 1'b1 & N1841;
  assign N1939 = 1'b1 & N1840;
  assign N1940 = 1'b1 & N1839;
  assign N1941 = 1'b1 & N1838;
  assign N1942 = 1'b1 & N1837;
  assign N1943 = 1'b1 & N1836;
  assign N1944 = 1'b1 & N1835;
  assign N1945 = 1'b1 & N1834;
  assign N1946 = 1'b1 & N1833;
  assign N1947 = 1'b1 & N1832;
  assign N1948 = 1'b1 & N1831;
  assign N1949 = 1'b1 & N1830;
  assign N1950 = 1'b1 & N1829;
  assign N1951 = 1'b1 & N1828;
  assign N1952 = 1'b1 & N1827;
  assign N1953 = 1'b1 & N1826;
  assign N2018 = ~mhpmcounter_we[2];
  assign N2019 = 1'b1 & csr_wdata_int[31];
  assign N2020 = 1'b1 & csr_wdata_int[30];
  assign N2021 = 1'b1 & csr_wdata_int[29];
  assign N2022 = 1'b1 & csr_wdata_int[28];
  assign N2023 = 1'b1 & csr_wdata_int[27];
  assign N2024 = 1'b1 & csr_wdata_int[26];
  assign N2025 = 1'b1 & csr_wdata_int[25];
  assign N2026 = 1'b1 & csr_wdata_int[24];
  assign N2027 = 1'b1 & csr_wdata_int[23];
  assign N2028 = 1'b1 & csr_wdata_int[22];
  assign N2029 = 1'b1 & csr_wdata_int[21];
  assign N2030 = 1'b1 & csr_wdata_int[20];
  assign N2031 = 1'b1 & csr_wdata_int[19];
  assign N2032 = 1'b1 & csr_wdata_int[18];
  assign N2033 = 1'b1 & csr_wdata_int[17];
  assign N2034 = 1'b1 & csr_wdata_int[16];
  assign N2035 = 1'b1 & csr_wdata_int[15];
  assign N2036 = 1'b1 & csr_wdata_int[14];
  assign N2037 = 1'b1 & csr_wdata_int[13];
  assign N2038 = 1'b1 & csr_wdata_int[12];
  assign N2039 = 1'b1 & csr_wdata_int[11];
  assign N2040 = 1'b1 & csr_wdata_int[10];
  assign N2041 = 1'b1 & csr_wdata_int[9];
  assign N2042 = 1'b1 & csr_wdata_int[8];
  assign N2043 = 1'b1 & csr_wdata_int[7];
  assign N2044 = 1'b1 & csr_wdata_int[6];
  assign N2045 = 1'b1 & csr_wdata_int[5];
  assign N2046 = 1'b1 & csr_wdata_int[4];
  assign N2047 = 1'b1 & csr_wdata_int[3];
  assign N2048 = 1'b1 & csr_wdata_int[2];
  assign N2049 = 1'b1 & csr_wdata_int[1];
  assign N2050 = 1'b1 & csr_wdata_int[0];
  assign N2051 = ~mhpmcounterh_we[2];
  assign N2052 = 1'b1 & csr_wdata_int[31];
  assign N2053 = 1'b1 & csr_wdata_int[30];
  assign N2054 = 1'b1 & csr_wdata_int[29];
  assign N2055 = 1'b1 & csr_wdata_int[28];
  assign N2056 = 1'b1 & csr_wdata_int[27];
  assign N2057 = 1'b1 & csr_wdata_int[26];
  assign N2058 = 1'b1 & csr_wdata_int[25];
  assign N2059 = 1'b1 & csr_wdata_int[24];
  assign N2060 = 1'b1 & csr_wdata_int[23];
  assign N2061 = 1'b1 & csr_wdata_int[22];
  assign N2062 = 1'b1 & csr_wdata_int[21];
  assign N2063 = 1'b1 & csr_wdata_int[20];
  assign N2064 = 1'b1 & csr_wdata_int[19];
  assign N2065 = 1'b1 & csr_wdata_int[18];
  assign N2066 = 1'b1 & csr_wdata_int[17];
  assign N2067 = 1'b1 & csr_wdata_int[16];
  assign N2068 = 1'b1 & csr_wdata_int[15];
  assign N2069 = 1'b1 & csr_wdata_int[14];
  assign N2070 = 1'b1 & csr_wdata_int[13];
  assign N2071 = 1'b1 & csr_wdata_int[12];
  assign N2072 = 1'b1 & csr_wdata_int[11];
  assign N2073 = 1'b1 & csr_wdata_int[10];
  assign N2074 = 1'b1 & csr_wdata_int[9];
  assign N2075 = 1'b1 & csr_wdata_int[8];
  assign N2076 = 1'b1 & csr_wdata_int[7];
  assign N2077 = 1'b1 & csr_wdata_int[6];
  assign N2078 = 1'b1 & csr_wdata_int[5];
  assign N2079 = 1'b1 & csr_wdata_int[4];
  assign N2080 = 1'b1 & csr_wdata_int[3];
  assign N2081 = 1'b1 & csr_wdata_int[2];
  assign N2082 = 1'b1 & csr_wdata_int[1];
  assign N2083 = 1'b1 & csr_wdata_int[0];
  assign N2116 = 1'b0 & N10708;
  assign N10708 = ~mcountinhibit[3];
  assign N2117 = ~N2116;
  assign N2182 = 1'b0 & N2181;
  assign N2183 = 1'b0 & N2180;
  assign N2184 = 1'b0 & N2179;
  assign N2185 = 1'b0 & N2178;
  assign N2186 = 1'b0 & N2177;
  assign N2187 = 1'b0 & N2176;
  assign N2188 = 1'b0 & N2175;
  assign N2189 = 1'b0 & N2174;
  assign N2190 = 1'b0 & N2173;
  assign N2191 = 1'b0 & N2172;
  assign N2192 = 1'b0 & N2171;
  assign N2193 = 1'b0 & N2170;
  assign N2194 = 1'b0 & N2169;
  assign N2195 = 1'b0 & N2168;
  assign N2196 = 1'b0 & N2167;
  assign N2197 = 1'b0 & N2166;
  assign N2198 = 1'b0 & N2165;
  assign N2199 = 1'b0 & N2164;
  assign N2200 = 1'b0 & N2163;
  assign N2201 = 1'b0 & N2162;
  assign N2202 = 1'b0 & N2161;
  assign N2203 = 1'b0 & N2160;
  assign N2204 = 1'b0 & N2159;
  assign N2205 = 1'b0 & N2158;
  assign N2206 = 1'b0 & N2157;
  assign N2207 = 1'b0 & N2156;
  assign N2208 = 1'b0 & N2155;
  assign N2209 = 1'b0 & N2154;
  assign N2210 = 1'b0 & N2153;
  assign N2211 = 1'b0 & N2152;
  assign N2212 = 1'b0 & N2151;
  assign N2213 = 1'b0 & N2150;
  assign N2214 = 1'b0 & N2149;
  assign N2215 = 1'b0 & N2148;
  assign N2216 = 1'b0 & N2147;
  assign N2217 = 1'b0 & N2146;
  assign N2218 = 1'b0 & N2145;
  assign N2219 = 1'b0 & N2144;
  assign N2220 = 1'b0 & N2143;
  assign N2221 = 1'b0 & N2142;
  assign N2222 = 1'b0 & N2141;
  assign N2223 = 1'b0 & N2140;
  assign N2224 = 1'b0 & N2139;
  assign N2225 = 1'b0 & N2138;
  assign N2226 = 1'b0 & N2137;
  assign N2227 = 1'b0 & N2136;
  assign N2228 = 1'b0 & N2135;
  assign N2229 = 1'b0 & N2134;
  assign N2230 = 1'b0 & N2133;
  assign N2231 = 1'b0 & N2132;
  assign N2232 = 1'b0 & N2131;
  assign N2233 = 1'b0 & N2130;
  assign N2234 = 1'b0 & N2129;
  assign N2235 = 1'b0 & N2128;
  assign N2236 = 1'b0 & N2127;
  assign N2237 = 1'b0 & N2126;
  assign N2238 = 1'b0 & N2125;
  assign N2239 = 1'b0 & N2124;
  assign N2240 = 1'b0 & N2123;
  assign N2241 = 1'b0 & N2122;
  assign N2242 = 1'b0 & N2121;
  assign N2243 = 1'b0 & N2120;
  assign N2244 = 1'b0 & N2119;
  assign N2245 = 1'b0 & N2118;
  assign N2310 = ~mhpmcounter_we[3];
  assign N2311 = 1'b0 & csr_wdata_int[31];
  assign N2312 = 1'b0 & csr_wdata_int[30];
  assign N2313 = 1'b0 & csr_wdata_int[29];
  assign N2314 = 1'b0 & csr_wdata_int[28];
  assign N2315 = 1'b0 & csr_wdata_int[27];
  assign N2316 = 1'b0 & csr_wdata_int[26];
  assign N2317 = 1'b0 & csr_wdata_int[25];
  assign N2318 = 1'b0 & csr_wdata_int[24];
  assign N2319 = 1'b0 & csr_wdata_int[23];
  assign N2320 = 1'b0 & csr_wdata_int[22];
  assign N2321 = 1'b0 & csr_wdata_int[21];
  assign N2322 = 1'b0 & csr_wdata_int[20];
  assign N2323 = 1'b0 & csr_wdata_int[19];
  assign N2324 = 1'b0 & csr_wdata_int[18];
  assign N2325 = 1'b0 & csr_wdata_int[17];
  assign N2326 = 1'b0 & csr_wdata_int[16];
  assign N2327 = 1'b0 & csr_wdata_int[15];
  assign N2328 = 1'b0 & csr_wdata_int[14];
  assign N2329 = 1'b0 & csr_wdata_int[13];
  assign N2330 = 1'b0 & csr_wdata_int[12];
  assign N2331 = 1'b0 & csr_wdata_int[11];
  assign N2332 = 1'b0 & csr_wdata_int[10];
  assign N2333 = 1'b0 & csr_wdata_int[9];
  assign N2334 = 1'b0 & csr_wdata_int[8];
  assign N2335 = 1'b0 & csr_wdata_int[7];
  assign N2336 = 1'b0 & csr_wdata_int[6];
  assign N2337 = 1'b0 & csr_wdata_int[5];
  assign N2338 = 1'b0 & csr_wdata_int[4];
  assign N2339 = 1'b0 & csr_wdata_int[3];
  assign N2340 = 1'b0 & csr_wdata_int[2];
  assign N2341 = 1'b0 & csr_wdata_int[1];
  assign N2342 = 1'b0 & csr_wdata_int[0];
  assign N2343 = ~mhpmcounterh_we[3];
  assign N2344 = 1'b0 & csr_wdata_int[31];
  assign N2345 = 1'b0 & csr_wdata_int[30];
  assign N2346 = 1'b0 & csr_wdata_int[29];
  assign N2347 = 1'b0 & csr_wdata_int[28];
  assign N2348 = 1'b0 & csr_wdata_int[27];
  assign N2349 = 1'b0 & csr_wdata_int[26];
  assign N2350 = 1'b0 & csr_wdata_int[25];
  assign N2351 = 1'b0 & csr_wdata_int[24];
  assign N2352 = 1'b0 & csr_wdata_int[23];
  assign N2353 = 1'b0 & csr_wdata_int[22];
  assign N2354 = 1'b0 & csr_wdata_int[21];
  assign N2355 = 1'b0 & csr_wdata_int[20];
  assign N2356 = 1'b0 & csr_wdata_int[19];
  assign N2357 = 1'b0 & csr_wdata_int[18];
  assign N2358 = 1'b0 & csr_wdata_int[17];
  assign N2359 = 1'b0 & csr_wdata_int[16];
  assign N2360 = 1'b0 & csr_wdata_int[15];
  assign N2361 = 1'b0 & csr_wdata_int[14];
  assign N2362 = 1'b0 & csr_wdata_int[13];
  assign N2363 = 1'b0 & csr_wdata_int[12];
  assign N2364 = 1'b0 & csr_wdata_int[11];
  assign N2365 = 1'b0 & csr_wdata_int[10];
  assign N2366 = 1'b0 & csr_wdata_int[9];
  assign N2367 = 1'b0 & csr_wdata_int[8];
  assign N2368 = 1'b0 & csr_wdata_int[7];
  assign N2369 = 1'b0 & csr_wdata_int[6];
  assign N2370 = 1'b0 & csr_wdata_int[5];
  assign N2371 = 1'b0 & csr_wdata_int[4];
  assign N2372 = 1'b0 & csr_wdata_int[3];
  assign N2373 = 1'b0 & csr_wdata_int[2];
  assign N2374 = 1'b0 & csr_wdata_int[1];
  assign N2375 = 1'b0 & csr_wdata_int[0];
  assign N2408 = 1'b0 & N10709;
  assign N10709 = ~mcountinhibit[4];
  assign N2409 = ~N2408;
  assign N2474 = 1'b0 & N2473;
  assign N2475 = 1'b0 & N2472;
  assign N2476 = 1'b0 & N2471;
  assign N2477 = 1'b0 & N2470;
  assign N2478 = 1'b0 & N2469;
  assign N2479 = 1'b0 & N2468;
  assign N2480 = 1'b0 & N2467;
  assign N2481 = 1'b0 & N2466;
  assign N2482 = 1'b0 & N2465;
  assign N2483 = 1'b0 & N2464;
  assign N2484 = 1'b0 & N2463;
  assign N2485 = 1'b0 & N2462;
  assign N2486 = 1'b0 & N2461;
  assign N2487 = 1'b0 & N2460;
  assign N2488 = 1'b0 & N2459;
  assign N2489 = 1'b0 & N2458;
  assign N2490 = 1'b0 & N2457;
  assign N2491 = 1'b0 & N2456;
  assign N2492 = 1'b0 & N2455;
  assign N2493 = 1'b0 & N2454;
  assign N2494 = 1'b0 & N2453;
  assign N2495 = 1'b0 & N2452;
  assign N2496 = 1'b0 & N2451;
  assign N2497 = 1'b0 & N2450;
  assign N2498 = 1'b0 & N2449;
  assign N2499 = 1'b0 & N2448;
  assign N2500 = 1'b0 & N2447;
  assign N2501 = 1'b0 & N2446;
  assign N2502 = 1'b0 & N2445;
  assign N2503 = 1'b0 & N2444;
  assign N2504 = 1'b0 & N2443;
  assign N2505 = 1'b0 & N2442;
  assign N2506 = 1'b0 & N2441;
  assign N2507 = 1'b0 & N2440;
  assign N2508 = 1'b0 & N2439;
  assign N2509 = 1'b0 & N2438;
  assign N2510 = 1'b0 & N2437;
  assign N2511 = 1'b0 & N2436;
  assign N2512 = 1'b0 & N2435;
  assign N2513 = 1'b0 & N2434;
  assign N2514 = 1'b0 & N2433;
  assign N2515 = 1'b0 & N2432;
  assign N2516 = 1'b0 & N2431;
  assign N2517 = 1'b0 & N2430;
  assign N2518 = 1'b0 & N2429;
  assign N2519 = 1'b0 & N2428;
  assign N2520 = 1'b0 & N2427;
  assign N2521 = 1'b0 & N2426;
  assign N2522 = 1'b0 & N2425;
  assign N2523 = 1'b0 & N2424;
  assign N2524 = 1'b0 & N2423;
  assign N2525 = 1'b0 & N2422;
  assign N2526 = 1'b0 & N2421;
  assign N2527 = 1'b0 & N2420;
  assign N2528 = 1'b0 & N2419;
  assign N2529 = 1'b0 & N2418;
  assign N2530 = 1'b0 & N2417;
  assign N2531 = 1'b0 & N2416;
  assign N2532 = 1'b0 & N2415;
  assign N2533 = 1'b0 & N2414;
  assign N2534 = 1'b0 & N2413;
  assign N2535 = 1'b0 & N2412;
  assign N2536 = 1'b0 & N2411;
  assign N2537 = 1'b0 & N2410;
  assign N2602 = ~mhpmcounter_we[4];
  assign N2603 = 1'b0 & csr_wdata_int[31];
  assign N2604 = 1'b0 & csr_wdata_int[30];
  assign N2605 = 1'b0 & csr_wdata_int[29];
  assign N2606 = 1'b0 & csr_wdata_int[28];
  assign N2607 = 1'b0 & csr_wdata_int[27];
  assign N2608 = 1'b0 & csr_wdata_int[26];
  assign N2609 = 1'b0 & csr_wdata_int[25];
  assign N2610 = 1'b0 & csr_wdata_int[24];
  assign N2611 = 1'b0 & csr_wdata_int[23];
  assign N2612 = 1'b0 & csr_wdata_int[22];
  assign N2613 = 1'b0 & csr_wdata_int[21];
  assign N2614 = 1'b0 & csr_wdata_int[20];
  assign N2615 = 1'b0 & csr_wdata_int[19];
  assign N2616 = 1'b0 & csr_wdata_int[18];
  assign N2617 = 1'b0 & csr_wdata_int[17];
  assign N2618 = 1'b0 & csr_wdata_int[16];
  assign N2619 = 1'b0 & csr_wdata_int[15];
  assign N2620 = 1'b0 & csr_wdata_int[14];
  assign N2621 = 1'b0 & csr_wdata_int[13];
  assign N2622 = 1'b0 & csr_wdata_int[12];
  assign N2623 = 1'b0 & csr_wdata_int[11];
  assign N2624 = 1'b0 & csr_wdata_int[10];
  assign N2625 = 1'b0 & csr_wdata_int[9];
  assign N2626 = 1'b0 & csr_wdata_int[8];
  assign N2627 = 1'b0 & csr_wdata_int[7];
  assign N2628 = 1'b0 & csr_wdata_int[6];
  assign N2629 = 1'b0 & csr_wdata_int[5];
  assign N2630 = 1'b0 & csr_wdata_int[4];
  assign N2631 = 1'b0 & csr_wdata_int[3];
  assign N2632 = 1'b0 & csr_wdata_int[2];
  assign N2633 = 1'b0 & csr_wdata_int[1];
  assign N2634 = 1'b0 & csr_wdata_int[0];
  assign N2635 = ~mhpmcounterh_we[4];
  assign N2636 = 1'b0 & csr_wdata_int[31];
  assign N2637 = 1'b0 & csr_wdata_int[30];
  assign N2638 = 1'b0 & csr_wdata_int[29];
  assign N2639 = 1'b0 & csr_wdata_int[28];
  assign N2640 = 1'b0 & csr_wdata_int[27];
  assign N2641 = 1'b0 & csr_wdata_int[26];
  assign N2642 = 1'b0 & csr_wdata_int[25];
  assign N2643 = 1'b0 & csr_wdata_int[24];
  assign N2644 = 1'b0 & csr_wdata_int[23];
  assign N2645 = 1'b0 & csr_wdata_int[22];
  assign N2646 = 1'b0 & csr_wdata_int[21];
  assign N2647 = 1'b0 & csr_wdata_int[20];
  assign N2648 = 1'b0 & csr_wdata_int[19];
  assign N2649 = 1'b0 & csr_wdata_int[18];
  assign N2650 = 1'b0 & csr_wdata_int[17];
  assign N2651 = 1'b0 & csr_wdata_int[16];
  assign N2652 = 1'b0 & csr_wdata_int[15];
  assign N2653 = 1'b0 & csr_wdata_int[14];
  assign N2654 = 1'b0 & csr_wdata_int[13];
  assign N2655 = 1'b0 & csr_wdata_int[12];
  assign N2656 = 1'b0 & csr_wdata_int[11];
  assign N2657 = 1'b0 & csr_wdata_int[10];
  assign N2658 = 1'b0 & csr_wdata_int[9];
  assign N2659 = 1'b0 & csr_wdata_int[8];
  assign N2660 = 1'b0 & csr_wdata_int[7];
  assign N2661 = 1'b0 & csr_wdata_int[6];
  assign N2662 = 1'b0 & csr_wdata_int[5];
  assign N2663 = 1'b0 & csr_wdata_int[4];
  assign N2664 = 1'b0 & csr_wdata_int[3];
  assign N2665 = 1'b0 & csr_wdata_int[2];
  assign N2666 = 1'b0 & csr_wdata_int[1];
  assign N2667 = 1'b0 & csr_wdata_int[0];
  assign N2700 = 1'b0 & N10710;
  assign N10710 = ~mcountinhibit[5];
  assign N2701 = ~N2700;
  assign N2766 = 1'b0 & N2765;
  assign N2767 = 1'b0 & N2764;
  assign N2768 = 1'b0 & N2763;
  assign N2769 = 1'b0 & N2762;
  assign N2770 = 1'b0 & N2761;
  assign N2771 = 1'b0 & N2760;
  assign N2772 = 1'b0 & N2759;
  assign N2773 = 1'b0 & N2758;
  assign N2774 = 1'b0 & N2757;
  assign N2775 = 1'b0 & N2756;
  assign N2776 = 1'b0 & N2755;
  assign N2777 = 1'b0 & N2754;
  assign N2778 = 1'b0 & N2753;
  assign N2779 = 1'b0 & N2752;
  assign N2780 = 1'b0 & N2751;
  assign N2781 = 1'b0 & N2750;
  assign N2782 = 1'b0 & N2749;
  assign N2783 = 1'b0 & N2748;
  assign N2784 = 1'b0 & N2747;
  assign N2785 = 1'b0 & N2746;
  assign N2786 = 1'b0 & N2745;
  assign N2787 = 1'b0 & N2744;
  assign N2788 = 1'b0 & N2743;
  assign N2789 = 1'b0 & N2742;
  assign N2790 = 1'b0 & N2741;
  assign N2791 = 1'b0 & N2740;
  assign N2792 = 1'b0 & N2739;
  assign N2793 = 1'b0 & N2738;
  assign N2794 = 1'b0 & N2737;
  assign N2795 = 1'b0 & N2736;
  assign N2796 = 1'b0 & N2735;
  assign N2797 = 1'b0 & N2734;
  assign N2798 = 1'b0 & N2733;
  assign N2799 = 1'b0 & N2732;
  assign N2800 = 1'b0 & N2731;
  assign N2801 = 1'b0 & N2730;
  assign N2802 = 1'b0 & N2729;
  assign N2803 = 1'b0 & N2728;
  assign N2804 = 1'b0 & N2727;
  assign N2805 = 1'b0 & N2726;
  assign N2806 = 1'b0 & N2725;
  assign N2807 = 1'b0 & N2724;
  assign N2808 = 1'b0 & N2723;
  assign N2809 = 1'b0 & N2722;
  assign N2810 = 1'b0 & N2721;
  assign N2811 = 1'b0 & N2720;
  assign N2812 = 1'b0 & N2719;
  assign N2813 = 1'b0 & N2718;
  assign N2814 = 1'b0 & N2717;
  assign N2815 = 1'b0 & N2716;
  assign N2816 = 1'b0 & N2715;
  assign N2817 = 1'b0 & N2714;
  assign N2818 = 1'b0 & N2713;
  assign N2819 = 1'b0 & N2712;
  assign N2820 = 1'b0 & N2711;
  assign N2821 = 1'b0 & N2710;
  assign N2822 = 1'b0 & N2709;
  assign N2823 = 1'b0 & N2708;
  assign N2824 = 1'b0 & N2707;
  assign N2825 = 1'b0 & N2706;
  assign N2826 = 1'b0 & N2705;
  assign N2827 = 1'b0 & N2704;
  assign N2828 = 1'b0 & N2703;
  assign N2829 = 1'b0 & N2702;
  assign N2894 = ~mhpmcounter_we[5];
  assign N2895 = 1'b0 & csr_wdata_int[31];
  assign N2896 = 1'b0 & csr_wdata_int[30];
  assign N2897 = 1'b0 & csr_wdata_int[29];
  assign N2898 = 1'b0 & csr_wdata_int[28];
  assign N2899 = 1'b0 & csr_wdata_int[27];
  assign N2900 = 1'b0 & csr_wdata_int[26];
  assign N2901 = 1'b0 & csr_wdata_int[25];
  assign N2902 = 1'b0 & csr_wdata_int[24];
  assign N2903 = 1'b0 & csr_wdata_int[23];
  assign N2904 = 1'b0 & csr_wdata_int[22];
  assign N2905 = 1'b0 & csr_wdata_int[21];
  assign N2906 = 1'b0 & csr_wdata_int[20];
  assign N2907 = 1'b0 & csr_wdata_int[19];
  assign N2908 = 1'b0 & csr_wdata_int[18];
  assign N2909 = 1'b0 & csr_wdata_int[17];
  assign N2910 = 1'b0 & csr_wdata_int[16];
  assign N2911 = 1'b0 & csr_wdata_int[15];
  assign N2912 = 1'b0 & csr_wdata_int[14];
  assign N2913 = 1'b0 & csr_wdata_int[13];
  assign N2914 = 1'b0 & csr_wdata_int[12];
  assign N2915 = 1'b0 & csr_wdata_int[11];
  assign N2916 = 1'b0 & csr_wdata_int[10];
  assign N2917 = 1'b0 & csr_wdata_int[9];
  assign N2918 = 1'b0 & csr_wdata_int[8];
  assign N2919 = 1'b0 & csr_wdata_int[7];
  assign N2920 = 1'b0 & csr_wdata_int[6];
  assign N2921 = 1'b0 & csr_wdata_int[5];
  assign N2922 = 1'b0 & csr_wdata_int[4];
  assign N2923 = 1'b0 & csr_wdata_int[3];
  assign N2924 = 1'b0 & csr_wdata_int[2];
  assign N2925 = 1'b0 & csr_wdata_int[1];
  assign N2926 = 1'b0 & csr_wdata_int[0];
  assign N2927 = ~mhpmcounterh_we[5];
  assign N2928 = 1'b0 & csr_wdata_int[31];
  assign N2929 = 1'b0 & csr_wdata_int[30];
  assign N2930 = 1'b0 & csr_wdata_int[29];
  assign N2931 = 1'b0 & csr_wdata_int[28];
  assign N2932 = 1'b0 & csr_wdata_int[27];
  assign N2933 = 1'b0 & csr_wdata_int[26];
  assign N2934 = 1'b0 & csr_wdata_int[25];
  assign N2935 = 1'b0 & csr_wdata_int[24];
  assign N2936 = 1'b0 & csr_wdata_int[23];
  assign N2937 = 1'b0 & csr_wdata_int[22];
  assign N2938 = 1'b0 & csr_wdata_int[21];
  assign N2939 = 1'b0 & csr_wdata_int[20];
  assign N2940 = 1'b0 & csr_wdata_int[19];
  assign N2941 = 1'b0 & csr_wdata_int[18];
  assign N2942 = 1'b0 & csr_wdata_int[17];
  assign N2943 = 1'b0 & csr_wdata_int[16];
  assign N2944 = 1'b0 & csr_wdata_int[15];
  assign N2945 = 1'b0 & csr_wdata_int[14];
  assign N2946 = 1'b0 & csr_wdata_int[13];
  assign N2947 = 1'b0 & csr_wdata_int[12];
  assign N2948 = 1'b0 & csr_wdata_int[11];
  assign N2949 = 1'b0 & csr_wdata_int[10];
  assign N2950 = 1'b0 & csr_wdata_int[9];
  assign N2951 = 1'b0 & csr_wdata_int[8];
  assign N2952 = 1'b0 & csr_wdata_int[7];
  assign N2953 = 1'b0 & csr_wdata_int[6];
  assign N2954 = 1'b0 & csr_wdata_int[5];
  assign N2955 = 1'b0 & csr_wdata_int[4];
  assign N2956 = 1'b0 & csr_wdata_int[3];
  assign N2957 = 1'b0 & csr_wdata_int[2];
  assign N2958 = 1'b0 & csr_wdata_int[1];
  assign N2959 = 1'b0 & csr_wdata_int[0];
  assign N2992 = 1'b0 & N10711;
  assign N10711 = ~mcountinhibit[6];
  assign N2993 = ~N2992;
  assign N3058 = 1'b0 & N3057;
  assign N3059 = 1'b0 & N3056;
  assign N3060 = 1'b0 & N3055;
  assign N3061 = 1'b0 & N3054;
  assign N3062 = 1'b0 & N3053;
  assign N3063 = 1'b0 & N3052;
  assign N3064 = 1'b0 & N3051;
  assign N3065 = 1'b0 & N3050;
  assign N3066 = 1'b0 & N3049;
  assign N3067 = 1'b0 & N3048;
  assign N3068 = 1'b0 & N3047;
  assign N3069 = 1'b0 & N3046;
  assign N3070 = 1'b0 & N3045;
  assign N3071 = 1'b0 & N3044;
  assign N3072 = 1'b0 & N3043;
  assign N3073 = 1'b0 & N3042;
  assign N3074 = 1'b0 & N3041;
  assign N3075 = 1'b0 & N3040;
  assign N3076 = 1'b0 & N3039;
  assign N3077 = 1'b0 & N3038;
  assign N3078 = 1'b0 & N3037;
  assign N3079 = 1'b0 & N3036;
  assign N3080 = 1'b0 & N3035;
  assign N3081 = 1'b0 & N3034;
  assign N3082 = 1'b0 & N3033;
  assign N3083 = 1'b0 & N3032;
  assign N3084 = 1'b0 & N3031;
  assign N3085 = 1'b0 & N3030;
  assign N3086 = 1'b0 & N3029;
  assign N3087 = 1'b0 & N3028;
  assign N3088 = 1'b0 & N3027;
  assign N3089 = 1'b0 & N3026;
  assign N3090 = 1'b0 & N3025;
  assign N3091 = 1'b0 & N3024;
  assign N3092 = 1'b0 & N3023;
  assign N3093 = 1'b0 & N3022;
  assign N3094 = 1'b0 & N3021;
  assign N3095 = 1'b0 & N3020;
  assign N3096 = 1'b0 & N3019;
  assign N3097 = 1'b0 & N3018;
  assign N3098 = 1'b0 & N3017;
  assign N3099 = 1'b0 & N3016;
  assign N3100 = 1'b0 & N3015;
  assign N3101 = 1'b0 & N3014;
  assign N3102 = 1'b0 & N3013;
  assign N3103 = 1'b0 & N3012;
  assign N3104 = 1'b0 & N3011;
  assign N3105 = 1'b0 & N3010;
  assign N3106 = 1'b0 & N3009;
  assign N3107 = 1'b0 & N3008;
  assign N3108 = 1'b0 & N3007;
  assign N3109 = 1'b0 & N3006;
  assign N3110 = 1'b0 & N3005;
  assign N3111 = 1'b0 & N3004;
  assign N3112 = 1'b0 & N3003;
  assign N3113 = 1'b0 & N3002;
  assign N3114 = 1'b0 & N3001;
  assign N3115 = 1'b0 & N3000;
  assign N3116 = 1'b0 & N2999;
  assign N3117 = 1'b0 & N2998;
  assign N3118 = 1'b0 & N2997;
  assign N3119 = 1'b0 & N2996;
  assign N3120 = 1'b0 & N2995;
  assign N3121 = 1'b0 & N2994;
  assign N3186 = ~mhpmcounter_we[6];
  assign N3187 = 1'b0 & csr_wdata_int[31];
  assign N3188 = 1'b0 & csr_wdata_int[30];
  assign N3189 = 1'b0 & csr_wdata_int[29];
  assign N3190 = 1'b0 & csr_wdata_int[28];
  assign N3191 = 1'b0 & csr_wdata_int[27];
  assign N3192 = 1'b0 & csr_wdata_int[26];
  assign N3193 = 1'b0 & csr_wdata_int[25];
  assign N3194 = 1'b0 & csr_wdata_int[24];
  assign N3195 = 1'b0 & csr_wdata_int[23];
  assign N3196 = 1'b0 & csr_wdata_int[22];
  assign N3197 = 1'b0 & csr_wdata_int[21];
  assign N3198 = 1'b0 & csr_wdata_int[20];
  assign N3199 = 1'b0 & csr_wdata_int[19];
  assign N3200 = 1'b0 & csr_wdata_int[18];
  assign N3201 = 1'b0 & csr_wdata_int[17];
  assign N3202 = 1'b0 & csr_wdata_int[16];
  assign N3203 = 1'b0 & csr_wdata_int[15];
  assign N3204 = 1'b0 & csr_wdata_int[14];
  assign N3205 = 1'b0 & csr_wdata_int[13];
  assign N3206 = 1'b0 & csr_wdata_int[12];
  assign N3207 = 1'b0 & csr_wdata_int[11];
  assign N3208 = 1'b0 & csr_wdata_int[10];
  assign N3209 = 1'b0 & csr_wdata_int[9];
  assign N3210 = 1'b0 & csr_wdata_int[8];
  assign N3211 = 1'b0 & csr_wdata_int[7];
  assign N3212 = 1'b0 & csr_wdata_int[6];
  assign N3213 = 1'b0 & csr_wdata_int[5];
  assign N3214 = 1'b0 & csr_wdata_int[4];
  assign N3215 = 1'b0 & csr_wdata_int[3];
  assign N3216 = 1'b0 & csr_wdata_int[2];
  assign N3217 = 1'b0 & csr_wdata_int[1];
  assign N3218 = 1'b0 & csr_wdata_int[0];
  assign N3219 = ~mhpmcounterh_we[6];
  assign N3220 = 1'b0 & csr_wdata_int[31];
  assign N3221 = 1'b0 & csr_wdata_int[30];
  assign N3222 = 1'b0 & csr_wdata_int[29];
  assign N3223 = 1'b0 & csr_wdata_int[28];
  assign N3224 = 1'b0 & csr_wdata_int[27];
  assign N3225 = 1'b0 & csr_wdata_int[26];
  assign N3226 = 1'b0 & csr_wdata_int[25];
  assign N3227 = 1'b0 & csr_wdata_int[24];
  assign N3228 = 1'b0 & csr_wdata_int[23];
  assign N3229 = 1'b0 & csr_wdata_int[22];
  assign N3230 = 1'b0 & csr_wdata_int[21];
  assign N3231 = 1'b0 & csr_wdata_int[20];
  assign N3232 = 1'b0 & csr_wdata_int[19];
  assign N3233 = 1'b0 & csr_wdata_int[18];
  assign N3234 = 1'b0 & csr_wdata_int[17];
  assign N3235 = 1'b0 & csr_wdata_int[16];
  assign N3236 = 1'b0 & csr_wdata_int[15];
  assign N3237 = 1'b0 & csr_wdata_int[14];
  assign N3238 = 1'b0 & csr_wdata_int[13];
  assign N3239 = 1'b0 & csr_wdata_int[12];
  assign N3240 = 1'b0 & csr_wdata_int[11];
  assign N3241 = 1'b0 & csr_wdata_int[10];
  assign N3242 = 1'b0 & csr_wdata_int[9];
  assign N3243 = 1'b0 & csr_wdata_int[8];
  assign N3244 = 1'b0 & csr_wdata_int[7];
  assign N3245 = 1'b0 & csr_wdata_int[6];
  assign N3246 = 1'b0 & csr_wdata_int[5];
  assign N3247 = 1'b0 & csr_wdata_int[4];
  assign N3248 = 1'b0 & csr_wdata_int[3];
  assign N3249 = 1'b0 & csr_wdata_int[2];
  assign N3250 = 1'b0 & csr_wdata_int[1];
  assign N3251 = 1'b0 & csr_wdata_int[0];
  assign N3284 = 1'b0 & N10712;
  assign N10712 = ~mcountinhibit[7];
  assign N3285 = ~N3284;
  assign N3350 = 1'b0 & N3349;
  assign N3351 = 1'b0 & N3348;
  assign N3352 = 1'b0 & N3347;
  assign N3353 = 1'b0 & N3346;
  assign N3354 = 1'b0 & N3345;
  assign N3355 = 1'b0 & N3344;
  assign N3356 = 1'b0 & N3343;
  assign N3357 = 1'b0 & N3342;
  assign N3358 = 1'b0 & N3341;
  assign N3359 = 1'b0 & N3340;
  assign N3360 = 1'b0 & N3339;
  assign N3361 = 1'b0 & N3338;
  assign N3362 = 1'b0 & N3337;
  assign N3363 = 1'b0 & N3336;
  assign N3364 = 1'b0 & N3335;
  assign N3365 = 1'b0 & N3334;
  assign N3366 = 1'b0 & N3333;
  assign N3367 = 1'b0 & N3332;
  assign N3368 = 1'b0 & N3331;
  assign N3369 = 1'b0 & N3330;
  assign N3370 = 1'b0 & N3329;
  assign N3371 = 1'b0 & N3328;
  assign N3372 = 1'b0 & N3327;
  assign N3373 = 1'b0 & N3326;
  assign N3374 = 1'b0 & N3325;
  assign N3375 = 1'b0 & N3324;
  assign N3376 = 1'b0 & N3323;
  assign N3377 = 1'b0 & N3322;
  assign N3378 = 1'b0 & N3321;
  assign N3379 = 1'b0 & N3320;
  assign N3380 = 1'b0 & N3319;
  assign N3381 = 1'b0 & N3318;
  assign N3382 = 1'b0 & N3317;
  assign N3383 = 1'b0 & N3316;
  assign N3384 = 1'b0 & N3315;
  assign N3385 = 1'b0 & N3314;
  assign N3386 = 1'b0 & N3313;
  assign N3387 = 1'b0 & N3312;
  assign N3388 = 1'b0 & N3311;
  assign N3389 = 1'b0 & N3310;
  assign N3390 = 1'b0 & N3309;
  assign N3391 = 1'b0 & N3308;
  assign N3392 = 1'b0 & N3307;
  assign N3393 = 1'b0 & N3306;
  assign N3394 = 1'b0 & N3305;
  assign N3395 = 1'b0 & N3304;
  assign N3396 = 1'b0 & N3303;
  assign N3397 = 1'b0 & N3302;
  assign N3398 = 1'b0 & N3301;
  assign N3399 = 1'b0 & N3300;
  assign N3400 = 1'b0 & N3299;
  assign N3401 = 1'b0 & N3298;
  assign N3402 = 1'b0 & N3297;
  assign N3403 = 1'b0 & N3296;
  assign N3404 = 1'b0 & N3295;
  assign N3405 = 1'b0 & N3294;
  assign N3406 = 1'b0 & N3293;
  assign N3407 = 1'b0 & N3292;
  assign N3408 = 1'b0 & N3291;
  assign N3409 = 1'b0 & N3290;
  assign N3410 = 1'b0 & N3289;
  assign N3411 = 1'b0 & N3288;
  assign N3412 = 1'b0 & N3287;
  assign N3413 = 1'b0 & N3286;
  assign N3478 = ~mhpmcounter_we[7];
  assign N3479 = 1'b0 & csr_wdata_int[31];
  assign N3480 = 1'b0 & csr_wdata_int[30];
  assign N3481 = 1'b0 & csr_wdata_int[29];
  assign N3482 = 1'b0 & csr_wdata_int[28];
  assign N3483 = 1'b0 & csr_wdata_int[27];
  assign N3484 = 1'b0 & csr_wdata_int[26];
  assign N3485 = 1'b0 & csr_wdata_int[25];
  assign N3486 = 1'b0 & csr_wdata_int[24];
  assign N3487 = 1'b0 & csr_wdata_int[23];
  assign N3488 = 1'b0 & csr_wdata_int[22];
  assign N3489 = 1'b0 & csr_wdata_int[21];
  assign N3490 = 1'b0 & csr_wdata_int[20];
  assign N3491 = 1'b0 & csr_wdata_int[19];
  assign N3492 = 1'b0 & csr_wdata_int[18];
  assign N3493 = 1'b0 & csr_wdata_int[17];
  assign N3494 = 1'b0 & csr_wdata_int[16];
  assign N3495 = 1'b0 & csr_wdata_int[15];
  assign N3496 = 1'b0 & csr_wdata_int[14];
  assign N3497 = 1'b0 & csr_wdata_int[13];
  assign N3498 = 1'b0 & csr_wdata_int[12];
  assign N3499 = 1'b0 & csr_wdata_int[11];
  assign N3500 = 1'b0 & csr_wdata_int[10];
  assign N3501 = 1'b0 & csr_wdata_int[9];
  assign N3502 = 1'b0 & csr_wdata_int[8];
  assign N3503 = 1'b0 & csr_wdata_int[7];
  assign N3504 = 1'b0 & csr_wdata_int[6];
  assign N3505 = 1'b0 & csr_wdata_int[5];
  assign N3506 = 1'b0 & csr_wdata_int[4];
  assign N3507 = 1'b0 & csr_wdata_int[3];
  assign N3508 = 1'b0 & csr_wdata_int[2];
  assign N3509 = 1'b0 & csr_wdata_int[1];
  assign N3510 = 1'b0 & csr_wdata_int[0];
  assign N3511 = ~mhpmcounterh_we[7];
  assign N3512 = 1'b0 & csr_wdata_int[31];
  assign N3513 = 1'b0 & csr_wdata_int[30];
  assign N3514 = 1'b0 & csr_wdata_int[29];
  assign N3515 = 1'b0 & csr_wdata_int[28];
  assign N3516 = 1'b0 & csr_wdata_int[27];
  assign N3517 = 1'b0 & csr_wdata_int[26];
  assign N3518 = 1'b0 & csr_wdata_int[25];
  assign N3519 = 1'b0 & csr_wdata_int[24];
  assign N3520 = 1'b0 & csr_wdata_int[23];
  assign N3521 = 1'b0 & csr_wdata_int[22];
  assign N3522 = 1'b0 & csr_wdata_int[21];
  assign N3523 = 1'b0 & csr_wdata_int[20];
  assign N3524 = 1'b0 & csr_wdata_int[19];
  assign N3525 = 1'b0 & csr_wdata_int[18];
  assign N3526 = 1'b0 & csr_wdata_int[17];
  assign N3527 = 1'b0 & csr_wdata_int[16];
  assign N3528 = 1'b0 & csr_wdata_int[15];
  assign N3529 = 1'b0 & csr_wdata_int[14];
  assign N3530 = 1'b0 & csr_wdata_int[13];
  assign N3531 = 1'b0 & csr_wdata_int[12];
  assign N3532 = 1'b0 & csr_wdata_int[11];
  assign N3533 = 1'b0 & csr_wdata_int[10];
  assign N3534 = 1'b0 & csr_wdata_int[9];
  assign N3535 = 1'b0 & csr_wdata_int[8];
  assign N3536 = 1'b0 & csr_wdata_int[7];
  assign N3537 = 1'b0 & csr_wdata_int[6];
  assign N3538 = 1'b0 & csr_wdata_int[5];
  assign N3539 = 1'b0 & csr_wdata_int[4];
  assign N3540 = 1'b0 & csr_wdata_int[3];
  assign N3541 = 1'b0 & csr_wdata_int[2];
  assign N3542 = 1'b0 & csr_wdata_int[1];
  assign N3543 = 1'b0 & csr_wdata_int[0];
  assign N3576 = 1'b0 & N10713;
  assign N10713 = ~mcountinhibit[8];
  assign N3577 = ~N3576;
  assign N3642 = 1'b0 & N3641;
  assign N3643 = 1'b0 & N3640;
  assign N3644 = 1'b0 & N3639;
  assign N3645 = 1'b0 & N3638;
  assign N3646 = 1'b0 & N3637;
  assign N3647 = 1'b0 & N3636;
  assign N3648 = 1'b0 & N3635;
  assign N3649 = 1'b0 & N3634;
  assign N3650 = 1'b0 & N3633;
  assign N3651 = 1'b0 & N3632;
  assign N3652 = 1'b0 & N3631;
  assign N3653 = 1'b0 & N3630;
  assign N3654 = 1'b0 & N3629;
  assign N3655 = 1'b0 & N3628;
  assign N3656 = 1'b0 & N3627;
  assign N3657 = 1'b0 & N3626;
  assign N3658 = 1'b0 & N3625;
  assign N3659 = 1'b0 & N3624;
  assign N3660 = 1'b0 & N3623;
  assign N3661 = 1'b0 & N3622;
  assign N3662 = 1'b0 & N3621;
  assign N3663 = 1'b0 & N3620;
  assign N3664 = 1'b0 & N3619;
  assign N3665 = 1'b0 & N3618;
  assign N3666 = 1'b0 & N3617;
  assign N3667 = 1'b0 & N3616;
  assign N3668 = 1'b0 & N3615;
  assign N3669 = 1'b0 & N3614;
  assign N3670 = 1'b0 & N3613;
  assign N3671 = 1'b0 & N3612;
  assign N3672 = 1'b0 & N3611;
  assign N3673 = 1'b0 & N3610;
  assign N3674 = 1'b0 & N3609;
  assign N3675 = 1'b0 & N3608;
  assign N3676 = 1'b0 & N3607;
  assign N3677 = 1'b0 & N3606;
  assign N3678 = 1'b0 & N3605;
  assign N3679 = 1'b0 & N3604;
  assign N3680 = 1'b0 & N3603;
  assign N3681 = 1'b0 & N3602;
  assign N3682 = 1'b0 & N3601;
  assign N3683 = 1'b0 & N3600;
  assign N3684 = 1'b0 & N3599;
  assign N3685 = 1'b0 & N3598;
  assign N3686 = 1'b0 & N3597;
  assign N3687 = 1'b0 & N3596;
  assign N3688 = 1'b0 & N3595;
  assign N3689 = 1'b0 & N3594;
  assign N3690 = 1'b0 & N3593;
  assign N3691 = 1'b0 & N3592;
  assign N3692 = 1'b0 & N3591;
  assign N3693 = 1'b0 & N3590;
  assign N3694 = 1'b0 & N3589;
  assign N3695 = 1'b0 & N3588;
  assign N3696 = 1'b0 & N3587;
  assign N3697 = 1'b0 & N3586;
  assign N3698 = 1'b0 & N3585;
  assign N3699 = 1'b0 & N3584;
  assign N3700 = 1'b0 & N3583;
  assign N3701 = 1'b0 & N3582;
  assign N3702 = 1'b0 & N3581;
  assign N3703 = 1'b0 & N3580;
  assign N3704 = 1'b0 & N3579;
  assign N3705 = 1'b0 & N3578;
  assign N3770 = ~mhpmcounter_we[8];
  assign N3771 = 1'b0 & csr_wdata_int[31];
  assign N3772 = 1'b0 & csr_wdata_int[30];
  assign N3773 = 1'b0 & csr_wdata_int[29];
  assign N3774 = 1'b0 & csr_wdata_int[28];
  assign N3775 = 1'b0 & csr_wdata_int[27];
  assign N3776 = 1'b0 & csr_wdata_int[26];
  assign N3777 = 1'b0 & csr_wdata_int[25];
  assign N3778 = 1'b0 & csr_wdata_int[24];
  assign N3779 = 1'b0 & csr_wdata_int[23];
  assign N3780 = 1'b0 & csr_wdata_int[22];
  assign N3781 = 1'b0 & csr_wdata_int[21];
  assign N3782 = 1'b0 & csr_wdata_int[20];
  assign N3783 = 1'b0 & csr_wdata_int[19];
  assign N3784 = 1'b0 & csr_wdata_int[18];
  assign N3785 = 1'b0 & csr_wdata_int[17];
  assign N3786 = 1'b0 & csr_wdata_int[16];
  assign N3787 = 1'b0 & csr_wdata_int[15];
  assign N3788 = 1'b0 & csr_wdata_int[14];
  assign N3789 = 1'b0 & csr_wdata_int[13];
  assign N3790 = 1'b0 & csr_wdata_int[12];
  assign N3791 = 1'b0 & csr_wdata_int[11];
  assign N3792 = 1'b0 & csr_wdata_int[10];
  assign N3793 = 1'b0 & csr_wdata_int[9];
  assign N3794 = 1'b0 & csr_wdata_int[8];
  assign N3795 = 1'b0 & csr_wdata_int[7];
  assign N3796 = 1'b0 & csr_wdata_int[6];
  assign N3797 = 1'b0 & csr_wdata_int[5];
  assign N3798 = 1'b0 & csr_wdata_int[4];
  assign N3799 = 1'b0 & csr_wdata_int[3];
  assign N3800 = 1'b0 & csr_wdata_int[2];
  assign N3801 = 1'b0 & csr_wdata_int[1];
  assign N3802 = 1'b0 & csr_wdata_int[0];
  assign N3803 = ~mhpmcounterh_we[8];
  assign N3804 = 1'b0 & csr_wdata_int[31];
  assign N3805 = 1'b0 & csr_wdata_int[30];
  assign N3806 = 1'b0 & csr_wdata_int[29];
  assign N3807 = 1'b0 & csr_wdata_int[28];
  assign N3808 = 1'b0 & csr_wdata_int[27];
  assign N3809 = 1'b0 & csr_wdata_int[26];
  assign N3810 = 1'b0 & csr_wdata_int[25];
  assign N3811 = 1'b0 & csr_wdata_int[24];
  assign N3812 = 1'b0 & csr_wdata_int[23];
  assign N3813 = 1'b0 & csr_wdata_int[22];
  assign N3814 = 1'b0 & csr_wdata_int[21];
  assign N3815 = 1'b0 & csr_wdata_int[20];
  assign N3816 = 1'b0 & csr_wdata_int[19];
  assign N3817 = 1'b0 & csr_wdata_int[18];
  assign N3818 = 1'b0 & csr_wdata_int[17];
  assign N3819 = 1'b0 & csr_wdata_int[16];
  assign N3820 = 1'b0 & csr_wdata_int[15];
  assign N3821 = 1'b0 & csr_wdata_int[14];
  assign N3822 = 1'b0 & csr_wdata_int[13];
  assign N3823 = 1'b0 & csr_wdata_int[12];
  assign N3824 = 1'b0 & csr_wdata_int[11];
  assign N3825 = 1'b0 & csr_wdata_int[10];
  assign N3826 = 1'b0 & csr_wdata_int[9];
  assign N3827 = 1'b0 & csr_wdata_int[8];
  assign N3828 = 1'b0 & csr_wdata_int[7];
  assign N3829 = 1'b0 & csr_wdata_int[6];
  assign N3830 = 1'b0 & csr_wdata_int[5];
  assign N3831 = 1'b0 & csr_wdata_int[4];
  assign N3832 = 1'b0 & csr_wdata_int[3];
  assign N3833 = 1'b0 & csr_wdata_int[2];
  assign N3834 = 1'b0 & csr_wdata_int[1];
  assign N3835 = 1'b0 & csr_wdata_int[0];
  assign N3868 = 1'b0 & N10714;
  assign N10714 = ~mcountinhibit[9];
  assign N3869 = ~N3868;
  assign N3934 = 1'b0 & N3933;
  assign N3935 = 1'b0 & N3932;
  assign N3936 = 1'b0 & N3931;
  assign N3937 = 1'b0 & N3930;
  assign N3938 = 1'b0 & N3929;
  assign N3939 = 1'b0 & N3928;
  assign N3940 = 1'b0 & N3927;
  assign N3941 = 1'b0 & N3926;
  assign N3942 = 1'b0 & N3925;
  assign N3943 = 1'b0 & N3924;
  assign N3944 = 1'b0 & N3923;
  assign N3945 = 1'b0 & N3922;
  assign N3946 = 1'b0 & N3921;
  assign N3947 = 1'b0 & N3920;
  assign N3948 = 1'b0 & N3919;
  assign N3949 = 1'b0 & N3918;
  assign N3950 = 1'b0 & N3917;
  assign N3951 = 1'b0 & N3916;
  assign N3952 = 1'b0 & N3915;
  assign N3953 = 1'b0 & N3914;
  assign N3954 = 1'b0 & N3913;
  assign N3955 = 1'b0 & N3912;
  assign N3956 = 1'b0 & N3911;
  assign N3957 = 1'b0 & N3910;
  assign N3958 = 1'b0 & N3909;
  assign N3959 = 1'b0 & N3908;
  assign N3960 = 1'b0 & N3907;
  assign N3961 = 1'b0 & N3906;
  assign N3962 = 1'b0 & N3905;
  assign N3963 = 1'b0 & N3904;
  assign N3964 = 1'b0 & N3903;
  assign N3965 = 1'b0 & N3902;
  assign N3966 = 1'b0 & N3901;
  assign N3967 = 1'b0 & N3900;
  assign N3968 = 1'b0 & N3899;
  assign N3969 = 1'b0 & N3898;
  assign N3970 = 1'b0 & N3897;
  assign N3971 = 1'b0 & N3896;
  assign N3972 = 1'b0 & N3895;
  assign N3973 = 1'b0 & N3894;
  assign N3974 = 1'b0 & N3893;
  assign N3975 = 1'b0 & N3892;
  assign N3976 = 1'b0 & N3891;
  assign N3977 = 1'b0 & N3890;
  assign N3978 = 1'b0 & N3889;
  assign N3979 = 1'b0 & N3888;
  assign N3980 = 1'b0 & N3887;
  assign N3981 = 1'b0 & N3886;
  assign N3982 = 1'b0 & N3885;
  assign N3983 = 1'b0 & N3884;
  assign N3984 = 1'b0 & N3883;
  assign N3985 = 1'b0 & N3882;
  assign N3986 = 1'b0 & N3881;
  assign N3987 = 1'b0 & N3880;
  assign N3988 = 1'b0 & N3879;
  assign N3989 = 1'b0 & N3878;
  assign N3990 = 1'b0 & N3877;
  assign N3991 = 1'b0 & N3876;
  assign N3992 = 1'b0 & N3875;
  assign N3993 = 1'b0 & N3874;
  assign N3994 = 1'b0 & N3873;
  assign N3995 = 1'b0 & N3872;
  assign N3996 = 1'b0 & N3871;
  assign N3997 = 1'b0 & N3870;
  assign N4062 = ~mhpmcounter_we[9];
  assign N4063 = 1'b0 & csr_wdata_int[31];
  assign N4064 = 1'b0 & csr_wdata_int[30];
  assign N4065 = 1'b0 & csr_wdata_int[29];
  assign N4066 = 1'b0 & csr_wdata_int[28];
  assign N4067 = 1'b0 & csr_wdata_int[27];
  assign N4068 = 1'b0 & csr_wdata_int[26];
  assign N4069 = 1'b0 & csr_wdata_int[25];
  assign N4070 = 1'b0 & csr_wdata_int[24];
  assign N4071 = 1'b0 & csr_wdata_int[23];
  assign N4072 = 1'b0 & csr_wdata_int[22];
  assign N4073 = 1'b0 & csr_wdata_int[21];
  assign N4074 = 1'b0 & csr_wdata_int[20];
  assign N4075 = 1'b0 & csr_wdata_int[19];
  assign N4076 = 1'b0 & csr_wdata_int[18];
  assign N4077 = 1'b0 & csr_wdata_int[17];
  assign N4078 = 1'b0 & csr_wdata_int[16];
  assign N4079 = 1'b0 & csr_wdata_int[15];
  assign N4080 = 1'b0 & csr_wdata_int[14];
  assign N4081 = 1'b0 & csr_wdata_int[13];
  assign N4082 = 1'b0 & csr_wdata_int[12];
  assign N4083 = 1'b0 & csr_wdata_int[11];
  assign N4084 = 1'b0 & csr_wdata_int[10];
  assign N4085 = 1'b0 & csr_wdata_int[9];
  assign N4086 = 1'b0 & csr_wdata_int[8];
  assign N4087 = 1'b0 & csr_wdata_int[7];
  assign N4088 = 1'b0 & csr_wdata_int[6];
  assign N4089 = 1'b0 & csr_wdata_int[5];
  assign N4090 = 1'b0 & csr_wdata_int[4];
  assign N4091 = 1'b0 & csr_wdata_int[3];
  assign N4092 = 1'b0 & csr_wdata_int[2];
  assign N4093 = 1'b0 & csr_wdata_int[1];
  assign N4094 = 1'b0 & csr_wdata_int[0];
  assign N4095 = ~mhpmcounterh_we[9];
  assign N4096 = 1'b0 & csr_wdata_int[31];
  assign N4097 = 1'b0 & csr_wdata_int[30];
  assign N4098 = 1'b0 & csr_wdata_int[29];
  assign N4099 = 1'b0 & csr_wdata_int[28];
  assign N4100 = 1'b0 & csr_wdata_int[27];
  assign N4101 = 1'b0 & csr_wdata_int[26];
  assign N4102 = 1'b0 & csr_wdata_int[25];
  assign N4103 = 1'b0 & csr_wdata_int[24];
  assign N4104 = 1'b0 & csr_wdata_int[23];
  assign N4105 = 1'b0 & csr_wdata_int[22];
  assign N4106 = 1'b0 & csr_wdata_int[21];
  assign N4107 = 1'b0 & csr_wdata_int[20];
  assign N4108 = 1'b0 & csr_wdata_int[19];
  assign N4109 = 1'b0 & csr_wdata_int[18];
  assign N4110 = 1'b0 & csr_wdata_int[17];
  assign N4111 = 1'b0 & csr_wdata_int[16];
  assign N4112 = 1'b0 & csr_wdata_int[15];
  assign N4113 = 1'b0 & csr_wdata_int[14];
  assign N4114 = 1'b0 & csr_wdata_int[13];
  assign N4115 = 1'b0 & csr_wdata_int[12];
  assign N4116 = 1'b0 & csr_wdata_int[11];
  assign N4117 = 1'b0 & csr_wdata_int[10];
  assign N4118 = 1'b0 & csr_wdata_int[9];
  assign N4119 = 1'b0 & csr_wdata_int[8];
  assign N4120 = 1'b0 & csr_wdata_int[7];
  assign N4121 = 1'b0 & csr_wdata_int[6];
  assign N4122 = 1'b0 & csr_wdata_int[5];
  assign N4123 = 1'b0 & csr_wdata_int[4];
  assign N4124 = 1'b0 & csr_wdata_int[3];
  assign N4125 = 1'b0 & csr_wdata_int[2];
  assign N4126 = 1'b0 & csr_wdata_int[1];
  assign N4127 = 1'b0 & csr_wdata_int[0];
  assign N4160 = 1'b0 & N10715;
  assign N10715 = ~mcountinhibit[10];
  assign N4161 = ~N4160;
  assign N4226 = 1'b0 & N4225;
  assign N4227 = 1'b0 & N4224;
  assign N4228 = 1'b0 & N4223;
  assign N4229 = 1'b0 & N4222;
  assign N4230 = 1'b0 & N4221;
  assign N4231 = 1'b0 & N4220;
  assign N4232 = 1'b0 & N4219;
  assign N4233 = 1'b0 & N4218;
  assign N4234 = 1'b0 & N4217;
  assign N4235 = 1'b0 & N4216;
  assign N4236 = 1'b0 & N4215;
  assign N4237 = 1'b0 & N4214;
  assign N4238 = 1'b0 & N4213;
  assign N4239 = 1'b0 & N4212;
  assign N4240 = 1'b0 & N4211;
  assign N4241 = 1'b0 & N4210;
  assign N4242 = 1'b0 & N4209;
  assign N4243 = 1'b0 & N4208;
  assign N4244 = 1'b0 & N4207;
  assign N4245 = 1'b0 & N4206;
  assign N4246 = 1'b0 & N4205;
  assign N4247 = 1'b0 & N4204;
  assign N4248 = 1'b0 & N4203;
  assign N4249 = 1'b0 & N4202;
  assign N4250 = 1'b0 & N4201;
  assign N4251 = 1'b0 & N4200;
  assign N4252 = 1'b0 & N4199;
  assign N4253 = 1'b0 & N4198;
  assign N4254 = 1'b0 & N4197;
  assign N4255 = 1'b0 & N4196;
  assign N4256 = 1'b0 & N4195;
  assign N4257 = 1'b0 & N4194;
  assign N4258 = 1'b0 & N4193;
  assign N4259 = 1'b0 & N4192;
  assign N4260 = 1'b0 & N4191;
  assign N4261 = 1'b0 & N4190;
  assign N4262 = 1'b0 & N4189;
  assign N4263 = 1'b0 & N4188;
  assign N4264 = 1'b0 & N4187;
  assign N4265 = 1'b0 & N4186;
  assign N4266 = 1'b0 & N4185;
  assign N4267 = 1'b0 & N4184;
  assign N4268 = 1'b0 & N4183;
  assign N4269 = 1'b0 & N4182;
  assign N4270 = 1'b0 & N4181;
  assign N4271 = 1'b0 & N4180;
  assign N4272 = 1'b0 & N4179;
  assign N4273 = 1'b0 & N4178;
  assign N4274 = 1'b0 & N4177;
  assign N4275 = 1'b0 & N4176;
  assign N4276 = 1'b0 & N4175;
  assign N4277 = 1'b0 & N4174;
  assign N4278 = 1'b0 & N4173;
  assign N4279 = 1'b0 & N4172;
  assign N4280 = 1'b0 & N4171;
  assign N4281 = 1'b0 & N4170;
  assign N4282 = 1'b0 & N4169;
  assign N4283 = 1'b0 & N4168;
  assign N4284 = 1'b0 & N4167;
  assign N4285 = 1'b0 & N4166;
  assign N4286 = 1'b0 & N4165;
  assign N4287 = 1'b0 & N4164;
  assign N4288 = 1'b0 & N4163;
  assign N4289 = 1'b0 & N4162;
  assign N4354 = ~mhpmcounter_we[10];
  assign N4355 = 1'b0 & csr_wdata_int[31];
  assign N4356 = 1'b0 & csr_wdata_int[30];
  assign N4357 = 1'b0 & csr_wdata_int[29];
  assign N4358 = 1'b0 & csr_wdata_int[28];
  assign N4359 = 1'b0 & csr_wdata_int[27];
  assign N4360 = 1'b0 & csr_wdata_int[26];
  assign N4361 = 1'b0 & csr_wdata_int[25];
  assign N4362 = 1'b0 & csr_wdata_int[24];
  assign N4363 = 1'b0 & csr_wdata_int[23];
  assign N4364 = 1'b0 & csr_wdata_int[22];
  assign N4365 = 1'b0 & csr_wdata_int[21];
  assign N4366 = 1'b0 & csr_wdata_int[20];
  assign N4367 = 1'b0 & csr_wdata_int[19];
  assign N4368 = 1'b0 & csr_wdata_int[18];
  assign N4369 = 1'b0 & csr_wdata_int[17];
  assign N4370 = 1'b0 & csr_wdata_int[16];
  assign N4371 = 1'b0 & csr_wdata_int[15];
  assign N4372 = 1'b0 & csr_wdata_int[14];
  assign N4373 = 1'b0 & csr_wdata_int[13];
  assign N4374 = 1'b0 & csr_wdata_int[12];
  assign N4375 = 1'b0 & csr_wdata_int[11];
  assign N4376 = 1'b0 & csr_wdata_int[10];
  assign N4377 = 1'b0 & csr_wdata_int[9];
  assign N4378 = 1'b0 & csr_wdata_int[8];
  assign N4379 = 1'b0 & csr_wdata_int[7];
  assign N4380 = 1'b0 & csr_wdata_int[6];
  assign N4381 = 1'b0 & csr_wdata_int[5];
  assign N4382 = 1'b0 & csr_wdata_int[4];
  assign N4383 = 1'b0 & csr_wdata_int[3];
  assign N4384 = 1'b0 & csr_wdata_int[2];
  assign N4385 = 1'b0 & csr_wdata_int[1];
  assign N4386 = 1'b0 & csr_wdata_int[0];
  assign N4387 = ~mhpmcounterh_we[10];
  assign N4388 = 1'b0 & csr_wdata_int[31];
  assign N4389 = 1'b0 & csr_wdata_int[30];
  assign N4390 = 1'b0 & csr_wdata_int[29];
  assign N4391 = 1'b0 & csr_wdata_int[28];
  assign N4392 = 1'b0 & csr_wdata_int[27];
  assign N4393 = 1'b0 & csr_wdata_int[26];
  assign N4394 = 1'b0 & csr_wdata_int[25];
  assign N4395 = 1'b0 & csr_wdata_int[24];
  assign N4396 = 1'b0 & csr_wdata_int[23];
  assign N4397 = 1'b0 & csr_wdata_int[22];
  assign N4398 = 1'b0 & csr_wdata_int[21];
  assign N4399 = 1'b0 & csr_wdata_int[20];
  assign N4400 = 1'b0 & csr_wdata_int[19];
  assign N4401 = 1'b0 & csr_wdata_int[18];
  assign N4402 = 1'b0 & csr_wdata_int[17];
  assign N4403 = 1'b0 & csr_wdata_int[16];
  assign N4404 = 1'b0 & csr_wdata_int[15];
  assign N4405 = 1'b0 & csr_wdata_int[14];
  assign N4406 = 1'b0 & csr_wdata_int[13];
  assign N4407 = 1'b0 & csr_wdata_int[12];
  assign N4408 = 1'b0 & csr_wdata_int[11];
  assign N4409 = 1'b0 & csr_wdata_int[10];
  assign N4410 = 1'b0 & csr_wdata_int[9];
  assign N4411 = 1'b0 & csr_wdata_int[8];
  assign N4412 = 1'b0 & csr_wdata_int[7];
  assign N4413 = 1'b0 & csr_wdata_int[6];
  assign N4414 = 1'b0 & csr_wdata_int[5];
  assign N4415 = 1'b0 & csr_wdata_int[4];
  assign N4416 = 1'b0 & csr_wdata_int[3];
  assign N4417 = 1'b0 & csr_wdata_int[2];
  assign N4418 = 1'b0 & csr_wdata_int[1];
  assign N4419 = 1'b0 & csr_wdata_int[0];
  assign N4452 = 1'b0 & N10716;
  assign N10716 = ~mcountinhibit[11];
  assign N4453 = ~N4452;
  assign N4518 = 1'b0 & N4517;
  assign N4519 = 1'b0 & N4516;
  assign N4520 = 1'b0 & N4515;
  assign N4521 = 1'b0 & N4514;
  assign N4522 = 1'b0 & N4513;
  assign N4523 = 1'b0 & N4512;
  assign N4524 = 1'b0 & N4511;
  assign N4525 = 1'b0 & N4510;
  assign N4526 = 1'b0 & N4509;
  assign N4527 = 1'b0 & N4508;
  assign N4528 = 1'b0 & N4507;
  assign N4529 = 1'b0 & N4506;
  assign N4530 = 1'b0 & N4505;
  assign N4531 = 1'b0 & N4504;
  assign N4532 = 1'b0 & N4503;
  assign N4533 = 1'b0 & N4502;
  assign N4534 = 1'b0 & N4501;
  assign N4535 = 1'b0 & N4500;
  assign N4536 = 1'b0 & N4499;
  assign N4537 = 1'b0 & N4498;
  assign N4538 = 1'b0 & N4497;
  assign N4539 = 1'b0 & N4496;
  assign N4540 = 1'b0 & N4495;
  assign N4541 = 1'b0 & N4494;
  assign N4542 = 1'b0 & N4493;
  assign N4543 = 1'b0 & N4492;
  assign N4544 = 1'b0 & N4491;
  assign N4545 = 1'b0 & N4490;
  assign N4546 = 1'b0 & N4489;
  assign N4547 = 1'b0 & N4488;
  assign N4548 = 1'b0 & N4487;
  assign N4549 = 1'b0 & N4486;
  assign N4550 = 1'b0 & N4485;
  assign N4551 = 1'b0 & N4484;
  assign N4552 = 1'b0 & N4483;
  assign N4553 = 1'b0 & N4482;
  assign N4554 = 1'b0 & N4481;
  assign N4555 = 1'b0 & N4480;
  assign N4556 = 1'b0 & N4479;
  assign N4557 = 1'b0 & N4478;
  assign N4558 = 1'b0 & N4477;
  assign N4559 = 1'b0 & N4476;
  assign N4560 = 1'b0 & N4475;
  assign N4561 = 1'b0 & N4474;
  assign N4562 = 1'b0 & N4473;
  assign N4563 = 1'b0 & N4472;
  assign N4564 = 1'b0 & N4471;
  assign N4565 = 1'b0 & N4470;
  assign N4566 = 1'b0 & N4469;
  assign N4567 = 1'b0 & N4468;
  assign N4568 = 1'b0 & N4467;
  assign N4569 = 1'b0 & N4466;
  assign N4570 = 1'b0 & N4465;
  assign N4571 = 1'b0 & N4464;
  assign N4572 = 1'b0 & N4463;
  assign N4573 = 1'b0 & N4462;
  assign N4574 = 1'b0 & N4461;
  assign N4575 = 1'b0 & N4460;
  assign N4576 = 1'b0 & N4459;
  assign N4577 = 1'b0 & N4458;
  assign N4578 = 1'b0 & N4457;
  assign N4579 = 1'b0 & N4456;
  assign N4580 = 1'b0 & N4455;
  assign N4581 = 1'b0 & N4454;
  assign N4646 = ~mhpmcounter_we[11];
  assign N4647 = 1'b0 & csr_wdata_int[31];
  assign N4648 = 1'b0 & csr_wdata_int[30];
  assign N4649 = 1'b0 & csr_wdata_int[29];
  assign N4650 = 1'b0 & csr_wdata_int[28];
  assign N4651 = 1'b0 & csr_wdata_int[27];
  assign N4652 = 1'b0 & csr_wdata_int[26];
  assign N4653 = 1'b0 & csr_wdata_int[25];
  assign N4654 = 1'b0 & csr_wdata_int[24];
  assign N4655 = 1'b0 & csr_wdata_int[23];
  assign N4656 = 1'b0 & csr_wdata_int[22];
  assign N4657 = 1'b0 & csr_wdata_int[21];
  assign N4658 = 1'b0 & csr_wdata_int[20];
  assign N4659 = 1'b0 & csr_wdata_int[19];
  assign N4660 = 1'b0 & csr_wdata_int[18];
  assign N4661 = 1'b0 & csr_wdata_int[17];
  assign N4662 = 1'b0 & csr_wdata_int[16];
  assign N4663 = 1'b0 & csr_wdata_int[15];
  assign N4664 = 1'b0 & csr_wdata_int[14];
  assign N4665 = 1'b0 & csr_wdata_int[13];
  assign N4666 = 1'b0 & csr_wdata_int[12];
  assign N4667 = 1'b0 & csr_wdata_int[11];
  assign N4668 = 1'b0 & csr_wdata_int[10];
  assign N4669 = 1'b0 & csr_wdata_int[9];
  assign N4670 = 1'b0 & csr_wdata_int[8];
  assign N4671 = 1'b0 & csr_wdata_int[7];
  assign N4672 = 1'b0 & csr_wdata_int[6];
  assign N4673 = 1'b0 & csr_wdata_int[5];
  assign N4674 = 1'b0 & csr_wdata_int[4];
  assign N4675 = 1'b0 & csr_wdata_int[3];
  assign N4676 = 1'b0 & csr_wdata_int[2];
  assign N4677 = 1'b0 & csr_wdata_int[1];
  assign N4678 = 1'b0 & csr_wdata_int[0];
  assign N4679 = ~mhpmcounterh_we[11];
  assign N4680 = 1'b0 & csr_wdata_int[31];
  assign N4681 = 1'b0 & csr_wdata_int[30];
  assign N4682 = 1'b0 & csr_wdata_int[29];
  assign N4683 = 1'b0 & csr_wdata_int[28];
  assign N4684 = 1'b0 & csr_wdata_int[27];
  assign N4685 = 1'b0 & csr_wdata_int[26];
  assign N4686 = 1'b0 & csr_wdata_int[25];
  assign N4687 = 1'b0 & csr_wdata_int[24];
  assign N4688 = 1'b0 & csr_wdata_int[23];
  assign N4689 = 1'b0 & csr_wdata_int[22];
  assign N4690 = 1'b0 & csr_wdata_int[21];
  assign N4691 = 1'b0 & csr_wdata_int[20];
  assign N4692 = 1'b0 & csr_wdata_int[19];
  assign N4693 = 1'b0 & csr_wdata_int[18];
  assign N4694 = 1'b0 & csr_wdata_int[17];
  assign N4695 = 1'b0 & csr_wdata_int[16];
  assign N4696 = 1'b0 & csr_wdata_int[15];
  assign N4697 = 1'b0 & csr_wdata_int[14];
  assign N4698 = 1'b0 & csr_wdata_int[13];
  assign N4699 = 1'b0 & csr_wdata_int[12];
  assign N4700 = 1'b0 & csr_wdata_int[11];
  assign N4701 = 1'b0 & csr_wdata_int[10];
  assign N4702 = 1'b0 & csr_wdata_int[9];
  assign N4703 = 1'b0 & csr_wdata_int[8];
  assign N4704 = 1'b0 & csr_wdata_int[7];
  assign N4705 = 1'b0 & csr_wdata_int[6];
  assign N4706 = 1'b0 & csr_wdata_int[5];
  assign N4707 = 1'b0 & csr_wdata_int[4];
  assign N4708 = 1'b0 & csr_wdata_int[3];
  assign N4709 = 1'b0 & csr_wdata_int[2];
  assign N4710 = 1'b0 & csr_wdata_int[1];
  assign N4711 = 1'b0 & csr_wdata_int[0];
  assign N4744 = 1'b0 & N10717;
  assign N10717 = ~mcountinhibit[12];
  assign N4745 = ~N4744;
  assign N4810 = 1'b0 & N4809;
  assign N4811 = 1'b0 & N4808;
  assign N4812 = 1'b0 & N4807;
  assign N4813 = 1'b0 & N4806;
  assign N4814 = 1'b0 & N4805;
  assign N4815 = 1'b0 & N4804;
  assign N4816 = 1'b0 & N4803;
  assign N4817 = 1'b0 & N4802;
  assign N4818 = 1'b0 & N4801;
  assign N4819 = 1'b0 & N4800;
  assign N4820 = 1'b0 & N4799;
  assign N4821 = 1'b0 & N4798;
  assign N4822 = 1'b0 & N4797;
  assign N4823 = 1'b0 & N4796;
  assign N4824 = 1'b0 & N4795;
  assign N4825 = 1'b0 & N4794;
  assign N4826 = 1'b0 & N4793;
  assign N4827 = 1'b0 & N4792;
  assign N4828 = 1'b0 & N4791;
  assign N4829 = 1'b0 & N4790;
  assign N4830 = 1'b0 & N4789;
  assign N4831 = 1'b0 & N4788;
  assign N4832 = 1'b0 & N4787;
  assign N4833 = 1'b0 & N4786;
  assign N4834 = 1'b0 & N4785;
  assign N4835 = 1'b0 & N4784;
  assign N4836 = 1'b0 & N4783;
  assign N4837 = 1'b0 & N4782;
  assign N4838 = 1'b0 & N4781;
  assign N4839 = 1'b0 & N4780;
  assign N4840 = 1'b0 & N4779;
  assign N4841 = 1'b0 & N4778;
  assign N4842 = 1'b0 & N4777;
  assign N4843 = 1'b0 & N4776;
  assign N4844 = 1'b0 & N4775;
  assign N4845 = 1'b0 & N4774;
  assign N4846 = 1'b0 & N4773;
  assign N4847 = 1'b0 & N4772;
  assign N4848 = 1'b0 & N4771;
  assign N4849 = 1'b0 & N4770;
  assign N4850 = 1'b0 & N4769;
  assign N4851 = 1'b0 & N4768;
  assign N4852 = 1'b0 & N4767;
  assign N4853 = 1'b0 & N4766;
  assign N4854 = 1'b0 & N4765;
  assign N4855 = 1'b0 & N4764;
  assign N4856 = 1'b0 & N4763;
  assign N4857 = 1'b0 & N4762;
  assign N4858 = 1'b0 & N4761;
  assign N4859 = 1'b0 & N4760;
  assign N4860 = 1'b0 & N4759;
  assign N4861 = 1'b0 & N4758;
  assign N4862 = 1'b0 & N4757;
  assign N4863 = 1'b0 & N4756;
  assign N4864 = 1'b0 & N4755;
  assign N4865 = 1'b0 & N4754;
  assign N4866 = 1'b0 & N4753;
  assign N4867 = 1'b0 & N4752;
  assign N4868 = 1'b0 & N4751;
  assign N4869 = 1'b0 & N4750;
  assign N4870 = 1'b0 & N4749;
  assign N4871 = 1'b0 & N4748;
  assign N4872 = 1'b0 & N4747;
  assign N4873 = 1'b0 & N4746;
  assign N4938 = ~mhpmcounter_we[12];
  assign N4939 = 1'b0 & csr_wdata_int[31];
  assign N4940 = 1'b0 & csr_wdata_int[30];
  assign N4941 = 1'b0 & csr_wdata_int[29];
  assign N4942 = 1'b0 & csr_wdata_int[28];
  assign N4943 = 1'b0 & csr_wdata_int[27];
  assign N4944 = 1'b0 & csr_wdata_int[26];
  assign N4945 = 1'b0 & csr_wdata_int[25];
  assign N4946 = 1'b0 & csr_wdata_int[24];
  assign N4947 = 1'b0 & csr_wdata_int[23];
  assign N4948 = 1'b0 & csr_wdata_int[22];
  assign N4949 = 1'b0 & csr_wdata_int[21];
  assign N4950 = 1'b0 & csr_wdata_int[20];
  assign N4951 = 1'b0 & csr_wdata_int[19];
  assign N4952 = 1'b0 & csr_wdata_int[18];
  assign N4953 = 1'b0 & csr_wdata_int[17];
  assign N4954 = 1'b0 & csr_wdata_int[16];
  assign N4955 = 1'b0 & csr_wdata_int[15];
  assign N4956 = 1'b0 & csr_wdata_int[14];
  assign N4957 = 1'b0 & csr_wdata_int[13];
  assign N4958 = 1'b0 & csr_wdata_int[12];
  assign N4959 = 1'b0 & csr_wdata_int[11];
  assign N4960 = 1'b0 & csr_wdata_int[10];
  assign N4961 = 1'b0 & csr_wdata_int[9];
  assign N4962 = 1'b0 & csr_wdata_int[8];
  assign N4963 = 1'b0 & csr_wdata_int[7];
  assign N4964 = 1'b0 & csr_wdata_int[6];
  assign N4965 = 1'b0 & csr_wdata_int[5];
  assign N4966 = 1'b0 & csr_wdata_int[4];
  assign N4967 = 1'b0 & csr_wdata_int[3];
  assign N4968 = 1'b0 & csr_wdata_int[2];
  assign N4969 = 1'b0 & csr_wdata_int[1];
  assign N4970 = 1'b0 & csr_wdata_int[0];
  assign N4971 = ~mhpmcounterh_we[12];
  assign N4972 = 1'b0 & csr_wdata_int[31];
  assign N4973 = 1'b0 & csr_wdata_int[30];
  assign N4974 = 1'b0 & csr_wdata_int[29];
  assign N4975 = 1'b0 & csr_wdata_int[28];
  assign N4976 = 1'b0 & csr_wdata_int[27];
  assign N4977 = 1'b0 & csr_wdata_int[26];
  assign N4978 = 1'b0 & csr_wdata_int[25];
  assign N4979 = 1'b0 & csr_wdata_int[24];
  assign N4980 = 1'b0 & csr_wdata_int[23];
  assign N4981 = 1'b0 & csr_wdata_int[22];
  assign N4982 = 1'b0 & csr_wdata_int[21];
  assign N4983 = 1'b0 & csr_wdata_int[20];
  assign N4984 = 1'b0 & csr_wdata_int[19];
  assign N4985 = 1'b0 & csr_wdata_int[18];
  assign N4986 = 1'b0 & csr_wdata_int[17];
  assign N4987 = 1'b0 & csr_wdata_int[16];
  assign N4988 = 1'b0 & csr_wdata_int[15];
  assign N4989 = 1'b0 & csr_wdata_int[14];
  assign N4990 = 1'b0 & csr_wdata_int[13];
  assign N4991 = 1'b0 & csr_wdata_int[12];
  assign N4992 = 1'b0 & csr_wdata_int[11];
  assign N4993 = 1'b0 & csr_wdata_int[10];
  assign N4994 = 1'b0 & csr_wdata_int[9];
  assign N4995 = 1'b0 & csr_wdata_int[8];
  assign N4996 = 1'b0 & csr_wdata_int[7];
  assign N4997 = 1'b0 & csr_wdata_int[6];
  assign N4998 = 1'b0 & csr_wdata_int[5];
  assign N4999 = 1'b0 & csr_wdata_int[4];
  assign N5000 = 1'b0 & csr_wdata_int[3];
  assign N5001 = 1'b0 & csr_wdata_int[2];
  assign N5002 = 1'b0 & csr_wdata_int[1];
  assign N5003 = 1'b0 & csr_wdata_int[0];
  assign N5036 = 1'b0 & N10718;
  assign N10718 = ~mcountinhibit[13];
  assign N5037 = ~N5036;
  assign N5102 = 1'b0 & N5101;
  assign N5103 = 1'b0 & N5100;
  assign N5104 = 1'b0 & N5099;
  assign N5105 = 1'b0 & N5098;
  assign N5106 = 1'b0 & N5097;
  assign N5107 = 1'b0 & N5096;
  assign N5108 = 1'b0 & N5095;
  assign N5109 = 1'b0 & N5094;
  assign N5110 = 1'b0 & N5093;
  assign N5111 = 1'b0 & N5092;
  assign N5112 = 1'b0 & N5091;
  assign N5113 = 1'b0 & N5090;
  assign N5114 = 1'b0 & N5089;
  assign N5115 = 1'b0 & N5088;
  assign N5116 = 1'b0 & N5087;
  assign N5117 = 1'b0 & N5086;
  assign N5118 = 1'b0 & N5085;
  assign N5119 = 1'b0 & N5084;
  assign N5120 = 1'b0 & N5083;
  assign N5121 = 1'b0 & N5082;
  assign N5122 = 1'b0 & N5081;
  assign N5123 = 1'b0 & N5080;
  assign N5124 = 1'b0 & N5079;
  assign N5125 = 1'b0 & N5078;
  assign N5126 = 1'b0 & N5077;
  assign N5127 = 1'b0 & N5076;
  assign N5128 = 1'b0 & N5075;
  assign N5129 = 1'b0 & N5074;
  assign N5130 = 1'b0 & N5073;
  assign N5131 = 1'b0 & N5072;
  assign N5132 = 1'b0 & N5071;
  assign N5133 = 1'b0 & N5070;
  assign N5134 = 1'b0 & N5069;
  assign N5135 = 1'b0 & N5068;
  assign N5136 = 1'b0 & N5067;
  assign N5137 = 1'b0 & N5066;
  assign N5138 = 1'b0 & N5065;
  assign N5139 = 1'b0 & N5064;
  assign N5140 = 1'b0 & N5063;
  assign N5141 = 1'b0 & N5062;
  assign N5142 = 1'b0 & N5061;
  assign N5143 = 1'b0 & N5060;
  assign N5144 = 1'b0 & N5059;
  assign N5145 = 1'b0 & N5058;
  assign N5146 = 1'b0 & N5057;
  assign N5147 = 1'b0 & N5056;
  assign N5148 = 1'b0 & N5055;
  assign N5149 = 1'b0 & N5054;
  assign N5150 = 1'b0 & N5053;
  assign N5151 = 1'b0 & N5052;
  assign N5152 = 1'b0 & N5051;
  assign N5153 = 1'b0 & N5050;
  assign N5154 = 1'b0 & N5049;
  assign N5155 = 1'b0 & N5048;
  assign N5156 = 1'b0 & N5047;
  assign N5157 = 1'b0 & N5046;
  assign N5158 = 1'b0 & N5045;
  assign N5159 = 1'b0 & N5044;
  assign N5160 = 1'b0 & N5043;
  assign N5161 = 1'b0 & N5042;
  assign N5162 = 1'b0 & N5041;
  assign N5163 = 1'b0 & N5040;
  assign N5164 = 1'b0 & N5039;
  assign N5165 = 1'b0 & N5038;
  assign N5230 = ~mhpmcounter_we[13];
  assign N5231 = 1'b0 & csr_wdata_int[31];
  assign N5232 = 1'b0 & csr_wdata_int[30];
  assign N5233 = 1'b0 & csr_wdata_int[29];
  assign N5234 = 1'b0 & csr_wdata_int[28];
  assign N5235 = 1'b0 & csr_wdata_int[27];
  assign N5236 = 1'b0 & csr_wdata_int[26];
  assign N5237 = 1'b0 & csr_wdata_int[25];
  assign N5238 = 1'b0 & csr_wdata_int[24];
  assign N5239 = 1'b0 & csr_wdata_int[23];
  assign N5240 = 1'b0 & csr_wdata_int[22];
  assign N5241 = 1'b0 & csr_wdata_int[21];
  assign N5242 = 1'b0 & csr_wdata_int[20];
  assign N5243 = 1'b0 & csr_wdata_int[19];
  assign N5244 = 1'b0 & csr_wdata_int[18];
  assign N5245 = 1'b0 & csr_wdata_int[17];
  assign N5246 = 1'b0 & csr_wdata_int[16];
  assign N5247 = 1'b0 & csr_wdata_int[15];
  assign N5248 = 1'b0 & csr_wdata_int[14];
  assign N5249 = 1'b0 & csr_wdata_int[13];
  assign N5250 = 1'b0 & csr_wdata_int[12];
  assign N5251 = 1'b0 & csr_wdata_int[11];
  assign N5252 = 1'b0 & csr_wdata_int[10];
  assign N5253 = 1'b0 & csr_wdata_int[9];
  assign N5254 = 1'b0 & csr_wdata_int[8];
  assign N5255 = 1'b0 & csr_wdata_int[7];
  assign N5256 = 1'b0 & csr_wdata_int[6];
  assign N5257 = 1'b0 & csr_wdata_int[5];
  assign N5258 = 1'b0 & csr_wdata_int[4];
  assign N5259 = 1'b0 & csr_wdata_int[3];
  assign N5260 = 1'b0 & csr_wdata_int[2];
  assign N5261 = 1'b0 & csr_wdata_int[1];
  assign N5262 = 1'b0 & csr_wdata_int[0];
  assign N5263 = ~mhpmcounterh_we[13];
  assign N5264 = 1'b0 & csr_wdata_int[31];
  assign N5265 = 1'b0 & csr_wdata_int[30];
  assign N5266 = 1'b0 & csr_wdata_int[29];
  assign N5267 = 1'b0 & csr_wdata_int[28];
  assign N5268 = 1'b0 & csr_wdata_int[27];
  assign N5269 = 1'b0 & csr_wdata_int[26];
  assign N5270 = 1'b0 & csr_wdata_int[25];
  assign N5271 = 1'b0 & csr_wdata_int[24];
  assign N5272 = 1'b0 & csr_wdata_int[23];
  assign N5273 = 1'b0 & csr_wdata_int[22];
  assign N5274 = 1'b0 & csr_wdata_int[21];
  assign N5275 = 1'b0 & csr_wdata_int[20];
  assign N5276 = 1'b0 & csr_wdata_int[19];
  assign N5277 = 1'b0 & csr_wdata_int[18];
  assign N5278 = 1'b0 & csr_wdata_int[17];
  assign N5279 = 1'b0 & csr_wdata_int[16];
  assign N5280 = 1'b0 & csr_wdata_int[15];
  assign N5281 = 1'b0 & csr_wdata_int[14];
  assign N5282 = 1'b0 & csr_wdata_int[13];
  assign N5283 = 1'b0 & csr_wdata_int[12];
  assign N5284 = 1'b0 & csr_wdata_int[11];
  assign N5285 = 1'b0 & csr_wdata_int[10];
  assign N5286 = 1'b0 & csr_wdata_int[9];
  assign N5287 = 1'b0 & csr_wdata_int[8];
  assign N5288 = 1'b0 & csr_wdata_int[7];
  assign N5289 = 1'b0 & csr_wdata_int[6];
  assign N5290 = 1'b0 & csr_wdata_int[5];
  assign N5291 = 1'b0 & csr_wdata_int[4];
  assign N5292 = 1'b0 & csr_wdata_int[3];
  assign N5293 = 1'b0 & csr_wdata_int[2];
  assign N5294 = 1'b0 & csr_wdata_int[1];
  assign N5295 = 1'b0 & csr_wdata_int[0];
  assign N5328 = 1'b0 & N10719;
  assign N10719 = ~mcountinhibit[14];
  assign N5329 = ~N5328;
  assign N5394 = 1'b0 & N5393;
  assign N5395 = 1'b0 & N5392;
  assign N5396 = 1'b0 & N5391;
  assign N5397 = 1'b0 & N5390;
  assign N5398 = 1'b0 & N5389;
  assign N5399 = 1'b0 & N5388;
  assign N5400 = 1'b0 & N5387;
  assign N5401 = 1'b0 & N5386;
  assign N5402 = 1'b0 & N5385;
  assign N5403 = 1'b0 & N5384;
  assign N5404 = 1'b0 & N5383;
  assign N5405 = 1'b0 & N5382;
  assign N5406 = 1'b0 & N5381;
  assign N5407 = 1'b0 & N5380;
  assign N5408 = 1'b0 & N5379;
  assign N5409 = 1'b0 & N5378;
  assign N5410 = 1'b0 & N5377;
  assign N5411 = 1'b0 & N5376;
  assign N5412 = 1'b0 & N5375;
  assign N5413 = 1'b0 & N5374;
  assign N5414 = 1'b0 & N5373;
  assign N5415 = 1'b0 & N5372;
  assign N5416 = 1'b0 & N5371;
  assign N5417 = 1'b0 & N5370;
  assign N5418 = 1'b0 & N5369;
  assign N5419 = 1'b0 & N5368;
  assign N5420 = 1'b0 & N5367;
  assign N5421 = 1'b0 & N5366;
  assign N5422 = 1'b0 & N5365;
  assign N5423 = 1'b0 & N5364;
  assign N5424 = 1'b0 & N5363;
  assign N5425 = 1'b0 & N5362;
  assign N5426 = 1'b0 & N5361;
  assign N5427 = 1'b0 & N5360;
  assign N5428 = 1'b0 & N5359;
  assign N5429 = 1'b0 & N5358;
  assign N5430 = 1'b0 & N5357;
  assign N5431 = 1'b0 & N5356;
  assign N5432 = 1'b0 & N5355;
  assign N5433 = 1'b0 & N5354;
  assign N5434 = 1'b0 & N5353;
  assign N5435 = 1'b0 & N5352;
  assign N5436 = 1'b0 & N5351;
  assign N5437 = 1'b0 & N5350;
  assign N5438 = 1'b0 & N5349;
  assign N5439 = 1'b0 & N5348;
  assign N5440 = 1'b0 & N5347;
  assign N5441 = 1'b0 & N5346;
  assign N5442 = 1'b0 & N5345;
  assign N5443 = 1'b0 & N5344;
  assign N5444 = 1'b0 & N5343;
  assign N5445 = 1'b0 & N5342;
  assign N5446 = 1'b0 & N5341;
  assign N5447 = 1'b0 & N5340;
  assign N5448 = 1'b0 & N5339;
  assign N5449 = 1'b0 & N5338;
  assign N5450 = 1'b0 & N5337;
  assign N5451 = 1'b0 & N5336;
  assign N5452 = 1'b0 & N5335;
  assign N5453 = 1'b0 & N5334;
  assign N5454 = 1'b0 & N5333;
  assign N5455 = 1'b0 & N5332;
  assign N5456 = 1'b0 & N5331;
  assign N5457 = 1'b0 & N5330;
  assign N5522 = ~mhpmcounter_we[14];
  assign N5523 = 1'b0 & csr_wdata_int[31];
  assign N5524 = 1'b0 & csr_wdata_int[30];
  assign N5525 = 1'b0 & csr_wdata_int[29];
  assign N5526 = 1'b0 & csr_wdata_int[28];
  assign N5527 = 1'b0 & csr_wdata_int[27];
  assign N5528 = 1'b0 & csr_wdata_int[26];
  assign N5529 = 1'b0 & csr_wdata_int[25];
  assign N5530 = 1'b0 & csr_wdata_int[24];
  assign N5531 = 1'b0 & csr_wdata_int[23];
  assign N5532 = 1'b0 & csr_wdata_int[22];
  assign N5533 = 1'b0 & csr_wdata_int[21];
  assign N5534 = 1'b0 & csr_wdata_int[20];
  assign N5535 = 1'b0 & csr_wdata_int[19];
  assign N5536 = 1'b0 & csr_wdata_int[18];
  assign N5537 = 1'b0 & csr_wdata_int[17];
  assign N5538 = 1'b0 & csr_wdata_int[16];
  assign N5539 = 1'b0 & csr_wdata_int[15];
  assign N5540 = 1'b0 & csr_wdata_int[14];
  assign N5541 = 1'b0 & csr_wdata_int[13];
  assign N5542 = 1'b0 & csr_wdata_int[12];
  assign N5543 = 1'b0 & csr_wdata_int[11];
  assign N5544 = 1'b0 & csr_wdata_int[10];
  assign N5545 = 1'b0 & csr_wdata_int[9];
  assign N5546 = 1'b0 & csr_wdata_int[8];
  assign N5547 = 1'b0 & csr_wdata_int[7];
  assign N5548 = 1'b0 & csr_wdata_int[6];
  assign N5549 = 1'b0 & csr_wdata_int[5];
  assign N5550 = 1'b0 & csr_wdata_int[4];
  assign N5551 = 1'b0 & csr_wdata_int[3];
  assign N5552 = 1'b0 & csr_wdata_int[2];
  assign N5553 = 1'b0 & csr_wdata_int[1];
  assign N5554 = 1'b0 & csr_wdata_int[0];
  assign N5555 = ~mhpmcounterh_we[14];
  assign N5556 = 1'b0 & csr_wdata_int[31];
  assign N5557 = 1'b0 & csr_wdata_int[30];
  assign N5558 = 1'b0 & csr_wdata_int[29];
  assign N5559 = 1'b0 & csr_wdata_int[28];
  assign N5560 = 1'b0 & csr_wdata_int[27];
  assign N5561 = 1'b0 & csr_wdata_int[26];
  assign N5562 = 1'b0 & csr_wdata_int[25];
  assign N5563 = 1'b0 & csr_wdata_int[24];
  assign N5564 = 1'b0 & csr_wdata_int[23];
  assign N5565 = 1'b0 & csr_wdata_int[22];
  assign N5566 = 1'b0 & csr_wdata_int[21];
  assign N5567 = 1'b0 & csr_wdata_int[20];
  assign N5568 = 1'b0 & csr_wdata_int[19];
  assign N5569 = 1'b0 & csr_wdata_int[18];
  assign N5570 = 1'b0 & csr_wdata_int[17];
  assign N5571 = 1'b0 & csr_wdata_int[16];
  assign N5572 = 1'b0 & csr_wdata_int[15];
  assign N5573 = 1'b0 & csr_wdata_int[14];
  assign N5574 = 1'b0 & csr_wdata_int[13];
  assign N5575 = 1'b0 & csr_wdata_int[12];
  assign N5576 = 1'b0 & csr_wdata_int[11];
  assign N5577 = 1'b0 & csr_wdata_int[10];
  assign N5578 = 1'b0 & csr_wdata_int[9];
  assign N5579 = 1'b0 & csr_wdata_int[8];
  assign N5580 = 1'b0 & csr_wdata_int[7];
  assign N5581 = 1'b0 & csr_wdata_int[6];
  assign N5582 = 1'b0 & csr_wdata_int[5];
  assign N5583 = 1'b0 & csr_wdata_int[4];
  assign N5584 = 1'b0 & csr_wdata_int[3];
  assign N5585 = 1'b0 & csr_wdata_int[2];
  assign N5586 = 1'b0 & csr_wdata_int[1];
  assign N5587 = 1'b0 & csr_wdata_int[0];
  assign N5620 = 1'b0 & N10720;
  assign N10720 = ~mcountinhibit[15];
  assign N5621 = ~N5620;
  assign N5686 = 1'b0 & N5685;
  assign N5687 = 1'b0 & N5684;
  assign N5688 = 1'b0 & N5683;
  assign N5689 = 1'b0 & N5682;
  assign N5690 = 1'b0 & N5681;
  assign N5691 = 1'b0 & N5680;
  assign N5692 = 1'b0 & N5679;
  assign N5693 = 1'b0 & N5678;
  assign N5694 = 1'b0 & N5677;
  assign N5695 = 1'b0 & N5676;
  assign N5696 = 1'b0 & N5675;
  assign N5697 = 1'b0 & N5674;
  assign N5698 = 1'b0 & N5673;
  assign N5699 = 1'b0 & N5672;
  assign N5700 = 1'b0 & N5671;
  assign N5701 = 1'b0 & N5670;
  assign N5702 = 1'b0 & N5669;
  assign N5703 = 1'b0 & N5668;
  assign N5704 = 1'b0 & N5667;
  assign N5705 = 1'b0 & N5666;
  assign N5706 = 1'b0 & N5665;
  assign N5707 = 1'b0 & N5664;
  assign N5708 = 1'b0 & N5663;
  assign N5709 = 1'b0 & N5662;
  assign N5710 = 1'b0 & N5661;
  assign N5711 = 1'b0 & N5660;
  assign N5712 = 1'b0 & N5659;
  assign N5713 = 1'b0 & N5658;
  assign N5714 = 1'b0 & N5657;
  assign N5715 = 1'b0 & N5656;
  assign N5716 = 1'b0 & N5655;
  assign N5717 = 1'b0 & N5654;
  assign N5718 = 1'b0 & N5653;
  assign N5719 = 1'b0 & N5652;
  assign N5720 = 1'b0 & N5651;
  assign N5721 = 1'b0 & N5650;
  assign N5722 = 1'b0 & N5649;
  assign N5723 = 1'b0 & N5648;
  assign N5724 = 1'b0 & N5647;
  assign N5725 = 1'b0 & N5646;
  assign N5726 = 1'b0 & N5645;
  assign N5727 = 1'b0 & N5644;
  assign N5728 = 1'b0 & N5643;
  assign N5729 = 1'b0 & N5642;
  assign N5730 = 1'b0 & N5641;
  assign N5731 = 1'b0 & N5640;
  assign N5732 = 1'b0 & N5639;
  assign N5733 = 1'b0 & N5638;
  assign N5734 = 1'b0 & N5637;
  assign N5735 = 1'b0 & N5636;
  assign N5736 = 1'b0 & N5635;
  assign N5737 = 1'b0 & N5634;
  assign N5738 = 1'b0 & N5633;
  assign N5739 = 1'b0 & N5632;
  assign N5740 = 1'b0 & N5631;
  assign N5741 = 1'b0 & N5630;
  assign N5742 = 1'b0 & N5629;
  assign N5743 = 1'b0 & N5628;
  assign N5744 = 1'b0 & N5627;
  assign N5745 = 1'b0 & N5626;
  assign N5746 = 1'b0 & N5625;
  assign N5747 = 1'b0 & N5624;
  assign N5748 = 1'b0 & N5623;
  assign N5749 = 1'b0 & N5622;
  assign N5814 = ~mhpmcounter_we[15];
  assign N5815 = 1'b0 & csr_wdata_int[31];
  assign N5816 = 1'b0 & csr_wdata_int[30];
  assign N5817 = 1'b0 & csr_wdata_int[29];
  assign N5818 = 1'b0 & csr_wdata_int[28];
  assign N5819 = 1'b0 & csr_wdata_int[27];
  assign N5820 = 1'b0 & csr_wdata_int[26];
  assign N5821 = 1'b0 & csr_wdata_int[25];
  assign N5822 = 1'b0 & csr_wdata_int[24];
  assign N5823 = 1'b0 & csr_wdata_int[23];
  assign N5824 = 1'b0 & csr_wdata_int[22];
  assign N5825 = 1'b0 & csr_wdata_int[21];
  assign N5826 = 1'b0 & csr_wdata_int[20];
  assign N5827 = 1'b0 & csr_wdata_int[19];
  assign N5828 = 1'b0 & csr_wdata_int[18];
  assign N5829 = 1'b0 & csr_wdata_int[17];
  assign N5830 = 1'b0 & csr_wdata_int[16];
  assign N5831 = 1'b0 & csr_wdata_int[15];
  assign N5832 = 1'b0 & csr_wdata_int[14];
  assign N5833 = 1'b0 & csr_wdata_int[13];
  assign N5834 = 1'b0 & csr_wdata_int[12];
  assign N5835 = 1'b0 & csr_wdata_int[11];
  assign N5836 = 1'b0 & csr_wdata_int[10];
  assign N5837 = 1'b0 & csr_wdata_int[9];
  assign N5838 = 1'b0 & csr_wdata_int[8];
  assign N5839 = 1'b0 & csr_wdata_int[7];
  assign N5840 = 1'b0 & csr_wdata_int[6];
  assign N5841 = 1'b0 & csr_wdata_int[5];
  assign N5842 = 1'b0 & csr_wdata_int[4];
  assign N5843 = 1'b0 & csr_wdata_int[3];
  assign N5844 = 1'b0 & csr_wdata_int[2];
  assign N5845 = 1'b0 & csr_wdata_int[1];
  assign N5846 = 1'b0 & csr_wdata_int[0];
  assign N5847 = ~mhpmcounterh_we[15];
  assign N5848 = 1'b0 & csr_wdata_int[31];
  assign N5849 = 1'b0 & csr_wdata_int[30];
  assign N5850 = 1'b0 & csr_wdata_int[29];
  assign N5851 = 1'b0 & csr_wdata_int[28];
  assign N5852 = 1'b0 & csr_wdata_int[27];
  assign N5853 = 1'b0 & csr_wdata_int[26];
  assign N5854 = 1'b0 & csr_wdata_int[25];
  assign N5855 = 1'b0 & csr_wdata_int[24];
  assign N5856 = 1'b0 & csr_wdata_int[23];
  assign N5857 = 1'b0 & csr_wdata_int[22];
  assign N5858 = 1'b0 & csr_wdata_int[21];
  assign N5859 = 1'b0 & csr_wdata_int[20];
  assign N5860 = 1'b0 & csr_wdata_int[19];
  assign N5861 = 1'b0 & csr_wdata_int[18];
  assign N5862 = 1'b0 & csr_wdata_int[17];
  assign N5863 = 1'b0 & csr_wdata_int[16];
  assign N5864 = 1'b0 & csr_wdata_int[15];
  assign N5865 = 1'b0 & csr_wdata_int[14];
  assign N5866 = 1'b0 & csr_wdata_int[13];
  assign N5867 = 1'b0 & csr_wdata_int[12];
  assign N5868 = 1'b0 & csr_wdata_int[11];
  assign N5869 = 1'b0 & csr_wdata_int[10];
  assign N5870 = 1'b0 & csr_wdata_int[9];
  assign N5871 = 1'b0 & csr_wdata_int[8];
  assign N5872 = 1'b0 & csr_wdata_int[7];
  assign N5873 = 1'b0 & csr_wdata_int[6];
  assign N5874 = 1'b0 & csr_wdata_int[5];
  assign N5875 = 1'b0 & csr_wdata_int[4];
  assign N5876 = 1'b0 & csr_wdata_int[3];
  assign N5877 = 1'b0 & csr_wdata_int[2];
  assign N5878 = 1'b0 & csr_wdata_int[1];
  assign N5879 = 1'b0 & csr_wdata_int[0];
  assign N5912 = 1'b0 & N10721;
  assign N10721 = ~mcountinhibit[16];
  assign N5913 = ~N5912;
  assign N5978 = 1'b0 & N5977;
  assign N5979 = 1'b0 & N5976;
  assign N5980 = 1'b0 & N5975;
  assign N5981 = 1'b0 & N5974;
  assign N5982 = 1'b0 & N5973;
  assign N5983 = 1'b0 & N5972;
  assign N5984 = 1'b0 & N5971;
  assign N5985 = 1'b0 & N5970;
  assign N5986 = 1'b0 & N5969;
  assign N5987 = 1'b0 & N5968;
  assign N5988 = 1'b0 & N5967;
  assign N5989 = 1'b0 & N5966;
  assign N5990 = 1'b0 & N5965;
  assign N5991 = 1'b0 & N5964;
  assign N5992 = 1'b0 & N5963;
  assign N5993 = 1'b0 & N5962;
  assign N5994 = 1'b0 & N5961;
  assign N5995 = 1'b0 & N5960;
  assign N5996 = 1'b0 & N5959;
  assign N5997 = 1'b0 & N5958;
  assign N5998 = 1'b0 & N5957;
  assign N5999 = 1'b0 & N5956;
  assign N6000 = 1'b0 & N5955;
  assign N6001 = 1'b0 & N5954;
  assign N6002 = 1'b0 & N5953;
  assign N6003 = 1'b0 & N5952;
  assign N6004 = 1'b0 & N5951;
  assign N6005 = 1'b0 & N5950;
  assign N6006 = 1'b0 & N5949;
  assign N6007 = 1'b0 & N5948;
  assign N6008 = 1'b0 & N5947;
  assign N6009 = 1'b0 & N5946;
  assign N6010 = 1'b0 & N5945;
  assign N6011 = 1'b0 & N5944;
  assign N6012 = 1'b0 & N5943;
  assign N6013 = 1'b0 & N5942;
  assign N6014 = 1'b0 & N5941;
  assign N6015 = 1'b0 & N5940;
  assign N6016 = 1'b0 & N5939;
  assign N6017 = 1'b0 & N5938;
  assign N6018 = 1'b0 & N5937;
  assign N6019 = 1'b0 & N5936;
  assign N6020 = 1'b0 & N5935;
  assign N6021 = 1'b0 & N5934;
  assign N6022 = 1'b0 & N5933;
  assign N6023 = 1'b0 & N5932;
  assign N6024 = 1'b0 & N5931;
  assign N6025 = 1'b0 & N5930;
  assign N6026 = 1'b0 & N5929;
  assign N6027 = 1'b0 & N5928;
  assign N6028 = 1'b0 & N5927;
  assign N6029 = 1'b0 & N5926;
  assign N6030 = 1'b0 & N5925;
  assign N6031 = 1'b0 & N5924;
  assign N6032 = 1'b0 & N5923;
  assign N6033 = 1'b0 & N5922;
  assign N6034 = 1'b0 & N5921;
  assign N6035 = 1'b0 & N5920;
  assign N6036 = 1'b0 & N5919;
  assign N6037 = 1'b0 & N5918;
  assign N6038 = 1'b0 & N5917;
  assign N6039 = 1'b0 & N5916;
  assign N6040 = 1'b0 & N5915;
  assign N6041 = 1'b0 & N5914;
  assign N6106 = ~mhpmcounter_we[16];
  assign N6107 = 1'b0 & csr_wdata_int[31];
  assign N6108 = 1'b0 & csr_wdata_int[30];
  assign N6109 = 1'b0 & csr_wdata_int[29];
  assign N6110 = 1'b0 & csr_wdata_int[28];
  assign N6111 = 1'b0 & csr_wdata_int[27];
  assign N6112 = 1'b0 & csr_wdata_int[26];
  assign N6113 = 1'b0 & csr_wdata_int[25];
  assign N6114 = 1'b0 & csr_wdata_int[24];
  assign N6115 = 1'b0 & csr_wdata_int[23];
  assign N6116 = 1'b0 & csr_wdata_int[22];
  assign N6117 = 1'b0 & csr_wdata_int[21];
  assign N6118 = 1'b0 & csr_wdata_int[20];
  assign N6119 = 1'b0 & csr_wdata_int[19];
  assign N6120 = 1'b0 & csr_wdata_int[18];
  assign N6121 = 1'b0 & csr_wdata_int[17];
  assign N6122 = 1'b0 & csr_wdata_int[16];
  assign N6123 = 1'b0 & csr_wdata_int[15];
  assign N6124 = 1'b0 & csr_wdata_int[14];
  assign N6125 = 1'b0 & csr_wdata_int[13];
  assign N6126 = 1'b0 & csr_wdata_int[12];
  assign N6127 = 1'b0 & csr_wdata_int[11];
  assign N6128 = 1'b0 & csr_wdata_int[10];
  assign N6129 = 1'b0 & csr_wdata_int[9];
  assign N6130 = 1'b0 & csr_wdata_int[8];
  assign N6131 = 1'b0 & csr_wdata_int[7];
  assign N6132 = 1'b0 & csr_wdata_int[6];
  assign N6133 = 1'b0 & csr_wdata_int[5];
  assign N6134 = 1'b0 & csr_wdata_int[4];
  assign N6135 = 1'b0 & csr_wdata_int[3];
  assign N6136 = 1'b0 & csr_wdata_int[2];
  assign N6137 = 1'b0 & csr_wdata_int[1];
  assign N6138 = 1'b0 & csr_wdata_int[0];
  assign N6139 = ~mhpmcounterh_we[16];
  assign N6140 = 1'b0 & csr_wdata_int[31];
  assign N6141 = 1'b0 & csr_wdata_int[30];
  assign N6142 = 1'b0 & csr_wdata_int[29];
  assign N6143 = 1'b0 & csr_wdata_int[28];
  assign N6144 = 1'b0 & csr_wdata_int[27];
  assign N6145 = 1'b0 & csr_wdata_int[26];
  assign N6146 = 1'b0 & csr_wdata_int[25];
  assign N6147 = 1'b0 & csr_wdata_int[24];
  assign N6148 = 1'b0 & csr_wdata_int[23];
  assign N6149 = 1'b0 & csr_wdata_int[22];
  assign N6150 = 1'b0 & csr_wdata_int[21];
  assign N6151 = 1'b0 & csr_wdata_int[20];
  assign N6152 = 1'b0 & csr_wdata_int[19];
  assign N6153 = 1'b0 & csr_wdata_int[18];
  assign N6154 = 1'b0 & csr_wdata_int[17];
  assign N6155 = 1'b0 & csr_wdata_int[16];
  assign N6156 = 1'b0 & csr_wdata_int[15];
  assign N6157 = 1'b0 & csr_wdata_int[14];
  assign N6158 = 1'b0 & csr_wdata_int[13];
  assign N6159 = 1'b0 & csr_wdata_int[12];
  assign N6160 = 1'b0 & csr_wdata_int[11];
  assign N6161 = 1'b0 & csr_wdata_int[10];
  assign N6162 = 1'b0 & csr_wdata_int[9];
  assign N6163 = 1'b0 & csr_wdata_int[8];
  assign N6164 = 1'b0 & csr_wdata_int[7];
  assign N6165 = 1'b0 & csr_wdata_int[6];
  assign N6166 = 1'b0 & csr_wdata_int[5];
  assign N6167 = 1'b0 & csr_wdata_int[4];
  assign N6168 = 1'b0 & csr_wdata_int[3];
  assign N6169 = 1'b0 & csr_wdata_int[2];
  assign N6170 = 1'b0 & csr_wdata_int[1];
  assign N6171 = 1'b0 & csr_wdata_int[0];
  assign N6204 = 1'b0 & N10722;
  assign N10722 = ~mcountinhibit[17];
  assign N6205 = ~N6204;
  assign N6270 = 1'b0 & N6269;
  assign N6271 = 1'b0 & N6268;
  assign N6272 = 1'b0 & N6267;
  assign N6273 = 1'b0 & N6266;
  assign N6274 = 1'b0 & N6265;
  assign N6275 = 1'b0 & N6264;
  assign N6276 = 1'b0 & N6263;
  assign N6277 = 1'b0 & N6262;
  assign N6278 = 1'b0 & N6261;
  assign N6279 = 1'b0 & N6260;
  assign N6280 = 1'b0 & N6259;
  assign N6281 = 1'b0 & N6258;
  assign N6282 = 1'b0 & N6257;
  assign N6283 = 1'b0 & N6256;
  assign N6284 = 1'b0 & N6255;
  assign N6285 = 1'b0 & N6254;
  assign N6286 = 1'b0 & N6253;
  assign N6287 = 1'b0 & N6252;
  assign N6288 = 1'b0 & N6251;
  assign N6289 = 1'b0 & N6250;
  assign N6290 = 1'b0 & N6249;
  assign N6291 = 1'b0 & N6248;
  assign N6292 = 1'b0 & N6247;
  assign N6293 = 1'b0 & N6246;
  assign N6294 = 1'b0 & N6245;
  assign N6295 = 1'b0 & N6244;
  assign N6296 = 1'b0 & N6243;
  assign N6297 = 1'b0 & N6242;
  assign N6298 = 1'b0 & N6241;
  assign N6299 = 1'b0 & N6240;
  assign N6300 = 1'b0 & N6239;
  assign N6301 = 1'b0 & N6238;
  assign N6302 = 1'b0 & N6237;
  assign N6303 = 1'b0 & N6236;
  assign N6304 = 1'b0 & N6235;
  assign N6305 = 1'b0 & N6234;
  assign N6306 = 1'b0 & N6233;
  assign N6307 = 1'b0 & N6232;
  assign N6308 = 1'b0 & N6231;
  assign N6309 = 1'b0 & N6230;
  assign N6310 = 1'b0 & N6229;
  assign N6311 = 1'b0 & N6228;
  assign N6312 = 1'b0 & N6227;
  assign N6313 = 1'b0 & N6226;
  assign N6314 = 1'b0 & N6225;
  assign N6315 = 1'b0 & N6224;
  assign N6316 = 1'b0 & N6223;
  assign N6317 = 1'b0 & N6222;
  assign N6318 = 1'b0 & N6221;
  assign N6319 = 1'b0 & N6220;
  assign N6320 = 1'b0 & N6219;
  assign N6321 = 1'b0 & N6218;
  assign N6322 = 1'b0 & N6217;
  assign N6323 = 1'b0 & N6216;
  assign N6324 = 1'b0 & N6215;
  assign N6325 = 1'b0 & N6214;
  assign N6326 = 1'b0 & N6213;
  assign N6327 = 1'b0 & N6212;
  assign N6328 = 1'b0 & N6211;
  assign N6329 = 1'b0 & N6210;
  assign N6330 = 1'b0 & N6209;
  assign N6331 = 1'b0 & N6208;
  assign N6332 = 1'b0 & N6207;
  assign N6333 = 1'b0 & N6206;
  assign N6398 = ~mhpmcounter_we[17];
  assign N6399 = 1'b0 & csr_wdata_int[31];
  assign N6400 = 1'b0 & csr_wdata_int[30];
  assign N6401 = 1'b0 & csr_wdata_int[29];
  assign N6402 = 1'b0 & csr_wdata_int[28];
  assign N6403 = 1'b0 & csr_wdata_int[27];
  assign N6404 = 1'b0 & csr_wdata_int[26];
  assign N6405 = 1'b0 & csr_wdata_int[25];
  assign N6406 = 1'b0 & csr_wdata_int[24];
  assign N6407 = 1'b0 & csr_wdata_int[23];
  assign N6408 = 1'b0 & csr_wdata_int[22];
  assign N6409 = 1'b0 & csr_wdata_int[21];
  assign N6410 = 1'b0 & csr_wdata_int[20];
  assign N6411 = 1'b0 & csr_wdata_int[19];
  assign N6412 = 1'b0 & csr_wdata_int[18];
  assign N6413 = 1'b0 & csr_wdata_int[17];
  assign N6414 = 1'b0 & csr_wdata_int[16];
  assign N6415 = 1'b0 & csr_wdata_int[15];
  assign N6416 = 1'b0 & csr_wdata_int[14];
  assign N6417 = 1'b0 & csr_wdata_int[13];
  assign N6418 = 1'b0 & csr_wdata_int[12];
  assign N6419 = 1'b0 & csr_wdata_int[11];
  assign N6420 = 1'b0 & csr_wdata_int[10];
  assign N6421 = 1'b0 & csr_wdata_int[9];
  assign N6422 = 1'b0 & csr_wdata_int[8];
  assign N6423 = 1'b0 & csr_wdata_int[7];
  assign N6424 = 1'b0 & csr_wdata_int[6];
  assign N6425 = 1'b0 & csr_wdata_int[5];
  assign N6426 = 1'b0 & csr_wdata_int[4];
  assign N6427 = 1'b0 & csr_wdata_int[3];
  assign N6428 = 1'b0 & csr_wdata_int[2];
  assign N6429 = 1'b0 & csr_wdata_int[1];
  assign N6430 = 1'b0 & csr_wdata_int[0];
  assign N6431 = ~mhpmcounterh_we[17];
  assign N6432 = 1'b0 & csr_wdata_int[31];
  assign N6433 = 1'b0 & csr_wdata_int[30];
  assign N6434 = 1'b0 & csr_wdata_int[29];
  assign N6435 = 1'b0 & csr_wdata_int[28];
  assign N6436 = 1'b0 & csr_wdata_int[27];
  assign N6437 = 1'b0 & csr_wdata_int[26];
  assign N6438 = 1'b0 & csr_wdata_int[25];
  assign N6439 = 1'b0 & csr_wdata_int[24];
  assign N6440 = 1'b0 & csr_wdata_int[23];
  assign N6441 = 1'b0 & csr_wdata_int[22];
  assign N6442 = 1'b0 & csr_wdata_int[21];
  assign N6443 = 1'b0 & csr_wdata_int[20];
  assign N6444 = 1'b0 & csr_wdata_int[19];
  assign N6445 = 1'b0 & csr_wdata_int[18];
  assign N6446 = 1'b0 & csr_wdata_int[17];
  assign N6447 = 1'b0 & csr_wdata_int[16];
  assign N6448 = 1'b0 & csr_wdata_int[15];
  assign N6449 = 1'b0 & csr_wdata_int[14];
  assign N6450 = 1'b0 & csr_wdata_int[13];
  assign N6451 = 1'b0 & csr_wdata_int[12];
  assign N6452 = 1'b0 & csr_wdata_int[11];
  assign N6453 = 1'b0 & csr_wdata_int[10];
  assign N6454 = 1'b0 & csr_wdata_int[9];
  assign N6455 = 1'b0 & csr_wdata_int[8];
  assign N6456 = 1'b0 & csr_wdata_int[7];
  assign N6457 = 1'b0 & csr_wdata_int[6];
  assign N6458 = 1'b0 & csr_wdata_int[5];
  assign N6459 = 1'b0 & csr_wdata_int[4];
  assign N6460 = 1'b0 & csr_wdata_int[3];
  assign N6461 = 1'b0 & csr_wdata_int[2];
  assign N6462 = 1'b0 & csr_wdata_int[1];
  assign N6463 = 1'b0 & csr_wdata_int[0];
  assign N6496 = 1'b0 & N10723;
  assign N10723 = ~mcountinhibit[18];
  assign N6497 = ~N6496;
  assign N6562 = 1'b0 & N6561;
  assign N6563 = 1'b0 & N6560;
  assign N6564 = 1'b0 & N6559;
  assign N6565 = 1'b0 & N6558;
  assign N6566 = 1'b0 & N6557;
  assign N6567 = 1'b0 & N6556;
  assign N6568 = 1'b0 & N6555;
  assign N6569 = 1'b0 & N6554;
  assign N6570 = 1'b0 & N6553;
  assign N6571 = 1'b0 & N6552;
  assign N6572 = 1'b0 & N6551;
  assign N6573 = 1'b0 & N6550;
  assign N6574 = 1'b0 & N6549;
  assign N6575 = 1'b0 & N6548;
  assign N6576 = 1'b0 & N6547;
  assign N6577 = 1'b0 & N6546;
  assign N6578 = 1'b0 & N6545;
  assign N6579 = 1'b0 & N6544;
  assign N6580 = 1'b0 & N6543;
  assign N6581 = 1'b0 & N6542;
  assign N6582 = 1'b0 & N6541;
  assign N6583 = 1'b0 & N6540;
  assign N6584 = 1'b0 & N6539;
  assign N6585 = 1'b0 & N6538;
  assign N6586 = 1'b0 & N6537;
  assign N6587 = 1'b0 & N6536;
  assign N6588 = 1'b0 & N6535;
  assign N6589 = 1'b0 & N6534;
  assign N6590 = 1'b0 & N6533;
  assign N6591 = 1'b0 & N6532;
  assign N6592 = 1'b0 & N6531;
  assign N6593 = 1'b0 & N6530;
  assign N6594 = 1'b0 & N6529;
  assign N6595 = 1'b0 & N6528;
  assign N6596 = 1'b0 & N6527;
  assign N6597 = 1'b0 & N6526;
  assign N6598 = 1'b0 & N6525;
  assign N6599 = 1'b0 & N6524;
  assign N6600 = 1'b0 & N6523;
  assign N6601 = 1'b0 & N6522;
  assign N6602 = 1'b0 & N6521;
  assign N6603 = 1'b0 & N6520;
  assign N6604 = 1'b0 & N6519;
  assign N6605 = 1'b0 & N6518;
  assign N6606 = 1'b0 & N6517;
  assign N6607 = 1'b0 & N6516;
  assign N6608 = 1'b0 & N6515;
  assign N6609 = 1'b0 & N6514;
  assign N6610 = 1'b0 & N6513;
  assign N6611 = 1'b0 & N6512;
  assign N6612 = 1'b0 & N6511;
  assign N6613 = 1'b0 & N6510;
  assign N6614 = 1'b0 & N6509;
  assign N6615 = 1'b0 & N6508;
  assign N6616 = 1'b0 & N6507;
  assign N6617 = 1'b0 & N6506;
  assign N6618 = 1'b0 & N6505;
  assign N6619 = 1'b0 & N6504;
  assign N6620 = 1'b0 & N6503;
  assign N6621 = 1'b0 & N6502;
  assign N6622 = 1'b0 & N6501;
  assign N6623 = 1'b0 & N6500;
  assign N6624 = 1'b0 & N6499;
  assign N6625 = 1'b0 & N6498;
  assign N6690 = ~mhpmcounter_we[18];
  assign N6691 = 1'b0 & csr_wdata_int[31];
  assign N6692 = 1'b0 & csr_wdata_int[30];
  assign N6693 = 1'b0 & csr_wdata_int[29];
  assign N6694 = 1'b0 & csr_wdata_int[28];
  assign N6695 = 1'b0 & csr_wdata_int[27];
  assign N6696 = 1'b0 & csr_wdata_int[26];
  assign N6697 = 1'b0 & csr_wdata_int[25];
  assign N6698 = 1'b0 & csr_wdata_int[24];
  assign N6699 = 1'b0 & csr_wdata_int[23];
  assign N6700 = 1'b0 & csr_wdata_int[22];
  assign N6701 = 1'b0 & csr_wdata_int[21];
  assign N6702 = 1'b0 & csr_wdata_int[20];
  assign N6703 = 1'b0 & csr_wdata_int[19];
  assign N6704 = 1'b0 & csr_wdata_int[18];
  assign N6705 = 1'b0 & csr_wdata_int[17];
  assign N6706 = 1'b0 & csr_wdata_int[16];
  assign N6707 = 1'b0 & csr_wdata_int[15];
  assign N6708 = 1'b0 & csr_wdata_int[14];
  assign N6709 = 1'b0 & csr_wdata_int[13];
  assign N6710 = 1'b0 & csr_wdata_int[12];
  assign N6711 = 1'b0 & csr_wdata_int[11];
  assign N6712 = 1'b0 & csr_wdata_int[10];
  assign N6713 = 1'b0 & csr_wdata_int[9];
  assign N6714 = 1'b0 & csr_wdata_int[8];
  assign N6715 = 1'b0 & csr_wdata_int[7];
  assign N6716 = 1'b0 & csr_wdata_int[6];
  assign N6717 = 1'b0 & csr_wdata_int[5];
  assign N6718 = 1'b0 & csr_wdata_int[4];
  assign N6719 = 1'b0 & csr_wdata_int[3];
  assign N6720 = 1'b0 & csr_wdata_int[2];
  assign N6721 = 1'b0 & csr_wdata_int[1];
  assign N6722 = 1'b0 & csr_wdata_int[0];
  assign N6723 = ~mhpmcounterh_we[18];
  assign N6724 = 1'b0 & csr_wdata_int[31];
  assign N6725 = 1'b0 & csr_wdata_int[30];
  assign N6726 = 1'b0 & csr_wdata_int[29];
  assign N6727 = 1'b0 & csr_wdata_int[28];
  assign N6728 = 1'b0 & csr_wdata_int[27];
  assign N6729 = 1'b0 & csr_wdata_int[26];
  assign N6730 = 1'b0 & csr_wdata_int[25];
  assign N6731 = 1'b0 & csr_wdata_int[24];
  assign N6732 = 1'b0 & csr_wdata_int[23];
  assign N6733 = 1'b0 & csr_wdata_int[22];
  assign N6734 = 1'b0 & csr_wdata_int[21];
  assign N6735 = 1'b0 & csr_wdata_int[20];
  assign N6736 = 1'b0 & csr_wdata_int[19];
  assign N6737 = 1'b0 & csr_wdata_int[18];
  assign N6738 = 1'b0 & csr_wdata_int[17];
  assign N6739 = 1'b0 & csr_wdata_int[16];
  assign N6740 = 1'b0 & csr_wdata_int[15];
  assign N6741 = 1'b0 & csr_wdata_int[14];
  assign N6742 = 1'b0 & csr_wdata_int[13];
  assign N6743 = 1'b0 & csr_wdata_int[12];
  assign N6744 = 1'b0 & csr_wdata_int[11];
  assign N6745 = 1'b0 & csr_wdata_int[10];
  assign N6746 = 1'b0 & csr_wdata_int[9];
  assign N6747 = 1'b0 & csr_wdata_int[8];
  assign N6748 = 1'b0 & csr_wdata_int[7];
  assign N6749 = 1'b0 & csr_wdata_int[6];
  assign N6750 = 1'b0 & csr_wdata_int[5];
  assign N6751 = 1'b0 & csr_wdata_int[4];
  assign N6752 = 1'b0 & csr_wdata_int[3];
  assign N6753 = 1'b0 & csr_wdata_int[2];
  assign N6754 = 1'b0 & csr_wdata_int[1];
  assign N6755 = 1'b0 & csr_wdata_int[0];
  assign N6788 = 1'b0 & N10724;
  assign N10724 = ~mcountinhibit[19];
  assign N6789 = ~N6788;
  assign N6854 = 1'b0 & N6853;
  assign N6855 = 1'b0 & N6852;
  assign N6856 = 1'b0 & N6851;
  assign N6857 = 1'b0 & N6850;
  assign N6858 = 1'b0 & N6849;
  assign N6859 = 1'b0 & N6848;
  assign N6860 = 1'b0 & N6847;
  assign N6861 = 1'b0 & N6846;
  assign N6862 = 1'b0 & N6845;
  assign N6863 = 1'b0 & N6844;
  assign N6864 = 1'b0 & N6843;
  assign N6865 = 1'b0 & N6842;
  assign N6866 = 1'b0 & N6841;
  assign N6867 = 1'b0 & N6840;
  assign N6868 = 1'b0 & N6839;
  assign N6869 = 1'b0 & N6838;
  assign N6870 = 1'b0 & N6837;
  assign N6871 = 1'b0 & N6836;
  assign N6872 = 1'b0 & N6835;
  assign N6873 = 1'b0 & N6834;
  assign N6874 = 1'b0 & N6833;
  assign N6875 = 1'b0 & N6832;
  assign N6876 = 1'b0 & N6831;
  assign N6877 = 1'b0 & N6830;
  assign N6878 = 1'b0 & N6829;
  assign N6879 = 1'b0 & N6828;
  assign N6880 = 1'b0 & N6827;
  assign N6881 = 1'b0 & N6826;
  assign N6882 = 1'b0 & N6825;
  assign N6883 = 1'b0 & N6824;
  assign N6884 = 1'b0 & N6823;
  assign N6885 = 1'b0 & N6822;
  assign N6886 = 1'b0 & N6821;
  assign N6887 = 1'b0 & N6820;
  assign N6888 = 1'b0 & N6819;
  assign N6889 = 1'b0 & N6818;
  assign N6890 = 1'b0 & N6817;
  assign N6891 = 1'b0 & N6816;
  assign N6892 = 1'b0 & N6815;
  assign N6893 = 1'b0 & N6814;
  assign N6894 = 1'b0 & N6813;
  assign N6895 = 1'b0 & N6812;
  assign N6896 = 1'b0 & N6811;
  assign N6897 = 1'b0 & N6810;
  assign N6898 = 1'b0 & N6809;
  assign N6899 = 1'b0 & N6808;
  assign N6900 = 1'b0 & N6807;
  assign N6901 = 1'b0 & N6806;
  assign N6902 = 1'b0 & N6805;
  assign N6903 = 1'b0 & N6804;
  assign N6904 = 1'b0 & N6803;
  assign N6905 = 1'b0 & N6802;
  assign N6906 = 1'b0 & N6801;
  assign N6907 = 1'b0 & N6800;
  assign N6908 = 1'b0 & N6799;
  assign N6909 = 1'b0 & N6798;
  assign N6910 = 1'b0 & N6797;
  assign N6911 = 1'b0 & N6796;
  assign N6912 = 1'b0 & N6795;
  assign N6913 = 1'b0 & N6794;
  assign N6914 = 1'b0 & N6793;
  assign N6915 = 1'b0 & N6792;
  assign N6916 = 1'b0 & N6791;
  assign N6917 = 1'b0 & N6790;
  assign N6982 = ~mhpmcounter_we[19];
  assign N6983 = 1'b0 & csr_wdata_int[31];
  assign N6984 = 1'b0 & csr_wdata_int[30];
  assign N6985 = 1'b0 & csr_wdata_int[29];
  assign N6986 = 1'b0 & csr_wdata_int[28];
  assign N6987 = 1'b0 & csr_wdata_int[27];
  assign N6988 = 1'b0 & csr_wdata_int[26];
  assign N6989 = 1'b0 & csr_wdata_int[25];
  assign N6990 = 1'b0 & csr_wdata_int[24];
  assign N6991 = 1'b0 & csr_wdata_int[23];
  assign N6992 = 1'b0 & csr_wdata_int[22];
  assign N6993 = 1'b0 & csr_wdata_int[21];
  assign N6994 = 1'b0 & csr_wdata_int[20];
  assign N6995 = 1'b0 & csr_wdata_int[19];
  assign N6996 = 1'b0 & csr_wdata_int[18];
  assign N6997 = 1'b0 & csr_wdata_int[17];
  assign N6998 = 1'b0 & csr_wdata_int[16];
  assign N6999 = 1'b0 & csr_wdata_int[15];
  assign N7000 = 1'b0 & csr_wdata_int[14];
  assign N7001 = 1'b0 & csr_wdata_int[13];
  assign N7002 = 1'b0 & csr_wdata_int[12];
  assign N7003 = 1'b0 & csr_wdata_int[11];
  assign N7004 = 1'b0 & csr_wdata_int[10];
  assign N7005 = 1'b0 & csr_wdata_int[9];
  assign N7006 = 1'b0 & csr_wdata_int[8];
  assign N7007 = 1'b0 & csr_wdata_int[7];
  assign N7008 = 1'b0 & csr_wdata_int[6];
  assign N7009 = 1'b0 & csr_wdata_int[5];
  assign N7010 = 1'b0 & csr_wdata_int[4];
  assign N7011 = 1'b0 & csr_wdata_int[3];
  assign N7012 = 1'b0 & csr_wdata_int[2];
  assign N7013 = 1'b0 & csr_wdata_int[1];
  assign N7014 = 1'b0 & csr_wdata_int[0];
  assign N7015 = ~mhpmcounterh_we[19];
  assign N7016 = 1'b0 & csr_wdata_int[31];
  assign N7017 = 1'b0 & csr_wdata_int[30];
  assign N7018 = 1'b0 & csr_wdata_int[29];
  assign N7019 = 1'b0 & csr_wdata_int[28];
  assign N7020 = 1'b0 & csr_wdata_int[27];
  assign N7021 = 1'b0 & csr_wdata_int[26];
  assign N7022 = 1'b0 & csr_wdata_int[25];
  assign N7023 = 1'b0 & csr_wdata_int[24];
  assign N7024 = 1'b0 & csr_wdata_int[23];
  assign N7025 = 1'b0 & csr_wdata_int[22];
  assign N7026 = 1'b0 & csr_wdata_int[21];
  assign N7027 = 1'b0 & csr_wdata_int[20];
  assign N7028 = 1'b0 & csr_wdata_int[19];
  assign N7029 = 1'b0 & csr_wdata_int[18];
  assign N7030 = 1'b0 & csr_wdata_int[17];
  assign N7031 = 1'b0 & csr_wdata_int[16];
  assign N7032 = 1'b0 & csr_wdata_int[15];
  assign N7033 = 1'b0 & csr_wdata_int[14];
  assign N7034 = 1'b0 & csr_wdata_int[13];
  assign N7035 = 1'b0 & csr_wdata_int[12];
  assign N7036 = 1'b0 & csr_wdata_int[11];
  assign N7037 = 1'b0 & csr_wdata_int[10];
  assign N7038 = 1'b0 & csr_wdata_int[9];
  assign N7039 = 1'b0 & csr_wdata_int[8];
  assign N7040 = 1'b0 & csr_wdata_int[7];
  assign N7041 = 1'b0 & csr_wdata_int[6];
  assign N7042 = 1'b0 & csr_wdata_int[5];
  assign N7043 = 1'b0 & csr_wdata_int[4];
  assign N7044 = 1'b0 & csr_wdata_int[3];
  assign N7045 = 1'b0 & csr_wdata_int[2];
  assign N7046 = 1'b0 & csr_wdata_int[1];
  assign N7047 = 1'b0 & csr_wdata_int[0];
  assign N7080 = 1'b0 & N10725;
  assign N10725 = ~mcountinhibit[20];
  assign N7081 = ~N7080;
  assign N7146 = 1'b0 & N7145;
  assign N7147 = 1'b0 & N7144;
  assign N7148 = 1'b0 & N7143;
  assign N7149 = 1'b0 & N7142;
  assign N7150 = 1'b0 & N7141;
  assign N7151 = 1'b0 & N7140;
  assign N7152 = 1'b0 & N7139;
  assign N7153 = 1'b0 & N7138;
  assign N7154 = 1'b0 & N7137;
  assign N7155 = 1'b0 & N7136;
  assign N7156 = 1'b0 & N7135;
  assign N7157 = 1'b0 & N7134;
  assign N7158 = 1'b0 & N7133;
  assign N7159 = 1'b0 & N7132;
  assign N7160 = 1'b0 & N7131;
  assign N7161 = 1'b0 & N7130;
  assign N7162 = 1'b0 & N7129;
  assign N7163 = 1'b0 & N7128;
  assign N7164 = 1'b0 & N7127;
  assign N7165 = 1'b0 & N7126;
  assign N7166 = 1'b0 & N7125;
  assign N7167 = 1'b0 & N7124;
  assign N7168 = 1'b0 & N7123;
  assign N7169 = 1'b0 & N7122;
  assign N7170 = 1'b0 & N7121;
  assign N7171 = 1'b0 & N7120;
  assign N7172 = 1'b0 & N7119;
  assign N7173 = 1'b0 & N7118;
  assign N7174 = 1'b0 & N7117;
  assign N7175 = 1'b0 & N7116;
  assign N7176 = 1'b0 & N7115;
  assign N7177 = 1'b0 & N7114;
  assign N7178 = 1'b0 & N7113;
  assign N7179 = 1'b0 & N7112;
  assign N7180 = 1'b0 & N7111;
  assign N7181 = 1'b0 & N7110;
  assign N7182 = 1'b0 & N7109;
  assign N7183 = 1'b0 & N7108;
  assign N7184 = 1'b0 & N7107;
  assign N7185 = 1'b0 & N7106;
  assign N7186 = 1'b0 & N7105;
  assign N7187 = 1'b0 & N7104;
  assign N7188 = 1'b0 & N7103;
  assign N7189 = 1'b0 & N7102;
  assign N7190 = 1'b0 & N7101;
  assign N7191 = 1'b0 & N7100;
  assign N7192 = 1'b0 & N7099;
  assign N7193 = 1'b0 & N7098;
  assign N7194 = 1'b0 & N7097;
  assign N7195 = 1'b0 & N7096;
  assign N7196 = 1'b0 & N7095;
  assign N7197 = 1'b0 & N7094;
  assign N7198 = 1'b0 & N7093;
  assign N7199 = 1'b0 & N7092;
  assign N7200 = 1'b0 & N7091;
  assign N7201 = 1'b0 & N7090;
  assign N7202 = 1'b0 & N7089;
  assign N7203 = 1'b0 & N7088;
  assign N7204 = 1'b0 & N7087;
  assign N7205 = 1'b0 & N7086;
  assign N7206 = 1'b0 & N7085;
  assign N7207 = 1'b0 & N7084;
  assign N7208 = 1'b0 & N7083;
  assign N7209 = 1'b0 & N7082;
  assign N7274 = ~mhpmcounter_we[20];
  assign N7275 = 1'b0 & csr_wdata_int[31];
  assign N7276 = 1'b0 & csr_wdata_int[30];
  assign N7277 = 1'b0 & csr_wdata_int[29];
  assign N7278 = 1'b0 & csr_wdata_int[28];
  assign N7279 = 1'b0 & csr_wdata_int[27];
  assign N7280 = 1'b0 & csr_wdata_int[26];
  assign N7281 = 1'b0 & csr_wdata_int[25];
  assign N7282 = 1'b0 & csr_wdata_int[24];
  assign N7283 = 1'b0 & csr_wdata_int[23];
  assign N7284 = 1'b0 & csr_wdata_int[22];
  assign N7285 = 1'b0 & csr_wdata_int[21];
  assign N7286 = 1'b0 & csr_wdata_int[20];
  assign N7287 = 1'b0 & csr_wdata_int[19];
  assign N7288 = 1'b0 & csr_wdata_int[18];
  assign N7289 = 1'b0 & csr_wdata_int[17];
  assign N7290 = 1'b0 & csr_wdata_int[16];
  assign N7291 = 1'b0 & csr_wdata_int[15];
  assign N7292 = 1'b0 & csr_wdata_int[14];
  assign N7293 = 1'b0 & csr_wdata_int[13];
  assign N7294 = 1'b0 & csr_wdata_int[12];
  assign N7295 = 1'b0 & csr_wdata_int[11];
  assign N7296 = 1'b0 & csr_wdata_int[10];
  assign N7297 = 1'b0 & csr_wdata_int[9];
  assign N7298 = 1'b0 & csr_wdata_int[8];
  assign N7299 = 1'b0 & csr_wdata_int[7];
  assign N7300 = 1'b0 & csr_wdata_int[6];
  assign N7301 = 1'b0 & csr_wdata_int[5];
  assign N7302 = 1'b0 & csr_wdata_int[4];
  assign N7303 = 1'b0 & csr_wdata_int[3];
  assign N7304 = 1'b0 & csr_wdata_int[2];
  assign N7305 = 1'b0 & csr_wdata_int[1];
  assign N7306 = 1'b0 & csr_wdata_int[0];
  assign N7307 = ~mhpmcounterh_we[20];
  assign N7308 = 1'b0 & csr_wdata_int[31];
  assign N7309 = 1'b0 & csr_wdata_int[30];
  assign N7310 = 1'b0 & csr_wdata_int[29];
  assign N7311 = 1'b0 & csr_wdata_int[28];
  assign N7312 = 1'b0 & csr_wdata_int[27];
  assign N7313 = 1'b0 & csr_wdata_int[26];
  assign N7314 = 1'b0 & csr_wdata_int[25];
  assign N7315 = 1'b0 & csr_wdata_int[24];
  assign N7316 = 1'b0 & csr_wdata_int[23];
  assign N7317 = 1'b0 & csr_wdata_int[22];
  assign N7318 = 1'b0 & csr_wdata_int[21];
  assign N7319 = 1'b0 & csr_wdata_int[20];
  assign N7320 = 1'b0 & csr_wdata_int[19];
  assign N7321 = 1'b0 & csr_wdata_int[18];
  assign N7322 = 1'b0 & csr_wdata_int[17];
  assign N7323 = 1'b0 & csr_wdata_int[16];
  assign N7324 = 1'b0 & csr_wdata_int[15];
  assign N7325 = 1'b0 & csr_wdata_int[14];
  assign N7326 = 1'b0 & csr_wdata_int[13];
  assign N7327 = 1'b0 & csr_wdata_int[12];
  assign N7328 = 1'b0 & csr_wdata_int[11];
  assign N7329 = 1'b0 & csr_wdata_int[10];
  assign N7330 = 1'b0 & csr_wdata_int[9];
  assign N7331 = 1'b0 & csr_wdata_int[8];
  assign N7332 = 1'b0 & csr_wdata_int[7];
  assign N7333 = 1'b0 & csr_wdata_int[6];
  assign N7334 = 1'b0 & csr_wdata_int[5];
  assign N7335 = 1'b0 & csr_wdata_int[4];
  assign N7336 = 1'b0 & csr_wdata_int[3];
  assign N7337 = 1'b0 & csr_wdata_int[2];
  assign N7338 = 1'b0 & csr_wdata_int[1];
  assign N7339 = 1'b0 & csr_wdata_int[0];
  assign N7372 = 1'b0 & N10726;
  assign N10726 = ~mcountinhibit[21];
  assign N7373 = ~N7372;
  assign N7438 = 1'b0 & N7437;
  assign N7439 = 1'b0 & N7436;
  assign N7440 = 1'b0 & N7435;
  assign N7441 = 1'b0 & N7434;
  assign N7442 = 1'b0 & N7433;
  assign N7443 = 1'b0 & N7432;
  assign N7444 = 1'b0 & N7431;
  assign N7445 = 1'b0 & N7430;
  assign N7446 = 1'b0 & N7429;
  assign N7447 = 1'b0 & N7428;
  assign N7448 = 1'b0 & N7427;
  assign N7449 = 1'b0 & N7426;
  assign N7450 = 1'b0 & N7425;
  assign N7451 = 1'b0 & N7424;
  assign N7452 = 1'b0 & N7423;
  assign N7453 = 1'b0 & N7422;
  assign N7454 = 1'b0 & N7421;
  assign N7455 = 1'b0 & N7420;
  assign N7456 = 1'b0 & N7419;
  assign N7457 = 1'b0 & N7418;
  assign N7458 = 1'b0 & N7417;
  assign N7459 = 1'b0 & N7416;
  assign N7460 = 1'b0 & N7415;
  assign N7461 = 1'b0 & N7414;
  assign N7462 = 1'b0 & N7413;
  assign N7463 = 1'b0 & N7412;
  assign N7464 = 1'b0 & N7411;
  assign N7465 = 1'b0 & N7410;
  assign N7466 = 1'b0 & N7409;
  assign N7467 = 1'b0 & N7408;
  assign N7468 = 1'b0 & N7407;
  assign N7469 = 1'b0 & N7406;
  assign N7470 = 1'b0 & N7405;
  assign N7471 = 1'b0 & N7404;
  assign N7472 = 1'b0 & N7403;
  assign N7473 = 1'b0 & N7402;
  assign N7474 = 1'b0 & N7401;
  assign N7475 = 1'b0 & N7400;
  assign N7476 = 1'b0 & N7399;
  assign N7477 = 1'b0 & N7398;
  assign N7478 = 1'b0 & N7397;
  assign N7479 = 1'b0 & N7396;
  assign N7480 = 1'b0 & N7395;
  assign N7481 = 1'b0 & N7394;
  assign N7482 = 1'b0 & N7393;
  assign N7483 = 1'b0 & N7392;
  assign N7484 = 1'b0 & N7391;
  assign N7485 = 1'b0 & N7390;
  assign N7486 = 1'b0 & N7389;
  assign N7487 = 1'b0 & N7388;
  assign N7488 = 1'b0 & N7387;
  assign N7489 = 1'b0 & N7386;
  assign N7490 = 1'b0 & N7385;
  assign N7491 = 1'b0 & N7384;
  assign N7492 = 1'b0 & N7383;
  assign N7493 = 1'b0 & N7382;
  assign N7494 = 1'b0 & N7381;
  assign N7495 = 1'b0 & N7380;
  assign N7496 = 1'b0 & N7379;
  assign N7497 = 1'b0 & N7378;
  assign N7498 = 1'b0 & N7377;
  assign N7499 = 1'b0 & N7376;
  assign N7500 = 1'b0 & N7375;
  assign N7501 = 1'b0 & N7374;
  assign N7566 = ~mhpmcounter_we[21];
  assign N7567 = 1'b0 & csr_wdata_int[31];
  assign N7568 = 1'b0 & csr_wdata_int[30];
  assign N7569 = 1'b0 & csr_wdata_int[29];
  assign N7570 = 1'b0 & csr_wdata_int[28];
  assign N7571 = 1'b0 & csr_wdata_int[27];
  assign N7572 = 1'b0 & csr_wdata_int[26];
  assign N7573 = 1'b0 & csr_wdata_int[25];
  assign N7574 = 1'b0 & csr_wdata_int[24];
  assign N7575 = 1'b0 & csr_wdata_int[23];
  assign N7576 = 1'b0 & csr_wdata_int[22];
  assign N7577 = 1'b0 & csr_wdata_int[21];
  assign N7578 = 1'b0 & csr_wdata_int[20];
  assign N7579 = 1'b0 & csr_wdata_int[19];
  assign N7580 = 1'b0 & csr_wdata_int[18];
  assign N7581 = 1'b0 & csr_wdata_int[17];
  assign N7582 = 1'b0 & csr_wdata_int[16];
  assign N7583 = 1'b0 & csr_wdata_int[15];
  assign N7584 = 1'b0 & csr_wdata_int[14];
  assign N7585 = 1'b0 & csr_wdata_int[13];
  assign N7586 = 1'b0 & csr_wdata_int[12];
  assign N7587 = 1'b0 & csr_wdata_int[11];
  assign N7588 = 1'b0 & csr_wdata_int[10];
  assign N7589 = 1'b0 & csr_wdata_int[9];
  assign N7590 = 1'b0 & csr_wdata_int[8];
  assign N7591 = 1'b0 & csr_wdata_int[7];
  assign N7592 = 1'b0 & csr_wdata_int[6];
  assign N7593 = 1'b0 & csr_wdata_int[5];
  assign N7594 = 1'b0 & csr_wdata_int[4];
  assign N7595 = 1'b0 & csr_wdata_int[3];
  assign N7596 = 1'b0 & csr_wdata_int[2];
  assign N7597 = 1'b0 & csr_wdata_int[1];
  assign N7598 = 1'b0 & csr_wdata_int[0];
  assign N7599 = ~mhpmcounterh_we[21];
  assign N7600 = 1'b0 & csr_wdata_int[31];
  assign N7601 = 1'b0 & csr_wdata_int[30];
  assign N7602 = 1'b0 & csr_wdata_int[29];
  assign N7603 = 1'b0 & csr_wdata_int[28];
  assign N7604 = 1'b0 & csr_wdata_int[27];
  assign N7605 = 1'b0 & csr_wdata_int[26];
  assign N7606 = 1'b0 & csr_wdata_int[25];
  assign N7607 = 1'b0 & csr_wdata_int[24];
  assign N7608 = 1'b0 & csr_wdata_int[23];
  assign N7609 = 1'b0 & csr_wdata_int[22];
  assign N7610 = 1'b0 & csr_wdata_int[21];
  assign N7611 = 1'b0 & csr_wdata_int[20];
  assign N7612 = 1'b0 & csr_wdata_int[19];
  assign N7613 = 1'b0 & csr_wdata_int[18];
  assign N7614 = 1'b0 & csr_wdata_int[17];
  assign N7615 = 1'b0 & csr_wdata_int[16];
  assign N7616 = 1'b0 & csr_wdata_int[15];
  assign N7617 = 1'b0 & csr_wdata_int[14];
  assign N7618 = 1'b0 & csr_wdata_int[13];
  assign N7619 = 1'b0 & csr_wdata_int[12];
  assign N7620 = 1'b0 & csr_wdata_int[11];
  assign N7621 = 1'b0 & csr_wdata_int[10];
  assign N7622 = 1'b0 & csr_wdata_int[9];
  assign N7623 = 1'b0 & csr_wdata_int[8];
  assign N7624 = 1'b0 & csr_wdata_int[7];
  assign N7625 = 1'b0 & csr_wdata_int[6];
  assign N7626 = 1'b0 & csr_wdata_int[5];
  assign N7627 = 1'b0 & csr_wdata_int[4];
  assign N7628 = 1'b0 & csr_wdata_int[3];
  assign N7629 = 1'b0 & csr_wdata_int[2];
  assign N7630 = 1'b0 & csr_wdata_int[1];
  assign N7631 = 1'b0 & csr_wdata_int[0];
  assign N7664 = 1'b0 & N10727;
  assign N10727 = ~mcountinhibit[22];
  assign N7665 = ~N7664;
  assign N7730 = 1'b0 & N7729;
  assign N7731 = 1'b0 & N7728;
  assign N7732 = 1'b0 & N7727;
  assign N7733 = 1'b0 & N7726;
  assign N7734 = 1'b0 & N7725;
  assign N7735 = 1'b0 & N7724;
  assign N7736 = 1'b0 & N7723;
  assign N7737 = 1'b0 & N7722;
  assign N7738 = 1'b0 & N7721;
  assign N7739 = 1'b0 & N7720;
  assign N7740 = 1'b0 & N7719;
  assign N7741 = 1'b0 & N7718;
  assign N7742 = 1'b0 & N7717;
  assign N7743 = 1'b0 & N7716;
  assign N7744 = 1'b0 & N7715;
  assign N7745 = 1'b0 & N7714;
  assign N7746 = 1'b0 & N7713;
  assign N7747 = 1'b0 & N7712;
  assign N7748 = 1'b0 & N7711;
  assign N7749 = 1'b0 & N7710;
  assign N7750 = 1'b0 & N7709;
  assign N7751 = 1'b0 & N7708;
  assign N7752 = 1'b0 & N7707;
  assign N7753 = 1'b0 & N7706;
  assign N7754 = 1'b0 & N7705;
  assign N7755 = 1'b0 & N7704;
  assign N7756 = 1'b0 & N7703;
  assign N7757 = 1'b0 & N7702;
  assign N7758 = 1'b0 & N7701;
  assign N7759 = 1'b0 & N7700;
  assign N7760 = 1'b0 & N7699;
  assign N7761 = 1'b0 & N7698;
  assign N7762 = 1'b0 & N7697;
  assign N7763 = 1'b0 & N7696;
  assign N7764 = 1'b0 & N7695;
  assign N7765 = 1'b0 & N7694;
  assign N7766 = 1'b0 & N7693;
  assign N7767 = 1'b0 & N7692;
  assign N7768 = 1'b0 & N7691;
  assign N7769 = 1'b0 & N7690;
  assign N7770 = 1'b0 & N7689;
  assign N7771 = 1'b0 & N7688;
  assign N7772 = 1'b0 & N7687;
  assign N7773 = 1'b0 & N7686;
  assign N7774 = 1'b0 & N7685;
  assign N7775 = 1'b0 & N7684;
  assign N7776 = 1'b0 & N7683;
  assign N7777 = 1'b0 & N7682;
  assign N7778 = 1'b0 & N7681;
  assign N7779 = 1'b0 & N7680;
  assign N7780 = 1'b0 & N7679;
  assign N7781 = 1'b0 & N7678;
  assign N7782 = 1'b0 & N7677;
  assign N7783 = 1'b0 & N7676;
  assign N7784 = 1'b0 & N7675;
  assign N7785 = 1'b0 & N7674;
  assign N7786 = 1'b0 & N7673;
  assign N7787 = 1'b0 & N7672;
  assign N7788 = 1'b0 & N7671;
  assign N7789 = 1'b0 & N7670;
  assign N7790 = 1'b0 & N7669;
  assign N7791 = 1'b0 & N7668;
  assign N7792 = 1'b0 & N7667;
  assign N7793 = 1'b0 & N7666;
  assign N7858 = ~mhpmcounter_we[22];
  assign N7859 = 1'b0 & csr_wdata_int[31];
  assign N7860 = 1'b0 & csr_wdata_int[30];
  assign N7861 = 1'b0 & csr_wdata_int[29];
  assign N7862 = 1'b0 & csr_wdata_int[28];
  assign N7863 = 1'b0 & csr_wdata_int[27];
  assign N7864 = 1'b0 & csr_wdata_int[26];
  assign N7865 = 1'b0 & csr_wdata_int[25];
  assign N7866 = 1'b0 & csr_wdata_int[24];
  assign N7867 = 1'b0 & csr_wdata_int[23];
  assign N7868 = 1'b0 & csr_wdata_int[22];
  assign N7869 = 1'b0 & csr_wdata_int[21];
  assign N7870 = 1'b0 & csr_wdata_int[20];
  assign N7871 = 1'b0 & csr_wdata_int[19];
  assign N7872 = 1'b0 & csr_wdata_int[18];
  assign N7873 = 1'b0 & csr_wdata_int[17];
  assign N7874 = 1'b0 & csr_wdata_int[16];
  assign N7875 = 1'b0 & csr_wdata_int[15];
  assign N7876 = 1'b0 & csr_wdata_int[14];
  assign N7877 = 1'b0 & csr_wdata_int[13];
  assign N7878 = 1'b0 & csr_wdata_int[12];
  assign N7879 = 1'b0 & csr_wdata_int[11];
  assign N7880 = 1'b0 & csr_wdata_int[10];
  assign N7881 = 1'b0 & csr_wdata_int[9];
  assign N7882 = 1'b0 & csr_wdata_int[8];
  assign N7883 = 1'b0 & csr_wdata_int[7];
  assign N7884 = 1'b0 & csr_wdata_int[6];
  assign N7885 = 1'b0 & csr_wdata_int[5];
  assign N7886 = 1'b0 & csr_wdata_int[4];
  assign N7887 = 1'b0 & csr_wdata_int[3];
  assign N7888 = 1'b0 & csr_wdata_int[2];
  assign N7889 = 1'b0 & csr_wdata_int[1];
  assign N7890 = 1'b0 & csr_wdata_int[0];
  assign N7891 = ~mhpmcounterh_we[22];
  assign N7892 = 1'b0 & csr_wdata_int[31];
  assign N7893 = 1'b0 & csr_wdata_int[30];
  assign N7894 = 1'b0 & csr_wdata_int[29];
  assign N7895 = 1'b0 & csr_wdata_int[28];
  assign N7896 = 1'b0 & csr_wdata_int[27];
  assign N7897 = 1'b0 & csr_wdata_int[26];
  assign N7898 = 1'b0 & csr_wdata_int[25];
  assign N7899 = 1'b0 & csr_wdata_int[24];
  assign N7900 = 1'b0 & csr_wdata_int[23];
  assign N7901 = 1'b0 & csr_wdata_int[22];
  assign N7902 = 1'b0 & csr_wdata_int[21];
  assign N7903 = 1'b0 & csr_wdata_int[20];
  assign N7904 = 1'b0 & csr_wdata_int[19];
  assign N7905 = 1'b0 & csr_wdata_int[18];
  assign N7906 = 1'b0 & csr_wdata_int[17];
  assign N7907 = 1'b0 & csr_wdata_int[16];
  assign N7908 = 1'b0 & csr_wdata_int[15];
  assign N7909 = 1'b0 & csr_wdata_int[14];
  assign N7910 = 1'b0 & csr_wdata_int[13];
  assign N7911 = 1'b0 & csr_wdata_int[12];
  assign N7912 = 1'b0 & csr_wdata_int[11];
  assign N7913 = 1'b0 & csr_wdata_int[10];
  assign N7914 = 1'b0 & csr_wdata_int[9];
  assign N7915 = 1'b0 & csr_wdata_int[8];
  assign N7916 = 1'b0 & csr_wdata_int[7];
  assign N7917 = 1'b0 & csr_wdata_int[6];
  assign N7918 = 1'b0 & csr_wdata_int[5];
  assign N7919 = 1'b0 & csr_wdata_int[4];
  assign N7920 = 1'b0 & csr_wdata_int[3];
  assign N7921 = 1'b0 & csr_wdata_int[2];
  assign N7922 = 1'b0 & csr_wdata_int[1];
  assign N7923 = 1'b0 & csr_wdata_int[0];
  assign N7956 = 1'b0 & N10728;
  assign N10728 = ~mcountinhibit[23];
  assign N7957 = ~N7956;
  assign N8022 = 1'b0 & N8021;
  assign N8023 = 1'b0 & N8020;
  assign N8024 = 1'b0 & N8019;
  assign N8025 = 1'b0 & N8018;
  assign N8026 = 1'b0 & N8017;
  assign N8027 = 1'b0 & N8016;
  assign N8028 = 1'b0 & N8015;
  assign N8029 = 1'b0 & N8014;
  assign N8030 = 1'b0 & N8013;
  assign N8031 = 1'b0 & N8012;
  assign N8032 = 1'b0 & N8011;
  assign N8033 = 1'b0 & N8010;
  assign N8034 = 1'b0 & N8009;
  assign N8035 = 1'b0 & N8008;
  assign N8036 = 1'b0 & N8007;
  assign N8037 = 1'b0 & N8006;
  assign N8038 = 1'b0 & N8005;
  assign N8039 = 1'b0 & N8004;
  assign N8040 = 1'b0 & N8003;
  assign N8041 = 1'b0 & N8002;
  assign N8042 = 1'b0 & N8001;
  assign N8043 = 1'b0 & N8000;
  assign N8044 = 1'b0 & N7999;
  assign N8045 = 1'b0 & N7998;
  assign N8046 = 1'b0 & N7997;
  assign N8047 = 1'b0 & N7996;
  assign N8048 = 1'b0 & N7995;
  assign N8049 = 1'b0 & N7994;
  assign N8050 = 1'b0 & N7993;
  assign N8051 = 1'b0 & N7992;
  assign N8052 = 1'b0 & N7991;
  assign N8053 = 1'b0 & N7990;
  assign N8054 = 1'b0 & N7989;
  assign N8055 = 1'b0 & N7988;
  assign N8056 = 1'b0 & N7987;
  assign N8057 = 1'b0 & N7986;
  assign N8058 = 1'b0 & N7985;
  assign N8059 = 1'b0 & N7984;
  assign N8060 = 1'b0 & N7983;
  assign N8061 = 1'b0 & N7982;
  assign N8062 = 1'b0 & N7981;
  assign N8063 = 1'b0 & N7980;
  assign N8064 = 1'b0 & N7979;
  assign N8065 = 1'b0 & N7978;
  assign N8066 = 1'b0 & N7977;
  assign N8067 = 1'b0 & N7976;
  assign N8068 = 1'b0 & N7975;
  assign N8069 = 1'b0 & N7974;
  assign N8070 = 1'b0 & N7973;
  assign N8071 = 1'b0 & N7972;
  assign N8072 = 1'b0 & N7971;
  assign N8073 = 1'b0 & N7970;
  assign N8074 = 1'b0 & N7969;
  assign N8075 = 1'b0 & N7968;
  assign N8076 = 1'b0 & N7967;
  assign N8077 = 1'b0 & N7966;
  assign N8078 = 1'b0 & N7965;
  assign N8079 = 1'b0 & N7964;
  assign N8080 = 1'b0 & N7963;
  assign N8081 = 1'b0 & N7962;
  assign N8082 = 1'b0 & N7961;
  assign N8083 = 1'b0 & N7960;
  assign N8084 = 1'b0 & N7959;
  assign N8085 = 1'b0 & N7958;
  assign N8150 = ~mhpmcounter_we[23];
  assign N8151 = 1'b0 & csr_wdata_int[31];
  assign N8152 = 1'b0 & csr_wdata_int[30];
  assign N8153 = 1'b0 & csr_wdata_int[29];
  assign N8154 = 1'b0 & csr_wdata_int[28];
  assign N8155 = 1'b0 & csr_wdata_int[27];
  assign N8156 = 1'b0 & csr_wdata_int[26];
  assign N8157 = 1'b0 & csr_wdata_int[25];
  assign N8158 = 1'b0 & csr_wdata_int[24];
  assign N8159 = 1'b0 & csr_wdata_int[23];
  assign N8160 = 1'b0 & csr_wdata_int[22];
  assign N8161 = 1'b0 & csr_wdata_int[21];
  assign N8162 = 1'b0 & csr_wdata_int[20];
  assign N8163 = 1'b0 & csr_wdata_int[19];
  assign N8164 = 1'b0 & csr_wdata_int[18];
  assign N8165 = 1'b0 & csr_wdata_int[17];
  assign N8166 = 1'b0 & csr_wdata_int[16];
  assign N8167 = 1'b0 & csr_wdata_int[15];
  assign N8168 = 1'b0 & csr_wdata_int[14];
  assign N8169 = 1'b0 & csr_wdata_int[13];
  assign N8170 = 1'b0 & csr_wdata_int[12];
  assign N8171 = 1'b0 & csr_wdata_int[11];
  assign N8172 = 1'b0 & csr_wdata_int[10];
  assign N8173 = 1'b0 & csr_wdata_int[9];
  assign N8174 = 1'b0 & csr_wdata_int[8];
  assign N8175 = 1'b0 & csr_wdata_int[7];
  assign N8176 = 1'b0 & csr_wdata_int[6];
  assign N8177 = 1'b0 & csr_wdata_int[5];
  assign N8178 = 1'b0 & csr_wdata_int[4];
  assign N8179 = 1'b0 & csr_wdata_int[3];
  assign N8180 = 1'b0 & csr_wdata_int[2];
  assign N8181 = 1'b0 & csr_wdata_int[1];
  assign N8182 = 1'b0 & csr_wdata_int[0];
  assign N8183 = ~mhpmcounterh_we[23];
  assign N8184 = 1'b0 & csr_wdata_int[31];
  assign N8185 = 1'b0 & csr_wdata_int[30];
  assign N8186 = 1'b0 & csr_wdata_int[29];
  assign N8187 = 1'b0 & csr_wdata_int[28];
  assign N8188 = 1'b0 & csr_wdata_int[27];
  assign N8189 = 1'b0 & csr_wdata_int[26];
  assign N8190 = 1'b0 & csr_wdata_int[25];
  assign N8191 = 1'b0 & csr_wdata_int[24];
  assign N8192 = 1'b0 & csr_wdata_int[23];
  assign N8193 = 1'b0 & csr_wdata_int[22];
  assign N8194 = 1'b0 & csr_wdata_int[21];
  assign N8195 = 1'b0 & csr_wdata_int[20];
  assign N8196 = 1'b0 & csr_wdata_int[19];
  assign N8197 = 1'b0 & csr_wdata_int[18];
  assign N8198 = 1'b0 & csr_wdata_int[17];
  assign N8199 = 1'b0 & csr_wdata_int[16];
  assign N8200 = 1'b0 & csr_wdata_int[15];
  assign N8201 = 1'b0 & csr_wdata_int[14];
  assign N8202 = 1'b0 & csr_wdata_int[13];
  assign N8203 = 1'b0 & csr_wdata_int[12];
  assign N8204 = 1'b0 & csr_wdata_int[11];
  assign N8205 = 1'b0 & csr_wdata_int[10];
  assign N8206 = 1'b0 & csr_wdata_int[9];
  assign N8207 = 1'b0 & csr_wdata_int[8];
  assign N8208 = 1'b0 & csr_wdata_int[7];
  assign N8209 = 1'b0 & csr_wdata_int[6];
  assign N8210 = 1'b0 & csr_wdata_int[5];
  assign N8211 = 1'b0 & csr_wdata_int[4];
  assign N8212 = 1'b0 & csr_wdata_int[3];
  assign N8213 = 1'b0 & csr_wdata_int[2];
  assign N8214 = 1'b0 & csr_wdata_int[1];
  assign N8215 = 1'b0 & csr_wdata_int[0];
  assign N8248 = 1'b0 & N10729;
  assign N10729 = ~mcountinhibit[24];
  assign N8249 = ~N8248;
  assign N8314 = 1'b0 & N8313;
  assign N8315 = 1'b0 & N8312;
  assign N8316 = 1'b0 & N8311;
  assign N8317 = 1'b0 & N8310;
  assign N8318 = 1'b0 & N8309;
  assign N8319 = 1'b0 & N8308;
  assign N8320 = 1'b0 & N8307;
  assign N8321 = 1'b0 & N8306;
  assign N8322 = 1'b0 & N8305;
  assign N8323 = 1'b0 & N8304;
  assign N8324 = 1'b0 & N8303;
  assign N8325 = 1'b0 & N8302;
  assign N8326 = 1'b0 & N8301;
  assign N8327 = 1'b0 & N8300;
  assign N8328 = 1'b0 & N8299;
  assign N8329 = 1'b0 & N8298;
  assign N8330 = 1'b0 & N8297;
  assign N8331 = 1'b0 & N8296;
  assign N8332 = 1'b0 & N8295;
  assign N8333 = 1'b0 & N8294;
  assign N8334 = 1'b0 & N8293;
  assign N8335 = 1'b0 & N8292;
  assign N8336 = 1'b0 & N8291;
  assign N8337 = 1'b0 & N8290;
  assign N8338 = 1'b0 & N8289;
  assign N8339 = 1'b0 & N8288;
  assign N8340 = 1'b0 & N8287;
  assign N8341 = 1'b0 & N8286;
  assign N8342 = 1'b0 & N8285;
  assign N8343 = 1'b0 & N8284;
  assign N8344 = 1'b0 & N8283;
  assign N8345 = 1'b0 & N8282;
  assign N8346 = 1'b0 & N8281;
  assign N8347 = 1'b0 & N8280;
  assign N8348 = 1'b0 & N8279;
  assign N8349 = 1'b0 & N8278;
  assign N8350 = 1'b0 & N8277;
  assign N8351 = 1'b0 & N8276;
  assign N8352 = 1'b0 & N8275;
  assign N8353 = 1'b0 & N8274;
  assign N8354 = 1'b0 & N8273;
  assign N8355 = 1'b0 & N8272;
  assign N8356 = 1'b0 & N8271;
  assign N8357 = 1'b0 & N8270;
  assign N8358 = 1'b0 & N8269;
  assign N8359 = 1'b0 & N8268;
  assign N8360 = 1'b0 & N8267;
  assign N8361 = 1'b0 & N8266;
  assign N8362 = 1'b0 & N8265;
  assign N8363 = 1'b0 & N8264;
  assign N8364 = 1'b0 & N8263;
  assign N8365 = 1'b0 & N8262;
  assign N8366 = 1'b0 & N8261;
  assign N8367 = 1'b0 & N8260;
  assign N8368 = 1'b0 & N8259;
  assign N8369 = 1'b0 & N8258;
  assign N8370 = 1'b0 & N8257;
  assign N8371 = 1'b0 & N8256;
  assign N8372 = 1'b0 & N8255;
  assign N8373 = 1'b0 & N8254;
  assign N8374 = 1'b0 & N8253;
  assign N8375 = 1'b0 & N8252;
  assign N8376 = 1'b0 & N8251;
  assign N8377 = 1'b0 & N8250;
  assign N8442 = ~mhpmcounter_we[24];
  assign N8443 = 1'b0 & csr_wdata_int[31];
  assign N8444 = 1'b0 & csr_wdata_int[30];
  assign N8445 = 1'b0 & csr_wdata_int[29];
  assign N8446 = 1'b0 & csr_wdata_int[28];
  assign N8447 = 1'b0 & csr_wdata_int[27];
  assign N8448 = 1'b0 & csr_wdata_int[26];
  assign N8449 = 1'b0 & csr_wdata_int[25];
  assign N8450 = 1'b0 & csr_wdata_int[24];
  assign N8451 = 1'b0 & csr_wdata_int[23];
  assign N8452 = 1'b0 & csr_wdata_int[22];
  assign N8453 = 1'b0 & csr_wdata_int[21];
  assign N8454 = 1'b0 & csr_wdata_int[20];
  assign N8455 = 1'b0 & csr_wdata_int[19];
  assign N8456 = 1'b0 & csr_wdata_int[18];
  assign N8457 = 1'b0 & csr_wdata_int[17];
  assign N8458 = 1'b0 & csr_wdata_int[16];
  assign N8459 = 1'b0 & csr_wdata_int[15];
  assign N8460 = 1'b0 & csr_wdata_int[14];
  assign N8461 = 1'b0 & csr_wdata_int[13];
  assign N8462 = 1'b0 & csr_wdata_int[12];
  assign N8463 = 1'b0 & csr_wdata_int[11];
  assign N8464 = 1'b0 & csr_wdata_int[10];
  assign N8465 = 1'b0 & csr_wdata_int[9];
  assign N8466 = 1'b0 & csr_wdata_int[8];
  assign N8467 = 1'b0 & csr_wdata_int[7];
  assign N8468 = 1'b0 & csr_wdata_int[6];
  assign N8469 = 1'b0 & csr_wdata_int[5];
  assign N8470 = 1'b0 & csr_wdata_int[4];
  assign N8471 = 1'b0 & csr_wdata_int[3];
  assign N8472 = 1'b0 & csr_wdata_int[2];
  assign N8473 = 1'b0 & csr_wdata_int[1];
  assign N8474 = 1'b0 & csr_wdata_int[0];
  assign N8475 = ~mhpmcounterh_we[24];
  assign N8476 = 1'b0 & csr_wdata_int[31];
  assign N8477 = 1'b0 & csr_wdata_int[30];
  assign N8478 = 1'b0 & csr_wdata_int[29];
  assign N8479 = 1'b0 & csr_wdata_int[28];
  assign N8480 = 1'b0 & csr_wdata_int[27];
  assign N8481 = 1'b0 & csr_wdata_int[26];
  assign N8482 = 1'b0 & csr_wdata_int[25];
  assign N8483 = 1'b0 & csr_wdata_int[24];
  assign N8484 = 1'b0 & csr_wdata_int[23];
  assign N8485 = 1'b0 & csr_wdata_int[22];
  assign N8486 = 1'b0 & csr_wdata_int[21];
  assign N8487 = 1'b0 & csr_wdata_int[20];
  assign N8488 = 1'b0 & csr_wdata_int[19];
  assign N8489 = 1'b0 & csr_wdata_int[18];
  assign N8490 = 1'b0 & csr_wdata_int[17];
  assign N8491 = 1'b0 & csr_wdata_int[16];
  assign N8492 = 1'b0 & csr_wdata_int[15];
  assign N8493 = 1'b0 & csr_wdata_int[14];
  assign N8494 = 1'b0 & csr_wdata_int[13];
  assign N8495 = 1'b0 & csr_wdata_int[12];
  assign N8496 = 1'b0 & csr_wdata_int[11];
  assign N8497 = 1'b0 & csr_wdata_int[10];
  assign N8498 = 1'b0 & csr_wdata_int[9];
  assign N8499 = 1'b0 & csr_wdata_int[8];
  assign N8500 = 1'b0 & csr_wdata_int[7];
  assign N8501 = 1'b0 & csr_wdata_int[6];
  assign N8502 = 1'b0 & csr_wdata_int[5];
  assign N8503 = 1'b0 & csr_wdata_int[4];
  assign N8504 = 1'b0 & csr_wdata_int[3];
  assign N8505 = 1'b0 & csr_wdata_int[2];
  assign N8506 = 1'b0 & csr_wdata_int[1];
  assign N8507 = 1'b0 & csr_wdata_int[0];
  assign N8540 = 1'b0 & N10730;
  assign N10730 = ~mcountinhibit[25];
  assign N8541 = ~N8540;
  assign N8606 = 1'b0 & N8605;
  assign N8607 = 1'b0 & N8604;
  assign N8608 = 1'b0 & N8603;
  assign N8609 = 1'b0 & N8602;
  assign N8610 = 1'b0 & N8601;
  assign N8611 = 1'b0 & N8600;
  assign N8612 = 1'b0 & N8599;
  assign N8613 = 1'b0 & N8598;
  assign N8614 = 1'b0 & N8597;
  assign N8615 = 1'b0 & N8596;
  assign N8616 = 1'b0 & N8595;
  assign N8617 = 1'b0 & N8594;
  assign N8618 = 1'b0 & N8593;
  assign N8619 = 1'b0 & N8592;
  assign N8620 = 1'b0 & N8591;
  assign N8621 = 1'b0 & N8590;
  assign N8622 = 1'b0 & N8589;
  assign N8623 = 1'b0 & N8588;
  assign N8624 = 1'b0 & N8587;
  assign N8625 = 1'b0 & N8586;
  assign N8626 = 1'b0 & N8585;
  assign N8627 = 1'b0 & N8584;
  assign N8628 = 1'b0 & N8583;
  assign N8629 = 1'b0 & N8582;
  assign N8630 = 1'b0 & N8581;
  assign N8631 = 1'b0 & N8580;
  assign N8632 = 1'b0 & N8579;
  assign N8633 = 1'b0 & N8578;
  assign N8634 = 1'b0 & N8577;
  assign N8635 = 1'b0 & N8576;
  assign N8636 = 1'b0 & N8575;
  assign N8637 = 1'b0 & N8574;
  assign N8638 = 1'b0 & N8573;
  assign N8639 = 1'b0 & N8572;
  assign N8640 = 1'b0 & N8571;
  assign N8641 = 1'b0 & N8570;
  assign N8642 = 1'b0 & N8569;
  assign N8643 = 1'b0 & N8568;
  assign N8644 = 1'b0 & N8567;
  assign N8645 = 1'b0 & N8566;
  assign N8646 = 1'b0 & N8565;
  assign N8647 = 1'b0 & N8564;
  assign N8648 = 1'b0 & N8563;
  assign N8649 = 1'b0 & N8562;
  assign N8650 = 1'b0 & N8561;
  assign N8651 = 1'b0 & N8560;
  assign N8652 = 1'b0 & N8559;
  assign N8653 = 1'b0 & N8558;
  assign N8654 = 1'b0 & N8557;
  assign N8655 = 1'b0 & N8556;
  assign N8656 = 1'b0 & N8555;
  assign N8657 = 1'b0 & N8554;
  assign N8658 = 1'b0 & N8553;
  assign N8659 = 1'b0 & N8552;
  assign N8660 = 1'b0 & N8551;
  assign N8661 = 1'b0 & N8550;
  assign N8662 = 1'b0 & N8549;
  assign N8663 = 1'b0 & N8548;
  assign N8664 = 1'b0 & N8547;
  assign N8665 = 1'b0 & N8546;
  assign N8666 = 1'b0 & N8545;
  assign N8667 = 1'b0 & N8544;
  assign N8668 = 1'b0 & N8543;
  assign N8669 = 1'b0 & N8542;
  assign N8734 = ~mhpmcounter_we[25];
  assign N8735 = 1'b0 & csr_wdata_int[31];
  assign N8736 = 1'b0 & csr_wdata_int[30];
  assign N8737 = 1'b0 & csr_wdata_int[29];
  assign N8738 = 1'b0 & csr_wdata_int[28];
  assign N8739 = 1'b0 & csr_wdata_int[27];
  assign N8740 = 1'b0 & csr_wdata_int[26];
  assign N8741 = 1'b0 & csr_wdata_int[25];
  assign N8742 = 1'b0 & csr_wdata_int[24];
  assign N8743 = 1'b0 & csr_wdata_int[23];
  assign N8744 = 1'b0 & csr_wdata_int[22];
  assign N8745 = 1'b0 & csr_wdata_int[21];
  assign N8746 = 1'b0 & csr_wdata_int[20];
  assign N8747 = 1'b0 & csr_wdata_int[19];
  assign N8748 = 1'b0 & csr_wdata_int[18];
  assign N8749 = 1'b0 & csr_wdata_int[17];
  assign N8750 = 1'b0 & csr_wdata_int[16];
  assign N8751 = 1'b0 & csr_wdata_int[15];
  assign N8752 = 1'b0 & csr_wdata_int[14];
  assign N8753 = 1'b0 & csr_wdata_int[13];
  assign N8754 = 1'b0 & csr_wdata_int[12];
  assign N8755 = 1'b0 & csr_wdata_int[11];
  assign N8756 = 1'b0 & csr_wdata_int[10];
  assign N8757 = 1'b0 & csr_wdata_int[9];
  assign N8758 = 1'b0 & csr_wdata_int[8];
  assign N8759 = 1'b0 & csr_wdata_int[7];
  assign N8760 = 1'b0 & csr_wdata_int[6];
  assign N8761 = 1'b0 & csr_wdata_int[5];
  assign N8762 = 1'b0 & csr_wdata_int[4];
  assign N8763 = 1'b0 & csr_wdata_int[3];
  assign N8764 = 1'b0 & csr_wdata_int[2];
  assign N8765 = 1'b0 & csr_wdata_int[1];
  assign N8766 = 1'b0 & csr_wdata_int[0];
  assign N8767 = ~mhpmcounterh_we[25];
  assign N8768 = 1'b0 & csr_wdata_int[31];
  assign N8769 = 1'b0 & csr_wdata_int[30];
  assign N8770 = 1'b0 & csr_wdata_int[29];
  assign N8771 = 1'b0 & csr_wdata_int[28];
  assign N8772 = 1'b0 & csr_wdata_int[27];
  assign N8773 = 1'b0 & csr_wdata_int[26];
  assign N8774 = 1'b0 & csr_wdata_int[25];
  assign N8775 = 1'b0 & csr_wdata_int[24];
  assign N8776 = 1'b0 & csr_wdata_int[23];
  assign N8777 = 1'b0 & csr_wdata_int[22];
  assign N8778 = 1'b0 & csr_wdata_int[21];
  assign N8779 = 1'b0 & csr_wdata_int[20];
  assign N8780 = 1'b0 & csr_wdata_int[19];
  assign N8781 = 1'b0 & csr_wdata_int[18];
  assign N8782 = 1'b0 & csr_wdata_int[17];
  assign N8783 = 1'b0 & csr_wdata_int[16];
  assign N8784 = 1'b0 & csr_wdata_int[15];
  assign N8785 = 1'b0 & csr_wdata_int[14];
  assign N8786 = 1'b0 & csr_wdata_int[13];
  assign N8787 = 1'b0 & csr_wdata_int[12];
  assign N8788 = 1'b0 & csr_wdata_int[11];
  assign N8789 = 1'b0 & csr_wdata_int[10];
  assign N8790 = 1'b0 & csr_wdata_int[9];
  assign N8791 = 1'b0 & csr_wdata_int[8];
  assign N8792 = 1'b0 & csr_wdata_int[7];
  assign N8793 = 1'b0 & csr_wdata_int[6];
  assign N8794 = 1'b0 & csr_wdata_int[5];
  assign N8795 = 1'b0 & csr_wdata_int[4];
  assign N8796 = 1'b0 & csr_wdata_int[3];
  assign N8797 = 1'b0 & csr_wdata_int[2];
  assign N8798 = 1'b0 & csr_wdata_int[1];
  assign N8799 = 1'b0 & csr_wdata_int[0];
  assign N8832 = 1'b0 & N10731;
  assign N10731 = ~mcountinhibit[26];
  assign N8833 = ~N8832;
  assign N8898 = 1'b0 & N8897;
  assign N8899 = 1'b0 & N8896;
  assign N8900 = 1'b0 & N8895;
  assign N8901 = 1'b0 & N8894;
  assign N8902 = 1'b0 & N8893;
  assign N8903 = 1'b0 & N8892;
  assign N8904 = 1'b0 & N8891;
  assign N8905 = 1'b0 & N8890;
  assign N8906 = 1'b0 & N8889;
  assign N8907 = 1'b0 & N8888;
  assign N8908 = 1'b0 & N8887;
  assign N8909 = 1'b0 & N8886;
  assign N8910 = 1'b0 & N8885;
  assign N8911 = 1'b0 & N8884;
  assign N8912 = 1'b0 & N8883;
  assign N8913 = 1'b0 & N8882;
  assign N8914 = 1'b0 & N8881;
  assign N8915 = 1'b0 & N8880;
  assign N8916 = 1'b0 & N8879;
  assign N8917 = 1'b0 & N8878;
  assign N8918 = 1'b0 & N8877;
  assign N8919 = 1'b0 & N8876;
  assign N8920 = 1'b0 & N8875;
  assign N8921 = 1'b0 & N8874;
  assign N8922 = 1'b0 & N8873;
  assign N8923 = 1'b0 & N8872;
  assign N8924 = 1'b0 & N8871;
  assign N8925 = 1'b0 & N8870;
  assign N8926 = 1'b0 & N8869;
  assign N8927 = 1'b0 & N8868;
  assign N8928 = 1'b0 & N8867;
  assign N8929 = 1'b0 & N8866;
  assign N8930 = 1'b0 & N8865;
  assign N8931 = 1'b0 & N8864;
  assign N8932 = 1'b0 & N8863;
  assign N8933 = 1'b0 & N8862;
  assign N8934 = 1'b0 & N8861;
  assign N8935 = 1'b0 & N8860;
  assign N8936 = 1'b0 & N8859;
  assign N8937 = 1'b0 & N8858;
  assign N8938 = 1'b0 & N8857;
  assign N8939 = 1'b0 & N8856;
  assign N8940 = 1'b0 & N8855;
  assign N8941 = 1'b0 & N8854;
  assign N8942 = 1'b0 & N8853;
  assign N8943 = 1'b0 & N8852;
  assign N8944 = 1'b0 & N8851;
  assign N8945 = 1'b0 & N8850;
  assign N8946 = 1'b0 & N8849;
  assign N8947 = 1'b0 & N8848;
  assign N8948 = 1'b0 & N8847;
  assign N8949 = 1'b0 & N8846;
  assign N8950 = 1'b0 & N8845;
  assign N8951 = 1'b0 & N8844;
  assign N8952 = 1'b0 & N8843;
  assign N8953 = 1'b0 & N8842;
  assign N8954 = 1'b0 & N8841;
  assign N8955 = 1'b0 & N8840;
  assign N8956 = 1'b0 & N8839;
  assign N8957 = 1'b0 & N8838;
  assign N8958 = 1'b0 & N8837;
  assign N8959 = 1'b0 & N8836;
  assign N8960 = 1'b0 & N8835;
  assign N8961 = 1'b0 & N8834;
  assign N9026 = ~mhpmcounter_we[26];
  assign N9027 = 1'b0 & csr_wdata_int[31];
  assign N9028 = 1'b0 & csr_wdata_int[30];
  assign N9029 = 1'b0 & csr_wdata_int[29];
  assign N9030 = 1'b0 & csr_wdata_int[28];
  assign N9031 = 1'b0 & csr_wdata_int[27];
  assign N9032 = 1'b0 & csr_wdata_int[26];
  assign N9033 = 1'b0 & csr_wdata_int[25];
  assign N9034 = 1'b0 & csr_wdata_int[24];
  assign N9035 = 1'b0 & csr_wdata_int[23];
  assign N9036 = 1'b0 & csr_wdata_int[22];
  assign N9037 = 1'b0 & csr_wdata_int[21];
  assign N9038 = 1'b0 & csr_wdata_int[20];
  assign N9039 = 1'b0 & csr_wdata_int[19];
  assign N9040 = 1'b0 & csr_wdata_int[18];
  assign N9041 = 1'b0 & csr_wdata_int[17];
  assign N9042 = 1'b0 & csr_wdata_int[16];
  assign N9043 = 1'b0 & csr_wdata_int[15];
  assign N9044 = 1'b0 & csr_wdata_int[14];
  assign N9045 = 1'b0 & csr_wdata_int[13];
  assign N9046 = 1'b0 & csr_wdata_int[12];
  assign N9047 = 1'b0 & csr_wdata_int[11];
  assign N9048 = 1'b0 & csr_wdata_int[10];
  assign N9049 = 1'b0 & csr_wdata_int[9];
  assign N9050 = 1'b0 & csr_wdata_int[8];
  assign N9051 = 1'b0 & csr_wdata_int[7];
  assign N9052 = 1'b0 & csr_wdata_int[6];
  assign N9053 = 1'b0 & csr_wdata_int[5];
  assign N9054 = 1'b0 & csr_wdata_int[4];
  assign N9055 = 1'b0 & csr_wdata_int[3];
  assign N9056 = 1'b0 & csr_wdata_int[2];
  assign N9057 = 1'b0 & csr_wdata_int[1];
  assign N9058 = 1'b0 & csr_wdata_int[0];
  assign N9059 = ~mhpmcounterh_we[26];
  assign N9060 = 1'b0 & csr_wdata_int[31];
  assign N9061 = 1'b0 & csr_wdata_int[30];
  assign N9062 = 1'b0 & csr_wdata_int[29];
  assign N9063 = 1'b0 & csr_wdata_int[28];
  assign N9064 = 1'b0 & csr_wdata_int[27];
  assign N9065 = 1'b0 & csr_wdata_int[26];
  assign N9066 = 1'b0 & csr_wdata_int[25];
  assign N9067 = 1'b0 & csr_wdata_int[24];
  assign N9068 = 1'b0 & csr_wdata_int[23];
  assign N9069 = 1'b0 & csr_wdata_int[22];
  assign N9070 = 1'b0 & csr_wdata_int[21];
  assign N9071 = 1'b0 & csr_wdata_int[20];
  assign N9072 = 1'b0 & csr_wdata_int[19];
  assign N9073 = 1'b0 & csr_wdata_int[18];
  assign N9074 = 1'b0 & csr_wdata_int[17];
  assign N9075 = 1'b0 & csr_wdata_int[16];
  assign N9076 = 1'b0 & csr_wdata_int[15];
  assign N9077 = 1'b0 & csr_wdata_int[14];
  assign N9078 = 1'b0 & csr_wdata_int[13];
  assign N9079 = 1'b0 & csr_wdata_int[12];
  assign N9080 = 1'b0 & csr_wdata_int[11];
  assign N9081 = 1'b0 & csr_wdata_int[10];
  assign N9082 = 1'b0 & csr_wdata_int[9];
  assign N9083 = 1'b0 & csr_wdata_int[8];
  assign N9084 = 1'b0 & csr_wdata_int[7];
  assign N9085 = 1'b0 & csr_wdata_int[6];
  assign N9086 = 1'b0 & csr_wdata_int[5];
  assign N9087 = 1'b0 & csr_wdata_int[4];
  assign N9088 = 1'b0 & csr_wdata_int[3];
  assign N9089 = 1'b0 & csr_wdata_int[2];
  assign N9090 = 1'b0 & csr_wdata_int[1];
  assign N9091 = 1'b0 & csr_wdata_int[0];
  assign N9124 = 1'b0 & N10732;
  assign N10732 = ~mcountinhibit[27];
  assign N9125 = ~N9124;
  assign N9190 = 1'b0 & N9189;
  assign N9191 = 1'b0 & N9188;
  assign N9192 = 1'b0 & N9187;
  assign N9193 = 1'b0 & N9186;
  assign N9194 = 1'b0 & N9185;
  assign N9195 = 1'b0 & N9184;
  assign N9196 = 1'b0 & N9183;
  assign N9197 = 1'b0 & N9182;
  assign N9198 = 1'b0 & N9181;
  assign N9199 = 1'b0 & N9180;
  assign N9200 = 1'b0 & N9179;
  assign N9201 = 1'b0 & N9178;
  assign N9202 = 1'b0 & N9177;
  assign N9203 = 1'b0 & N9176;
  assign N9204 = 1'b0 & N9175;
  assign N9205 = 1'b0 & N9174;
  assign N9206 = 1'b0 & N9173;
  assign N9207 = 1'b0 & N9172;
  assign N9208 = 1'b0 & N9171;
  assign N9209 = 1'b0 & N9170;
  assign N9210 = 1'b0 & N9169;
  assign N9211 = 1'b0 & N9168;
  assign N9212 = 1'b0 & N9167;
  assign N9213 = 1'b0 & N9166;
  assign N9214 = 1'b0 & N9165;
  assign N9215 = 1'b0 & N9164;
  assign N9216 = 1'b0 & N9163;
  assign N9217 = 1'b0 & N9162;
  assign N9218 = 1'b0 & N9161;
  assign N9219 = 1'b0 & N9160;
  assign N9220 = 1'b0 & N9159;
  assign N9221 = 1'b0 & N9158;
  assign N9222 = 1'b0 & N9157;
  assign N9223 = 1'b0 & N9156;
  assign N9224 = 1'b0 & N9155;
  assign N9225 = 1'b0 & N9154;
  assign N9226 = 1'b0 & N9153;
  assign N9227 = 1'b0 & N9152;
  assign N9228 = 1'b0 & N9151;
  assign N9229 = 1'b0 & N9150;
  assign N9230 = 1'b0 & N9149;
  assign N9231 = 1'b0 & N9148;
  assign N9232 = 1'b0 & N9147;
  assign N9233 = 1'b0 & N9146;
  assign N9234 = 1'b0 & N9145;
  assign N9235 = 1'b0 & N9144;
  assign N9236 = 1'b0 & N9143;
  assign N9237 = 1'b0 & N9142;
  assign N9238 = 1'b0 & N9141;
  assign N9239 = 1'b0 & N9140;
  assign N9240 = 1'b0 & N9139;
  assign N9241 = 1'b0 & N9138;
  assign N9242 = 1'b0 & N9137;
  assign N9243 = 1'b0 & N9136;
  assign N9244 = 1'b0 & N9135;
  assign N9245 = 1'b0 & N9134;
  assign N9246 = 1'b0 & N9133;
  assign N9247 = 1'b0 & N9132;
  assign N9248 = 1'b0 & N9131;
  assign N9249 = 1'b0 & N9130;
  assign N9250 = 1'b0 & N9129;
  assign N9251 = 1'b0 & N9128;
  assign N9252 = 1'b0 & N9127;
  assign N9253 = 1'b0 & N9126;
  assign N9318 = ~mhpmcounter_we[27];
  assign N9319 = 1'b0 & csr_wdata_int[31];
  assign N9320 = 1'b0 & csr_wdata_int[30];
  assign N9321 = 1'b0 & csr_wdata_int[29];
  assign N9322 = 1'b0 & csr_wdata_int[28];
  assign N9323 = 1'b0 & csr_wdata_int[27];
  assign N9324 = 1'b0 & csr_wdata_int[26];
  assign N9325 = 1'b0 & csr_wdata_int[25];
  assign N9326 = 1'b0 & csr_wdata_int[24];
  assign N9327 = 1'b0 & csr_wdata_int[23];
  assign N9328 = 1'b0 & csr_wdata_int[22];
  assign N9329 = 1'b0 & csr_wdata_int[21];
  assign N9330 = 1'b0 & csr_wdata_int[20];
  assign N9331 = 1'b0 & csr_wdata_int[19];
  assign N9332 = 1'b0 & csr_wdata_int[18];
  assign N9333 = 1'b0 & csr_wdata_int[17];
  assign N9334 = 1'b0 & csr_wdata_int[16];
  assign N9335 = 1'b0 & csr_wdata_int[15];
  assign N9336 = 1'b0 & csr_wdata_int[14];
  assign N9337 = 1'b0 & csr_wdata_int[13];
  assign N9338 = 1'b0 & csr_wdata_int[12];
  assign N9339 = 1'b0 & csr_wdata_int[11];
  assign N9340 = 1'b0 & csr_wdata_int[10];
  assign N9341 = 1'b0 & csr_wdata_int[9];
  assign N9342 = 1'b0 & csr_wdata_int[8];
  assign N9343 = 1'b0 & csr_wdata_int[7];
  assign N9344 = 1'b0 & csr_wdata_int[6];
  assign N9345 = 1'b0 & csr_wdata_int[5];
  assign N9346 = 1'b0 & csr_wdata_int[4];
  assign N9347 = 1'b0 & csr_wdata_int[3];
  assign N9348 = 1'b0 & csr_wdata_int[2];
  assign N9349 = 1'b0 & csr_wdata_int[1];
  assign N9350 = 1'b0 & csr_wdata_int[0];
  assign N9351 = ~mhpmcounterh_we[27];
  assign N9352 = 1'b0 & csr_wdata_int[31];
  assign N9353 = 1'b0 & csr_wdata_int[30];
  assign N9354 = 1'b0 & csr_wdata_int[29];
  assign N9355 = 1'b0 & csr_wdata_int[28];
  assign N9356 = 1'b0 & csr_wdata_int[27];
  assign N9357 = 1'b0 & csr_wdata_int[26];
  assign N9358 = 1'b0 & csr_wdata_int[25];
  assign N9359 = 1'b0 & csr_wdata_int[24];
  assign N9360 = 1'b0 & csr_wdata_int[23];
  assign N9361 = 1'b0 & csr_wdata_int[22];
  assign N9362 = 1'b0 & csr_wdata_int[21];
  assign N9363 = 1'b0 & csr_wdata_int[20];
  assign N9364 = 1'b0 & csr_wdata_int[19];
  assign N9365 = 1'b0 & csr_wdata_int[18];
  assign N9366 = 1'b0 & csr_wdata_int[17];
  assign N9367 = 1'b0 & csr_wdata_int[16];
  assign N9368 = 1'b0 & csr_wdata_int[15];
  assign N9369 = 1'b0 & csr_wdata_int[14];
  assign N9370 = 1'b0 & csr_wdata_int[13];
  assign N9371 = 1'b0 & csr_wdata_int[12];
  assign N9372 = 1'b0 & csr_wdata_int[11];
  assign N9373 = 1'b0 & csr_wdata_int[10];
  assign N9374 = 1'b0 & csr_wdata_int[9];
  assign N9375 = 1'b0 & csr_wdata_int[8];
  assign N9376 = 1'b0 & csr_wdata_int[7];
  assign N9377 = 1'b0 & csr_wdata_int[6];
  assign N9378 = 1'b0 & csr_wdata_int[5];
  assign N9379 = 1'b0 & csr_wdata_int[4];
  assign N9380 = 1'b0 & csr_wdata_int[3];
  assign N9381 = 1'b0 & csr_wdata_int[2];
  assign N9382 = 1'b0 & csr_wdata_int[1];
  assign N9383 = 1'b0 & csr_wdata_int[0];
  assign N9416 = 1'b0 & N10733;
  assign N10733 = ~mcountinhibit[28];
  assign N9417 = ~N9416;
  assign N9482 = 1'b0 & N9481;
  assign N9483 = 1'b0 & N9480;
  assign N9484 = 1'b0 & N9479;
  assign N9485 = 1'b0 & N9478;
  assign N9486 = 1'b0 & N9477;
  assign N9487 = 1'b0 & N9476;
  assign N9488 = 1'b0 & N9475;
  assign N9489 = 1'b0 & N9474;
  assign N9490 = 1'b0 & N9473;
  assign N9491 = 1'b0 & N9472;
  assign N9492 = 1'b0 & N9471;
  assign N9493 = 1'b0 & N9470;
  assign N9494 = 1'b0 & N9469;
  assign N9495 = 1'b0 & N9468;
  assign N9496 = 1'b0 & N9467;
  assign N9497 = 1'b0 & N9466;
  assign N9498 = 1'b0 & N9465;
  assign N9499 = 1'b0 & N9464;
  assign N9500 = 1'b0 & N9463;
  assign N9501 = 1'b0 & N9462;
  assign N9502 = 1'b0 & N9461;
  assign N9503 = 1'b0 & N9460;
  assign N9504 = 1'b0 & N9459;
  assign N9505 = 1'b0 & N9458;
  assign N9506 = 1'b0 & N9457;
  assign N9507 = 1'b0 & N9456;
  assign N9508 = 1'b0 & N9455;
  assign N9509 = 1'b0 & N9454;
  assign N9510 = 1'b0 & N9453;
  assign N9511 = 1'b0 & N9452;
  assign N9512 = 1'b0 & N9451;
  assign N9513 = 1'b0 & N9450;
  assign N9514 = 1'b0 & N9449;
  assign N9515 = 1'b0 & N9448;
  assign N9516 = 1'b0 & N9447;
  assign N9517 = 1'b0 & N9446;
  assign N9518 = 1'b0 & N9445;
  assign N9519 = 1'b0 & N9444;
  assign N9520 = 1'b0 & N9443;
  assign N9521 = 1'b0 & N9442;
  assign N9522 = 1'b0 & N9441;
  assign N9523 = 1'b0 & N9440;
  assign N9524 = 1'b0 & N9439;
  assign N9525 = 1'b0 & N9438;
  assign N9526 = 1'b0 & N9437;
  assign N9527 = 1'b0 & N9436;
  assign N9528 = 1'b0 & N9435;
  assign N9529 = 1'b0 & N9434;
  assign N9530 = 1'b0 & N9433;
  assign N9531 = 1'b0 & N9432;
  assign N9532 = 1'b0 & N9431;
  assign N9533 = 1'b0 & N9430;
  assign N9534 = 1'b0 & N9429;
  assign N9535 = 1'b0 & N9428;
  assign N9536 = 1'b0 & N9427;
  assign N9537 = 1'b0 & N9426;
  assign N9538 = 1'b0 & N9425;
  assign N9539 = 1'b0 & N9424;
  assign N9540 = 1'b0 & N9423;
  assign N9541 = 1'b0 & N9422;
  assign N9542 = 1'b0 & N9421;
  assign N9543 = 1'b0 & N9420;
  assign N9544 = 1'b0 & N9419;
  assign N9545 = 1'b0 & N9418;
  assign N9610 = ~mhpmcounter_we[28];
  assign N9611 = 1'b0 & csr_wdata_int[31];
  assign N9612 = 1'b0 & csr_wdata_int[30];
  assign N9613 = 1'b0 & csr_wdata_int[29];
  assign N9614 = 1'b0 & csr_wdata_int[28];
  assign N9615 = 1'b0 & csr_wdata_int[27];
  assign N9616 = 1'b0 & csr_wdata_int[26];
  assign N9617 = 1'b0 & csr_wdata_int[25];
  assign N9618 = 1'b0 & csr_wdata_int[24];
  assign N9619 = 1'b0 & csr_wdata_int[23];
  assign N9620 = 1'b0 & csr_wdata_int[22];
  assign N9621 = 1'b0 & csr_wdata_int[21];
  assign N9622 = 1'b0 & csr_wdata_int[20];
  assign N9623 = 1'b0 & csr_wdata_int[19];
  assign N9624 = 1'b0 & csr_wdata_int[18];
  assign N9625 = 1'b0 & csr_wdata_int[17];
  assign N9626 = 1'b0 & csr_wdata_int[16];
  assign N9627 = 1'b0 & csr_wdata_int[15];
  assign N9628 = 1'b0 & csr_wdata_int[14];
  assign N9629 = 1'b0 & csr_wdata_int[13];
  assign N9630 = 1'b0 & csr_wdata_int[12];
  assign N9631 = 1'b0 & csr_wdata_int[11];
  assign N9632 = 1'b0 & csr_wdata_int[10];
  assign N9633 = 1'b0 & csr_wdata_int[9];
  assign N9634 = 1'b0 & csr_wdata_int[8];
  assign N9635 = 1'b0 & csr_wdata_int[7];
  assign N9636 = 1'b0 & csr_wdata_int[6];
  assign N9637 = 1'b0 & csr_wdata_int[5];
  assign N9638 = 1'b0 & csr_wdata_int[4];
  assign N9639 = 1'b0 & csr_wdata_int[3];
  assign N9640 = 1'b0 & csr_wdata_int[2];
  assign N9641 = 1'b0 & csr_wdata_int[1];
  assign N9642 = 1'b0 & csr_wdata_int[0];
  assign N9643 = ~mhpmcounterh_we[28];
  assign N9644 = 1'b0 & csr_wdata_int[31];
  assign N9645 = 1'b0 & csr_wdata_int[30];
  assign N9646 = 1'b0 & csr_wdata_int[29];
  assign N9647 = 1'b0 & csr_wdata_int[28];
  assign N9648 = 1'b0 & csr_wdata_int[27];
  assign N9649 = 1'b0 & csr_wdata_int[26];
  assign N9650 = 1'b0 & csr_wdata_int[25];
  assign N9651 = 1'b0 & csr_wdata_int[24];
  assign N9652 = 1'b0 & csr_wdata_int[23];
  assign N9653 = 1'b0 & csr_wdata_int[22];
  assign N9654 = 1'b0 & csr_wdata_int[21];
  assign N9655 = 1'b0 & csr_wdata_int[20];
  assign N9656 = 1'b0 & csr_wdata_int[19];
  assign N9657 = 1'b0 & csr_wdata_int[18];
  assign N9658 = 1'b0 & csr_wdata_int[17];
  assign N9659 = 1'b0 & csr_wdata_int[16];
  assign N9660 = 1'b0 & csr_wdata_int[15];
  assign N9661 = 1'b0 & csr_wdata_int[14];
  assign N9662 = 1'b0 & csr_wdata_int[13];
  assign N9663 = 1'b0 & csr_wdata_int[12];
  assign N9664 = 1'b0 & csr_wdata_int[11];
  assign N9665 = 1'b0 & csr_wdata_int[10];
  assign N9666 = 1'b0 & csr_wdata_int[9];
  assign N9667 = 1'b0 & csr_wdata_int[8];
  assign N9668 = 1'b0 & csr_wdata_int[7];
  assign N9669 = 1'b0 & csr_wdata_int[6];
  assign N9670 = 1'b0 & csr_wdata_int[5];
  assign N9671 = 1'b0 & csr_wdata_int[4];
  assign N9672 = 1'b0 & csr_wdata_int[3];
  assign N9673 = 1'b0 & csr_wdata_int[2];
  assign N9674 = 1'b0 & csr_wdata_int[1];
  assign N9675 = 1'b0 & csr_wdata_int[0];
  assign N9708 = 1'b0 & N10734;
  assign N10734 = ~mcountinhibit[29];
  assign N9709 = ~N9708;
  assign N9774 = 1'b0 & N9773;
  assign N9775 = 1'b0 & N9772;
  assign N9776 = 1'b0 & N9771;
  assign N9777 = 1'b0 & N9770;
  assign N9778 = 1'b0 & N9769;
  assign N9779 = 1'b0 & N9768;
  assign N9780 = 1'b0 & N9767;
  assign N9781 = 1'b0 & N9766;
  assign N9782 = 1'b0 & N9765;
  assign N9783 = 1'b0 & N9764;
  assign N9784 = 1'b0 & N9763;
  assign N9785 = 1'b0 & N9762;
  assign N9786 = 1'b0 & N9761;
  assign N9787 = 1'b0 & N9760;
  assign N9788 = 1'b0 & N9759;
  assign N9789 = 1'b0 & N9758;
  assign N9790 = 1'b0 & N9757;
  assign N9791 = 1'b0 & N9756;
  assign N9792 = 1'b0 & N9755;
  assign N9793 = 1'b0 & N9754;
  assign N9794 = 1'b0 & N9753;
  assign N9795 = 1'b0 & N9752;
  assign N9796 = 1'b0 & N9751;
  assign N9797 = 1'b0 & N9750;
  assign N9798 = 1'b0 & N9749;
  assign N9799 = 1'b0 & N9748;
  assign N9800 = 1'b0 & N9747;
  assign N9801 = 1'b0 & N9746;
  assign N9802 = 1'b0 & N9745;
  assign N9803 = 1'b0 & N9744;
  assign N9804 = 1'b0 & N9743;
  assign N9805 = 1'b0 & N9742;
  assign N9806 = 1'b0 & N9741;
  assign N9807 = 1'b0 & N9740;
  assign N9808 = 1'b0 & N9739;
  assign N9809 = 1'b0 & N9738;
  assign N9810 = 1'b0 & N9737;
  assign N9811 = 1'b0 & N9736;
  assign N9812 = 1'b0 & N9735;
  assign N9813 = 1'b0 & N9734;
  assign N9814 = 1'b0 & N9733;
  assign N9815 = 1'b0 & N9732;
  assign N9816 = 1'b0 & N9731;
  assign N9817 = 1'b0 & N9730;
  assign N9818 = 1'b0 & N9729;
  assign N9819 = 1'b0 & N9728;
  assign N9820 = 1'b0 & N9727;
  assign N9821 = 1'b0 & N9726;
  assign N9822 = 1'b0 & N9725;
  assign N9823 = 1'b0 & N9724;
  assign N9824 = 1'b0 & N9723;
  assign N9825 = 1'b0 & N9722;
  assign N9826 = 1'b0 & N9721;
  assign N9827 = 1'b0 & N9720;
  assign N9828 = 1'b0 & N9719;
  assign N9829 = 1'b0 & N9718;
  assign N9830 = 1'b0 & N9717;
  assign N9831 = 1'b0 & N9716;
  assign N9832 = 1'b0 & N9715;
  assign N9833 = 1'b0 & N9714;
  assign N9834 = 1'b0 & N9713;
  assign N9835 = 1'b0 & N9712;
  assign N9836 = 1'b0 & N9711;
  assign N9837 = 1'b0 & N9710;
  assign N9902 = ~mhpmcounter_we[29];
  assign N9903 = 1'b0 & csr_wdata_int[31];
  assign N9904 = 1'b0 & csr_wdata_int[30];
  assign N9905 = 1'b0 & csr_wdata_int[29];
  assign N9906 = 1'b0 & csr_wdata_int[28];
  assign N9907 = 1'b0 & csr_wdata_int[27];
  assign N9908 = 1'b0 & csr_wdata_int[26];
  assign N9909 = 1'b0 & csr_wdata_int[25];
  assign N9910 = 1'b0 & csr_wdata_int[24];
  assign N9911 = 1'b0 & csr_wdata_int[23];
  assign N9912 = 1'b0 & csr_wdata_int[22];
  assign N9913 = 1'b0 & csr_wdata_int[21];
  assign N9914 = 1'b0 & csr_wdata_int[20];
  assign N9915 = 1'b0 & csr_wdata_int[19];
  assign N9916 = 1'b0 & csr_wdata_int[18];
  assign N9917 = 1'b0 & csr_wdata_int[17];
  assign N9918 = 1'b0 & csr_wdata_int[16];
  assign N9919 = 1'b0 & csr_wdata_int[15];
  assign N9920 = 1'b0 & csr_wdata_int[14];
  assign N9921 = 1'b0 & csr_wdata_int[13];
  assign N9922 = 1'b0 & csr_wdata_int[12];
  assign N9923 = 1'b0 & csr_wdata_int[11];
  assign N9924 = 1'b0 & csr_wdata_int[10];
  assign N9925 = 1'b0 & csr_wdata_int[9];
  assign N9926 = 1'b0 & csr_wdata_int[8];
  assign N9927 = 1'b0 & csr_wdata_int[7];
  assign N9928 = 1'b0 & csr_wdata_int[6];
  assign N9929 = 1'b0 & csr_wdata_int[5];
  assign N9930 = 1'b0 & csr_wdata_int[4];
  assign N9931 = 1'b0 & csr_wdata_int[3];
  assign N9932 = 1'b0 & csr_wdata_int[2];
  assign N9933 = 1'b0 & csr_wdata_int[1];
  assign N9934 = 1'b0 & csr_wdata_int[0];
  assign N9935 = ~mhpmcounterh_we[29];
  assign N9936 = 1'b0 & csr_wdata_int[31];
  assign N9937 = 1'b0 & csr_wdata_int[30];
  assign N9938 = 1'b0 & csr_wdata_int[29];
  assign N9939 = 1'b0 & csr_wdata_int[28];
  assign N9940 = 1'b0 & csr_wdata_int[27];
  assign N9941 = 1'b0 & csr_wdata_int[26];
  assign N9942 = 1'b0 & csr_wdata_int[25];
  assign N9943 = 1'b0 & csr_wdata_int[24];
  assign N9944 = 1'b0 & csr_wdata_int[23];
  assign N9945 = 1'b0 & csr_wdata_int[22];
  assign N9946 = 1'b0 & csr_wdata_int[21];
  assign N9947 = 1'b0 & csr_wdata_int[20];
  assign N9948 = 1'b0 & csr_wdata_int[19];
  assign N9949 = 1'b0 & csr_wdata_int[18];
  assign N9950 = 1'b0 & csr_wdata_int[17];
  assign N9951 = 1'b0 & csr_wdata_int[16];
  assign N9952 = 1'b0 & csr_wdata_int[15];
  assign N9953 = 1'b0 & csr_wdata_int[14];
  assign N9954 = 1'b0 & csr_wdata_int[13];
  assign N9955 = 1'b0 & csr_wdata_int[12];
  assign N9956 = 1'b0 & csr_wdata_int[11];
  assign N9957 = 1'b0 & csr_wdata_int[10];
  assign N9958 = 1'b0 & csr_wdata_int[9];
  assign N9959 = 1'b0 & csr_wdata_int[8];
  assign N9960 = 1'b0 & csr_wdata_int[7];
  assign N9961 = 1'b0 & csr_wdata_int[6];
  assign N9962 = 1'b0 & csr_wdata_int[5];
  assign N9963 = 1'b0 & csr_wdata_int[4];
  assign N9964 = 1'b0 & csr_wdata_int[3];
  assign N9965 = 1'b0 & csr_wdata_int[2];
  assign N9966 = 1'b0 & csr_wdata_int[1];
  assign N9967 = 1'b0 & csr_wdata_int[0];
  assign N10000 = 1'b0 & N10735;
  assign N10735 = ~mcountinhibit[30];
  assign N10001 = ~N10000;
  assign N10066 = 1'b0 & N10065;
  assign N10067 = 1'b0 & N10064;
  assign N10068 = 1'b0 & N10063;
  assign N10069 = 1'b0 & N10062;
  assign N10070 = 1'b0 & N10061;
  assign N10071 = 1'b0 & N10060;
  assign N10072 = 1'b0 & N10059;
  assign N10073 = 1'b0 & N10058;
  assign N10074 = 1'b0 & N10057;
  assign N10075 = 1'b0 & N10056;
  assign N10076 = 1'b0 & N10055;
  assign N10077 = 1'b0 & N10054;
  assign N10078 = 1'b0 & N10053;
  assign N10079 = 1'b0 & N10052;
  assign N10080 = 1'b0 & N10051;
  assign N10081 = 1'b0 & N10050;
  assign N10082 = 1'b0 & N10049;
  assign N10083 = 1'b0 & N10048;
  assign N10084 = 1'b0 & N10047;
  assign N10085 = 1'b0 & N10046;
  assign N10086 = 1'b0 & N10045;
  assign N10087 = 1'b0 & N10044;
  assign N10088 = 1'b0 & N10043;
  assign N10089 = 1'b0 & N10042;
  assign N10090 = 1'b0 & N10041;
  assign N10091 = 1'b0 & N10040;
  assign N10092 = 1'b0 & N10039;
  assign N10093 = 1'b0 & N10038;
  assign N10094 = 1'b0 & N10037;
  assign N10095 = 1'b0 & N10036;
  assign N10096 = 1'b0 & N10035;
  assign N10097 = 1'b0 & N10034;
  assign N10098 = 1'b0 & N10033;
  assign N10099 = 1'b0 & N10032;
  assign N10100 = 1'b0 & N10031;
  assign N10101 = 1'b0 & N10030;
  assign N10102 = 1'b0 & N10029;
  assign N10103 = 1'b0 & N10028;
  assign N10104 = 1'b0 & N10027;
  assign N10105 = 1'b0 & N10026;
  assign N10106 = 1'b0 & N10025;
  assign N10107 = 1'b0 & N10024;
  assign N10108 = 1'b0 & N10023;
  assign N10109 = 1'b0 & N10022;
  assign N10110 = 1'b0 & N10021;
  assign N10111 = 1'b0 & N10020;
  assign N10112 = 1'b0 & N10019;
  assign N10113 = 1'b0 & N10018;
  assign N10114 = 1'b0 & N10017;
  assign N10115 = 1'b0 & N10016;
  assign N10116 = 1'b0 & N10015;
  assign N10117 = 1'b0 & N10014;
  assign N10118 = 1'b0 & N10013;
  assign N10119 = 1'b0 & N10012;
  assign N10120 = 1'b0 & N10011;
  assign N10121 = 1'b0 & N10010;
  assign N10122 = 1'b0 & N10009;
  assign N10123 = 1'b0 & N10008;
  assign N10124 = 1'b0 & N10007;
  assign N10125 = 1'b0 & N10006;
  assign N10126 = 1'b0 & N10005;
  assign N10127 = 1'b0 & N10004;
  assign N10128 = 1'b0 & N10003;
  assign N10129 = 1'b0 & N10002;
  assign N10194 = ~mhpmcounter_we[30];
  assign N10195 = 1'b0 & csr_wdata_int[31];
  assign N10196 = 1'b0 & csr_wdata_int[30];
  assign N10197 = 1'b0 & csr_wdata_int[29];
  assign N10198 = 1'b0 & csr_wdata_int[28];
  assign N10199 = 1'b0 & csr_wdata_int[27];
  assign N10200 = 1'b0 & csr_wdata_int[26];
  assign N10201 = 1'b0 & csr_wdata_int[25];
  assign N10202 = 1'b0 & csr_wdata_int[24];
  assign N10203 = 1'b0 & csr_wdata_int[23];
  assign N10204 = 1'b0 & csr_wdata_int[22];
  assign N10205 = 1'b0 & csr_wdata_int[21];
  assign N10206 = 1'b0 & csr_wdata_int[20];
  assign N10207 = 1'b0 & csr_wdata_int[19];
  assign N10208 = 1'b0 & csr_wdata_int[18];
  assign N10209 = 1'b0 & csr_wdata_int[17];
  assign N10210 = 1'b0 & csr_wdata_int[16];
  assign N10211 = 1'b0 & csr_wdata_int[15];
  assign N10212 = 1'b0 & csr_wdata_int[14];
  assign N10213 = 1'b0 & csr_wdata_int[13];
  assign N10214 = 1'b0 & csr_wdata_int[12];
  assign N10215 = 1'b0 & csr_wdata_int[11];
  assign N10216 = 1'b0 & csr_wdata_int[10];
  assign N10217 = 1'b0 & csr_wdata_int[9];
  assign N10218 = 1'b0 & csr_wdata_int[8];
  assign N10219 = 1'b0 & csr_wdata_int[7];
  assign N10220 = 1'b0 & csr_wdata_int[6];
  assign N10221 = 1'b0 & csr_wdata_int[5];
  assign N10222 = 1'b0 & csr_wdata_int[4];
  assign N10223 = 1'b0 & csr_wdata_int[3];
  assign N10224 = 1'b0 & csr_wdata_int[2];
  assign N10225 = 1'b0 & csr_wdata_int[1];
  assign N10226 = 1'b0 & csr_wdata_int[0];
  assign N10227 = ~mhpmcounterh_we[30];
  assign N10228 = 1'b0 & csr_wdata_int[31];
  assign N10229 = 1'b0 & csr_wdata_int[30];
  assign N10230 = 1'b0 & csr_wdata_int[29];
  assign N10231 = 1'b0 & csr_wdata_int[28];
  assign N10232 = 1'b0 & csr_wdata_int[27];
  assign N10233 = 1'b0 & csr_wdata_int[26];
  assign N10234 = 1'b0 & csr_wdata_int[25];
  assign N10235 = 1'b0 & csr_wdata_int[24];
  assign N10236 = 1'b0 & csr_wdata_int[23];
  assign N10237 = 1'b0 & csr_wdata_int[22];
  assign N10238 = 1'b0 & csr_wdata_int[21];
  assign N10239 = 1'b0 & csr_wdata_int[20];
  assign N10240 = 1'b0 & csr_wdata_int[19];
  assign N10241 = 1'b0 & csr_wdata_int[18];
  assign N10242 = 1'b0 & csr_wdata_int[17];
  assign N10243 = 1'b0 & csr_wdata_int[16];
  assign N10244 = 1'b0 & csr_wdata_int[15];
  assign N10245 = 1'b0 & csr_wdata_int[14];
  assign N10246 = 1'b0 & csr_wdata_int[13];
  assign N10247 = 1'b0 & csr_wdata_int[12];
  assign N10248 = 1'b0 & csr_wdata_int[11];
  assign N10249 = 1'b0 & csr_wdata_int[10];
  assign N10250 = 1'b0 & csr_wdata_int[9];
  assign N10251 = 1'b0 & csr_wdata_int[8];
  assign N10252 = 1'b0 & csr_wdata_int[7];
  assign N10253 = 1'b0 & csr_wdata_int[6];
  assign N10254 = 1'b0 & csr_wdata_int[5];
  assign N10255 = 1'b0 & csr_wdata_int[4];
  assign N10256 = 1'b0 & csr_wdata_int[3];
  assign N10257 = 1'b0 & csr_wdata_int[2];
  assign N10258 = 1'b0 & csr_wdata_int[1];
  assign N10259 = 1'b0 & csr_wdata_int[0];
  assign N10292 = 1'b0 & N10736;
  assign N10736 = ~mcountinhibit[31];
  assign N10293 = ~N10292;
  assign N10358 = 1'b0 & N10357;
  assign N10359 = 1'b0 & N10356;
  assign N10360 = 1'b0 & N10355;
  assign N10361 = 1'b0 & N10354;
  assign N10362 = 1'b0 & N10353;
  assign N10363 = 1'b0 & N10352;
  assign N10364 = 1'b0 & N10351;
  assign N10365 = 1'b0 & N10350;
  assign N10366 = 1'b0 & N10349;
  assign N10367 = 1'b0 & N10348;
  assign N10368 = 1'b0 & N10347;
  assign N10369 = 1'b0 & N10346;
  assign N10370 = 1'b0 & N10345;
  assign N10371 = 1'b0 & N10344;
  assign N10372 = 1'b0 & N10343;
  assign N10373 = 1'b0 & N10342;
  assign N10374 = 1'b0 & N10341;
  assign N10375 = 1'b0 & N10340;
  assign N10376 = 1'b0 & N10339;
  assign N10377 = 1'b0 & N10338;
  assign N10378 = 1'b0 & N10337;
  assign N10379 = 1'b0 & N10336;
  assign N10380 = 1'b0 & N10335;
  assign N10381 = 1'b0 & N10334;
  assign N10382 = 1'b0 & N10333;
  assign N10383 = 1'b0 & N10332;
  assign N10384 = 1'b0 & N10331;
  assign N10385 = 1'b0 & N10330;
  assign N10386 = 1'b0 & N10329;
  assign N10387 = 1'b0 & N10328;
  assign N10388 = 1'b0 & N10327;
  assign N10389 = 1'b0 & N10326;
  assign N10390 = 1'b0 & N10325;
  assign N10391 = 1'b0 & N10324;
  assign N10392 = 1'b0 & N10323;
  assign N10393 = 1'b0 & N10322;
  assign N10394 = 1'b0 & N10321;
  assign N10395 = 1'b0 & N10320;
  assign N10396 = 1'b0 & N10319;
  assign N10397 = 1'b0 & N10318;
  assign N10398 = 1'b0 & N10317;
  assign N10399 = 1'b0 & N10316;
  assign N10400 = 1'b0 & N10315;
  assign N10401 = 1'b0 & N10314;
  assign N10402 = 1'b0 & N10313;
  assign N10403 = 1'b0 & N10312;
  assign N10404 = 1'b0 & N10311;
  assign N10405 = 1'b0 & N10310;
  assign N10406 = 1'b0 & N10309;
  assign N10407 = 1'b0 & N10308;
  assign N10408 = 1'b0 & N10307;
  assign N10409 = 1'b0 & N10306;
  assign N10410 = 1'b0 & N10305;
  assign N10411 = 1'b0 & N10304;
  assign N10412 = 1'b0 & N10303;
  assign N10413 = 1'b0 & N10302;
  assign N10414 = 1'b0 & N10301;
  assign N10415 = 1'b0 & N10300;
  assign N10416 = 1'b0 & N10299;
  assign N10417 = 1'b0 & N10298;
  assign N10418 = 1'b0 & N10297;
  assign N10419 = 1'b0 & N10296;
  assign N10420 = 1'b0 & N10295;
  assign N10421 = 1'b0 & N10294;
  assign N10486 = ~mhpmcounter_we[31];
  assign N10487 = 1'b0 & csr_wdata_int[31];
  assign N10488 = 1'b0 & csr_wdata_int[30];
  assign N10489 = 1'b0 & csr_wdata_int[29];
  assign N10490 = 1'b0 & csr_wdata_int[28];
  assign N10491 = 1'b0 & csr_wdata_int[27];
  assign N10492 = 1'b0 & csr_wdata_int[26];
  assign N10493 = 1'b0 & csr_wdata_int[25];
  assign N10494 = 1'b0 & csr_wdata_int[24];
  assign N10495 = 1'b0 & csr_wdata_int[23];
  assign N10496 = 1'b0 & csr_wdata_int[22];
  assign N10497 = 1'b0 & csr_wdata_int[21];
  assign N10498 = 1'b0 & csr_wdata_int[20];
  assign N10499 = 1'b0 & csr_wdata_int[19];
  assign N10500 = 1'b0 & csr_wdata_int[18];
  assign N10501 = 1'b0 & csr_wdata_int[17];
  assign N10502 = 1'b0 & csr_wdata_int[16];
  assign N10503 = 1'b0 & csr_wdata_int[15];
  assign N10504 = 1'b0 & csr_wdata_int[14];
  assign N10505 = 1'b0 & csr_wdata_int[13];
  assign N10506 = 1'b0 & csr_wdata_int[12];
  assign N10507 = 1'b0 & csr_wdata_int[11];
  assign N10508 = 1'b0 & csr_wdata_int[10];
  assign N10509 = 1'b0 & csr_wdata_int[9];
  assign N10510 = 1'b0 & csr_wdata_int[8];
  assign N10511 = 1'b0 & csr_wdata_int[7];
  assign N10512 = 1'b0 & csr_wdata_int[6];
  assign N10513 = 1'b0 & csr_wdata_int[5];
  assign N10514 = 1'b0 & csr_wdata_int[4];
  assign N10515 = 1'b0 & csr_wdata_int[3];
  assign N10516 = 1'b0 & csr_wdata_int[2];
  assign N10517 = 1'b0 & csr_wdata_int[1];
  assign N10518 = 1'b0 & csr_wdata_int[0];
  assign N10519 = ~mhpmcounterh_we[31];
  assign N10520 = 1'b0 & csr_wdata_int[31];
  assign N10521 = 1'b0 & csr_wdata_int[30];
  assign N10522 = 1'b0 & csr_wdata_int[29];
  assign N10523 = 1'b0 & csr_wdata_int[28];
  assign N10524 = 1'b0 & csr_wdata_int[27];
  assign N10525 = 1'b0 & csr_wdata_int[26];
  assign N10526 = 1'b0 & csr_wdata_int[25];
  assign N10527 = 1'b0 & csr_wdata_int[24];
  assign N10528 = 1'b0 & csr_wdata_int[23];
  assign N10529 = 1'b0 & csr_wdata_int[22];
  assign N10530 = 1'b0 & csr_wdata_int[21];
  assign N10531 = 1'b0 & csr_wdata_int[20];
  assign N10532 = 1'b0 & csr_wdata_int[19];
  assign N10533 = 1'b0 & csr_wdata_int[18];
  assign N10534 = 1'b0 & csr_wdata_int[17];
  assign N10535 = 1'b0 & csr_wdata_int[16];
  assign N10536 = 1'b0 & csr_wdata_int[15];
  assign N10537 = 1'b0 & csr_wdata_int[14];
  assign N10538 = 1'b0 & csr_wdata_int[13];
  assign N10539 = 1'b0 & csr_wdata_int[12];
  assign N10540 = 1'b0 & csr_wdata_int[11];
  assign N10541 = 1'b0 & csr_wdata_int[10];
  assign N10542 = 1'b0 & csr_wdata_int[9];
  assign N10543 = 1'b0 & csr_wdata_int[8];
  assign N10544 = 1'b0 & csr_wdata_int[7];
  assign N10545 = 1'b0 & csr_wdata_int[6];
  assign N10546 = 1'b0 & csr_wdata_int[5];
  assign N10547 = 1'b0 & csr_wdata_int[4];
  assign N10548 = 1'b0 & csr_wdata_int[3];
  assign N10549 = 1'b0 & csr_wdata_int[2];
  assign N10550 = 1'b0 & csr_wdata_int[1];
  assign N10551 = 1'b0 & csr_wdata_int[0];
  assign N10584 = N409 | N411;
  assign N10585 = N10584 | N413;
  assign N10586 = N10585 | N415;
  assign N10587 = N10586 | N421;
  assign N10588 = N10587 | N423;
  assign N10589 = N10588 | N427;
  assign N10590 = N10589 | N429;
  assign N10591 = N10590 | N447;
  assign N10592 = N10591 | N449;
  assign N10593 = N10592 | N453;
  assign N10594 = N10593 | N458;
  assign N10595 = N10594 | N470;
  assign N10596 = ~N10595;
  assign N10597 = N409 | N413;
  assign N10598 = N10597 | N415;
  assign N10599 = N10598 | N421;
  assign N10600 = N10599 | N423;
  assign N10601 = N10600 | N427;
  assign N10602 = N10601 | N429;
  assign N10603 = N10602 | N440;
  assign N10604 = N10603 | N447;
  assign N10605 = N10604 | N449;
  assign N10606 = N10605 | N453;
  assign N10607 = N10606 | N458;
  assign N10608 = N10607 | N470;
  assign N10609 = ~N10608;
  assign N10610 = N10589 | N440;
  assign N10611 = N10610 | N447;
  assign N10612 = N10611 | N449;
  assign N10613 = N10612 | N453;
  assign N10614 = N10613 | N458;
  assign N10615 = N10614 | N470;
  assign N10616 = ~N10615;

endmodule



module ibex_core
(
  clk_i,
  rst_ni,
  test_en_i,
  core_id_i,
  cluster_id_i,
  boot_addr_i,
  instr_req_o,
  instr_gnt_i,
  instr_rvalid_i,
  instr_addr_o,
  instr_rdata_i,
  data_req_o,
  data_gnt_i,
  data_rvalid_i,
  data_we_o,
  data_be_o,
  data_addr_o,
  data_wdata_o,
  data_rdata_i,
  data_err_i,
  irq_i,
  irq_id_i,
  irq_ack_o,
  irq_id_o,
  debug_req_i,
  fetch_enable_i
);

  input [3:0] core_id_i;
  input [5:0] cluster_id_i;
  input [31:0] boot_addr_i;
  output [31:0] instr_addr_o;
  input [31:0] instr_rdata_i;
  output [3:0] data_be_o;
  output [31:0] data_addr_o;
  output [31:0] data_wdata_o;
  input [31:0] data_rdata_i;
  input [4:0] irq_id_i;
  output [4:0] irq_id_o;
  input clk_i;
  input rst_ni;
  input test_en_i;
  input instr_gnt_i;
  input instr_rvalid_i;
  input data_gnt_i;
  input data_rvalid_i;
  input data_err_i;
  input irq_i;
  input debug_req_i;
  input fetch_enable_i;
  output instr_req_o;
  output data_req_o;
  output data_we_o;
  output irq_ack_o;
  wire [31:0] instr_addr_o,data_addr_o,data_wdata_o,instr_rdata_id,pc_if,pc_id,jump_target_ex,
  csr_mepc,csr_depc,csr_mtvec,alu_operand_a_ex,alu_operand_b_ex,
  multdiv_operand_a_ex,multdiv_operand_b_ex,csr_mtval,data_wdata_ex,lsu_addr_last,regfile_wdata_lsu,
  regfile_wdata_ex,csr_rdata,alu_adder_result_ex;
  wire [3:0] data_be_o;
  wire [4:0] irq_id_o,alu_operator_ex;
  wire instr_req_o,data_req_o,data_we_o,irq_ack_o,N0,N1,N2,N3,if_busy,ctrl_busy,
  lsu_busy,core_busy_int,N4,core_ctrl_firstfetch,N5,core_busy,clock_en,clk,instr_req_int,
  instr_valid_id,instr_new_id,instr_is_compressed_id,illegal_c_insn_id,
  instr_valid_clear,pc_set,id_in_ready,perf_imiss,illegal_insn_id,branch_decision,ex_valid,
  lsu_data_valid,mult_en_ex,div_en_ex,csr_access,csr_save_if,csr_save_id,
  csr_restore_mret_id,csr_restore_dret_id,csr_save_cause,illegal_csr_insn_id,data_req_ex,
  data_we_ex,data_sign_ext_ex,lsu_addr_incr_req,lsu_load_err,lsu_store_err,
  m_irq_enable,debug_csr_save,debug_single_step,debug_ebreakm,perf_jump,perf_branch,
  perf_tbranch,instr_ret,instr_ret_compressed,N6,N7,perf_load,perf_store,N8,N9,N10,N11,N12;
  wire [15:0] instr_rdata_c_id;
  wire [2:0] pc_mux_id,debug_cause;
  wire [1:0] exc_pc_mux_id,multdiv_operator_ex,multdiv_signed_mode_ex,csr_op,data_type_ex,
  data_reg_offset_ex;
  wire [5:0] exc_cause;
  wire [11:0] csr_addr;
  reg core_busy_q;

  always @(posedge clk_i or posedge N4) begin
    if(N4) begin
      core_busy_q <= 1'b0;
    end else if(1'b1) begin
      core_busy_q <= core_busy_int;
    end 
  end


  prim_clock_gating
  core_clock_gate_i
  (
    .clk_i(clk_i),
    .en_i(clock_en),
    .test_en_i(test_en_i),
    .clk_o(clk)
  );


  ibex_if_stage_1a110800_1a110808
  if_stage_i
  (
    .clk_i(clk),
    .rst_ni(rst_ni),
    .boot_addr_i(boot_addr_i),
    .req_i(instr_req_int),
    .instr_req_o(instr_req_o),
    .instr_addr_o(instr_addr_o),
    .instr_gnt_i(instr_gnt_i),
    .instr_rvalid_i(instr_rvalid_i),
    .instr_rdata_i(instr_rdata_i),
    .instr_valid_id_o(instr_valid_id),
    .instr_new_id_o(instr_new_id),
    .instr_rdata_id_o(instr_rdata_id),
    .instr_rdata_c_id_o(instr_rdata_c_id),
    .instr_is_compressed_id_o(instr_is_compressed_id),
    .illegal_c_insn_id_o(illegal_c_insn_id),
    .pc_if_o(pc_if),
    .pc_id_o(pc_id),
    .instr_valid_clear_i(instr_valid_clear),
    .pc_set_i(pc_set),
    .csr_mepc_i(csr_mepc),
    .csr_depc_i(csr_depc),
    .pc_mux_i(pc_mux_id),
    .exc_pc_mux_i(exc_pc_mux_id),
    .exc_cause(exc_cause),
    .jump_target_ex_i(jump_target_ex),
    .csr_mtvec_o(csr_mtvec),
    .id_in_ready_i(id_in_ready),
    .if_busy_o(if_busy),
    .perf_imiss_o(perf_imiss)
  );


  ibex_id_stage_0_1
  id_stage_i
  (
    .clk_i(clk),
    .rst_ni(rst_ni),
    .test_en_i(test_en_i),
    .fetch_enable_i(fetch_enable_i),
    .ctrl_busy_o(ctrl_busy),
    .core_ctrl_firstfetch_o(core_ctrl_firstfetch),
    .illegal_insn_o(illegal_insn_id),
    .instr_valid_i(instr_valid_id),
    .instr_new_i(instr_new_id),
    .instr_rdata_i(instr_rdata_id),
    .instr_rdata_c_i(instr_rdata_c_id),
    .instr_is_compressed_i(instr_is_compressed_id),
    .instr_req_o(instr_req_int),
    .instr_valid_clear_o(instr_valid_clear),
    .id_in_ready_o(id_in_ready),
    .branch_decision_i(branch_decision),
    .pc_set_o(pc_set),
    .pc_mux_o(pc_mux_id),
    .exc_pc_mux_o(exc_pc_mux_id),
    .illegal_c_insn_i(illegal_c_insn_id),
    .pc_id_i(pc_id),
    .ex_valid_i(ex_valid),
    .lsu_valid_i(lsu_data_valid),
    .alu_operator_ex_o(alu_operator_ex),
    .alu_operand_a_ex_o(alu_operand_a_ex),
    .alu_operand_b_ex_o(alu_operand_b_ex),
    .mult_en_ex_o(mult_en_ex),
    .div_en_ex_o(div_en_ex),
    .multdiv_operator_ex_o(multdiv_operator_ex),
    .multdiv_signed_mode_ex_o(multdiv_signed_mode_ex),
    .multdiv_operand_a_ex_o(multdiv_operand_a_ex),
    .multdiv_operand_b_ex_o(multdiv_operand_b_ex),
    .csr_access_o(csr_access),
    .csr_op_o(csr_op),
    .csr_save_if_o(csr_save_if),
    .csr_save_id_o(csr_save_id),
    .csr_restore_mret_id_o(csr_restore_mret_id),
    .csr_restore_dret_id_o(csr_restore_dret_id),
    .csr_save_cause_o(csr_save_cause),
    .csr_mtval_o(csr_mtval),
    .illegal_csr_insn_i(illegal_csr_insn_id),
    .data_req_ex_o(data_req_ex),
    .data_we_ex_o(data_we_ex),
    .data_type_ex_o(data_type_ex),
    .data_sign_ext_ex_o(data_sign_ext_ex),
    .data_reg_offset_ex_o(data_reg_offset_ex),
    .data_wdata_ex_o(data_wdata_ex),
    .lsu_addr_incr_req_i(lsu_addr_incr_req),
    .lsu_addr_last_i(lsu_addr_last),
    .irq_i(irq_i),
    .irq_id_i(irq_id_i),
    .m_irq_enable_i(m_irq_enable),
    .irq_ack_o(irq_ack_o),
    .irq_id_o(irq_id_o),
    .exc_cause_o(exc_cause),
    .lsu_load_err_i(lsu_load_err),
    .lsu_store_err_i(lsu_store_err),
    .debug_cause_o(debug_cause),
    .debug_csr_save_o(debug_csr_save),
    .debug_req_i(debug_req_i),
    .debug_single_step_i(debug_single_step),
    .debug_ebreakm_i(debug_ebreakm),
    .regfile_wdata_lsu_i(regfile_wdata_lsu),
    .regfile_wdata_ex_i(regfile_wdata_ex),
    .csr_rdata_i(csr_rdata),
    .perf_jump_o(perf_jump),
    .perf_branch_o(perf_branch),
    .perf_tbranch_o(perf_tbranch),
    .instr_ret_o(instr_ret),
    .instr_ret_compressed_o(instr_ret_compressed)
  );


  ibex_ex_block_1
  ex_block_i
  (
    .clk_i(clk),
    .rst_ni(rst_ni),
    .alu_operator_i(alu_operator_ex),
    .alu_operand_a_i(alu_operand_a_ex),
    .alu_operand_b_i(alu_operand_b_ex),
    .multdiv_operator_i(multdiv_operator_ex),
    .mult_en_i(mult_en_ex),
    .div_en_i(div_en_ex),
    .multdiv_signed_mode_i(multdiv_signed_mode_ex),
    .multdiv_operand_a_i(multdiv_operand_a_ex),
    .multdiv_operand_b_i(multdiv_operand_b_ex),
    .alu_adder_result_ex_o(alu_adder_result_ex),
    .regfile_wdata_ex_o(regfile_wdata_ex),
    .jump_target_o(jump_target_ex),
    .branch_decision_o(branch_decision),
    .ex_valid_o(ex_valid)
  );


  ibex_load_store_unit
  load_store_unit_i
  (
    .clk_i(clk),
    .rst_ni(rst_ni),
    .data_req_o(data_req_o),
    .data_gnt_i(data_gnt_i),
    .data_rvalid_i(data_rvalid_i),
    .data_err_i(data_err_i),
    .data_addr_o(data_addr_o),
    .data_we_o(data_we_o),
    .data_be_o(data_be_o),
    .data_wdata_o(data_wdata_o),
    .data_rdata_i(data_rdata_i),
    .data_we_ex_i(data_we_ex),
    .data_type_ex_i(data_type_ex),
    .data_wdata_ex_i(data_wdata_ex),
    .data_reg_offset_ex_i(data_reg_offset_ex),
    .data_sign_ext_ex_i(data_sign_ext_ex),
    .data_rdata_ex_o(regfile_wdata_lsu),
    .data_req_ex_i(data_req_ex),
    .adder_result_ex_i(alu_adder_result_ex),
    .addr_incr_req_o(lsu_addr_incr_req),
    .addr_last_o(lsu_addr_last),
    .data_valid_o(lsu_data_valid),
    .load_err_o(lsu_load_err),
    .store_err_o(lsu_store_err),
    .busy_o(lsu_busy)
  );


  ibex_cs_registers_00000000_00000028_0_1
  cs_registers_i
  (
    .clk_i(clk),
    .rst_ni(rst_ni),
    .core_id_i(core_id_i),
    .cluster_id_i(cluster_id_i),
    .csr_access_i(csr_access),
    .csr_addr_i(csr_addr),
    .csr_wdata_i(alu_operand_a_ex),
    .csr_op_i(csr_op),
    .csr_rdata_o(csr_rdata),
    .m_irq_enable_o(m_irq_enable),
    .csr_mepc_o(csr_mepc),
    .debug_cause_i(debug_cause),
    .debug_csr_save_i(debug_csr_save),
    .csr_depc_o(csr_depc),
    .debug_single_step_o(debug_single_step),
    .debug_ebreakm_o(debug_ebreakm),
    .pc_if_i(pc_if),
    .pc_id_i(pc_id),
    .csr_save_if_i(csr_save_if),
    .csr_save_id_i(csr_save_id),
    .csr_restore_mret_i(csr_restore_mret_id),
    .csr_restore_dret_i(csr_restore_dret_id),
    .csr_save_cause_i(csr_save_cause),
    .csr_mtvec_i(csr_mtvec),
    .csr_mcause_i(exc_cause),
    .csr_mtval_i(csr_mtval),
    .illegal_csr_insn_o(illegal_csr_insn_id),
    .instr_new_id_i(instr_new_id),
    .instr_ret_i(instr_ret),
    .instr_ret_compressed_i(instr_ret_compressed),
    .imiss_i(perf_imiss),
    .pc_set_i(pc_set),
    .jump_i(perf_jump),
    .branch_i(perf_branch),
    .branch_taken_i(perf_tbranch),
    .mem_load_i(perf_load),
    .mem_store_i(perf_store),
    .lsu_busy_i(lsu_busy)
  );

  assign core_busy = (N0)? 1'b1 : 
                     (N1)? core_busy_q : 1'b0;
  assign N0 = core_ctrl_firstfetch;
  assign N1 = N5;
  assign csr_addr = (N2)? alu_operand_b_ex[11:0] : 
                    (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N2 = N7;
  assign N3 = N6;
  assign core_busy_int = N8 | lsu_busy;
  assign N8 = if_busy | ctrl_busy;
  assign N4 = ~rst_ni;
  assign N5 = ~core_ctrl_firstfetch;
  assign clock_en = N9 | debug_req_i;
  assign N9 = core_busy | irq_i;
  assign N6 = ~csr_access;
  assign N7 = csr_access;
  assign perf_load = N10 & N11;
  assign N10 = data_req_o & data_gnt_i;
  assign N11 = ~data_we_o;
  assign perf_store = N12 & data_we_o;
  assign N12 = data_req_o & data_gnt_i;

endmodule

