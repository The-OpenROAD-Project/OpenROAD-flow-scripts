VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram130_2x576
  FOREIGN fakeram130_2x576 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 589.570 BY 169.400 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 23.500 1.000 24.500 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 28.300 1.000 29.300 ;
    END
  END w_mask_in[1]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 35.500 1.000 36.500 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 40.300 1.000 41.300 ;
    END
  END rd_out[1]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 47.500 1.000 48.500 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 52.300 1.000 53.300 ;
    END
  END wd_in[1]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 59.500 1.000 60.500 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 64.300 1.000 65.300 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 69.100 1.000 70.100 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 73.900 1.000 74.900 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 78.700 1.000 79.700 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 83.500 1.000 84.500 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 88.300 1.000 89.300 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 93.100 1.000 94.100 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 97.900 1.000 98.900 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 102.700 1.000 103.700 ;
    END
  END addr_in[9]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 109.900 1.000 110.900 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 114.700 1.000 115.700 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 119.500 1.000 120.500 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
      RECT 22.000 24.000 26.000 145.400 ;
      RECT 60.400 24.000 64.400 145.400 ;
      RECT 98.800 24.000 102.800 145.400 ;
      RECT 137.200 24.000 141.200 145.400 ;
      RECT 175.600 24.000 179.600 145.400 ;
      RECT 214.000 24.000 218.000 145.400 ;
      RECT 252.400 24.000 256.400 145.400 ;
      RECT 290.800 24.000 294.800 145.400 ;
      RECT 329.200 24.000 333.200 145.400 ;
      RECT 367.600 24.000 371.600 145.400 ;
      RECT 406.000 24.000 410.000 145.400 ;
      RECT 444.400 24.000 448.400 145.400 ;
      RECT 482.800 24.000 486.800 145.400 ;
      RECT 521.200 24.000 525.200 145.400 ;
      RECT 559.600 24.000 563.600 145.400 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
      RECT 41.200 24.000 45.200 145.400 ;
      RECT 79.600 24.000 83.600 145.400 ;
      RECT 118.000 24.000 122.000 145.400 ;
      RECT 156.400 24.000 160.400 145.400 ;
      RECT 194.800 24.000 198.800 145.400 ;
      RECT 233.200 24.000 237.200 145.400 ;
      RECT 271.600 24.000 275.600 145.400 ;
      RECT 310.000 24.000 314.000 145.400 ;
      RECT 348.400 24.000 352.400 145.400 ;
      RECT 386.800 24.000 390.800 145.400 ;
      RECT 425.200 24.000 429.200 145.400 ;
      RECT 463.600 24.000 467.600 145.400 ;
      RECT 502.000 24.000 506.000 145.400 ;
      RECT 540.400 24.000 544.400 145.400 ;
    END
  END VDD
  OBS
    LAYER met1 ;
    RECT 0 0 589.570 169.400 ;
    LAYER met2 ;
    RECT 0 0 589.570 169.400 ;
    LAYER met3 ;
    RECT 1.000 0 589.570 169.400 ;
    RECT 0 0.000 1.000 23.500 ;
    RECT 0 24.500 1.000 28.300 ;
    RECT 0 29.300 1.000 35.500 ;
    RECT 0 36.500 1.000 40.300 ;
    RECT 0 41.300 1.000 47.500 ;
    RECT 0 48.500 1.000 52.300 ;
    RECT 0 53.300 1.000 59.500 ;
    RECT 0 60.500 1.000 64.300 ;
    RECT 0 65.300 1.000 69.100 ;
    RECT 0 70.100 1.000 73.900 ;
    RECT 0 74.900 1.000 78.700 ;
    RECT 0 79.700 1.000 83.500 ;
    RECT 0 84.500 1.000 88.300 ;
    RECT 0 89.300 1.000 93.100 ;
    RECT 0 94.100 1.000 97.900 ;
    RECT 0 98.900 1.000 102.700 ;
    RECT 0 103.700 1.000 109.900 ;
    RECT 0 110.900 1.000 114.700 ;
    RECT 0 115.700 1.000 119.500 ;
    RECT 0 120.500 1.000 169.400 ;
    LAYER met4 ;
    RECT 0 0 589.570 24.000 ;
    RECT 0 145.400 589.570 169.400 ;
    RECT 0.000 24.000 22.000 145.400 ;
    RECT 26.000 24.000 41.200 145.400 ;
    RECT 45.200 24.000 60.400 145.400 ;
    RECT 64.400 24.000 79.600 145.400 ;
    RECT 83.600 24.000 98.800 145.400 ;
    RECT 102.800 24.000 118.000 145.400 ;
    RECT 122.000 24.000 137.200 145.400 ;
    RECT 141.200 24.000 156.400 145.400 ;
    RECT 160.400 24.000 175.600 145.400 ;
    RECT 179.600 24.000 194.800 145.400 ;
    RECT 198.800 24.000 214.000 145.400 ;
    RECT 218.000 24.000 233.200 145.400 ;
    RECT 237.200 24.000 252.400 145.400 ;
    RECT 256.400 24.000 271.600 145.400 ;
    RECT 275.600 24.000 290.800 145.400 ;
    RECT 294.800 24.000 310.000 145.400 ;
    RECT 314.000 24.000 329.200 145.400 ;
    RECT 333.200 24.000 348.400 145.400 ;
    RECT 352.400 24.000 367.600 145.400 ;
    RECT 371.600 24.000 386.800 145.400 ;
    RECT 390.800 24.000 406.000 145.400 ;
    RECT 410.000 24.000 425.200 145.400 ;
    RECT 429.200 24.000 444.400 145.400 ;
    RECT 448.400 24.000 463.600 145.400 ;
    RECT 467.600 24.000 482.800 145.400 ;
    RECT 486.800 24.000 502.000 145.400 ;
    RECT 506.000 24.000 521.200 145.400 ;
    RECT 525.200 24.000 540.400 145.400 ;
    RECT 544.400 24.000 559.600 145.400 ;
    RECT 563.600 24.000 589.570 145.400 ;
    LAYER OVERLAP ;
    RECT 0 0 589.570 169.400 ;
  END
END fakeram130_2x576

END LIBRARY
