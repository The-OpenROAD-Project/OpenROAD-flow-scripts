VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_64x96
  FOREIGN fakeram45_64x96 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 54.530 BY 77.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.400 0.070 1.470 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.540 0.070 1.610 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.680 0.070 1.750 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.820 0.070 1.890 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.960 0.070 2.030 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.100 0.070 2.170 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.240 0.070 2.310 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.380 0.070 2.450 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.520 0.070 2.590 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.660 0.070 2.730 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.800 0.070 2.870 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.940 0.070 3.010 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.080 0.070 3.150 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.220 0.070 3.290 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.360 0.070 3.430 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.500 0.070 3.570 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.640 0.070 3.710 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.780 0.070 3.850 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.920 0.070 3.990 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.060 0.070 4.130 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.200 0.070 4.270 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.340 0.070 4.410 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.480 0.070 4.550 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.620 0.070 4.690 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.760 0.070 4.830 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.900 0.070 4.970 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.040 0.070 5.110 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.180 0.070 5.250 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.320 0.070 5.390 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.460 0.070 5.530 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.600 0.070 5.670 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.740 0.070 5.810 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.880 0.070 5.950 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.020 0.070 6.090 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.160 0.070 6.230 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.300 0.070 6.370 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.440 0.070 6.510 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.580 0.070 6.650 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.720 0.070 6.790 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.860 0.070 6.930 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.000 0.070 7.070 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.140 0.070 7.210 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.280 0.070 7.350 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.420 0.070 7.490 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.560 0.070 7.630 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.700 0.070 7.770 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.840 0.070 7.910 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.980 0.070 8.050 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.120 0.070 8.190 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.260 0.070 8.330 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.400 0.070 8.470 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.540 0.070 8.610 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.680 0.070 8.750 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.820 0.070 8.890 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.960 0.070 9.030 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.100 0.070 9.170 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.240 0.070 9.310 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.380 0.070 9.450 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.520 0.070 9.590 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.660 0.070 9.730 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.800 0.070 9.870 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.940 0.070 10.010 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.080 0.070 10.150 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.220 0.070 10.290 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.360 0.070 10.430 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.500 0.070 10.570 ;
    END
  END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.640 0.070 10.710 ;
    END
  END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.780 0.070 10.850 ;
    END
  END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.920 0.070 10.990 ;
    END
  END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.060 0.070 11.130 ;
    END
  END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.200 0.070 11.270 ;
    END
  END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.340 0.070 11.410 ;
    END
  END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.480 0.070 11.550 ;
    END
  END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.620 0.070 11.690 ;
    END
  END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.760 0.070 11.830 ;
    END
  END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.900 0.070 11.970 ;
    END
  END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.040 0.070 12.110 ;
    END
  END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.180 0.070 12.250 ;
    END
  END w_mask_in[77]
  PIN w_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.320 0.070 12.390 ;
    END
  END w_mask_in[78]
  PIN w_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.460 0.070 12.530 ;
    END
  END w_mask_in[79]
  PIN w_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.600 0.070 12.670 ;
    END
  END w_mask_in[80]
  PIN w_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.740 0.070 12.810 ;
    END
  END w_mask_in[81]
  PIN w_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.880 0.070 12.950 ;
    END
  END w_mask_in[82]
  PIN w_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.020 0.070 13.090 ;
    END
  END w_mask_in[83]
  PIN w_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.160 0.070 13.230 ;
    END
  END w_mask_in[84]
  PIN w_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.300 0.070 13.370 ;
    END
  END w_mask_in[85]
  PIN w_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.440 0.070 13.510 ;
    END
  END w_mask_in[86]
  PIN w_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.580 0.070 13.650 ;
    END
  END w_mask_in[87]
  PIN w_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.720 0.070 13.790 ;
    END
  END w_mask_in[88]
  PIN w_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.860 0.070 13.930 ;
    END
  END w_mask_in[89]
  PIN w_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.000 0.070 14.070 ;
    END
  END w_mask_in[90]
  PIN w_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.140 0.070 14.210 ;
    END
  END w_mask_in[91]
  PIN w_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.280 0.070 14.350 ;
    END
  END w_mask_in[92]
  PIN w_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.420 0.070 14.490 ;
    END
  END w_mask_in[93]
  PIN w_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.560 0.070 14.630 ;
    END
  END w_mask_in[94]
  PIN w_mask_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.700 0.070 14.770 ;
    END
  END w_mask_in[95]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.820 0.070 22.890 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.960 0.070 23.030 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.100 0.070 23.170 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.240 0.070 23.310 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.380 0.070 23.450 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.520 0.070 23.590 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.660 0.070 23.730 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.800 0.070 23.870 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.940 0.070 24.010 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.080 0.070 24.150 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.220 0.070 24.290 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.360 0.070 24.430 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.500 0.070 24.570 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.640 0.070 24.710 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.780 0.070 24.850 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.920 0.070 24.990 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.060 0.070 25.130 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.200 0.070 25.270 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.340 0.070 25.410 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.480 0.070 25.550 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.620 0.070 25.690 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.760 0.070 25.830 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.900 0.070 25.970 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.040 0.070 26.110 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.180 0.070 26.250 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.320 0.070 26.390 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.460 0.070 26.530 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.600 0.070 26.670 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.740 0.070 26.810 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.880 0.070 26.950 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.020 0.070 27.090 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.160 0.070 27.230 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.300 0.070 27.370 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.440 0.070 27.510 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.580 0.070 27.650 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.720 0.070 27.790 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.860 0.070 27.930 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.000 0.070 28.070 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.140 0.070 28.210 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.280 0.070 28.350 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.420 0.070 28.490 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.560 0.070 28.630 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.700 0.070 28.770 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.840 0.070 28.910 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.980 0.070 29.050 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.120 0.070 29.190 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.260 0.070 29.330 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.400 0.070 29.470 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.540 0.070 29.610 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.680 0.070 29.750 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.820 0.070 29.890 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.960 0.070 30.030 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.100 0.070 30.170 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.240 0.070 30.310 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.380 0.070 30.450 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.520 0.070 30.590 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.660 0.070 30.730 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.800 0.070 30.870 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.940 0.070 31.010 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.080 0.070 31.150 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.220 0.070 31.290 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.360 0.070 31.430 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.500 0.070 31.570 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.640 0.070 31.710 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.780 0.070 31.850 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.920 0.070 31.990 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.060 0.070 32.130 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.200 0.070 32.270 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.340 0.070 32.410 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.480 0.070 32.550 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.620 0.070 32.690 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.760 0.070 32.830 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.900 0.070 32.970 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.040 0.070 33.110 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.180 0.070 33.250 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.320 0.070 33.390 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.460 0.070 33.530 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.600 0.070 33.670 ;
    END
  END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.740 0.070 33.810 ;
    END
  END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.880 0.070 33.950 ;
    END
  END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.020 0.070 34.090 ;
    END
  END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.160 0.070 34.230 ;
    END
  END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.300 0.070 34.370 ;
    END
  END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.440 0.070 34.510 ;
    END
  END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.580 0.070 34.650 ;
    END
  END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.720 0.070 34.790 ;
    END
  END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.860 0.070 34.930 ;
    END
  END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.000 0.070 35.070 ;
    END
  END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.140 0.070 35.210 ;
    END
  END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.280 0.070 35.350 ;
    END
  END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.420 0.070 35.490 ;
    END
  END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.560 0.070 35.630 ;
    END
  END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.700 0.070 35.770 ;
    END
  END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.840 0.070 35.910 ;
    END
  END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.980 0.070 36.050 ;
    END
  END rd_out[94]
  PIN rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.120 0.070 36.190 ;
    END
  END rd_out[95]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.240 0.070 44.310 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.380 0.070 44.450 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.520 0.070 44.590 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.660 0.070 44.730 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.800 0.070 44.870 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.940 0.070 45.010 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.080 0.070 45.150 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.220 0.070 45.290 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.360 0.070 45.430 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.500 0.070 45.570 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.640 0.070 45.710 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.780 0.070 45.850 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.920 0.070 45.990 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.060 0.070 46.130 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.200 0.070 46.270 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.340 0.070 46.410 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.480 0.070 46.550 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.620 0.070 46.690 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.760 0.070 46.830 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.900 0.070 46.970 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.040 0.070 47.110 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.180 0.070 47.250 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.320 0.070 47.390 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.460 0.070 47.530 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.600 0.070 47.670 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.740 0.070 47.810 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.880 0.070 47.950 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.020 0.070 48.090 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.160 0.070 48.230 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.300 0.070 48.370 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.440 0.070 48.510 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.580 0.070 48.650 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.720 0.070 48.790 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.860 0.070 48.930 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.000 0.070 49.070 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.140 0.070 49.210 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.280 0.070 49.350 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.420 0.070 49.490 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.560 0.070 49.630 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.700 0.070 49.770 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.840 0.070 49.910 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.980 0.070 50.050 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.120 0.070 50.190 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.260 0.070 50.330 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.400 0.070 50.470 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.540 0.070 50.610 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.680 0.070 50.750 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.820 0.070 50.890 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.960 0.070 51.030 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.100 0.070 51.170 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.240 0.070 51.310 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.380 0.070 51.450 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.520 0.070 51.590 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.660 0.070 51.730 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.800 0.070 51.870 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.940 0.070 52.010 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.080 0.070 52.150 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.220 0.070 52.290 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.360 0.070 52.430 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.500 0.070 52.570 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.640 0.070 52.710 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.780 0.070 52.850 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.920 0.070 52.990 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.060 0.070 53.130 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.200 0.070 53.270 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.340 0.070 53.410 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.480 0.070 53.550 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.620 0.070 53.690 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.760 0.070 53.830 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.900 0.070 53.970 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.040 0.070 54.110 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.180 0.070 54.250 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.320 0.070 54.390 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.460 0.070 54.530 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.600 0.070 54.670 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.740 0.070 54.810 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.880 0.070 54.950 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.020 0.070 55.090 ;
    END
  END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.160 0.070 55.230 ;
    END
  END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.300 0.070 55.370 ;
    END
  END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.440 0.070 55.510 ;
    END
  END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.580 0.070 55.650 ;
    END
  END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.720 0.070 55.790 ;
    END
  END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.860 0.070 55.930 ;
    END
  END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.000 0.070 56.070 ;
    END
  END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.140 0.070 56.210 ;
    END
  END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.280 0.070 56.350 ;
    END
  END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.420 0.070 56.490 ;
    END
  END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.560 0.070 56.630 ;
    END
  END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.700 0.070 56.770 ;
    END
  END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.840 0.070 56.910 ;
    END
  END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.980 0.070 57.050 ;
    END
  END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.120 0.070 57.190 ;
    END
  END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.260 0.070 57.330 ;
    END
  END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.400 0.070 57.470 ;
    END
  END wd_in[94]
  PIN wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.540 0.070 57.610 ;
    END
  END wd_in[95]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.660 0.070 65.730 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.800 0.070 65.870 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.940 0.070 66.010 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.080 0.070 66.150 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.220 0.070 66.290 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.360 0.070 66.430 ;
    END
  END addr_in[5]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.480 0.070 74.550 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.620 0.070 74.690 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.760 0.070 74.830 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 75.600 ;
      RECT 3.500 1.400 3.780 75.600 ;
      RECT 5.740 1.400 6.020 75.600 ;
      RECT 7.980 1.400 8.260 75.600 ;
      RECT 10.220 1.400 10.500 75.600 ;
      RECT 12.460 1.400 12.740 75.600 ;
      RECT 14.700 1.400 14.980 75.600 ;
      RECT 16.940 1.400 17.220 75.600 ;
      RECT 19.180 1.400 19.460 75.600 ;
      RECT 21.420 1.400 21.700 75.600 ;
      RECT 23.660 1.400 23.940 75.600 ;
      RECT 25.900 1.400 26.180 75.600 ;
      RECT 28.140 1.400 28.420 75.600 ;
      RECT 30.380 1.400 30.660 75.600 ;
      RECT 32.620 1.400 32.900 75.600 ;
      RECT 34.860 1.400 35.140 75.600 ;
      RECT 37.100 1.400 37.380 75.600 ;
      RECT 39.340 1.400 39.620 75.600 ;
      RECT 41.580 1.400 41.860 75.600 ;
      RECT 43.820 1.400 44.100 75.600 ;
      RECT 46.060 1.400 46.340 75.600 ;
      RECT 48.300 1.400 48.580 75.600 ;
      RECT 50.540 1.400 50.820 75.600 ;
      RECT 52.780 1.400 53.060 75.600 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 75.600 ;
      RECT 4.620 1.400 4.900 75.600 ;
      RECT 6.860 1.400 7.140 75.600 ;
      RECT 9.100 1.400 9.380 75.600 ;
      RECT 11.340 1.400 11.620 75.600 ;
      RECT 13.580 1.400 13.860 75.600 ;
      RECT 15.820 1.400 16.100 75.600 ;
      RECT 18.060 1.400 18.340 75.600 ;
      RECT 20.300 1.400 20.580 75.600 ;
      RECT 22.540 1.400 22.820 75.600 ;
      RECT 24.780 1.400 25.060 75.600 ;
      RECT 27.020 1.400 27.300 75.600 ;
      RECT 29.260 1.400 29.540 75.600 ;
      RECT 31.500 1.400 31.780 75.600 ;
      RECT 33.740 1.400 34.020 75.600 ;
      RECT 35.980 1.400 36.260 75.600 ;
      RECT 38.220 1.400 38.500 75.600 ;
      RECT 40.460 1.400 40.740 75.600 ;
      RECT 42.700 1.400 42.980 75.600 ;
      RECT 44.940 1.400 45.220 75.600 ;
      RECT 47.180 1.400 47.460 75.600 ;
      RECT 49.420 1.400 49.700 75.600 ;
      RECT 51.660 1.400 51.940 75.600 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 54.530 77.000 ;
    LAYER metal2 ;
    RECT 0 0 54.530 77.000 ;
    LAYER metal3 ;
    RECT 0.070 0 54.530 77.000 ;
    RECT 0 0.000 0.070 1.400 ;
    RECT 0 1.470 0.070 1.540 ;
    RECT 0 1.610 0.070 1.680 ;
    RECT 0 1.750 0.070 1.820 ;
    RECT 0 1.890 0.070 1.960 ;
    RECT 0 2.030 0.070 2.100 ;
    RECT 0 2.170 0.070 2.240 ;
    RECT 0 2.310 0.070 2.380 ;
    RECT 0 2.450 0.070 2.520 ;
    RECT 0 2.590 0.070 2.660 ;
    RECT 0 2.730 0.070 2.800 ;
    RECT 0 2.870 0.070 2.940 ;
    RECT 0 3.010 0.070 3.080 ;
    RECT 0 3.150 0.070 3.220 ;
    RECT 0 3.290 0.070 3.360 ;
    RECT 0 3.430 0.070 3.500 ;
    RECT 0 3.570 0.070 3.640 ;
    RECT 0 3.710 0.070 3.780 ;
    RECT 0 3.850 0.070 3.920 ;
    RECT 0 3.990 0.070 4.060 ;
    RECT 0 4.130 0.070 4.200 ;
    RECT 0 4.270 0.070 4.340 ;
    RECT 0 4.410 0.070 4.480 ;
    RECT 0 4.550 0.070 4.620 ;
    RECT 0 4.690 0.070 4.760 ;
    RECT 0 4.830 0.070 4.900 ;
    RECT 0 4.970 0.070 5.040 ;
    RECT 0 5.110 0.070 5.180 ;
    RECT 0 5.250 0.070 5.320 ;
    RECT 0 5.390 0.070 5.460 ;
    RECT 0 5.530 0.070 5.600 ;
    RECT 0 5.670 0.070 5.740 ;
    RECT 0 5.810 0.070 5.880 ;
    RECT 0 5.950 0.070 6.020 ;
    RECT 0 6.090 0.070 6.160 ;
    RECT 0 6.230 0.070 6.300 ;
    RECT 0 6.370 0.070 6.440 ;
    RECT 0 6.510 0.070 6.580 ;
    RECT 0 6.650 0.070 6.720 ;
    RECT 0 6.790 0.070 6.860 ;
    RECT 0 6.930 0.070 7.000 ;
    RECT 0 7.070 0.070 7.140 ;
    RECT 0 7.210 0.070 7.280 ;
    RECT 0 7.350 0.070 7.420 ;
    RECT 0 7.490 0.070 7.560 ;
    RECT 0 7.630 0.070 7.700 ;
    RECT 0 7.770 0.070 7.840 ;
    RECT 0 7.910 0.070 7.980 ;
    RECT 0 8.050 0.070 8.120 ;
    RECT 0 8.190 0.070 8.260 ;
    RECT 0 8.330 0.070 8.400 ;
    RECT 0 8.470 0.070 8.540 ;
    RECT 0 8.610 0.070 8.680 ;
    RECT 0 8.750 0.070 8.820 ;
    RECT 0 8.890 0.070 8.960 ;
    RECT 0 9.030 0.070 9.100 ;
    RECT 0 9.170 0.070 9.240 ;
    RECT 0 9.310 0.070 9.380 ;
    RECT 0 9.450 0.070 9.520 ;
    RECT 0 9.590 0.070 9.660 ;
    RECT 0 9.730 0.070 9.800 ;
    RECT 0 9.870 0.070 9.940 ;
    RECT 0 10.010 0.070 10.080 ;
    RECT 0 10.150 0.070 10.220 ;
    RECT 0 10.290 0.070 10.360 ;
    RECT 0 10.430 0.070 10.500 ;
    RECT 0 10.570 0.070 10.640 ;
    RECT 0 10.710 0.070 10.780 ;
    RECT 0 10.850 0.070 10.920 ;
    RECT 0 10.990 0.070 11.060 ;
    RECT 0 11.130 0.070 11.200 ;
    RECT 0 11.270 0.070 11.340 ;
    RECT 0 11.410 0.070 11.480 ;
    RECT 0 11.550 0.070 11.620 ;
    RECT 0 11.690 0.070 11.760 ;
    RECT 0 11.830 0.070 11.900 ;
    RECT 0 11.970 0.070 12.040 ;
    RECT 0 12.110 0.070 12.180 ;
    RECT 0 12.250 0.070 12.320 ;
    RECT 0 12.390 0.070 12.460 ;
    RECT 0 12.530 0.070 12.600 ;
    RECT 0 12.670 0.070 12.740 ;
    RECT 0 12.810 0.070 12.880 ;
    RECT 0 12.950 0.070 13.020 ;
    RECT 0 13.090 0.070 13.160 ;
    RECT 0 13.230 0.070 13.300 ;
    RECT 0 13.370 0.070 13.440 ;
    RECT 0 13.510 0.070 13.580 ;
    RECT 0 13.650 0.070 13.720 ;
    RECT 0 13.790 0.070 13.860 ;
    RECT 0 13.930 0.070 14.000 ;
    RECT 0 14.070 0.070 14.140 ;
    RECT 0 14.210 0.070 14.280 ;
    RECT 0 14.350 0.070 14.420 ;
    RECT 0 14.490 0.070 14.560 ;
    RECT 0 14.630 0.070 14.700 ;
    RECT 0 14.770 0.070 22.820 ;
    RECT 0 22.890 0.070 22.960 ;
    RECT 0 23.030 0.070 23.100 ;
    RECT 0 23.170 0.070 23.240 ;
    RECT 0 23.310 0.070 23.380 ;
    RECT 0 23.450 0.070 23.520 ;
    RECT 0 23.590 0.070 23.660 ;
    RECT 0 23.730 0.070 23.800 ;
    RECT 0 23.870 0.070 23.940 ;
    RECT 0 24.010 0.070 24.080 ;
    RECT 0 24.150 0.070 24.220 ;
    RECT 0 24.290 0.070 24.360 ;
    RECT 0 24.430 0.070 24.500 ;
    RECT 0 24.570 0.070 24.640 ;
    RECT 0 24.710 0.070 24.780 ;
    RECT 0 24.850 0.070 24.920 ;
    RECT 0 24.990 0.070 25.060 ;
    RECT 0 25.130 0.070 25.200 ;
    RECT 0 25.270 0.070 25.340 ;
    RECT 0 25.410 0.070 25.480 ;
    RECT 0 25.550 0.070 25.620 ;
    RECT 0 25.690 0.070 25.760 ;
    RECT 0 25.830 0.070 25.900 ;
    RECT 0 25.970 0.070 26.040 ;
    RECT 0 26.110 0.070 26.180 ;
    RECT 0 26.250 0.070 26.320 ;
    RECT 0 26.390 0.070 26.460 ;
    RECT 0 26.530 0.070 26.600 ;
    RECT 0 26.670 0.070 26.740 ;
    RECT 0 26.810 0.070 26.880 ;
    RECT 0 26.950 0.070 27.020 ;
    RECT 0 27.090 0.070 27.160 ;
    RECT 0 27.230 0.070 27.300 ;
    RECT 0 27.370 0.070 27.440 ;
    RECT 0 27.510 0.070 27.580 ;
    RECT 0 27.650 0.070 27.720 ;
    RECT 0 27.790 0.070 27.860 ;
    RECT 0 27.930 0.070 28.000 ;
    RECT 0 28.070 0.070 28.140 ;
    RECT 0 28.210 0.070 28.280 ;
    RECT 0 28.350 0.070 28.420 ;
    RECT 0 28.490 0.070 28.560 ;
    RECT 0 28.630 0.070 28.700 ;
    RECT 0 28.770 0.070 28.840 ;
    RECT 0 28.910 0.070 28.980 ;
    RECT 0 29.050 0.070 29.120 ;
    RECT 0 29.190 0.070 29.260 ;
    RECT 0 29.330 0.070 29.400 ;
    RECT 0 29.470 0.070 29.540 ;
    RECT 0 29.610 0.070 29.680 ;
    RECT 0 29.750 0.070 29.820 ;
    RECT 0 29.890 0.070 29.960 ;
    RECT 0 30.030 0.070 30.100 ;
    RECT 0 30.170 0.070 30.240 ;
    RECT 0 30.310 0.070 30.380 ;
    RECT 0 30.450 0.070 30.520 ;
    RECT 0 30.590 0.070 30.660 ;
    RECT 0 30.730 0.070 30.800 ;
    RECT 0 30.870 0.070 30.940 ;
    RECT 0 31.010 0.070 31.080 ;
    RECT 0 31.150 0.070 31.220 ;
    RECT 0 31.290 0.070 31.360 ;
    RECT 0 31.430 0.070 31.500 ;
    RECT 0 31.570 0.070 31.640 ;
    RECT 0 31.710 0.070 31.780 ;
    RECT 0 31.850 0.070 31.920 ;
    RECT 0 31.990 0.070 32.060 ;
    RECT 0 32.130 0.070 32.200 ;
    RECT 0 32.270 0.070 32.340 ;
    RECT 0 32.410 0.070 32.480 ;
    RECT 0 32.550 0.070 32.620 ;
    RECT 0 32.690 0.070 32.760 ;
    RECT 0 32.830 0.070 32.900 ;
    RECT 0 32.970 0.070 33.040 ;
    RECT 0 33.110 0.070 33.180 ;
    RECT 0 33.250 0.070 33.320 ;
    RECT 0 33.390 0.070 33.460 ;
    RECT 0 33.530 0.070 33.600 ;
    RECT 0 33.670 0.070 33.740 ;
    RECT 0 33.810 0.070 33.880 ;
    RECT 0 33.950 0.070 34.020 ;
    RECT 0 34.090 0.070 34.160 ;
    RECT 0 34.230 0.070 34.300 ;
    RECT 0 34.370 0.070 34.440 ;
    RECT 0 34.510 0.070 34.580 ;
    RECT 0 34.650 0.070 34.720 ;
    RECT 0 34.790 0.070 34.860 ;
    RECT 0 34.930 0.070 35.000 ;
    RECT 0 35.070 0.070 35.140 ;
    RECT 0 35.210 0.070 35.280 ;
    RECT 0 35.350 0.070 35.420 ;
    RECT 0 35.490 0.070 35.560 ;
    RECT 0 35.630 0.070 35.700 ;
    RECT 0 35.770 0.070 35.840 ;
    RECT 0 35.910 0.070 35.980 ;
    RECT 0 36.050 0.070 36.120 ;
    RECT 0 36.190 0.070 44.240 ;
    RECT 0 44.310 0.070 44.380 ;
    RECT 0 44.450 0.070 44.520 ;
    RECT 0 44.590 0.070 44.660 ;
    RECT 0 44.730 0.070 44.800 ;
    RECT 0 44.870 0.070 44.940 ;
    RECT 0 45.010 0.070 45.080 ;
    RECT 0 45.150 0.070 45.220 ;
    RECT 0 45.290 0.070 45.360 ;
    RECT 0 45.430 0.070 45.500 ;
    RECT 0 45.570 0.070 45.640 ;
    RECT 0 45.710 0.070 45.780 ;
    RECT 0 45.850 0.070 45.920 ;
    RECT 0 45.990 0.070 46.060 ;
    RECT 0 46.130 0.070 46.200 ;
    RECT 0 46.270 0.070 46.340 ;
    RECT 0 46.410 0.070 46.480 ;
    RECT 0 46.550 0.070 46.620 ;
    RECT 0 46.690 0.070 46.760 ;
    RECT 0 46.830 0.070 46.900 ;
    RECT 0 46.970 0.070 47.040 ;
    RECT 0 47.110 0.070 47.180 ;
    RECT 0 47.250 0.070 47.320 ;
    RECT 0 47.390 0.070 47.460 ;
    RECT 0 47.530 0.070 47.600 ;
    RECT 0 47.670 0.070 47.740 ;
    RECT 0 47.810 0.070 47.880 ;
    RECT 0 47.950 0.070 48.020 ;
    RECT 0 48.090 0.070 48.160 ;
    RECT 0 48.230 0.070 48.300 ;
    RECT 0 48.370 0.070 48.440 ;
    RECT 0 48.510 0.070 48.580 ;
    RECT 0 48.650 0.070 48.720 ;
    RECT 0 48.790 0.070 48.860 ;
    RECT 0 48.930 0.070 49.000 ;
    RECT 0 49.070 0.070 49.140 ;
    RECT 0 49.210 0.070 49.280 ;
    RECT 0 49.350 0.070 49.420 ;
    RECT 0 49.490 0.070 49.560 ;
    RECT 0 49.630 0.070 49.700 ;
    RECT 0 49.770 0.070 49.840 ;
    RECT 0 49.910 0.070 49.980 ;
    RECT 0 50.050 0.070 50.120 ;
    RECT 0 50.190 0.070 50.260 ;
    RECT 0 50.330 0.070 50.400 ;
    RECT 0 50.470 0.070 50.540 ;
    RECT 0 50.610 0.070 50.680 ;
    RECT 0 50.750 0.070 50.820 ;
    RECT 0 50.890 0.070 50.960 ;
    RECT 0 51.030 0.070 51.100 ;
    RECT 0 51.170 0.070 51.240 ;
    RECT 0 51.310 0.070 51.380 ;
    RECT 0 51.450 0.070 51.520 ;
    RECT 0 51.590 0.070 51.660 ;
    RECT 0 51.730 0.070 51.800 ;
    RECT 0 51.870 0.070 51.940 ;
    RECT 0 52.010 0.070 52.080 ;
    RECT 0 52.150 0.070 52.220 ;
    RECT 0 52.290 0.070 52.360 ;
    RECT 0 52.430 0.070 52.500 ;
    RECT 0 52.570 0.070 52.640 ;
    RECT 0 52.710 0.070 52.780 ;
    RECT 0 52.850 0.070 52.920 ;
    RECT 0 52.990 0.070 53.060 ;
    RECT 0 53.130 0.070 53.200 ;
    RECT 0 53.270 0.070 53.340 ;
    RECT 0 53.410 0.070 53.480 ;
    RECT 0 53.550 0.070 53.620 ;
    RECT 0 53.690 0.070 53.760 ;
    RECT 0 53.830 0.070 53.900 ;
    RECT 0 53.970 0.070 54.040 ;
    RECT 0 54.110 0.070 54.180 ;
    RECT 0 54.250 0.070 54.320 ;
    RECT 0 54.390 0.070 54.460 ;
    RECT 0 54.530 0.070 54.600 ;
    RECT 0 54.670 0.070 54.740 ;
    RECT 0 54.810 0.070 54.880 ;
    RECT 0 54.950 0.070 55.020 ;
    RECT 0 55.090 0.070 55.160 ;
    RECT 0 55.230 0.070 55.300 ;
    RECT 0 55.370 0.070 55.440 ;
    RECT 0 55.510 0.070 55.580 ;
    RECT 0 55.650 0.070 55.720 ;
    RECT 0 55.790 0.070 55.860 ;
    RECT 0 55.930 0.070 56.000 ;
    RECT 0 56.070 0.070 56.140 ;
    RECT 0 56.210 0.070 56.280 ;
    RECT 0 56.350 0.070 56.420 ;
    RECT 0 56.490 0.070 56.560 ;
    RECT 0 56.630 0.070 56.700 ;
    RECT 0 56.770 0.070 56.840 ;
    RECT 0 56.910 0.070 56.980 ;
    RECT 0 57.050 0.070 57.120 ;
    RECT 0 57.190 0.070 57.260 ;
    RECT 0 57.330 0.070 57.400 ;
    RECT 0 57.470 0.070 57.540 ;
    RECT 0 57.610 0.070 65.660 ;
    RECT 0 65.730 0.070 65.800 ;
    RECT 0 65.870 0.070 65.940 ;
    RECT 0 66.010 0.070 66.080 ;
    RECT 0 66.150 0.070 66.220 ;
    RECT 0 66.290 0.070 66.360 ;
    RECT 0 66.430 0.070 74.480 ;
    RECT 0 74.550 0.070 74.620 ;
    RECT 0 74.690 0.070 74.760 ;
    RECT 0 74.830 0.070 77.000 ;
    LAYER metal4 ;
    RECT 0 0 54.530 1.400 ;
    RECT 0 75.600 54.530 77.000 ;
    RECT 0.000 1.400 1.260 75.600 ;
    RECT 1.540 1.400 2.380 75.600 ;
    RECT 2.660 1.400 3.500 75.600 ;
    RECT 3.780 1.400 4.620 75.600 ;
    RECT 4.900 1.400 5.740 75.600 ;
    RECT 6.020 1.400 6.860 75.600 ;
    RECT 7.140 1.400 7.980 75.600 ;
    RECT 8.260 1.400 9.100 75.600 ;
    RECT 9.380 1.400 10.220 75.600 ;
    RECT 10.500 1.400 11.340 75.600 ;
    RECT 11.620 1.400 12.460 75.600 ;
    RECT 12.740 1.400 13.580 75.600 ;
    RECT 13.860 1.400 14.700 75.600 ;
    RECT 14.980 1.400 15.820 75.600 ;
    RECT 16.100 1.400 16.940 75.600 ;
    RECT 17.220 1.400 18.060 75.600 ;
    RECT 18.340 1.400 19.180 75.600 ;
    RECT 19.460 1.400 20.300 75.600 ;
    RECT 20.580 1.400 21.420 75.600 ;
    RECT 21.700 1.400 22.540 75.600 ;
    RECT 22.820 1.400 23.660 75.600 ;
    RECT 23.940 1.400 24.780 75.600 ;
    RECT 25.060 1.400 25.900 75.600 ;
    RECT 26.180 1.400 27.020 75.600 ;
    RECT 27.300 1.400 28.140 75.600 ;
    RECT 28.420 1.400 29.260 75.600 ;
    RECT 29.540 1.400 30.380 75.600 ;
    RECT 30.660 1.400 31.500 75.600 ;
    RECT 31.780 1.400 32.620 75.600 ;
    RECT 32.900 1.400 33.740 75.600 ;
    RECT 34.020 1.400 34.860 75.600 ;
    RECT 35.140 1.400 35.980 75.600 ;
    RECT 36.260 1.400 37.100 75.600 ;
    RECT 37.380 1.400 38.220 75.600 ;
    RECT 38.500 1.400 39.340 75.600 ;
    RECT 39.620 1.400 40.460 75.600 ;
    RECT 40.740 1.400 41.580 75.600 ;
    RECT 41.860 1.400 42.700 75.600 ;
    RECT 42.980 1.400 43.820 75.600 ;
    RECT 44.100 1.400 44.940 75.600 ;
    RECT 45.220 1.400 46.060 75.600 ;
    RECT 46.340 1.400 47.180 75.600 ;
    RECT 47.460 1.400 48.300 75.600 ;
    RECT 48.580 1.400 49.420 75.600 ;
    RECT 49.700 1.400 50.540 75.600 ;
    RECT 50.820 1.400 51.660 75.600 ;
    RECT 51.940 1.400 52.780 75.600 ;
    RECT 53.060 1.400 54.530 75.600 ;
    LAYER OVERLAP ;
    RECT 0 0 54.530 77.000 ;
  END
END fakeram45_64x96

END LIBRARY
