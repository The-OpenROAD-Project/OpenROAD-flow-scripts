module MuxTest_width_16_inputs_8_outputs_8_pipeline_5( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [2:0]  io_selects_0_0, // @[:@6.4]
  input  [2:0]  io_selects_0_1, // @[:@6.4]
  input  [2:0]  io_selects_1_0, // @[:@6.4]
  input  [2:0]  io_selects_1_1, // @[:@6.4]
  input  [2:0]  io_selects_2_0, // @[:@6.4]
  input  [2:0]  io_selects_2_1, // @[:@6.4]
  input  [2:0]  io_selects_3_0, // @[:@6.4]
  input  [2:0]  io_selects_3_1, // @[:@6.4]
  input  [2:0]  io_selects_4_0, // @[:@6.4]
  input  [2:0]  io_selects_4_1, // @[:@6.4]
  input  [2:0]  io_selects_5_0, // @[:@6.4]
  input  [2:0]  io_selects_5_1, // @[:@6.4]
  input  [2:0]  io_selects_6_0, // @[:@6.4]
  input  [2:0]  io_selects_6_1, // @[:@6.4]
  input  [2:0]  io_selects_7_0, // @[:@6.4]
  input  [2:0]  io_selects_7_1, // @[:@6.4]
  input  [2:0]  io_operation_0, // @[:@6.4]
  input  [2:0]  io_operation_1, // @[:@6.4]
  input  [2:0]  io_operation_2, // @[:@6.4]
  input  [2:0]  io_operation_3, // @[:@6.4]
  input  [2:0]  io_operation_4, // @[:@6.4]
  input  [2:0]  io_operation_5, // @[:@6.4]
  input  [2:0]  io_operation_6, // @[:@6.4]
  input  [2:0]  io_operation_7, // @[:@6.4]
  input  [15:0] io_inputs_0, // @[:@6.4]
  input  [15:0] io_inputs_1, // @[:@6.4]
  input  [15:0] io_inputs_2, // @[:@6.4]
  input  [15:0] io_inputs_3, // @[:@6.4]
  input  [15:0] io_inputs_4, // @[:@6.4]
  input  [15:0] io_inputs_5, // @[:@6.4]
  input  [15:0] io_inputs_6, // @[:@6.4]
  input  [15:0] io_inputs_7, // @[:@6.4]
  output [15:0] io_outputs_0, // @[:@6.4]
  output [15:0] io_outputs_1, // @[:@6.4]
  output [15:0] io_outputs_2, // @[:@6.4]
  output [15:0] io_outputs_3, // @[:@6.4]
  output [15:0] io_outputs_4, // @[:@6.4]
  output [15:0] io_outputs_5, // @[:@6.4]
  output [15:0] io_outputs_6, // @[:@6.4]
  output [15:0] io_outputs_7 // @[:@6.4]
);
  wire [15:0] _GEN_1; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  wire [15:0] _GEN_2; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  wire [15:0] _GEN_3; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  wire [15:0] _GEN_4; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  wire [15:0] _GEN_5; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  wire [15:0] _GEN_6; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  wire [15:0] _GEN_7; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  wire [15:0] _GEN_9; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  wire [15:0] _GEN_10; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  wire [15:0] _GEN_11; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  wire [15:0] _GEN_12; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  wire [15:0] _GEN_13; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  wire [15:0] _GEN_14; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  wire [15:0] _GEN_15; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  wire [16:0] _T_402; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  wire [15:0] _T_403; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@9.4]
  wire [31:0] _T_405; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 33:58:@10.4]
  wire [15:0] _T_407; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 34:56:@11.4]
  wire  _T_408; // @[Mux.scala 46:19:@12.4]
  wire [15:0] _T_409; // @[Mux.scala 46:16:@13.4]
  wire  _T_410; // @[Mux.scala 46:19:@14.4]
  wire [31:0] _T_411; // @[Mux.scala 46:16:@15.4]
  wire  _T_412; // @[Mux.scala 46:19:@16.4]
  wire [31:0] _T_413; // @[Mux.scala 46:16:@17.4]
  wire  _T_414; // @[Mux.scala 46:19:@18.4]
  wire [15:0] _GEN_17; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  wire [15:0] _GEN_18; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  wire [15:0] _GEN_19; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  wire [15:0] _GEN_20; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  wire [15:0] _GEN_21; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  wire [15:0] _GEN_22; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  wire [15:0] _GEN_23; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  wire [15:0] _GEN_25; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  wire [15:0] _GEN_26; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  wire [15:0] _GEN_27; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  wire [15:0] _GEN_28; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  wire [15:0] _GEN_29; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  wire [15:0] _GEN_30; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  wire [15:0] _GEN_31; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  wire [16:0] _T_419; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  wire [15:0] _T_420; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@21.4]
  wire [31:0] _T_422; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 33:58:@22.4]
  wire [15:0] _T_424; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 34:56:@23.4]
  wire  _T_425; // @[Mux.scala 46:19:@24.4]
  wire [15:0] _T_426; // @[Mux.scala 46:16:@25.4]
  wire  _T_427; // @[Mux.scala 46:19:@26.4]
  wire [31:0] _T_428; // @[Mux.scala 46:16:@27.4]
  wire  _T_429; // @[Mux.scala 46:19:@28.4]
  wire [31:0] _T_430; // @[Mux.scala 46:16:@29.4]
  wire  _T_431; // @[Mux.scala 46:19:@30.4]
  wire [15:0] _GEN_33; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  wire [15:0] _GEN_34; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  wire [15:0] _GEN_35; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  wire [15:0] _GEN_36; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  wire [15:0] _GEN_37; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  wire [15:0] _GEN_38; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  wire [15:0] _GEN_39; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  wire [15:0] _GEN_41; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  wire [15:0] _GEN_42; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  wire [15:0] _GEN_43; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  wire [15:0] _GEN_44; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  wire [15:0] _GEN_45; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  wire [15:0] _GEN_46; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  wire [15:0] _GEN_47; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  wire [16:0] _T_436; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  wire [15:0] _T_437; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@33.4]
  wire [31:0] _T_439; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 33:58:@34.4]
  wire [15:0] _T_441; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 34:56:@35.4]
  wire  _T_442; // @[Mux.scala 46:19:@36.4]
  wire [15:0] _T_443; // @[Mux.scala 46:16:@37.4]
  wire  _T_444; // @[Mux.scala 46:19:@38.4]
  wire [31:0] _T_445; // @[Mux.scala 46:16:@39.4]
  wire  _T_446; // @[Mux.scala 46:19:@40.4]
  wire [31:0] _T_447; // @[Mux.scala 46:16:@41.4]
  wire  _T_448; // @[Mux.scala 46:19:@42.4]
  wire [15:0] _GEN_49; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  wire [15:0] _GEN_50; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  wire [15:0] _GEN_51; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  wire [15:0] _GEN_52; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  wire [15:0] _GEN_53; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  wire [15:0] _GEN_54; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  wire [15:0] _GEN_55; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  wire [15:0] _GEN_57; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  wire [15:0] _GEN_58; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  wire [15:0] _GEN_59; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  wire [15:0] _GEN_60; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  wire [15:0] _GEN_61; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  wire [15:0] _GEN_62; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  wire [15:0] _GEN_63; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  wire [16:0] _T_453; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  wire [15:0] _T_454; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@45.4]
  wire [31:0] _T_456; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 33:58:@46.4]
  wire [15:0] _T_458; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 34:56:@47.4]
  wire  _T_459; // @[Mux.scala 46:19:@48.4]
  wire [15:0] _T_460; // @[Mux.scala 46:16:@49.4]
  wire  _T_461; // @[Mux.scala 46:19:@50.4]
  wire [31:0] _T_462; // @[Mux.scala 46:16:@51.4]
  wire  _T_463; // @[Mux.scala 46:19:@52.4]
  wire [31:0] _T_464; // @[Mux.scala 46:16:@53.4]
  wire  _T_465; // @[Mux.scala 46:19:@54.4]
  wire [15:0] _GEN_65; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  wire [15:0] _GEN_66; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  wire [15:0] _GEN_67; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  wire [15:0] _GEN_68; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  wire [15:0] _GEN_69; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  wire [15:0] _GEN_70; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  wire [15:0] _GEN_71; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  wire [15:0] _GEN_73; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  wire [15:0] _GEN_74; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  wire [15:0] _GEN_75; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  wire [15:0] _GEN_76; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  wire [15:0] _GEN_77; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  wire [15:0] _GEN_78; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  wire [15:0] _GEN_79; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  wire [16:0] _T_470; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  wire [15:0] _T_471; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@57.4]
  wire [31:0] _T_473; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 33:58:@58.4]
  wire [15:0] _T_475; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 34:56:@59.4]
  wire  _T_476; // @[Mux.scala 46:19:@60.4]
  wire [15:0] _T_477; // @[Mux.scala 46:16:@61.4]
  wire  _T_478; // @[Mux.scala 46:19:@62.4]
  wire [31:0] _T_479; // @[Mux.scala 46:16:@63.4]
  wire  _T_480; // @[Mux.scala 46:19:@64.4]
  wire [31:0] _T_481; // @[Mux.scala 46:16:@65.4]
  wire  _T_482; // @[Mux.scala 46:19:@66.4]
  wire [15:0] _GEN_81; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  wire [15:0] _GEN_82; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  wire [15:0] _GEN_83; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  wire [15:0] _GEN_84; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  wire [15:0] _GEN_85; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  wire [15:0] _GEN_86; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  wire [15:0] _GEN_87; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  wire [15:0] _GEN_89; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  wire [15:0] _GEN_90; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  wire [15:0] _GEN_91; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  wire [15:0] _GEN_92; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  wire [15:0] _GEN_93; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  wire [15:0] _GEN_94; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  wire [15:0] _GEN_95; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  wire [16:0] _T_487; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  wire [15:0] _T_488; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@69.4]
  wire [31:0] _T_490; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 33:58:@70.4]
  wire [15:0] _T_492; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 34:56:@71.4]
  wire  _T_493; // @[Mux.scala 46:19:@72.4]
  wire [15:0] _T_494; // @[Mux.scala 46:16:@73.4]
  wire  _T_495; // @[Mux.scala 46:19:@74.4]
  wire [31:0] _T_496; // @[Mux.scala 46:16:@75.4]
  wire  _T_497; // @[Mux.scala 46:19:@76.4]
  wire [31:0] _T_498; // @[Mux.scala 46:16:@77.4]
  wire  _T_499; // @[Mux.scala 46:19:@78.4]
  wire [15:0] _GEN_97; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  wire [15:0] _GEN_98; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  wire [15:0] _GEN_99; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  wire [15:0] _GEN_100; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  wire [15:0] _GEN_101; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  wire [15:0] _GEN_102; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  wire [15:0] _GEN_103; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  wire [15:0] _GEN_105; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  wire [15:0] _GEN_106; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  wire [15:0] _GEN_107; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  wire [15:0] _GEN_108; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  wire [15:0] _GEN_109; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  wire [15:0] _GEN_110; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  wire [15:0] _GEN_111; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  wire [16:0] _T_504; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  wire [15:0] _T_505; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@81.4]
  wire [31:0] _T_507; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 33:58:@82.4]
  wire [15:0] _T_509; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 34:56:@83.4]
  wire  _T_510; // @[Mux.scala 46:19:@84.4]
  wire [15:0] _T_511; // @[Mux.scala 46:16:@85.4]
  wire  _T_512; // @[Mux.scala 46:19:@86.4]
  wire [31:0] _T_513; // @[Mux.scala 46:16:@87.4]
  wire  _T_514; // @[Mux.scala 46:19:@88.4]
  wire [31:0] _T_515; // @[Mux.scala 46:16:@89.4]
  wire  _T_516; // @[Mux.scala 46:19:@90.4]
  wire [15:0] _GEN_113; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  wire [15:0] _GEN_114; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  wire [15:0] _GEN_115; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  wire [15:0] _GEN_116; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  wire [15:0] _GEN_117; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  wire [15:0] _GEN_118; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  wire [15:0] _GEN_119; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  wire [15:0] _GEN_121; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  wire [15:0] _GEN_122; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  wire [15:0] _GEN_123; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  wire [15:0] _GEN_124; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  wire [15:0] _GEN_125; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  wire [15:0] _GEN_126; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  wire [15:0] _GEN_127; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  wire [16:0] _T_521; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  wire [15:0] _T_522; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@93.4]
  wire [31:0] _T_524; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 33:58:@94.4]
  wire [15:0] _T_526; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 34:56:@95.4]
  wire  _T_527; // @[Mux.scala 46:19:@96.4]
  wire [15:0] _T_528; // @[Mux.scala 46:16:@97.4]
  wire  _T_529; // @[Mux.scala 46:19:@98.4]
  wire [31:0] _T_530; // @[Mux.scala 46:16:@99.4]
  wire  _T_531; // @[Mux.scala 46:19:@100.4]
  wire [31:0] _T_532; // @[Mux.scala 46:16:@101.4]
  wire  _T_533; // @[Mux.scala 46:19:@102.4]
  reg [31:0] _T_537; // @[Reg.scala 11:16:@104.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_539; // @[Reg.scala 11:16:@108.4]
  reg [31:0] _RAND_1;
  reg [31:0] _T_541; // @[Reg.scala 11:16:@112.4]
  reg [31:0] _RAND_2;
  reg [31:0] _T_543; // @[Reg.scala 11:16:@116.4]
  reg [31:0] _RAND_3;
  reg [31:0] _T_545; // @[Reg.scala 11:16:@120.4]
  reg [31:0] _RAND_4;
  reg [31:0] _T_548; // @[Reg.scala 11:16:@124.4]
  reg [31:0] _RAND_5;
  reg [31:0] _T_550; // @[Reg.scala 11:16:@128.4]
  reg [31:0] _RAND_6;
  reg [31:0] _T_552; // @[Reg.scala 11:16:@132.4]
  reg [31:0] _RAND_7;
  reg [31:0] _T_554; // @[Reg.scala 11:16:@136.4]
  reg [31:0] _RAND_8;
  reg [31:0] _T_556; // @[Reg.scala 11:16:@140.4]
  reg [31:0] _RAND_9;
  reg [31:0] _T_559; // @[Reg.scala 11:16:@144.4]
  reg [31:0] _RAND_10;
  reg [31:0] _T_561; // @[Reg.scala 11:16:@148.4]
  reg [31:0] _RAND_11;
  reg [31:0] _T_563; // @[Reg.scala 11:16:@152.4]
  reg [31:0] _RAND_12;
  reg [31:0] _T_565; // @[Reg.scala 11:16:@156.4]
  reg [31:0] _RAND_13;
  reg [31:0] _T_567; // @[Reg.scala 11:16:@160.4]
  reg [31:0] _RAND_14;
  reg [31:0] _T_570; // @[Reg.scala 11:16:@164.4]
  reg [31:0] _RAND_15;
  reg [31:0] _T_572; // @[Reg.scala 11:16:@168.4]
  reg [31:0] _RAND_16;
  reg [31:0] _T_574; // @[Reg.scala 11:16:@172.4]
  reg [31:0] _RAND_17;
  reg [31:0] _T_576; // @[Reg.scala 11:16:@176.4]
  reg [31:0] _RAND_18;
  reg [31:0] _T_578; // @[Reg.scala 11:16:@180.4]
  reg [31:0] _RAND_19;
  reg [31:0] _T_581; // @[Reg.scala 11:16:@184.4]
  reg [31:0] _RAND_20;
  reg [31:0] _T_583; // @[Reg.scala 11:16:@188.4]
  reg [31:0] _RAND_21;
  reg [31:0] _T_585; // @[Reg.scala 11:16:@192.4]
  reg [31:0] _RAND_22;
  reg [31:0] _T_587; // @[Reg.scala 11:16:@196.4]
  reg [31:0] _RAND_23;
  reg [31:0] _T_589; // @[Reg.scala 11:16:@200.4]
  reg [31:0] _RAND_24;
  reg [31:0] _T_592; // @[Reg.scala 11:16:@204.4]
  reg [31:0] _RAND_25;
  reg [31:0] _T_594; // @[Reg.scala 11:16:@208.4]
  reg [31:0] _RAND_26;
  reg [31:0] _T_596; // @[Reg.scala 11:16:@212.4]
  reg [31:0] _RAND_27;
  reg [31:0] _T_598; // @[Reg.scala 11:16:@216.4]
  reg [31:0] _RAND_28;
  reg [31:0] _T_600; // @[Reg.scala 11:16:@220.4]
  reg [31:0] _RAND_29;
  reg [31:0] _T_603; // @[Reg.scala 11:16:@224.4]
  reg [31:0] _RAND_30;
  reg [31:0] _T_605; // @[Reg.scala 11:16:@228.4]
  reg [31:0] _RAND_31;
  reg [31:0] _T_607; // @[Reg.scala 11:16:@232.4]
  reg [31:0] _RAND_32;
  reg [31:0] _T_609; // @[Reg.scala 11:16:@236.4]
  reg [31:0] _RAND_33;
  reg [31:0] _T_611; // @[Reg.scala 11:16:@240.4]
  reg [31:0] _RAND_34;
  reg [31:0] _T_614; // @[Reg.scala 11:16:@244.4]
  reg [31:0] _RAND_35;
  reg [31:0] _T_616; // @[Reg.scala 11:16:@248.4]
  reg [31:0] _RAND_36;
  reg [31:0] _T_618; // @[Reg.scala 11:16:@252.4]
  reg [31:0] _RAND_37;
  reg [31:0] _T_620; // @[Reg.scala 11:16:@256.4]
  reg [31:0] _RAND_38;
  reg [31:0] _T_622; // @[Reg.scala 11:16:@260.4]
  reg [31:0] _RAND_39;
  assign _GEN_1 = 3'h1 == io_selects_0_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_2 = 3'h2 == io_selects_0_0 ? io_inputs_2 : _GEN_1; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_3 = 3'h3 == io_selects_0_0 ? io_inputs_3 : _GEN_2; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_4 = 3'h4 == io_selects_0_0 ? io_inputs_4 : _GEN_3; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_5 = 3'h5 == io_selects_0_0 ? io_inputs_5 : _GEN_4; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_6 = 3'h6 == io_selects_0_0 ? io_inputs_6 : _GEN_5; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_7 = 3'h7 == io_selects_0_0 ? io_inputs_7 : _GEN_6; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_9 = 3'h1 == io_selects_0_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_10 = 3'h2 == io_selects_0_1 ? io_inputs_2 : _GEN_9; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_11 = 3'h3 == io_selects_0_1 ? io_inputs_3 : _GEN_10; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_12 = 3'h4 == io_selects_0_1 ? io_inputs_4 : _GEN_11; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_13 = 3'h5 == io_selects_0_1 ? io_inputs_5 : _GEN_12; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_14 = 3'h6 == io_selects_0_1 ? io_inputs_6 : _GEN_13; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_15 = 3'h7 == io_selects_0_1 ? io_inputs_7 : _GEN_14; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  assign _T_402 = _GEN_7 + _GEN_15; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@8.4]
  assign _T_403 = _GEN_7 + _GEN_15; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@9.4]
  assign _T_405 = _GEN_7 * _GEN_15; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 33:58:@10.4]
  assign _T_407 = _GEN_7 / _GEN_15; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 34:56:@11.4]
  assign _T_408 = 3'h3 == io_operation_0; // @[Mux.scala 46:19:@12.4]
  assign _T_409 = _T_408 ? _T_407 : 16'h0; // @[Mux.scala 46:16:@13.4]
  assign _T_410 = 3'h2 == io_operation_0; // @[Mux.scala 46:19:@14.4]
  assign _T_411 = _T_410 ? _T_405 : {{16'd0}, _T_409}; // @[Mux.scala 46:16:@15.4]
  assign _T_412 = 3'h1 == io_operation_0; // @[Mux.scala 46:19:@16.4]
  assign _T_413 = _T_412 ? {{16'd0}, _T_403} : _T_411; // @[Mux.scala 46:16:@17.4]
  assign _T_414 = 3'h0 == io_operation_0; // @[Mux.scala 46:19:@18.4]
  assign _GEN_17 = 3'h1 == io_selects_1_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_18 = 3'h2 == io_selects_1_0 ? io_inputs_2 : _GEN_17; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_19 = 3'h3 == io_selects_1_0 ? io_inputs_3 : _GEN_18; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_20 = 3'h4 == io_selects_1_0 ? io_inputs_4 : _GEN_19; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_21 = 3'h5 == io_selects_1_0 ? io_inputs_5 : _GEN_20; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_22 = 3'h6 == io_selects_1_0 ? io_inputs_6 : _GEN_21; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_23 = 3'h7 == io_selects_1_0 ? io_inputs_7 : _GEN_22; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_25 = 3'h1 == io_selects_1_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_26 = 3'h2 == io_selects_1_1 ? io_inputs_2 : _GEN_25; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_27 = 3'h3 == io_selects_1_1 ? io_inputs_3 : _GEN_26; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_28 = 3'h4 == io_selects_1_1 ? io_inputs_4 : _GEN_27; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_29 = 3'h5 == io_selects_1_1 ? io_inputs_5 : _GEN_28; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_30 = 3'h6 == io_selects_1_1 ? io_inputs_6 : _GEN_29; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_31 = 3'h7 == io_selects_1_1 ? io_inputs_7 : _GEN_30; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  assign _T_419 = _GEN_23 + _GEN_31; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@20.4]
  assign _T_420 = _GEN_23 + _GEN_31; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@21.4]
  assign _T_422 = _GEN_23 * _GEN_31; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 33:58:@22.4]
  assign _T_424 = _GEN_23 / _GEN_31; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 34:56:@23.4]
  assign _T_425 = 3'h3 == io_operation_1; // @[Mux.scala 46:19:@24.4]
  assign _T_426 = _T_425 ? _T_424 : 16'h0; // @[Mux.scala 46:16:@25.4]
  assign _T_427 = 3'h2 == io_operation_1; // @[Mux.scala 46:19:@26.4]
  assign _T_428 = _T_427 ? _T_422 : {{16'd0}, _T_426}; // @[Mux.scala 46:16:@27.4]
  assign _T_429 = 3'h1 == io_operation_1; // @[Mux.scala 46:19:@28.4]
  assign _T_430 = _T_429 ? {{16'd0}, _T_420} : _T_428; // @[Mux.scala 46:16:@29.4]
  assign _T_431 = 3'h0 == io_operation_1; // @[Mux.scala 46:19:@30.4]
  assign _GEN_33 = 3'h1 == io_selects_2_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_34 = 3'h2 == io_selects_2_0 ? io_inputs_2 : _GEN_33; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_35 = 3'h3 == io_selects_2_0 ? io_inputs_3 : _GEN_34; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_36 = 3'h4 == io_selects_2_0 ? io_inputs_4 : _GEN_35; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_37 = 3'h5 == io_selects_2_0 ? io_inputs_5 : _GEN_36; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_38 = 3'h6 == io_selects_2_0 ? io_inputs_6 : _GEN_37; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_39 = 3'h7 == io_selects_2_0 ? io_inputs_7 : _GEN_38; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_41 = 3'h1 == io_selects_2_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_42 = 3'h2 == io_selects_2_1 ? io_inputs_2 : _GEN_41; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_43 = 3'h3 == io_selects_2_1 ? io_inputs_3 : _GEN_42; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_44 = 3'h4 == io_selects_2_1 ? io_inputs_4 : _GEN_43; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_45 = 3'h5 == io_selects_2_1 ? io_inputs_5 : _GEN_44; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_46 = 3'h6 == io_selects_2_1 ? io_inputs_6 : _GEN_45; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_47 = 3'h7 == io_selects_2_1 ? io_inputs_7 : _GEN_46; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  assign _T_436 = _GEN_39 + _GEN_47; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@32.4]
  assign _T_437 = _GEN_39 + _GEN_47; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@33.4]
  assign _T_439 = _GEN_39 * _GEN_47; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 33:58:@34.4]
  assign _T_441 = _GEN_39 / _GEN_47; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 34:56:@35.4]
  assign _T_442 = 3'h3 == io_operation_2; // @[Mux.scala 46:19:@36.4]
  assign _T_443 = _T_442 ? _T_441 : 16'h0; // @[Mux.scala 46:16:@37.4]
  assign _T_444 = 3'h2 == io_operation_2; // @[Mux.scala 46:19:@38.4]
  assign _T_445 = _T_444 ? _T_439 : {{16'd0}, _T_443}; // @[Mux.scala 46:16:@39.4]
  assign _T_446 = 3'h1 == io_operation_2; // @[Mux.scala 46:19:@40.4]
  assign _T_447 = _T_446 ? {{16'd0}, _T_437} : _T_445; // @[Mux.scala 46:16:@41.4]
  assign _T_448 = 3'h0 == io_operation_2; // @[Mux.scala 46:19:@42.4]
  assign _GEN_49 = 3'h1 == io_selects_3_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_50 = 3'h2 == io_selects_3_0 ? io_inputs_2 : _GEN_49; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_51 = 3'h3 == io_selects_3_0 ? io_inputs_3 : _GEN_50; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_52 = 3'h4 == io_selects_3_0 ? io_inputs_4 : _GEN_51; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_53 = 3'h5 == io_selects_3_0 ? io_inputs_5 : _GEN_52; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_54 = 3'h6 == io_selects_3_0 ? io_inputs_6 : _GEN_53; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_55 = 3'h7 == io_selects_3_0 ? io_inputs_7 : _GEN_54; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_57 = 3'h1 == io_selects_3_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_58 = 3'h2 == io_selects_3_1 ? io_inputs_2 : _GEN_57; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_59 = 3'h3 == io_selects_3_1 ? io_inputs_3 : _GEN_58; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_60 = 3'h4 == io_selects_3_1 ? io_inputs_4 : _GEN_59; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_61 = 3'h5 == io_selects_3_1 ? io_inputs_5 : _GEN_60; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_62 = 3'h6 == io_selects_3_1 ? io_inputs_6 : _GEN_61; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_63 = 3'h7 == io_selects_3_1 ? io_inputs_7 : _GEN_62; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  assign _T_453 = _GEN_55 + _GEN_63; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@44.4]
  assign _T_454 = _GEN_55 + _GEN_63; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@45.4]
  assign _T_456 = _GEN_55 * _GEN_63; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 33:58:@46.4]
  assign _T_458 = _GEN_55 / _GEN_63; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 34:56:@47.4]
  assign _T_459 = 3'h3 == io_operation_3; // @[Mux.scala 46:19:@48.4]
  assign _T_460 = _T_459 ? _T_458 : 16'h0; // @[Mux.scala 46:16:@49.4]
  assign _T_461 = 3'h2 == io_operation_3; // @[Mux.scala 46:19:@50.4]
  assign _T_462 = _T_461 ? _T_456 : {{16'd0}, _T_460}; // @[Mux.scala 46:16:@51.4]
  assign _T_463 = 3'h1 == io_operation_3; // @[Mux.scala 46:19:@52.4]
  assign _T_464 = _T_463 ? {{16'd0}, _T_454} : _T_462; // @[Mux.scala 46:16:@53.4]
  assign _T_465 = 3'h0 == io_operation_3; // @[Mux.scala 46:19:@54.4]
  assign _GEN_65 = 3'h1 == io_selects_4_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_66 = 3'h2 == io_selects_4_0 ? io_inputs_2 : _GEN_65; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_67 = 3'h3 == io_selects_4_0 ? io_inputs_3 : _GEN_66; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_68 = 3'h4 == io_selects_4_0 ? io_inputs_4 : _GEN_67; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_69 = 3'h5 == io_selects_4_0 ? io_inputs_5 : _GEN_68; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_70 = 3'h6 == io_selects_4_0 ? io_inputs_6 : _GEN_69; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_71 = 3'h7 == io_selects_4_0 ? io_inputs_7 : _GEN_70; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_73 = 3'h1 == io_selects_4_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_74 = 3'h2 == io_selects_4_1 ? io_inputs_2 : _GEN_73; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_75 = 3'h3 == io_selects_4_1 ? io_inputs_3 : _GEN_74; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_76 = 3'h4 == io_selects_4_1 ? io_inputs_4 : _GEN_75; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_77 = 3'h5 == io_selects_4_1 ? io_inputs_5 : _GEN_76; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_78 = 3'h6 == io_selects_4_1 ? io_inputs_6 : _GEN_77; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_79 = 3'h7 == io_selects_4_1 ? io_inputs_7 : _GEN_78; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  assign _T_470 = _GEN_71 + _GEN_79; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@56.4]
  assign _T_471 = _GEN_71 + _GEN_79; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@57.4]
  assign _T_473 = _GEN_71 * _GEN_79; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 33:58:@58.4]
  assign _T_475 = _GEN_71 / _GEN_79; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 34:56:@59.4]
  assign _T_476 = 3'h3 == io_operation_4; // @[Mux.scala 46:19:@60.4]
  assign _T_477 = _T_476 ? _T_475 : 16'h0; // @[Mux.scala 46:16:@61.4]
  assign _T_478 = 3'h2 == io_operation_4; // @[Mux.scala 46:19:@62.4]
  assign _T_479 = _T_478 ? _T_473 : {{16'd0}, _T_477}; // @[Mux.scala 46:16:@63.4]
  assign _T_480 = 3'h1 == io_operation_4; // @[Mux.scala 46:19:@64.4]
  assign _T_481 = _T_480 ? {{16'd0}, _T_471} : _T_479; // @[Mux.scala 46:16:@65.4]
  assign _T_482 = 3'h0 == io_operation_4; // @[Mux.scala 46:19:@66.4]
  assign _GEN_81 = 3'h1 == io_selects_5_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_82 = 3'h2 == io_selects_5_0 ? io_inputs_2 : _GEN_81; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_83 = 3'h3 == io_selects_5_0 ? io_inputs_3 : _GEN_82; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_84 = 3'h4 == io_selects_5_0 ? io_inputs_4 : _GEN_83; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_85 = 3'h5 == io_selects_5_0 ? io_inputs_5 : _GEN_84; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_86 = 3'h6 == io_selects_5_0 ? io_inputs_6 : _GEN_85; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_87 = 3'h7 == io_selects_5_0 ? io_inputs_7 : _GEN_86; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_89 = 3'h1 == io_selects_5_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_90 = 3'h2 == io_selects_5_1 ? io_inputs_2 : _GEN_89; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_91 = 3'h3 == io_selects_5_1 ? io_inputs_3 : _GEN_90; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_92 = 3'h4 == io_selects_5_1 ? io_inputs_4 : _GEN_91; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_93 = 3'h5 == io_selects_5_1 ? io_inputs_5 : _GEN_92; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_94 = 3'h6 == io_selects_5_1 ? io_inputs_6 : _GEN_93; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_95 = 3'h7 == io_selects_5_1 ? io_inputs_7 : _GEN_94; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  assign _T_487 = _GEN_87 + _GEN_95; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@68.4]
  assign _T_488 = _GEN_87 + _GEN_95; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@69.4]
  assign _T_490 = _GEN_87 * _GEN_95; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 33:58:@70.4]
  assign _T_492 = _GEN_87 / _GEN_95; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 34:56:@71.4]
  assign _T_493 = 3'h3 == io_operation_5; // @[Mux.scala 46:19:@72.4]
  assign _T_494 = _T_493 ? _T_492 : 16'h0; // @[Mux.scala 46:16:@73.4]
  assign _T_495 = 3'h2 == io_operation_5; // @[Mux.scala 46:19:@74.4]
  assign _T_496 = _T_495 ? _T_490 : {{16'd0}, _T_494}; // @[Mux.scala 46:16:@75.4]
  assign _T_497 = 3'h1 == io_operation_5; // @[Mux.scala 46:19:@76.4]
  assign _T_498 = _T_497 ? {{16'd0}, _T_488} : _T_496; // @[Mux.scala 46:16:@77.4]
  assign _T_499 = 3'h0 == io_operation_5; // @[Mux.scala 46:19:@78.4]
  assign _GEN_97 = 3'h1 == io_selects_6_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_98 = 3'h2 == io_selects_6_0 ? io_inputs_2 : _GEN_97; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_99 = 3'h3 == io_selects_6_0 ? io_inputs_3 : _GEN_98; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_100 = 3'h4 == io_selects_6_0 ? io_inputs_4 : _GEN_99; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_101 = 3'h5 == io_selects_6_0 ? io_inputs_5 : _GEN_100; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_102 = 3'h6 == io_selects_6_0 ? io_inputs_6 : _GEN_101; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_103 = 3'h7 == io_selects_6_0 ? io_inputs_7 : _GEN_102; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_105 = 3'h1 == io_selects_6_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_106 = 3'h2 == io_selects_6_1 ? io_inputs_2 : _GEN_105; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_107 = 3'h3 == io_selects_6_1 ? io_inputs_3 : _GEN_106; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_108 = 3'h4 == io_selects_6_1 ? io_inputs_4 : _GEN_107; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_109 = 3'h5 == io_selects_6_1 ? io_inputs_5 : _GEN_108; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_110 = 3'h6 == io_selects_6_1 ? io_inputs_6 : _GEN_109; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_111 = 3'h7 == io_selects_6_1 ? io_inputs_7 : _GEN_110; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  assign _T_504 = _GEN_103 + _GEN_111; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@80.4]
  assign _T_505 = _GEN_103 + _GEN_111; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@81.4]
  assign _T_507 = _GEN_103 * _GEN_111; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 33:58:@82.4]
  assign _T_509 = _GEN_103 / _GEN_111; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 34:56:@83.4]
  assign _T_510 = 3'h3 == io_operation_6; // @[Mux.scala 46:19:@84.4]
  assign _T_511 = _T_510 ? _T_509 : 16'h0; // @[Mux.scala 46:16:@85.4]
  assign _T_512 = 3'h2 == io_operation_6; // @[Mux.scala 46:19:@86.4]
  assign _T_513 = _T_512 ? _T_507 : {{16'd0}, _T_511}; // @[Mux.scala 46:16:@87.4]
  assign _T_514 = 3'h1 == io_operation_6; // @[Mux.scala 46:19:@88.4]
  assign _T_515 = _T_514 ? {{16'd0}, _T_505} : _T_513; // @[Mux.scala 46:16:@89.4]
  assign _T_516 = 3'h0 == io_operation_6; // @[Mux.scala 46:19:@90.4]
  assign _GEN_113 = 3'h1 == io_selects_7_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_114 = 3'h2 == io_selects_7_0 ? io_inputs_2 : _GEN_113; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_115 = 3'h3 == io_selects_7_0 ? io_inputs_3 : _GEN_114; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_116 = 3'h4 == io_selects_7_0 ? io_inputs_4 : _GEN_115; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_117 = 3'h5 == io_selects_7_0 ? io_inputs_5 : _GEN_116; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_118 = 3'h6 == io_selects_7_0 ? io_inputs_6 : _GEN_117; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_119 = 3'h7 == io_selects_7_0 ? io_inputs_7 : _GEN_118; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_121 = 3'h1 == io_selects_7_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_122 = 3'h2 == io_selects_7_1 ? io_inputs_2 : _GEN_121; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_123 = 3'h3 == io_selects_7_1 ? io_inputs_3 : _GEN_122; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_124 = 3'h4 == io_selects_7_1 ? io_inputs_4 : _GEN_123; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_125 = 3'h5 == io_selects_7_1 ? io_inputs_5 : _GEN_124; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_126 = 3'h6 == io_selects_7_1 ? io_inputs_6 : _GEN_125; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_127 = 3'h7 == io_selects_7_1 ? io_inputs_7 : _GEN_126; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  assign _T_521 = _GEN_119 + _GEN_127; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@92.4]
  assign _T_522 = _GEN_119 + _GEN_127; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 32:53:@93.4]
  assign _T_524 = _GEN_119 * _GEN_127; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 33:58:@94.4]
  assign _T_526 = _GEN_119 / _GEN_127; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 34:56:@95.4]
  assign _T_527 = 3'h3 == io_operation_7; // @[Mux.scala 46:19:@96.4]
  assign _T_528 = _T_527 ? _T_526 : 16'h0; // @[Mux.scala 46:16:@97.4]
  assign _T_529 = 3'h2 == io_operation_7; // @[Mux.scala 46:19:@98.4]
  assign _T_530 = _T_529 ? _T_524 : {{16'd0}, _T_528}; // @[Mux.scala 46:16:@99.4]
  assign _T_531 = 3'h1 == io_operation_7; // @[Mux.scala 46:19:@100.4]
  assign _T_532 = _T_531 ? {{16'd0}, _T_522} : _T_530; // @[Mux.scala 46:16:@101.4]
  assign _T_533 = 3'h0 == io_operation_7; // @[Mux.scala 46:19:@102.4]
  assign io_outputs_0 = _T_545[15:0]; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 23:14:@264.4]
  assign io_outputs_1 = _T_556[15:0]; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 23:14:@265.4]
  assign io_outputs_2 = _T_567[15:0]; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 23:14:@266.4]
  assign io_outputs_3 = _T_578[15:0]; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 23:14:@267.4]
  assign io_outputs_4 = _T_589[15:0]; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 23:14:@268.4]
  assign io_outputs_5 = _T_600[15:0]; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 23:14:@269.4]
  assign io_outputs_6 = _T_611[15:0]; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 23:14:@270.4]
  assign io_outputs_7 = _T_622[15:0]; // @[MuxTest_width_16_inputs_8_outputs_8_pipeline_5s.scala 23:14:@271.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_537 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_539 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_541 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_543 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_545 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_548 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_550 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_552 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_554 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_556 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_559 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_561 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_563 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_565 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_567 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_570 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_572 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_574 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_576 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_578 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_581 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_583 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_585 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_587 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_589 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_592 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_594 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_596 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_598 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_600 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_603 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_605 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_607 = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_609 = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_611 = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_614 = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_616 = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_618 = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_620 = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_622 = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_414) begin
      _T_537 <= {{16'd0}, _GEN_7};
    end else begin
      _T_537 <= _T_413;
    end
    _T_539 <= _T_537;
    _T_541 <= _T_539;
    _T_543 <= _T_541;
    _T_545 <= _T_543;
    if (_T_431) begin
      _T_548 <= {{16'd0}, _GEN_23};
    end else begin
      _T_548 <= _T_430;
    end
    _T_550 <= _T_548;
    _T_552 <= _T_550;
    _T_554 <= _T_552;
    _T_556 <= _T_554;
    if (_T_448) begin
      _T_559 <= {{16'd0}, _GEN_39};
    end else begin
      _T_559 <= _T_447;
    end
    _T_561 <= _T_559;
    _T_563 <= _T_561;
    _T_565 <= _T_563;
    _T_567 <= _T_565;
    if (_T_465) begin
      _T_570 <= {{16'd0}, _GEN_55};
    end else begin
      _T_570 <= _T_464;
    end
    _T_572 <= _T_570;
    _T_574 <= _T_572;
    _T_576 <= _T_574;
    _T_578 <= _T_576;
    if (_T_482) begin
      _T_581 <= {{16'd0}, _GEN_71};
    end else begin
      _T_581 <= _T_481;
    end
    _T_583 <= _T_581;
    _T_585 <= _T_583;
    _T_587 <= _T_585;
    _T_589 <= _T_587;
    if (_T_499) begin
      _T_592 <= {{16'd0}, _GEN_87};
    end else begin
      _T_592 <= _T_498;
    end
    _T_594 <= _T_592;
    _T_596 <= _T_594;
    _T_598 <= _T_596;
    _T_600 <= _T_598;
    if (_T_516) begin
      _T_603 <= {{16'd0}, _GEN_103};
    end else begin
      _T_603 <= _T_515;
    end
    _T_605 <= _T_603;
    _T_607 <= _T_605;
    _T_609 <= _T_607;
    _T_611 <= _T_609;
    if (_T_533) begin
      _T_614 <= {{16'd0}, _GEN_119};
    end else begin
      _T_614 <= _T_532;
    end
    _T_616 <= _T_614;
    _T_618 <= _T_616;
    _T_620 <= _T_618;
    _T_622 <= _T_620;
  end
endmodule
