VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_128x256
  FOREIGN fakeram45_128x256 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 151.810 BY 154.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.400 0.070 1.470 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.540 0.070 1.610 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.680 0.070 1.750 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.820 0.070 1.890 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.960 0.070 2.030 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.100 0.070 2.170 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.240 0.070 2.310 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.380 0.070 2.450 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.520 0.070 2.590 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.660 0.070 2.730 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.800 0.070 2.870 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.940 0.070 3.010 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.080 0.070 3.150 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.220 0.070 3.290 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.360 0.070 3.430 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.500 0.070 3.570 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.640 0.070 3.710 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.780 0.070 3.850 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.920 0.070 3.990 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.060 0.070 4.130 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.200 0.070 4.270 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.340 0.070 4.410 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.480 0.070 4.550 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.620 0.070 4.690 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.760 0.070 4.830 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.900 0.070 4.970 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.040 0.070 5.110 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.180 0.070 5.250 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.320 0.070 5.390 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.460 0.070 5.530 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.600 0.070 5.670 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.740 0.070 5.810 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.880 0.070 5.950 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.020 0.070 6.090 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.160 0.070 6.230 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.300 0.070 6.370 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.440 0.070 6.510 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.580 0.070 6.650 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.720 0.070 6.790 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.860 0.070 6.930 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.000 0.070 7.070 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.140 0.070 7.210 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.280 0.070 7.350 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.420 0.070 7.490 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.560 0.070 7.630 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.700 0.070 7.770 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.840 0.070 7.910 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.980 0.070 8.050 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.120 0.070 8.190 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.260 0.070 8.330 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.400 0.070 8.470 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.540 0.070 8.610 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.680 0.070 8.750 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.820 0.070 8.890 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.960 0.070 9.030 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.100 0.070 9.170 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.240 0.070 9.310 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.380 0.070 9.450 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.520 0.070 9.590 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.660 0.070 9.730 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.800 0.070 9.870 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.940 0.070 10.010 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.080 0.070 10.150 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.220 0.070 10.290 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.360 0.070 10.430 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.500 0.070 10.570 ;
    END
  END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.640 0.070 10.710 ;
    END
  END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.780 0.070 10.850 ;
    END
  END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.920 0.070 10.990 ;
    END
  END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.060 0.070 11.130 ;
    END
  END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.200 0.070 11.270 ;
    END
  END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.340 0.070 11.410 ;
    END
  END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.480 0.070 11.550 ;
    END
  END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.620 0.070 11.690 ;
    END
  END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.760 0.070 11.830 ;
    END
  END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.900 0.070 11.970 ;
    END
  END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.040 0.070 12.110 ;
    END
  END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.180 0.070 12.250 ;
    END
  END w_mask_in[77]
  PIN w_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.320 0.070 12.390 ;
    END
  END w_mask_in[78]
  PIN w_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.460 0.070 12.530 ;
    END
  END w_mask_in[79]
  PIN w_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.600 0.070 12.670 ;
    END
  END w_mask_in[80]
  PIN w_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.740 0.070 12.810 ;
    END
  END w_mask_in[81]
  PIN w_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.880 0.070 12.950 ;
    END
  END w_mask_in[82]
  PIN w_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.020 0.070 13.090 ;
    END
  END w_mask_in[83]
  PIN w_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.160 0.070 13.230 ;
    END
  END w_mask_in[84]
  PIN w_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.300 0.070 13.370 ;
    END
  END w_mask_in[85]
  PIN w_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.440 0.070 13.510 ;
    END
  END w_mask_in[86]
  PIN w_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.580 0.070 13.650 ;
    END
  END w_mask_in[87]
  PIN w_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.720 0.070 13.790 ;
    END
  END w_mask_in[88]
  PIN w_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.860 0.070 13.930 ;
    END
  END w_mask_in[89]
  PIN w_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.000 0.070 14.070 ;
    END
  END w_mask_in[90]
  PIN w_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.140 0.070 14.210 ;
    END
  END w_mask_in[91]
  PIN w_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.280 0.070 14.350 ;
    END
  END w_mask_in[92]
  PIN w_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.420 0.070 14.490 ;
    END
  END w_mask_in[93]
  PIN w_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.560 0.070 14.630 ;
    END
  END w_mask_in[94]
  PIN w_mask_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.700 0.070 14.770 ;
    END
  END w_mask_in[95]
  PIN w_mask_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.840 0.070 14.910 ;
    END
  END w_mask_in[96]
  PIN w_mask_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.980 0.070 15.050 ;
    END
  END w_mask_in[97]
  PIN w_mask_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.120 0.070 15.190 ;
    END
  END w_mask_in[98]
  PIN w_mask_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.260 0.070 15.330 ;
    END
  END w_mask_in[99]
  PIN w_mask_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.400 0.070 15.470 ;
    END
  END w_mask_in[100]
  PIN w_mask_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.540 0.070 15.610 ;
    END
  END w_mask_in[101]
  PIN w_mask_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.680 0.070 15.750 ;
    END
  END w_mask_in[102]
  PIN w_mask_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.820 0.070 15.890 ;
    END
  END w_mask_in[103]
  PIN w_mask_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.960 0.070 16.030 ;
    END
  END w_mask_in[104]
  PIN w_mask_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.100 0.070 16.170 ;
    END
  END w_mask_in[105]
  PIN w_mask_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.240 0.070 16.310 ;
    END
  END w_mask_in[106]
  PIN w_mask_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.380 0.070 16.450 ;
    END
  END w_mask_in[107]
  PIN w_mask_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.520 0.070 16.590 ;
    END
  END w_mask_in[108]
  PIN w_mask_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.660 0.070 16.730 ;
    END
  END w_mask_in[109]
  PIN w_mask_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.800 0.070 16.870 ;
    END
  END w_mask_in[110]
  PIN w_mask_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.940 0.070 17.010 ;
    END
  END w_mask_in[111]
  PIN w_mask_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.080 0.070 17.150 ;
    END
  END w_mask_in[112]
  PIN w_mask_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.220 0.070 17.290 ;
    END
  END w_mask_in[113]
  PIN w_mask_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.360 0.070 17.430 ;
    END
  END w_mask_in[114]
  PIN w_mask_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.500 0.070 17.570 ;
    END
  END w_mask_in[115]
  PIN w_mask_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.640 0.070 17.710 ;
    END
  END w_mask_in[116]
  PIN w_mask_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.780 0.070 17.850 ;
    END
  END w_mask_in[117]
  PIN w_mask_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.920 0.070 17.990 ;
    END
  END w_mask_in[118]
  PIN w_mask_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.060 0.070 18.130 ;
    END
  END w_mask_in[119]
  PIN w_mask_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.200 0.070 18.270 ;
    END
  END w_mask_in[120]
  PIN w_mask_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.340 0.070 18.410 ;
    END
  END w_mask_in[121]
  PIN w_mask_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.480 0.070 18.550 ;
    END
  END w_mask_in[122]
  PIN w_mask_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.620 0.070 18.690 ;
    END
  END w_mask_in[123]
  PIN w_mask_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.760 0.070 18.830 ;
    END
  END w_mask_in[124]
  PIN w_mask_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.900 0.070 18.970 ;
    END
  END w_mask_in[125]
  PIN w_mask_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.040 0.070 19.110 ;
    END
  END w_mask_in[126]
  PIN w_mask_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.180 0.070 19.250 ;
    END
  END w_mask_in[127]
  PIN w_mask_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.320 0.070 19.390 ;
    END
  END w_mask_in[128]
  PIN w_mask_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.460 0.070 19.530 ;
    END
  END w_mask_in[129]
  PIN w_mask_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.600 0.070 19.670 ;
    END
  END w_mask_in[130]
  PIN w_mask_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.740 0.070 19.810 ;
    END
  END w_mask_in[131]
  PIN w_mask_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.880 0.070 19.950 ;
    END
  END w_mask_in[132]
  PIN w_mask_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.020 0.070 20.090 ;
    END
  END w_mask_in[133]
  PIN w_mask_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.160 0.070 20.230 ;
    END
  END w_mask_in[134]
  PIN w_mask_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.300 0.070 20.370 ;
    END
  END w_mask_in[135]
  PIN w_mask_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.440 0.070 20.510 ;
    END
  END w_mask_in[136]
  PIN w_mask_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.580 0.070 20.650 ;
    END
  END w_mask_in[137]
  PIN w_mask_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.720 0.070 20.790 ;
    END
  END w_mask_in[138]
  PIN w_mask_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.860 0.070 20.930 ;
    END
  END w_mask_in[139]
  PIN w_mask_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.000 0.070 21.070 ;
    END
  END w_mask_in[140]
  PIN w_mask_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.140 0.070 21.210 ;
    END
  END w_mask_in[141]
  PIN w_mask_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.280 0.070 21.350 ;
    END
  END w_mask_in[142]
  PIN w_mask_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.420 0.070 21.490 ;
    END
  END w_mask_in[143]
  PIN w_mask_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.560 0.070 21.630 ;
    END
  END w_mask_in[144]
  PIN w_mask_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.700 0.070 21.770 ;
    END
  END w_mask_in[145]
  PIN w_mask_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.840 0.070 21.910 ;
    END
  END w_mask_in[146]
  PIN w_mask_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.980 0.070 22.050 ;
    END
  END w_mask_in[147]
  PIN w_mask_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.120 0.070 22.190 ;
    END
  END w_mask_in[148]
  PIN w_mask_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.260 0.070 22.330 ;
    END
  END w_mask_in[149]
  PIN w_mask_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.400 0.070 22.470 ;
    END
  END w_mask_in[150]
  PIN w_mask_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.540 0.070 22.610 ;
    END
  END w_mask_in[151]
  PIN w_mask_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.680 0.070 22.750 ;
    END
  END w_mask_in[152]
  PIN w_mask_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.820 0.070 22.890 ;
    END
  END w_mask_in[153]
  PIN w_mask_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.960 0.070 23.030 ;
    END
  END w_mask_in[154]
  PIN w_mask_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.100 0.070 23.170 ;
    END
  END w_mask_in[155]
  PIN w_mask_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.240 0.070 23.310 ;
    END
  END w_mask_in[156]
  PIN w_mask_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.380 0.070 23.450 ;
    END
  END w_mask_in[157]
  PIN w_mask_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.520 0.070 23.590 ;
    END
  END w_mask_in[158]
  PIN w_mask_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.660 0.070 23.730 ;
    END
  END w_mask_in[159]
  PIN w_mask_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.800 0.070 23.870 ;
    END
  END w_mask_in[160]
  PIN w_mask_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.940 0.070 24.010 ;
    END
  END w_mask_in[161]
  PIN w_mask_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.080 0.070 24.150 ;
    END
  END w_mask_in[162]
  PIN w_mask_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.220 0.070 24.290 ;
    END
  END w_mask_in[163]
  PIN w_mask_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.360 0.070 24.430 ;
    END
  END w_mask_in[164]
  PIN w_mask_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.500 0.070 24.570 ;
    END
  END w_mask_in[165]
  PIN w_mask_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.640 0.070 24.710 ;
    END
  END w_mask_in[166]
  PIN w_mask_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.780 0.070 24.850 ;
    END
  END w_mask_in[167]
  PIN w_mask_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.920 0.070 24.990 ;
    END
  END w_mask_in[168]
  PIN w_mask_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.060 0.070 25.130 ;
    END
  END w_mask_in[169]
  PIN w_mask_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.200 0.070 25.270 ;
    END
  END w_mask_in[170]
  PIN w_mask_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.340 0.070 25.410 ;
    END
  END w_mask_in[171]
  PIN w_mask_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.480 0.070 25.550 ;
    END
  END w_mask_in[172]
  PIN w_mask_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.620 0.070 25.690 ;
    END
  END w_mask_in[173]
  PIN w_mask_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.760 0.070 25.830 ;
    END
  END w_mask_in[174]
  PIN w_mask_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.900 0.070 25.970 ;
    END
  END w_mask_in[175]
  PIN w_mask_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.040 0.070 26.110 ;
    END
  END w_mask_in[176]
  PIN w_mask_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.180 0.070 26.250 ;
    END
  END w_mask_in[177]
  PIN w_mask_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.320 0.070 26.390 ;
    END
  END w_mask_in[178]
  PIN w_mask_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.460 0.070 26.530 ;
    END
  END w_mask_in[179]
  PIN w_mask_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.600 0.070 26.670 ;
    END
  END w_mask_in[180]
  PIN w_mask_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.740 0.070 26.810 ;
    END
  END w_mask_in[181]
  PIN w_mask_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.880 0.070 26.950 ;
    END
  END w_mask_in[182]
  PIN w_mask_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.020 0.070 27.090 ;
    END
  END w_mask_in[183]
  PIN w_mask_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.160 0.070 27.230 ;
    END
  END w_mask_in[184]
  PIN w_mask_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.300 0.070 27.370 ;
    END
  END w_mask_in[185]
  PIN w_mask_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.440 0.070 27.510 ;
    END
  END w_mask_in[186]
  PIN w_mask_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.580 0.070 27.650 ;
    END
  END w_mask_in[187]
  PIN w_mask_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.720 0.070 27.790 ;
    END
  END w_mask_in[188]
  PIN w_mask_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.860 0.070 27.930 ;
    END
  END w_mask_in[189]
  PIN w_mask_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.000 0.070 28.070 ;
    END
  END w_mask_in[190]
  PIN w_mask_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.140 0.070 28.210 ;
    END
  END w_mask_in[191]
  PIN w_mask_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.280 0.070 28.350 ;
    END
  END w_mask_in[192]
  PIN w_mask_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.420 0.070 28.490 ;
    END
  END w_mask_in[193]
  PIN w_mask_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.560 0.070 28.630 ;
    END
  END w_mask_in[194]
  PIN w_mask_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.700 0.070 28.770 ;
    END
  END w_mask_in[195]
  PIN w_mask_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.840 0.070 28.910 ;
    END
  END w_mask_in[196]
  PIN w_mask_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.980 0.070 29.050 ;
    END
  END w_mask_in[197]
  PIN w_mask_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.120 0.070 29.190 ;
    END
  END w_mask_in[198]
  PIN w_mask_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.260 0.070 29.330 ;
    END
  END w_mask_in[199]
  PIN w_mask_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.400 0.070 29.470 ;
    END
  END w_mask_in[200]
  PIN w_mask_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.540 0.070 29.610 ;
    END
  END w_mask_in[201]
  PIN w_mask_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.680 0.070 29.750 ;
    END
  END w_mask_in[202]
  PIN w_mask_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.820 0.070 29.890 ;
    END
  END w_mask_in[203]
  PIN w_mask_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.960 0.070 30.030 ;
    END
  END w_mask_in[204]
  PIN w_mask_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.100 0.070 30.170 ;
    END
  END w_mask_in[205]
  PIN w_mask_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.240 0.070 30.310 ;
    END
  END w_mask_in[206]
  PIN w_mask_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.380 0.070 30.450 ;
    END
  END w_mask_in[207]
  PIN w_mask_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.520 0.070 30.590 ;
    END
  END w_mask_in[208]
  PIN w_mask_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.660 0.070 30.730 ;
    END
  END w_mask_in[209]
  PIN w_mask_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.800 0.070 30.870 ;
    END
  END w_mask_in[210]
  PIN w_mask_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.940 0.070 31.010 ;
    END
  END w_mask_in[211]
  PIN w_mask_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.080 0.070 31.150 ;
    END
  END w_mask_in[212]
  PIN w_mask_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.220 0.070 31.290 ;
    END
  END w_mask_in[213]
  PIN w_mask_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.360 0.070 31.430 ;
    END
  END w_mask_in[214]
  PIN w_mask_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.500 0.070 31.570 ;
    END
  END w_mask_in[215]
  PIN w_mask_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.640 0.070 31.710 ;
    END
  END w_mask_in[216]
  PIN w_mask_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.780 0.070 31.850 ;
    END
  END w_mask_in[217]
  PIN w_mask_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.920 0.070 31.990 ;
    END
  END w_mask_in[218]
  PIN w_mask_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.060 0.070 32.130 ;
    END
  END w_mask_in[219]
  PIN w_mask_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.200 0.070 32.270 ;
    END
  END w_mask_in[220]
  PIN w_mask_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.340 0.070 32.410 ;
    END
  END w_mask_in[221]
  PIN w_mask_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.480 0.070 32.550 ;
    END
  END w_mask_in[222]
  PIN w_mask_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.620 0.070 32.690 ;
    END
  END w_mask_in[223]
  PIN w_mask_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.760 0.070 32.830 ;
    END
  END w_mask_in[224]
  PIN w_mask_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.900 0.070 32.970 ;
    END
  END w_mask_in[225]
  PIN w_mask_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.040 0.070 33.110 ;
    END
  END w_mask_in[226]
  PIN w_mask_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.180 0.070 33.250 ;
    END
  END w_mask_in[227]
  PIN w_mask_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.320 0.070 33.390 ;
    END
  END w_mask_in[228]
  PIN w_mask_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.460 0.070 33.530 ;
    END
  END w_mask_in[229]
  PIN w_mask_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.600 0.070 33.670 ;
    END
  END w_mask_in[230]
  PIN w_mask_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.740 0.070 33.810 ;
    END
  END w_mask_in[231]
  PIN w_mask_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.880 0.070 33.950 ;
    END
  END w_mask_in[232]
  PIN w_mask_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.020 0.070 34.090 ;
    END
  END w_mask_in[233]
  PIN w_mask_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.160 0.070 34.230 ;
    END
  END w_mask_in[234]
  PIN w_mask_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.300 0.070 34.370 ;
    END
  END w_mask_in[235]
  PIN w_mask_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.440 0.070 34.510 ;
    END
  END w_mask_in[236]
  PIN w_mask_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.580 0.070 34.650 ;
    END
  END w_mask_in[237]
  PIN w_mask_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.720 0.070 34.790 ;
    END
  END w_mask_in[238]
  PIN w_mask_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.860 0.070 34.930 ;
    END
  END w_mask_in[239]
  PIN w_mask_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.000 0.070 35.070 ;
    END
  END w_mask_in[240]
  PIN w_mask_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.140 0.070 35.210 ;
    END
  END w_mask_in[241]
  PIN w_mask_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.280 0.070 35.350 ;
    END
  END w_mask_in[242]
  PIN w_mask_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.420 0.070 35.490 ;
    END
  END w_mask_in[243]
  PIN w_mask_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.560 0.070 35.630 ;
    END
  END w_mask_in[244]
  PIN w_mask_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.700 0.070 35.770 ;
    END
  END w_mask_in[245]
  PIN w_mask_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.840 0.070 35.910 ;
    END
  END w_mask_in[246]
  PIN w_mask_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.980 0.070 36.050 ;
    END
  END w_mask_in[247]
  PIN w_mask_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.120 0.070 36.190 ;
    END
  END w_mask_in[248]
  PIN w_mask_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.260 0.070 36.330 ;
    END
  END w_mask_in[249]
  PIN w_mask_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.400 0.070 36.470 ;
    END
  END w_mask_in[250]
  PIN w_mask_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.540 0.070 36.610 ;
    END
  END w_mask_in[251]
  PIN w_mask_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.680 0.070 36.750 ;
    END
  END w_mask_in[252]
  PIN w_mask_in[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.820 0.070 36.890 ;
    END
  END w_mask_in[253]
  PIN w_mask_in[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.960 0.070 37.030 ;
    END
  END w_mask_in[254]
  PIN w_mask_in[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.100 0.070 37.170 ;
    END
  END w_mask_in[255]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.600 0.070 47.670 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.740 0.070 47.810 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.880 0.070 47.950 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.020 0.070 48.090 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.160 0.070 48.230 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.300 0.070 48.370 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.440 0.070 48.510 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.580 0.070 48.650 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.720 0.070 48.790 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.860 0.070 48.930 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.000 0.070 49.070 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.140 0.070 49.210 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.280 0.070 49.350 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.420 0.070 49.490 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.560 0.070 49.630 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.700 0.070 49.770 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.840 0.070 49.910 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.980 0.070 50.050 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.120 0.070 50.190 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.260 0.070 50.330 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.400 0.070 50.470 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.540 0.070 50.610 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.680 0.070 50.750 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.820 0.070 50.890 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.960 0.070 51.030 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.100 0.070 51.170 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.240 0.070 51.310 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.380 0.070 51.450 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.520 0.070 51.590 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.660 0.070 51.730 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.800 0.070 51.870 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.940 0.070 52.010 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.080 0.070 52.150 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.220 0.070 52.290 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.360 0.070 52.430 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.500 0.070 52.570 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.640 0.070 52.710 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.780 0.070 52.850 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.920 0.070 52.990 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.060 0.070 53.130 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.200 0.070 53.270 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.340 0.070 53.410 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.480 0.070 53.550 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.620 0.070 53.690 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.760 0.070 53.830 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.900 0.070 53.970 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.040 0.070 54.110 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.180 0.070 54.250 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.320 0.070 54.390 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.460 0.070 54.530 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.600 0.070 54.670 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.740 0.070 54.810 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.880 0.070 54.950 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.020 0.070 55.090 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.160 0.070 55.230 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.300 0.070 55.370 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.440 0.070 55.510 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.580 0.070 55.650 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.720 0.070 55.790 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.860 0.070 55.930 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.000 0.070 56.070 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.140 0.070 56.210 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.280 0.070 56.350 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.420 0.070 56.490 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.560 0.070 56.630 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.700 0.070 56.770 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.840 0.070 56.910 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.980 0.070 57.050 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.120 0.070 57.190 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.260 0.070 57.330 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.400 0.070 57.470 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.540 0.070 57.610 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.680 0.070 57.750 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.820 0.070 57.890 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.960 0.070 58.030 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.100 0.070 58.170 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.240 0.070 58.310 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.380 0.070 58.450 ;
    END
  END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.520 0.070 58.590 ;
    END
  END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.660 0.070 58.730 ;
    END
  END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.800 0.070 58.870 ;
    END
  END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.940 0.070 59.010 ;
    END
  END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.080 0.070 59.150 ;
    END
  END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.220 0.070 59.290 ;
    END
  END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.360 0.070 59.430 ;
    END
  END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.500 0.070 59.570 ;
    END
  END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.640 0.070 59.710 ;
    END
  END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.780 0.070 59.850 ;
    END
  END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.920 0.070 59.990 ;
    END
  END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.060 0.070 60.130 ;
    END
  END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.200 0.070 60.270 ;
    END
  END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.340 0.070 60.410 ;
    END
  END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.480 0.070 60.550 ;
    END
  END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.620 0.070 60.690 ;
    END
  END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.760 0.070 60.830 ;
    END
  END rd_out[94]
  PIN rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.900 0.070 60.970 ;
    END
  END rd_out[95]
  PIN rd_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.040 0.070 61.110 ;
    END
  END rd_out[96]
  PIN rd_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.180 0.070 61.250 ;
    END
  END rd_out[97]
  PIN rd_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.320 0.070 61.390 ;
    END
  END rd_out[98]
  PIN rd_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.460 0.070 61.530 ;
    END
  END rd_out[99]
  PIN rd_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.600 0.070 61.670 ;
    END
  END rd_out[100]
  PIN rd_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.740 0.070 61.810 ;
    END
  END rd_out[101]
  PIN rd_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.880 0.070 61.950 ;
    END
  END rd_out[102]
  PIN rd_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.020 0.070 62.090 ;
    END
  END rd_out[103]
  PIN rd_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.160 0.070 62.230 ;
    END
  END rd_out[104]
  PIN rd_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.300 0.070 62.370 ;
    END
  END rd_out[105]
  PIN rd_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.440 0.070 62.510 ;
    END
  END rd_out[106]
  PIN rd_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.580 0.070 62.650 ;
    END
  END rd_out[107]
  PIN rd_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.720 0.070 62.790 ;
    END
  END rd_out[108]
  PIN rd_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.860 0.070 62.930 ;
    END
  END rd_out[109]
  PIN rd_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.000 0.070 63.070 ;
    END
  END rd_out[110]
  PIN rd_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.140 0.070 63.210 ;
    END
  END rd_out[111]
  PIN rd_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.280 0.070 63.350 ;
    END
  END rd_out[112]
  PIN rd_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.420 0.070 63.490 ;
    END
  END rd_out[113]
  PIN rd_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.560 0.070 63.630 ;
    END
  END rd_out[114]
  PIN rd_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.700 0.070 63.770 ;
    END
  END rd_out[115]
  PIN rd_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.840 0.070 63.910 ;
    END
  END rd_out[116]
  PIN rd_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.980 0.070 64.050 ;
    END
  END rd_out[117]
  PIN rd_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.120 0.070 64.190 ;
    END
  END rd_out[118]
  PIN rd_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.260 0.070 64.330 ;
    END
  END rd_out[119]
  PIN rd_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.400 0.070 64.470 ;
    END
  END rd_out[120]
  PIN rd_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.540 0.070 64.610 ;
    END
  END rd_out[121]
  PIN rd_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.680 0.070 64.750 ;
    END
  END rd_out[122]
  PIN rd_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.820 0.070 64.890 ;
    END
  END rd_out[123]
  PIN rd_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.960 0.070 65.030 ;
    END
  END rd_out[124]
  PIN rd_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.100 0.070 65.170 ;
    END
  END rd_out[125]
  PIN rd_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.240 0.070 65.310 ;
    END
  END rd_out[126]
  PIN rd_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.380 0.070 65.450 ;
    END
  END rd_out[127]
  PIN rd_out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.520 0.070 65.590 ;
    END
  END rd_out[128]
  PIN rd_out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.660 0.070 65.730 ;
    END
  END rd_out[129]
  PIN rd_out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.800 0.070 65.870 ;
    END
  END rd_out[130]
  PIN rd_out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.940 0.070 66.010 ;
    END
  END rd_out[131]
  PIN rd_out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.080 0.070 66.150 ;
    END
  END rd_out[132]
  PIN rd_out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.220 0.070 66.290 ;
    END
  END rd_out[133]
  PIN rd_out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.360 0.070 66.430 ;
    END
  END rd_out[134]
  PIN rd_out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.500 0.070 66.570 ;
    END
  END rd_out[135]
  PIN rd_out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.640 0.070 66.710 ;
    END
  END rd_out[136]
  PIN rd_out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.780 0.070 66.850 ;
    END
  END rd_out[137]
  PIN rd_out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.920 0.070 66.990 ;
    END
  END rd_out[138]
  PIN rd_out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.060 0.070 67.130 ;
    END
  END rd_out[139]
  PIN rd_out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.200 0.070 67.270 ;
    END
  END rd_out[140]
  PIN rd_out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.340 0.070 67.410 ;
    END
  END rd_out[141]
  PIN rd_out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.480 0.070 67.550 ;
    END
  END rd_out[142]
  PIN rd_out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.620 0.070 67.690 ;
    END
  END rd_out[143]
  PIN rd_out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.760 0.070 67.830 ;
    END
  END rd_out[144]
  PIN rd_out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.900 0.070 67.970 ;
    END
  END rd_out[145]
  PIN rd_out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.040 0.070 68.110 ;
    END
  END rd_out[146]
  PIN rd_out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.180 0.070 68.250 ;
    END
  END rd_out[147]
  PIN rd_out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.320 0.070 68.390 ;
    END
  END rd_out[148]
  PIN rd_out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.460 0.070 68.530 ;
    END
  END rd_out[149]
  PIN rd_out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.600 0.070 68.670 ;
    END
  END rd_out[150]
  PIN rd_out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.740 0.070 68.810 ;
    END
  END rd_out[151]
  PIN rd_out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.880 0.070 68.950 ;
    END
  END rd_out[152]
  PIN rd_out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.020 0.070 69.090 ;
    END
  END rd_out[153]
  PIN rd_out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.160 0.070 69.230 ;
    END
  END rd_out[154]
  PIN rd_out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.300 0.070 69.370 ;
    END
  END rd_out[155]
  PIN rd_out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.440 0.070 69.510 ;
    END
  END rd_out[156]
  PIN rd_out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.580 0.070 69.650 ;
    END
  END rd_out[157]
  PIN rd_out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.720 0.070 69.790 ;
    END
  END rd_out[158]
  PIN rd_out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.860 0.070 69.930 ;
    END
  END rd_out[159]
  PIN rd_out[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.000 0.070 70.070 ;
    END
  END rd_out[160]
  PIN rd_out[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.140 0.070 70.210 ;
    END
  END rd_out[161]
  PIN rd_out[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.280 0.070 70.350 ;
    END
  END rd_out[162]
  PIN rd_out[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.420 0.070 70.490 ;
    END
  END rd_out[163]
  PIN rd_out[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.560 0.070 70.630 ;
    END
  END rd_out[164]
  PIN rd_out[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.700 0.070 70.770 ;
    END
  END rd_out[165]
  PIN rd_out[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.840 0.070 70.910 ;
    END
  END rd_out[166]
  PIN rd_out[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.980 0.070 71.050 ;
    END
  END rd_out[167]
  PIN rd_out[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.120 0.070 71.190 ;
    END
  END rd_out[168]
  PIN rd_out[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.260 0.070 71.330 ;
    END
  END rd_out[169]
  PIN rd_out[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.400 0.070 71.470 ;
    END
  END rd_out[170]
  PIN rd_out[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.540 0.070 71.610 ;
    END
  END rd_out[171]
  PIN rd_out[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.680 0.070 71.750 ;
    END
  END rd_out[172]
  PIN rd_out[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.820 0.070 71.890 ;
    END
  END rd_out[173]
  PIN rd_out[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.960 0.070 72.030 ;
    END
  END rd_out[174]
  PIN rd_out[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.100 0.070 72.170 ;
    END
  END rd_out[175]
  PIN rd_out[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.240 0.070 72.310 ;
    END
  END rd_out[176]
  PIN rd_out[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.380 0.070 72.450 ;
    END
  END rd_out[177]
  PIN rd_out[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.520 0.070 72.590 ;
    END
  END rd_out[178]
  PIN rd_out[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.660 0.070 72.730 ;
    END
  END rd_out[179]
  PIN rd_out[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.800 0.070 72.870 ;
    END
  END rd_out[180]
  PIN rd_out[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.940 0.070 73.010 ;
    END
  END rd_out[181]
  PIN rd_out[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.080 0.070 73.150 ;
    END
  END rd_out[182]
  PIN rd_out[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.220 0.070 73.290 ;
    END
  END rd_out[183]
  PIN rd_out[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.360 0.070 73.430 ;
    END
  END rd_out[184]
  PIN rd_out[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.500 0.070 73.570 ;
    END
  END rd_out[185]
  PIN rd_out[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.640 0.070 73.710 ;
    END
  END rd_out[186]
  PIN rd_out[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.780 0.070 73.850 ;
    END
  END rd_out[187]
  PIN rd_out[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.920 0.070 73.990 ;
    END
  END rd_out[188]
  PIN rd_out[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.060 0.070 74.130 ;
    END
  END rd_out[189]
  PIN rd_out[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.200 0.070 74.270 ;
    END
  END rd_out[190]
  PIN rd_out[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.340 0.070 74.410 ;
    END
  END rd_out[191]
  PIN rd_out[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.480 0.070 74.550 ;
    END
  END rd_out[192]
  PIN rd_out[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.620 0.070 74.690 ;
    END
  END rd_out[193]
  PIN rd_out[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.760 0.070 74.830 ;
    END
  END rd_out[194]
  PIN rd_out[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.900 0.070 74.970 ;
    END
  END rd_out[195]
  PIN rd_out[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.040 0.070 75.110 ;
    END
  END rd_out[196]
  PIN rd_out[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.180 0.070 75.250 ;
    END
  END rd_out[197]
  PIN rd_out[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.320 0.070 75.390 ;
    END
  END rd_out[198]
  PIN rd_out[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.460 0.070 75.530 ;
    END
  END rd_out[199]
  PIN rd_out[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.600 0.070 75.670 ;
    END
  END rd_out[200]
  PIN rd_out[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.740 0.070 75.810 ;
    END
  END rd_out[201]
  PIN rd_out[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.880 0.070 75.950 ;
    END
  END rd_out[202]
  PIN rd_out[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.020 0.070 76.090 ;
    END
  END rd_out[203]
  PIN rd_out[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.160 0.070 76.230 ;
    END
  END rd_out[204]
  PIN rd_out[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.300 0.070 76.370 ;
    END
  END rd_out[205]
  PIN rd_out[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.440 0.070 76.510 ;
    END
  END rd_out[206]
  PIN rd_out[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.580 0.070 76.650 ;
    END
  END rd_out[207]
  PIN rd_out[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.720 0.070 76.790 ;
    END
  END rd_out[208]
  PIN rd_out[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.860 0.070 76.930 ;
    END
  END rd_out[209]
  PIN rd_out[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.000 0.070 77.070 ;
    END
  END rd_out[210]
  PIN rd_out[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.140 0.070 77.210 ;
    END
  END rd_out[211]
  PIN rd_out[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.280 0.070 77.350 ;
    END
  END rd_out[212]
  PIN rd_out[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.420 0.070 77.490 ;
    END
  END rd_out[213]
  PIN rd_out[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.560 0.070 77.630 ;
    END
  END rd_out[214]
  PIN rd_out[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.700 0.070 77.770 ;
    END
  END rd_out[215]
  PIN rd_out[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.840 0.070 77.910 ;
    END
  END rd_out[216]
  PIN rd_out[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.980 0.070 78.050 ;
    END
  END rd_out[217]
  PIN rd_out[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.120 0.070 78.190 ;
    END
  END rd_out[218]
  PIN rd_out[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.260 0.070 78.330 ;
    END
  END rd_out[219]
  PIN rd_out[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.400 0.070 78.470 ;
    END
  END rd_out[220]
  PIN rd_out[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.540 0.070 78.610 ;
    END
  END rd_out[221]
  PIN rd_out[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.680 0.070 78.750 ;
    END
  END rd_out[222]
  PIN rd_out[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.820 0.070 78.890 ;
    END
  END rd_out[223]
  PIN rd_out[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.960 0.070 79.030 ;
    END
  END rd_out[224]
  PIN rd_out[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.100 0.070 79.170 ;
    END
  END rd_out[225]
  PIN rd_out[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.240 0.070 79.310 ;
    END
  END rd_out[226]
  PIN rd_out[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.380 0.070 79.450 ;
    END
  END rd_out[227]
  PIN rd_out[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.520 0.070 79.590 ;
    END
  END rd_out[228]
  PIN rd_out[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.660 0.070 79.730 ;
    END
  END rd_out[229]
  PIN rd_out[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.800 0.070 79.870 ;
    END
  END rd_out[230]
  PIN rd_out[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.940 0.070 80.010 ;
    END
  END rd_out[231]
  PIN rd_out[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.080 0.070 80.150 ;
    END
  END rd_out[232]
  PIN rd_out[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.220 0.070 80.290 ;
    END
  END rd_out[233]
  PIN rd_out[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.360 0.070 80.430 ;
    END
  END rd_out[234]
  PIN rd_out[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.500 0.070 80.570 ;
    END
  END rd_out[235]
  PIN rd_out[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.640 0.070 80.710 ;
    END
  END rd_out[236]
  PIN rd_out[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.780 0.070 80.850 ;
    END
  END rd_out[237]
  PIN rd_out[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.920 0.070 80.990 ;
    END
  END rd_out[238]
  PIN rd_out[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.060 0.070 81.130 ;
    END
  END rd_out[239]
  PIN rd_out[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.200 0.070 81.270 ;
    END
  END rd_out[240]
  PIN rd_out[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.340 0.070 81.410 ;
    END
  END rd_out[241]
  PIN rd_out[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.480 0.070 81.550 ;
    END
  END rd_out[242]
  PIN rd_out[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.620 0.070 81.690 ;
    END
  END rd_out[243]
  PIN rd_out[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.760 0.070 81.830 ;
    END
  END rd_out[244]
  PIN rd_out[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.900 0.070 81.970 ;
    END
  END rd_out[245]
  PIN rd_out[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.040 0.070 82.110 ;
    END
  END rd_out[246]
  PIN rd_out[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.180 0.070 82.250 ;
    END
  END rd_out[247]
  PIN rd_out[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.320 0.070 82.390 ;
    END
  END rd_out[248]
  PIN rd_out[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.460 0.070 82.530 ;
    END
  END rd_out[249]
  PIN rd_out[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.600 0.070 82.670 ;
    END
  END rd_out[250]
  PIN rd_out[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.740 0.070 82.810 ;
    END
  END rd_out[251]
  PIN rd_out[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.880 0.070 82.950 ;
    END
  END rd_out[252]
  PIN rd_out[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.020 0.070 83.090 ;
    END
  END rd_out[253]
  PIN rd_out[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.160 0.070 83.230 ;
    END
  END rd_out[254]
  PIN rd_out[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.300 0.070 83.370 ;
    END
  END rd_out[255]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.800 0.070 93.870 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.940 0.070 94.010 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.080 0.070 94.150 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.220 0.070 94.290 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.360 0.070 94.430 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.500 0.070 94.570 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.640 0.070 94.710 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.780 0.070 94.850 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.920 0.070 94.990 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.060 0.070 95.130 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.200 0.070 95.270 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.340 0.070 95.410 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.480 0.070 95.550 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.620 0.070 95.690 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.760 0.070 95.830 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.900 0.070 95.970 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.040 0.070 96.110 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.180 0.070 96.250 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.320 0.070 96.390 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.460 0.070 96.530 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.600 0.070 96.670 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.740 0.070 96.810 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.880 0.070 96.950 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.020 0.070 97.090 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.160 0.070 97.230 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.300 0.070 97.370 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.440 0.070 97.510 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.580 0.070 97.650 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.720 0.070 97.790 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.860 0.070 97.930 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.000 0.070 98.070 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.140 0.070 98.210 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.280 0.070 98.350 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.420 0.070 98.490 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.560 0.070 98.630 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.700 0.070 98.770 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.840 0.070 98.910 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.980 0.070 99.050 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.120 0.070 99.190 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.260 0.070 99.330 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.400 0.070 99.470 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.540 0.070 99.610 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.680 0.070 99.750 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.820 0.070 99.890 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.960 0.070 100.030 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.100 0.070 100.170 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.240 0.070 100.310 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.380 0.070 100.450 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.520 0.070 100.590 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.660 0.070 100.730 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.800 0.070 100.870 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.940 0.070 101.010 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.080 0.070 101.150 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.220 0.070 101.290 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.360 0.070 101.430 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.500 0.070 101.570 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.640 0.070 101.710 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.780 0.070 101.850 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.920 0.070 101.990 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.060 0.070 102.130 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.200 0.070 102.270 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.340 0.070 102.410 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.480 0.070 102.550 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.620 0.070 102.690 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.760 0.070 102.830 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.900 0.070 102.970 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.040 0.070 103.110 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.180 0.070 103.250 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.320 0.070 103.390 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.460 0.070 103.530 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.600 0.070 103.670 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.740 0.070 103.810 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.880 0.070 103.950 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.020 0.070 104.090 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.160 0.070 104.230 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.300 0.070 104.370 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.440 0.070 104.510 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.580 0.070 104.650 ;
    END
  END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.720 0.070 104.790 ;
    END
  END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.860 0.070 104.930 ;
    END
  END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.000 0.070 105.070 ;
    END
  END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.140 0.070 105.210 ;
    END
  END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.280 0.070 105.350 ;
    END
  END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.420 0.070 105.490 ;
    END
  END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.560 0.070 105.630 ;
    END
  END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.700 0.070 105.770 ;
    END
  END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.840 0.070 105.910 ;
    END
  END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.980 0.070 106.050 ;
    END
  END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.120 0.070 106.190 ;
    END
  END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.260 0.070 106.330 ;
    END
  END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.400 0.070 106.470 ;
    END
  END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.540 0.070 106.610 ;
    END
  END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.680 0.070 106.750 ;
    END
  END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.820 0.070 106.890 ;
    END
  END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.960 0.070 107.030 ;
    END
  END wd_in[94]
  PIN wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.100 0.070 107.170 ;
    END
  END wd_in[95]
  PIN wd_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.240 0.070 107.310 ;
    END
  END wd_in[96]
  PIN wd_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.380 0.070 107.450 ;
    END
  END wd_in[97]
  PIN wd_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.520 0.070 107.590 ;
    END
  END wd_in[98]
  PIN wd_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.660 0.070 107.730 ;
    END
  END wd_in[99]
  PIN wd_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.800 0.070 107.870 ;
    END
  END wd_in[100]
  PIN wd_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.940 0.070 108.010 ;
    END
  END wd_in[101]
  PIN wd_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.080 0.070 108.150 ;
    END
  END wd_in[102]
  PIN wd_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.220 0.070 108.290 ;
    END
  END wd_in[103]
  PIN wd_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.360 0.070 108.430 ;
    END
  END wd_in[104]
  PIN wd_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.500 0.070 108.570 ;
    END
  END wd_in[105]
  PIN wd_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.640 0.070 108.710 ;
    END
  END wd_in[106]
  PIN wd_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.780 0.070 108.850 ;
    END
  END wd_in[107]
  PIN wd_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.920 0.070 108.990 ;
    END
  END wd_in[108]
  PIN wd_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.060 0.070 109.130 ;
    END
  END wd_in[109]
  PIN wd_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.200 0.070 109.270 ;
    END
  END wd_in[110]
  PIN wd_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.340 0.070 109.410 ;
    END
  END wd_in[111]
  PIN wd_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.480 0.070 109.550 ;
    END
  END wd_in[112]
  PIN wd_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.620 0.070 109.690 ;
    END
  END wd_in[113]
  PIN wd_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.760 0.070 109.830 ;
    END
  END wd_in[114]
  PIN wd_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.900 0.070 109.970 ;
    END
  END wd_in[115]
  PIN wd_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.040 0.070 110.110 ;
    END
  END wd_in[116]
  PIN wd_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.180 0.070 110.250 ;
    END
  END wd_in[117]
  PIN wd_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.320 0.070 110.390 ;
    END
  END wd_in[118]
  PIN wd_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.460 0.070 110.530 ;
    END
  END wd_in[119]
  PIN wd_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.600 0.070 110.670 ;
    END
  END wd_in[120]
  PIN wd_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.740 0.070 110.810 ;
    END
  END wd_in[121]
  PIN wd_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.880 0.070 110.950 ;
    END
  END wd_in[122]
  PIN wd_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.020 0.070 111.090 ;
    END
  END wd_in[123]
  PIN wd_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.160 0.070 111.230 ;
    END
  END wd_in[124]
  PIN wd_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.300 0.070 111.370 ;
    END
  END wd_in[125]
  PIN wd_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.440 0.070 111.510 ;
    END
  END wd_in[126]
  PIN wd_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.580 0.070 111.650 ;
    END
  END wd_in[127]
  PIN wd_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.720 0.070 111.790 ;
    END
  END wd_in[128]
  PIN wd_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.860 0.070 111.930 ;
    END
  END wd_in[129]
  PIN wd_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.000 0.070 112.070 ;
    END
  END wd_in[130]
  PIN wd_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.140 0.070 112.210 ;
    END
  END wd_in[131]
  PIN wd_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.280 0.070 112.350 ;
    END
  END wd_in[132]
  PIN wd_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.420 0.070 112.490 ;
    END
  END wd_in[133]
  PIN wd_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.560 0.070 112.630 ;
    END
  END wd_in[134]
  PIN wd_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.700 0.070 112.770 ;
    END
  END wd_in[135]
  PIN wd_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.840 0.070 112.910 ;
    END
  END wd_in[136]
  PIN wd_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.980 0.070 113.050 ;
    END
  END wd_in[137]
  PIN wd_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.120 0.070 113.190 ;
    END
  END wd_in[138]
  PIN wd_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.260 0.070 113.330 ;
    END
  END wd_in[139]
  PIN wd_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.400 0.070 113.470 ;
    END
  END wd_in[140]
  PIN wd_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.540 0.070 113.610 ;
    END
  END wd_in[141]
  PIN wd_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.680 0.070 113.750 ;
    END
  END wd_in[142]
  PIN wd_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.820 0.070 113.890 ;
    END
  END wd_in[143]
  PIN wd_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.960 0.070 114.030 ;
    END
  END wd_in[144]
  PIN wd_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.100 0.070 114.170 ;
    END
  END wd_in[145]
  PIN wd_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.240 0.070 114.310 ;
    END
  END wd_in[146]
  PIN wd_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.380 0.070 114.450 ;
    END
  END wd_in[147]
  PIN wd_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.520 0.070 114.590 ;
    END
  END wd_in[148]
  PIN wd_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.660 0.070 114.730 ;
    END
  END wd_in[149]
  PIN wd_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.800 0.070 114.870 ;
    END
  END wd_in[150]
  PIN wd_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.940 0.070 115.010 ;
    END
  END wd_in[151]
  PIN wd_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.080 0.070 115.150 ;
    END
  END wd_in[152]
  PIN wd_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.220 0.070 115.290 ;
    END
  END wd_in[153]
  PIN wd_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.360 0.070 115.430 ;
    END
  END wd_in[154]
  PIN wd_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.500 0.070 115.570 ;
    END
  END wd_in[155]
  PIN wd_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.640 0.070 115.710 ;
    END
  END wd_in[156]
  PIN wd_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.780 0.070 115.850 ;
    END
  END wd_in[157]
  PIN wd_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.920 0.070 115.990 ;
    END
  END wd_in[158]
  PIN wd_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.060 0.070 116.130 ;
    END
  END wd_in[159]
  PIN wd_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.200 0.070 116.270 ;
    END
  END wd_in[160]
  PIN wd_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.340 0.070 116.410 ;
    END
  END wd_in[161]
  PIN wd_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.480 0.070 116.550 ;
    END
  END wd_in[162]
  PIN wd_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.620 0.070 116.690 ;
    END
  END wd_in[163]
  PIN wd_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.760 0.070 116.830 ;
    END
  END wd_in[164]
  PIN wd_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.900 0.070 116.970 ;
    END
  END wd_in[165]
  PIN wd_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.040 0.070 117.110 ;
    END
  END wd_in[166]
  PIN wd_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.180 0.070 117.250 ;
    END
  END wd_in[167]
  PIN wd_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.320 0.070 117.390 ;
    END
  END wd_in[168]
  PIN wd_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.460 0.070 117.530 ;
    END
  END wd_in[169]
  PIN wd_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.600 0.070 117.670 ;
    END
  END wd_in[170]
  PIN wd_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.740 0.070 117.810 ;
    END
  END wd_in[171]
  PIN wd_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.880 0.070 117.950 ;
    END
  END wd_in[172]
  PIN wd_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.020 0.070 118.090 ;
    END
  END wd_in[173]
  PIN wd_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.160 0.070 118.230 ;
    END
  END wd_in[174]
  PIN wd_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.300 0.070 118.370 ;
    END
  END wd_in[175]
  PIN wd_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.440 0.070 118.510 ;
    END
  END wd_in[176]
  PIN wd_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.580 0.070 118.650 ;
    END
  END wd_in[177]
  PIN wd_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.720 0.070 118.790 ;
    END
  END wd_in[178]
  PIN wd_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.860 0.070 118.930 ;
    END
  END wd_in[179]
  PIN wd_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.000 0.070 119.070 ;
    END
  END wd_in[180]
  PIN wd_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.140 0.070 119.210 ;
    END
  END wd_in[181]
  PIN wd_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.280 0.070 119.350 ;
    END
  END wd_in[182]
  PIN wd_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.420 0.070 119.490 ;
    END
  END wd_in[183]
  PIN wd_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.560 0.070 119.630 ;
    END
  END wd_in[184]
  PIN wd_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.700 0.070 119.770 ;
    END
  END wd_in[185]
  PIN wd_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.840 0.070 119.910 ;
    END
  END wd_in[186]
  PIN wd_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.980 0.070 120.050 ;
    END
  END wd_in[187]
  PIN wd_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.120 0.070 120.190 ;
    END
  END wd_in[188]
  PIN wd_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.260 0.070 120.330 ;
    END
  END wd_in[189]
  PIN wd_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.400 0.070 120.470 ;
    END
  END wd_in[190]
  PIN wd_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.540 0.070 120.610 ;
    END
  END wd_in[191]
  PIN wd_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.680 0.070 120.750 ;
    END
  END wd_in[192]
  PIN wd_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.820 0.070 120.890 ;
    END
  END wd_in[193]
  PIN wd_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.960 0.070 121.030 ;
    END
  END wd_in[194]
  PIN wd_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.100 0.070 121.170 ;
    END
  END wd_in[195]
  PIN wd_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.240 0.070 121.310 ;
    END
  END wd_in[196]
  PIN wd_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.380 0.070 121.450 ;
    END
  END wd_in[197]
  PIN wd_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.520 0.070 121.590 ;
    END
  END wd_in[198]
  PIN wd_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.660 0.070 121.730 ;
    END
  END wd_in[199]
  PIN wd_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.800 0.070 121.870 ;
    END
  END wd_in[200]
  PIN wd_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.940 0.070 122.010 ;
    END
  END wd_in[201]
  PIN wd_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.080 0.070 122.150 ;
    END
  END wd_in[202]
  PIN wd_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.220 0.070 122.290 ;
    END
  END wd_in[203]
  PIN wd_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.360 0.070 122.430 ;
    END
  END wd_in[204]
  PIN wd_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.500 0.070 122.570 ;
    END
  END wd_in[205]
  PIN wd_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.640 0.070 122.710 ;
    END
  END wd_in[206]
  PIN wd_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.780 0.070 122.850 ;
    END
  END wd_in[207]
  PIN wd_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.920 0.070 122.990 ;
    END
  END wd_in[208]
  PIN wd_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.060 0.070 123.130 ;
    END
  END wd_in[209]
  PIN wd_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.200 0.070 123.270 ;
    END
  END wd_in[210]
  PIN wd_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.340 0.070 123.410 ;
    END
  END wd_in[211]
  PIN wd_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.480 0.070 123.550 ;
    END
  END wd_in[212]
  PIN wd_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.620 0.070 123.690 ;
    END
  END wd_in[213]
  PIN wd_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.760 0.070 123.830 ;
    END
  END wd_in[214]
  PIN wd_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.900 0.070 123.970 ;
    END
  END wd_in[215]
  PIN wd_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.040 0.070 124.110 ;
    END
  END wd_in[216]
  PIN wd_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.180 0.070 124.250 ;
    END
  END wd_in[217]
  PIN wd_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.320 0.070 124.390 ;
    END
  END wd_in[218]
  PIN wd_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.460 0.070 124.530 ;
    END
  END wd_in[219]
  PIN wd_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.600 0.070 124.670 ;
    END
  END wd_in[220]
  PIN wd_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.740 0.070 124.810 ;
    END
  END wd_in[221]
  PIN wd_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.880 0.070 124.950 ;
    END
  END wd_in[222]
  PIN wd_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.020 0.070 125.090 ;
    END
  END wd_in[223]
  PIN wd_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.160 0.070 125.230 ;
    END
  END wd_in[224]
  PIN wd_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.300 0.070 125.370 ;
    END
  END wd_in[225]
  PIN wd_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.440 0.070 125.510 ;
    END
  END wd_in[226]
  PIN wd_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.580 0.070 125.650 ;
    END
  END wd_in[227]
  PIN wd_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.720 0.070 125.790 ;
    END
  END wd_in[228]
  PIN wd_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.860 0.070 125.930 ;
    END
  END wd_in[229]
  PIN wd_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.000 0.070 126.070 ;
    END
  END wd_in[230]
  PIN wd_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.140 0.070 126.210 ;
    END
  END wd_in[231]
  PIN wd_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.280 0.070 126.350 ;
    END
  END wd_in[232]
  PIN wd_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.420 0.070 126.490 ;
    END
  END wd_in[233]
  PIN wd_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.560 0.070 126.630 ;
    END
  END wd_in[234]
  PIN wd_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.700 0.070 126.770 ;
    END
  END wd_in[235]
  PIN wd_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.840 0.070 126.910 ;
    END
  END wd_in[236]
  PIN wd_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.980 0.070 127.050 ;
    END
  END wd_in[237]
  PIN wd_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.120 0.070 127.190 ;
    END
  END wd_in[238]
  PIN wd_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.260 0.070 127.330 ;
    END
  END wd_in[239]
  PIN wd_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.400 0.070 127.470 ;
    END
  END wd_in[240]
  PIN wd_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.540 0.070 127.610 ;
    END
  END wd_in[241]
  PIN wd_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.680 0.070 127.750 ;
    END
  END wd_in[242]
  PIN wd_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.820 0.070 127.890 ;
    END
  END wd_in[243]
  PIN wd_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.960 0.070 128.030 ;
    END
  END wd_in[244]
  PIN wd_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.100 0.070 128.170 ;
    END
  END wd_in[245]
  PIN wd_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.240 0.070 128.310 ;
    END
  END wd_in[246]
  PIN wd_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.380 0.070 128.450 ;
    END
  END wd_in[247]
  PIN wd_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.520 0.070 128.590 ;
    END
  END wd_in[248]
  PIN wd_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.660 0.070 128.730 ;
    END
  END wd_in[249]
  PIN wd_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.800 0.070 128.870 ;
    END
  END wd_in[250]
  PIN wd_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.940 0.070 129.010 ;
    END
  END wd_in[251]
  PIN wd_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.080 0.070 129.150 ;
    END
  END wd_in[252]
  PIN wd_in[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.220 0.070 129.290 ;
    END
  END wd_in[253]
  PIN wd_in[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.360 0.070 129.430 ;
    END
  END wd_in[254]
  PIN wd_in[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.500 0.070 129.570 ;
    END
  END wd_in[255]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.000 0.070 140.070 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.140 0.070 140.210 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.280 0.070 140.350 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.420 0.070 140.490 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.560 0.070 140.630 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.700 0.070 140.770 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.840 0.070 140.910 ;
    END
  END addr_in[6]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.340 0.070 151.410 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.480 0.070 151.550 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.620 0.070 151.690 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 152.600 ;
      RECT 3.500 1.400 3.780 152.600 ;
      RECT 5.740 1.400 6.020 152.600 ;
      RECT 7.980 1.400 8.260 152.600 ;
      RECT 10.220 1.400 10.500 152.600 ;
      RECT 12.460 1.400 12.740 152.600 ;
      RECT 14.700 1.400 14.980 152.600 ;
      RECT 16.940 1.400 17.220 152.600 ;
      RECT 19.180 1.400 19.460 152.600 ;
      RECT 21.420 1.400 21.700 152.600 ;
      RECT 23.660 1.400 23.940 152.600 ;
      RECT 25.900 1.400 26.180 152.600 ;
      RECT 28.140 1.400 28.420 152.600 ;
      RECT 30.380 1.400 30.660 152.600 ;
      RECT 32.620 1.400 32.900 152.600 ;
      RECT 34.860 1.400 35.140 152.600 ;
      RECT 37.100 1.400 37.380 152.600 ;
      RECT 39.340 1.400 39.620 152.600 ;
      RECT 41.580 1.400 41.860 152.600 ;
      RECT 43.820 1.400 44.100 152.600 ;
      RECT 46.060 1.400 46.340 152.600 ;
      RECT 48.300 1.400 48.580 152.600 ;
      RECT 50.540 1.400 50.820 152.600 ;
      RECT 52.780 1.400 53.060 152.600 ;
      RECT 55.020 1.400 55.300 152.600 ;
      RECT 57.260 1.400 57.540 152.600 ;
      RECT 59.500 1.400 59.780 152.600 ;
      RECT 61.740 1.400 62.020 152.600 ;
      RECT 63.980 1.400 64.260 152.600 ;
      RECT 66.220 1.400 66.500 152.600 ;
      RECT 68.460 1.400 68.740 152.600 ;
      RECT 70.700 1.400 70.980 152.600 ;
      RECT 72.940 1.400 73.220 152.600 ;
      RECT 75.180 1.400 75.460 152.600 ;
      RECT 77.420 1.400 77.700 152.600 ;
      RECT 79.660 1.400 79.940 152.600 ;
      RECT 81.900 1.400 82.180 152.600 ;
      RECT 84.140 1.400 84.420 152.600 ;
      RECT 86.380 1.400 86.660 152.600 ;
      RECT 88.620 1.400 88.900 152.600 ;
      RECT 90.860 1.400 91.140 152.600 ;
      RECT 93.100 1.400 93.380 152.600 ;
      RECT 95.340 1.400 95.620 152.600 ;
      RECT 97.580 1.400 97.860 152.600 ;
      RECT 99.820 1.400 100.100 152.600 ;
      RECT 102.060 1.400 102.340 152.600 ;
      RECT 104.300 1.400 104.580 152.600 ;
      RECT 106.540 1.400 106.820 152.600 ;
      RECT 108.780 1.400 109.060 152.600 ;
      RECT 111.020 1.400 111.300 152.600 ;
      RECT 113.260 1.400 113.540 152.600 ;
      RECT 115.500 1.400 115.780 152.600 ;
      RECT 117.740 1.400 118.020 152.600 ;
      RECT 119.980 1.400 120.260 152.600 ;
      RECT 122.220 1.400 122.500 152.600 ;
      RECT 124.460 1.400 124.740 152.600 ;
      RECT 126.700 1.400 126.980 152.600 ;
      RECT 128.940 1.400 129.220 152.600 ;
      RECT 131.180 1.400 131.460 152.600 ;
      RECT 133.420 1.400 133.700 152.600 ;
      RECT 135.660 1.400 135.940 152.600 ;
      RECT 137.900 1.400 138.180 152.600 ;
      RECT 140.140 1.400 140.420 152.600 ;
      RECT 142.380 1.400 142.660 152.600 ;
      RECT 144.620 1.400 144.900 152.600 ;
      RECT 146.860 1.400 147.140 152.600 ;
      RECT 149.100 1.400 149.380 152.600 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 152.600 ;
      RECT 4.620 1.400 4.900 152.600 ;
      RECT 6.860 1.400 7.140 152.600 ;
      RECT 9.100 1.400 9.380 152.600 ;
      RECT 11.340 1.400 11.620 152.600 ;
      RECT 13.580 1.400 13.860 152.600 ;
      RECT 15.820 1.400 16.100 152.600 ;
      RECT 18.060 1.400 18.340 152.600 ;
      RECT 20.300 1.400 20.580 152.600 ;
      RECT 22.540 1.400 22.820 152.600 ;
      RECT 24.780 1.400 25.060 152.600 ;
      RECT 27.020 1.400 27.300 152.600 ;
      RECT 29.260 1.400 29.540 152.600 ;
      RECT 31.500 1.400 31.780 152.600 ;
      RECT 33.740 1.400 34.020 152.600 ;
      RECT 35.980 1.400 36.260 152.600 ;
      RECT 38.220 1.400 38.500 152.600 ;
      RECT 40.460 1.400 40.740 152.600 ;
      RECT 42.700 1.400 42.980 152.600 ;
      RECT 44.940 1.400 45.220 152.600 ;
      RECT 47.180 1.400 47.460 152.600 ;
      RECT 49.420 1.400 49.700 152.600 ;
      RECT 51.660 1.400 51.940 152.600 ;
      RECT 53.900 1.400 54.180 152.600 ;
      RECT 56.140 1.400 56.420 152.600 ;
      RECT 58.380 1.400 58.660 152.600 ;
      RECT 60.620 1.400 60.900 152.600 ;
      RECT 62.860 1.400 63.140 152.600 ;
      RECT 65.100 1.400 65.380 152.600 ;
      RECT 67.340 1.400 67.620 152.600 ;
      RECT 69.580 1.400 69.860 152.600 ;
      RECT 71.820 1.400 72.100 152.600 ;
      RECT 74.060 1.400 74.340 152.600 ;
      RECT 76.300 1.400 76.580 152.600 ;
      RECT 78.540 1.400 78.820 152.600 ;
      RECT 80.780 1.400 81.060 152.600 ;
      RECT 83.020 1.400 83.300 152.600 ;
      RECT 85.260 1.400 85.540 152.600 ;
      RECT 87.500 1.400 87.780 152.600 ;
      RECT 89.740 1.400 90.020 152.600 ;
      RECT 91.980 1.400 92.260 152.600 ;
      RECT 94.220 1.400 94.500 152.600 ;
      RECT 96.460 1.400 96.740 152.600 ;
      RECT 98.700 1.400 98.980 152.600 ;
      RECT 100.940 1.400 101.220 152.600 ;
      RECT 103.180 1.400 103.460 152.600 ;
      RECT 105.420 1.400 105.700 152.600 ;
      RECT 107.660 1.400 107.940 152.600 ;
      RECT 109.900 1.400 110.180 152.600 ;
      RECT 112.140 1.400 112.420 152.600 ;
      RECT 114.380 1.400 114.660 152.600 ;
      RECT 116.620 1.400 116.900 152.600 ;
      RECT 118.860 1.400 119.140 152.600 ;
      RECT 121.100 1.400 121.380 152.600 ;
      RECT 123.340 1.400 123.620 152.600 ;
      RECT 125.580 1.400 125.860 152.600 ;
      RECT 127.820 1.400 128.100 152.600 ;
      RECT 130.060 1.400 130.340 152.600 ;
      RECT 132.300 1.400 132.580 152.600 ;
      RECT 134.540 1.400 134.820 152.600 ;
      RECT 136.780 1.400 137.060 152.600 ;
      RECT 139.020 1.400 139.300 152.600 ;
      RECT 141.260 1.400 141.540 152.600 ;
      RECT 143.500 1.400 143.780 152.600 ;
      RECT 145.740 1.400 146.020 152.600 ;
      RECT 147.980 1.400 148.260 152.600 ;
      RECT 150.220 1.400 150.500 152.600 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 151.810 154.000 ;
    LAYER metal2 ;
    RECT 0 0 151.810 154.000 ;
    LAYER metal3 ;
    RECT 0.070 0 151.810 154.000 ;
    RECT 0 0.000 0.070 1.400 ;
    RECT 0 1.470 0.070 1.540 ;
    RECT 0 1.610 0.070 1.680 ;
    RECT 0 1.750 0.070 1.820 ;
    RECT 0 1.890 0.070 1.960 ;
    RECT 0 2.030 0.070 2.100 ;
    RECT 0 2.170 0.070 2.240 ;
    RECT 0 2.310 0.070 2.380 ;
    RECT 0 2.450 0.070 2.520 ;
    RECT 0 2.590 0.070 2.660 ;
    RECT 0 2.730 0.070 2.800 ;
    RECT 0 2.870 0.070 2.940 ;
    RECT 0 3.010 0.070 3.080 ;
    RECT 0 3.150 0.070 3.220 ;
    RECT 0 3.290 0.070 3.360 ;
    RECT 0 3.430 0.070 3.500 ;
    RECT 0 3.570 0.070 3.640 ;
    RECT 0 3.710 0.070 3.780 ;
    RECT 0 3.850 0.070 3.920 ;
    RECT 0 3.990 0.070 4.060 ;
    RECT 0 4.130 0.070 4.200 ;
    RECT 0 4.270 0.070 4.340 ;
    RECT 0 4.410 0.070 4.480 ;
    RECT 0 4.550 0.070 4.620 ;
    RECT 0 4.690 0.070 4.760 ;
    RECT 0 4.830 0.070 4.900 ;
    RECT 0 4.970 0.070 5.040 ;
    RECT 0 5.110 0.070 5.180 ;
    RECT 0 5.250 0.070 5.320 ;
    RECT 0 5.390 0.070 5.460 ;
    RECT 0 5.530 0.070 5.600 ;
    RECT 0 5.670 0.070 5.740 ;
    RECT 0 5.810 0.070 5.880 ;
    RECT 0 5.950 0.070 6.020 ;
    RECT 0 6.090 0.070 6.160 ;
    RECT 0 6.230 0.070 6.300 ;
    RECT 0 6.370 0.070 6.440 ;
    RECT 0 6.510 0.070 6.580 ;
    RECT 0 6.650 0.070 6.720 ;
    RECT 0 6.790 0.070 6.860 ;
    RECT 0 6.930 0.070 7.000 ;
    RECT 0 7.070 0.070 7.140 ;
    RECT 0 7.210 0.070 7.280 ;
    RECT 0 7.350 0.070 7.420 ;
    RECT 0 7.490 0.070 7.560 ;
    RECT 0 7.630 0.070 7.700 ;
    RECT 0 7.770 0.070 7.840 ;
    RECT 0 7.910 0.070 7.980 ;
    RECT 0 8.050 0.070 8.120 ;
    RECT 0 8.190 0.070 8.260 ;
    RECT 0 8.330 0.070 8.400 ;
    RECT 0 8.470 0.070 8.540 ;
    RECT 0 8.610 0.070 8.680 ;
    RECT 0 8.750 0.070 8.820 ;
    RECT 0 8.890 0.070 8.960 ;
    RECT 0 9.030 0.070 9.100 ;
    RECT 0 9.170 0.070 9.240 ;
    RECT 0 9.310 0.070 9.380 ;
    RECT 0 9.450 0.070 9.520 ;
    RECT 0 9.590 0.070 9.660 ;
    RECT 0 9.730 0.070 9.800 ;
    RECT 0 9.870 0.070 9.940 ;
    RECT 0 10.010 0.070 10.080 ;
    RECT 0 10.150 0.070 10.220 ;
    RECT 0 10.290 0.070 10.360 ;
    RECT 0 10.430 0.070 10.500 ;
    RECT 0 10.570 0.070 10.640 ;
    RECT 0 10.710 0.070 10.780 ;
    RECT 0 10.850 0.070 10.920 ;
    RECT 0 10.990 0.070 11.060 ;
    RECT 0 11.130 0.070 11.200 ;
    RECT 0 11.270 0.070 11.340 ;
    RECT 0 11.410 0.070 11.480 ;
    RECT 0 11.550 0.070 11.620 ;
    RECT 0 11.690 0.070 11.760 ;
    RECT 0 11.830 0.070 11.900 ;
    RECT 0 11.970 0.070 12.040 ;
    RECT 0 12.110 0.070 12.180 ;
    RECT 0 12.250 0.070 12.320 ;
    RECT 0 12.390 0.070 12.460 ;
    RECT 0 12.530 0.070 12.600 ;
    RECT 0 12.670 0.070 12.740 ;
    RECT 0 12.810 0.070 12.880 ;
    RECT 0 12.950 0.070 13.020 ;
    RECT 0 13.090 0.070 13.160 ;
    RECT 0 13.230 0.070 13.300 ;
    RECT 0 13.370 0.070 13.440 ;
    RECT 0 13.510 0.070 13.580 ;
    RECT 0 13.650 0.070 13.720 ;
    RECT 0 13.790 0.070 13.860 ;
    RECT 0 13.930 0.070 14.000 ;
    RECT 0 14.070 0.070 14.140 ;
    RECT 0 14.210 0.070 14.280 ;
    RECT 0 14.350 0.070 14.420 ;
    RECT 0 14.490 0.070 14.560 ;
    RECT 0 14.630 0.070 14.700 ;
    RECT 0 14.770 0.070 14.840 ;
    RECT 0 14.910 0.070 14.980 ;
    RECT 0 15.050 0.070 15.120 ;
    RECT 0 15.190 0.070 15.260 ;
    RECT 0 15.330 0.070 15.400 ;
    RECT 0 15.470 0.070 15.540 ;
    RECT 0 15.610 0.070 15.680 ;
    RECT 0 15.750 0.070 15.820 ;
    RECT 0 15.890 0.070 15.960 ;
    RECT 0 16.030 0.070 16.100 ;
    RECT 0 16.170 0.070 16.240 ;
    RECT 0 16.310 0.070 16.380 ;
    RECT 0 16.450 0.070 16.520 ;
    RECT 0 16.590 0.070 16.660 ;
    RECT 0 16.730 0.070 16.800 ;
    RECT 0 16.870 0.070 16.940 ;
    RECT 0 17.010 0.070 17.080 ;
    RECT 0 17.150 0.070 17.220 ;
    RECT 0 17.290 0.070 17.360 ;
    RECT 0 17.430 0.070 17.500 ;
    RECT 0 17.570 0.070 17.640 ;
    RECT 0 17.710 0.070 17.780 ;
    RECT 0 17.850 0.070 17.920 ;
    RECT 0 17.990 0.070 18.060 ;
    RECT 0 18.130 0.070 18.200 ;
    RECT 0 18.270 0.070 18.340 ;
    RECT 0 18.410 0.070 18.480 ;
    RECT 0 18.550 0.070 18.620 ;
    RECT 0 18.690 0.070 18.760 ;
    RECT 0 18.830 0.070 18.900 ;
    RECT 0 18.970 0.070 19.040 ;
    RECT 0 19.110 0.070 19.180 ;
    RECT 0 19.250 0.070 19.320 ;
    RECT 0 19.390 0.070 19.460 ;
    RECT 0 19.530 0.070 19.600 ;
    RECT 0 19.670 0.070 19.740 ;
    RECT 0 19.810 0.070 19.880 ;
    RECT 0 19.950 0.070 20.020 ;
    RECT 0 20.090 0.070 20.160 ;
    RECT 0 20.230 0.070 20.300 ;
    RECT 0 20.370 0.070 20.440 ;
    RECT 0 20.510 0.070 20.580 ;
    RECT 0 20.650 0.070 20.720 ;
    RECT 0 20.790 0.070 20.860 ;
    RECT 0 20.930 0.070 21.000 ;
    RECT 0 21.070 0.070 21.140 ;
    RECT 0 21.210 0.070 21.280 ;
    RECT 0 21.350 0.070 21.420 ;
    RECT 0 21.490 0.070 21.560 ;
    RECT 0 21.630 0.070 21.700 ;
    RECT 0 21.770 0.070 21.840 ;
    RECT 0 21.910 0.070 21.980 ;
    RECT 0 22.050 0.070 22.120 ;
    RECT 0 22.190 0.070 22.260 ;
    RECT 0 22.330 0.070 22.400 ;
    RECT 0 22.470 0.070 22.540 ;
    RECT 0 22.610 0.070 22.680 ;
    RECT 0 22.750 0.070 22.820 ;
    RECT 0 22.890 0.070 22.960 ;
    RECT 0 23.030 0.070 23.100 ;
    RECT 0 23.170 0.070 23.240 ;
    RECT 0 23.310 0.070 23.380 ;
    RECT 0 23.450 0.070 23.520 ;
    RECT 0 23.590 0.070 23.660 ;
    RECT 0 23.730 0.070 23.800 ;
    RECT 0 23.870 0.070 23.940 ;
    RECT 0 24.010 0.070 24.080 ;
    RECT 0 24.150 0.070 24.220 ;
    RECT 0 24.290 0.070 24.360 ;
    RECT 0 24.430 0.070 24.500 ;
    RECT 0 24.570 0.070 24.640 ;
    RECT 0 24.710 0.070 24.780 ;
    RECT 0 24.850 0.070 24.920 ;
    RECT 0 24.990 0.070 25.060 ;
    RECT 0 25.130 0.070 25.200 ;
    RECT 0 25.270 0.070 25.340 ;
    RECT 0 25.410 0.070 25.480 ;
    RECT 0 25.550 0.070 25.620 ;
    RECT 0 25.690 0.070 25.760 ;
    RECT 0 25.830 0.070 25.900 ;
    RECT 0 25.970 0.070 26.040 ;
    RECT 0 26.110 0.070 26.180 ;
    RECT 0 26.250 0.070 26.320 ;
    RECT 0 26.390 0.070 26.460 ;
    RECT 0 26.530 0.070 26.600 ;
    RECT 0 26.670 0.070 26.740 ;
    RECT 0 26.810 0.070 26.880 ;
    RECT 0 26.950 0.070 27.020 ;
    RECT 0 27.090 0.070 27.160 ;
    RECT 0 27.230 0.070 27.300 ;
    RECT 0 27.370 0.070 27.440 ;
    RECT 0 27.510 0.070 27.580 ;
    RECT 0 27.650 0.070 27.720 ;
    RECT 0 27.790 0.070 27.860 ;
    RECT 0 27.930 0.070 28.000 ;
    RECT 0 28.070 0.070 28.140 ;
    RECT 0 28.210 0.070 28.280 ;
    RECT 0 28.350 0.070 28.420 ;
    RECT 0 28.490 0.070 28.560 ;
    RECT 0 28.630 0.070 28.700 ;
    RECT 0 28.770 0.070 28.840 ;
    RECT 0 28.910 0.070 28.980 ;
    RECT 0 29.050 0.070 29.120 ;
    RECT 0 29.190 0.070 29.260 ;
    RECT 0 29.330 0.070 29.400 ;
    RECT 0 29.470 0.070 29.540 ;
    RECT 0 29.610 0.070 29.680 ;
    RECT 0 29.750 0.070 29.820 ;
    RECT 0 29.890 0.070 29.960 ;
    RECT 0 30.030 0.070 30.100 ;
    RECT 0 30.170 0.070 30.240 ;
    RECT 0 30.310 0.070 30.380 ;
    RECT 0 30.450 0.070 30.520 ;
    RECT 0 30.590 0.070 30.660 ;
    RECT 0 30.730 0.070 30.800 ;
    RECT 0 30.870 0.070 30.940 ;
    RECT 0 31.010 0.070 31.080 ;
    RECT 0 31.150 0.070 31.220 ;
    RECT 0 31.290 0.070 31.360 ;
    RECT 0 31.430 0.070 31.500 ;
    RECT 0 31.570 0.070 31.640 ;
    RECT 0 31.710 0.070 31.780 ;
    RECT 0 31.850 0.070 31.920 ;
    RECT 0 31.990 0.070 32.060 ;
    RECT 0 32.130 0.070 32.200 ;
    RECT 0 32.270 0.070 32.340 ;
    RECT 0 32.410 0.070 32.480 ;
    RECT 0 32.550 0.070 32.620 ;
    RECT 0 32.690 0.070 32.760 ;
    RECT 0 32.830 0.070 32.900 ;
    RECT 0 32.970 0.070 33.040 ;
    RECT 0 33.110 0.070 33.180 ;
    RECT 0 33.250 0.070 33.320 ;
    RECT 0 33.390 0.070 33.460 ;
    RECT 0 33.530 0.070 33.600 ;
    RECT 0 33.670 0.070 33.740 ;
    RECT 0 33.810 0.070 33.880 ;
    RECT 0 33.950 0.070 34.020 ;
    RECT 0 34.090 0.070 34.160 ;
    RECT 0 34.230 0.070 34.300 ;
    RECT 0 34.370 0.070 34.440 ;
    RECT 0 34.510 0.070 34.580 ;
    RECT 0 34.650 0.070 34.720 ;
    RECT 0 34.790 0.070 34.860 ;
    RECT 0 34.930 0.070 35.000 ;
    RECT 0 35.070 0.070 35.140 ;
    RECT 0 35.210 0.070 35.280 ;
    RECT 0 35.350 0.070 35.420 ;
    RECT 0 35.490 0.070 35.560 ;
    RECT 0 35.630 0.070 35.700 ;
    RECT 0 35.770 0.070 35.840 ;
    RECT 0 35.910 0.070 35.980 ;
    RECT 0 36.050 0.070 36.120 ;
    RECT 0 36.190 0.070 36.260 ;
    RECT 0 36.330 0.070 36.400 ;
    RECT 0 36.470 0.070 36.540 ;
    RECT 0 36.610 0.070 36.680 ;
    RECT 0 36.750 0.070 36.820 ;
    RECT 0 36.890 0.070 36.960 ;
    RECT 0 37.030 0.070 37.100 ;
    RECT 0 37.170 0.070 47.600 ;
    RECT 0 47.670 0.070 47.740 ;
    RECT 0 47.810 0.070 47.880 ;
    RECT 0 47.950 0.070 48.020 ;
    RECT 0 48.090 0.070 48.160 ;
    RECT 0 48.230 0.070 48.300 ;
    RECT 0 48.370 0.070 48.440 ;
    RECT 0 48.510 0.070 48.580 ;
    RECT 0 48.650 0.070 48.720 ;
    RECT 0 48.790 0.070 48.860 ;
    RECT 0 48.930 0.070 49.000 ;
    RECT 0 49.070 0.070 49.140 ;
    RECT 0 49.210 0.070 49.280 ;
    RECT 0 49.350 0.070 49.420 ;
    RECT 0 49.490 0.070 49.560 ;
    RECT 0 49.630 0.070 49.700 ;
    RECT 0 49.770 0.070 49.840 ;
    RECT 0 49.910 0.070 49.980 ;
    RECT 0 50.050 0.070 50.120 ;
    RECT 0 50.190 0.070 50.260 ;
    RECT 0 50.330 0.070 50.400 ;
    RECT 0 50.470 0.070 50.540 ;
    RECT 0 50.610 0.070 50.680 ;
    RECT 0 50.750 0.070 50.820 ;
    RECT 0 50.890 0.070 50.960 ;
    RECT 0 51.030 0.070 51.100 ;
    RECT 0 51.170 0.070 51.240 ;
    RECT 0 51.310 0.070 51.380 ;
    RECT 0 51.450 0.070 51.520 ;
    RECT 0 51.590 0.070 51.660 ;
    RECT 0 51.730 0.070 51.800 ;
    RECT 0 51.870 0.070 51.940 ;
    RECT 0 52.010 0.070 52.080 ;
    RECT 0 52.150 0.070 52.220 ;
    RECT 0 52.290 0.070 52.360 ;
    RECT 0 52.430 0.070 52.500 ;
    RECT 0 52.570 0.070 52.640 ;
    RECT 0 52.710 0.070 52.780 ;
    RECT 0 52.850 0.070 52.920 ;
    RECT 0 52.990 0.070 53.060 ;
    RECT 0 53.130 0.070 53.200 ;
    RECT 0 53.270 0.070 53.340 ;
    RECT 0 53.410 0.070 53.480 ;
    RECT 0 53.550 0.070 53.620 ;
    RECT 0 53.690 0.070 53.760 ;
    RECT 0 53.830 0.070 53.900 ;
    RECT 0 53.970 0.070 54.040 ;
    RECT 0 54.110 0.070 54.180 ;
    RECT 0 54.250 0.070 54.320 ;
    RECT 0 54.390 0.070 54.460 ;
    RECT 0 54.530 0.070 54.600 ;
    RECT 0 54.670 0.070 54.740 ;
    RECT 0 54.810 0.070 54.880 ;
    RECT 0 54.950 0.070 55.020 ;
    RECT 0 55.090 0.070 55.160 ;
    RECT 0 55.230 0.070 55.300 ;
    RECT 0 55.370 0.070 55.440 ;
    RECT 0 55.510 0.070 55.580 ;
    RECT 0 55.650 0.070 55.720 ;
    RECT 0 55.790 0.070 55.860 ;
    RECT 0 55.930 0.070 56.000 ;
    RECT 0 56.070 0.070 56.140 ;
    RECT 0 56.210 0.070 56.280 ;
    RECT 0 56.350 0.070 56.420 ;
    RECT 0 56.490 0.070 56.560 ;
    RECT 0 56.630 0.070 56.700 ;
    RECT 0 56.770 0.070 56.840 ;
    RECT 0 56.910 0.070 56.980 ;
    RECT 0 57.050 0.070 57.120 ;
    RECT 0 57.190 0.070 57.260 ;
    RECT 0 57.330 0.070 57.400 ;
    RECT 0 57.470 0.070 57.540 ;
    RECT 0 57.610 0.070 57.680 ;
    RECT 0 57.750 0.070 57.820 ;
    RECT 0 57.890 0.070 57.960 ;
    RECT 0 58.030 0.070 58.100 ;
    RECT 0 58.170 0.070 58.240 ;
    RECT 0 58.310 0.070 58.380 ;
    RECT 0 58.450 0.070 58.520 ;
    RECT 0 58.590 0.070 58.660 ;
    RECT 0 58.730 0.070 58.800 ;
    RECT 0 58.870 0.070 58.940 ;
    RECT 0 59.010 0.070 59.080 ;
    RECT 0 59.150 0.070 59.220 ;
    RECT 0 59.290 0.070 59.360 ;
    RECT 0 59.430 0.070 59.500 ;
    RECT 0 59.570 0.070 59.640 ;
    RECT 0 59.710 0.070 59.780 ;
    RECT 0 59.850 0.070 59.920 ;
    RECT 0 59.990 0.070 60.060 ;
    RECT 0 60.130 0.070 60.200 ;
    RECT 0 60.270 0.070 60.340 ;
    RECT 0 60.410 0.070 60.480 ;
    RECT 0 60.550 0.070 60.620 ;
    RECT 0 60.690 0.070 60.760 ;
    RECT 0 60.830 0.070 60.900 ;
    RECT 0 60.970 0.070 61.040 ;
    RECT 0 61.110 0.070 61.180 ;
    RECT 0 61.250 0.070 61.320 ;
    RECT 0 61.390 0.070 61.460 ;
    RECT 0 61.530 0.070 61.600 ;
    RECT 0 61.670 0.070 61.740 ;
    RECT 0 61.810 0.070 61.880 ;
    RECT 0 61.950 0.070 62.020 ;
    RECT 0 62.090 0.070 62.160 ;
    RECT 0 62.230 0.070 62.300 ;
    RECT 0 62.370 0.070 62.440 ;
    RECT 0 62.510 0.070 62.580 ;
    RECT 0 62.650 0.070 62.720 ;
    RECT 0 62.790 0.070 62.860 ;
    RECT 0 62.930 0.070 63.000 ;
    RECT 0 63.070 0.070 63.140 ;
    RECT 0 63.210 0.070 63.280 ;
    RECT 0 63.350 0.070 63.420 ;
    RECT 0 63.490 0.070 63.560 ;
    RECT 0 63.630 0.070 63.700 ;
    RECT 0 63.770 0.070 63.840 ;
    RECT 0 63.910 0.070 63.980 ;
    RECT 0 64.050 0.070 64.120 ;
    RECT 0 64.190 0.070 64.260 ;
    RECT 0 64.330 0.070 64.400 ;
    RECT 0 64.470 0.070 64.540 ;
    RECT 0 64.610 0.070 64.680 ;
    RECT 0 64.750 0.070 64.820 ;
    RECT 0 64.890 0.070 64.960 ;
    RECT 0 65.030 0.070 65.100 ;
    RECT 0 65.170 0.070 65.240 ;
    RECT 0 65.310 0.070 65.380 ;
    RECT 0 65.450 0.070 65.520 ;
    RECT 0 65.590 0.070 65.660 ;
    RECT 0 65.730 0.070 65.800 ;
    RECT 0 65.870 0.070 65.940 ;
    RECT 0 66.010 0.070 66.080 ;
    RECT 0 66.150 0.070 66.220 ;
    RECT 0 66.290 0.070 66.360 ;
    RECT 0 66.430 0.070 66.500 ;
    RECT 0 66.570 0.070 66.640 ;
    RECT 0 66.710 0.070 66.780 ;
    RECT 0 66.850 0.070 66.920 ;
    RECT 0 66.990 0.070 67.060 ;
    RECT 0 67.130 0.070 67.200 ;
    RECT 0 67.270 0.070 67.340 ;
    RECT 0 67.410 0.070 67.480 ;
    RECT 0 67.550 0.070 67.620 ;
    RECT 0 67.690 0.070 67.760 ;
    RECT 0 67.830 0.070 67.900 ;
    RECT 0 67.970 0.070 68.040 ;
    RECT 0 68.110 0.070 68.180 ;
    RECT 0 68.250 0.070 68.320 ;
    RECT 0 68.390 0.070 68.460 ;
    RECT 0 68.530 0.070 68.600 ;
    RECT 0 68.670 0.070 68.740 ;
    RECT 0 68.810 0.070 68.880 ;
    RECT 0 68.950 0.070 69.020 ;
    RECT 0 69.090 0.070 69.160 ;
    RECT 0 69.230 0.070 69.300 ;
    RECT 0 69.370 0.070 69.440 ;
    RECT 0 69.510 0.070 69.580 ;
    RECT 0 69.650 0.070 69.720 ;
    RECT 0 69.790 0.070 69.860 ;
    RECT 0 69.930 0.070 70.000 ;
    RECT 0 70.070 0.070 70.140 ;
    RECT 0 70.210 0.070 70.280 ;
    RECT 0 70.350 0.070 70.420 ;
    RECT 0 70.490 0.070 70.560 ;
    RECT 0 70.630 0.070 70.700 ;
    RECT 0 70.770 0.070 70.840 ;
    RECT 0 70.910 0.070 70.980 ;
    RECT 0 71.050 0.070 71.120 ;
    RECT 0 71.190 0.070 71.260 ;
    RECT 0 71.330 0.070 71.400 ;
    RECT 0 71.470 0.070 71.540 ;
    RECT 0 71.610 0.070 71.680 ;
    RECT 0 71.750 0.070 71.820 ;
    RECT 0 71.890 0.070 71.960 ;
    RECT 0 72.030 0.070 72.100 ;
    RECT 0 72.170 0.070 72.240 ;
    RECT 0 72.310 0.070 72.380 ;
    RECT 0 72.450 0.070 72.520 ;
    RECT 0 72.590 0.070 72.660 ;
    RECT 0 72.730 0.070 72.800 ;
    RECT 0 72.870 0.070 72.940 ;
    RECT 0 73.010 0.070 73.080 ;
    RECT 0 73.150 0.070 73.220 ;
    RECT 0 73.290 0.070 73.360 ;
    RECT 0 73.430 0.070 73.500 ;
    RECT 0 73.570 0.070 73.640 ;
    RECT 0 73.710 0.070 73.780 ;
    RECT 0 73.850 0.070 73.920 ;
    RECT 0 73.990 0.070 74.060 ;
    RECT 0 74.130 0.070 74.200 ;
    RECT 0 74.270 0.070 74.340 ;
    RECT 0 74.410 0.070 74.480 ;
    RECT 0 74.550 0.070 74.620 ;
    RECT 0 74.690 0.070 74.760 ;
    RECT 0 74.830 0.070 74.900 ;
    RECT 0 74.970 0.070 75.040 ;
    RECT 0 75.110 0.070 75.180 ;
    RECT 0 75.250 0.070 75.320 ;
    RECT 0 75.390 0.070 75.460 ;
    RECT 0 75.530 0.070 75.600 ;
    RECT 0 75.670 0.070 75.740 ;
    RECT 0 75.810 0.070 75.880 ;
    RECT 0 75.950 0.070 76.020 ;
    RECT 0 76.090 0.070 76.160 ;
    RECT 0 76.230 0.070 76.300 ;
    RECT 0 76.370 0.070 76.440 ;
    RECT 0 76.510 0.070 76.580 ;
    RECT 0 76.650 0.070 76.720 ;
    RECT 0 76.790 0.070 76.860 ;
    RECT 0 76.930 0.070 77.000 ;
    RECT 0 77.070 0.070 77.140 ;
    RECT 0 77.210 0.070 77.280 ;
    RECT 0 77.350 0.070 77.420 ;
    RECT 0 77.490 0.070 77.560 ;
    RECT 0 77.630 0.070 77.700 ;
    RECT 0 77.770 0.070 77.840 ;
    RECT 0 77.910 0.070 77.980 ;
    RECT 0 78.050 0.070 78.120 ;
    RECT 0 78.190 0.070 78.260 ;
    RECT 0 78.330 0.070 78.400 ;
    RECT 0 78.470 0.070 78.540 ;
    RECT 0 78.610 0.070 78.680 ;
    RECT 0 78.750 0.070 78.820 ;
    RECT 0 78.890 0.070 78.960 ;
    RECT 0 79.030 0.070 79.100 ;
    RECT 0 79.170 0.070 79.240 ;
    RECT 0 79.310 0.070 79.380 ;
    RECT 0 79.450 0.070 79.520 ;
    RECT 0 79.590 0.070 79.660 ;
    RECT 0 79.730 0.070 79.800 ;
    RECT 0 79.870 0.070 79.940 ;
    RECT 0 80.010 0.070 80.080 ;
    RECT 0 80.150 0.070 80.220 ;
    RECT 0 80.290 0.070 80.360 ;
    RECT 0 80.430 0.070 80.500 ;
    RECT 0 80.570 0.070 80.640 ;
    RECT 0 80.710 0.070 80.780 ;
    RECT 0 80.850 0.070 80.920 ;
    RECT 0 80.990 0.070 81.060 ;
    RECT 0 81.130 0.070 81.200 ;
    RECT 0 81.270 0.070 81.340 ;
    RECT 0 81.410 0.070 81.480 ;
    RECT 0 81.550 0.070 81.620 ;
    RECT 0 81.690 0.070 81.760 ;
    RECT 0 81.830 0.070 81.900 ;
    RECT 0 81.970 0.070 82.040 ;
    RECT 0 82.110 0.070 82.180 ;
    RECT 0 82.250 0.070 82.320 ;
    RECT 0 82.390 0.070 82.460 ;
    RECT 0 82.530 0.070 82.600 ;
    RECT 0 82.670 0.070 82.740 ;
    RECT 0 82.810 0.070 82.880 ;
    RECT 0 82.950 0.070 83.020 ;
    RECT 0 83.090 0.070 83.160 ;
    RECT 0 83.230 0.070 83.300 ;
    RECT 0 83.370 0.070 93.800 ;
    RECT 0 93.870 0.070 93.940 ;
    RECT 0 94.010 0.070 94.080 ;
    RECT 0 94.150 0.070 94.220 ;
    RECT 0 94.290 0.070 94.360 ;
    RECT 0 94.430 0.070 94.500 ;
    RECT 0 94.570 0.070 94.640 ;
    RECT 0 94.710 0.070 94.780 ;
    RECT 0 94.850 0.070 94.920 ;
    RECT 0 94.990 0.070 95.060 ;
    RECT 0 95.130 0.070 95.200 ;
    RECT 0 95.270 0.070 95.340 ;
    RECT 0 95.410 0.070 95.480 ;
    RECT 0 95.550 0.070 95.620 ;
    RECT 0 95.690 0.070 95.760 ;
    RECT 0 95.830 0.070 95.900 ;
    RECT 0 95.970 0.070 96.040 ;
    RECT 0 96.110 0.070 96.180 ;
    RECT 0 96.250 0.070 96.320 ;
    RECT 0 96.390 0.070 96.460 ;
    RECT 0 96.530 0.070 96.600 ;
    RECT 0 96.670 0.070 96.740 ;
    RECT 0 96.810 0.070 96.880 ;
    RECT 0 96.950 0.070 97.020 ;
    RECT 0 97.090 0.070 97.160 ;
    RECT 0 97.230 0.070 97.300 ;
    RECT 0 97.370 0.070 97.440 ;
    RECT 0 97.510 0.070 97.580 ;
    RECT 0 97.650 0.070 97.720 ;
    RECT 0 97.790 0.070 97.860 ;
    RECT 0 97.930 0.070 98.000 ;
    RECT 0 98.070 0.070 98.140 ;
    RECT 0 98.210 0.070 98.280 ;
    RECT 0 98.350 0.070 98.420 ;
    RECT 0 98.490 0.070 98.560 ;
    RECT 0 98.630 0.070 98.700 ;
    RECT 0 98.770 0.070 98.840 ;
    RECT 0 98.910 0.070 98.980 ;
    RECT 0 99.050 0.070 99.120 ;
    RECT 0 99.190 0.070 99.260 ;
    RECT 0 99.330 0.070 99.400 ;
    RECT 0 99.470 0.070 99.540 ;
    RECT 0 99.610 0.070 99.680 ;
    RECT 0 99.750 0.070 99.820 ;
    RECT 0 99.890 0.070 99.960 ;
    RECT 0 100.030 0.070 100.100 ;
    RECT 0 100.170 0.070 100.240 ;
    RECT 0 100.310 0.070 100.380 ;
    RECT 0 100.450 0.070 100.520 ;
    RECT 0 100.590 0.070 100.660 ;
    RECT 0 100.730 0.070 100.800 ;
    RECT 0 100.870 0.070 100.940 ;
    RECT 0 101.010 0.070 101.080 ;
    RECT 0 101.150 0.070 101.220 ;
    RECT 0 101.290 0.070 101.360 ;
    RECT 0 101.430 0.070 101.500 ;
    RECT 0 101.570 0.070 101.640 ;
    RECT 0 101.710 0.070 101.780 ;
    RECT 0 101.850 0.070 101.920 ;
    RECT 0 101.990 0.070 102.060 ;
    RECT 0 102.130 0.070 102.200 ;
    RECT 0 102.270 0.070 102.340 ;
    RECT 0 102.410 0.070 102.480 ;
    RECT 0 102.550 0.070 102.620 ;
    RECT 0 102.690 0.070 102.760 ;
    RECT 0 102.830 0.070 102.900 ;
    RECT 0 102.970 0.070 103.040 ;
    RECT 0 103.110 0.070 103.180 ;
    RECT 0 103.250 0.070 103.320 ;
    RECT 0 103.390 0.070 103.460 ;
    RECT 0 103.530 0.070 103.600 ;
    RECT 0 103.670 0.070 103.740 ;
    RECT 0 103.810 0.070 103.880 ;
    RECT 0 103.950 0.070 104.020 ;
    RECT 0 104.090 0.070 104.160 ;
    RECT 0 104.230 0.070 104.300 ;
    RECT 0 104.370 0.070 104.440 ;
    RECT 0 104.510 0.070 104.580 ;
    RECT 0 104.650 0.070 104.720 ;
    RECT 0 104.790 0.070 104.860 ;
    RECT 0 104.930 0.070 105.000 ;
    RECT 0 105.070 0.070 105.140 ;
    RECT 0 105.210 0.070 105.280 ;
    RECT 0 105.350 0.070 105.420 ;
    RECT 0 105.490 0.070 105.560 ;
    RECT 0 105.630 0.070 105.700 ;
    RECT 0 105.770 0.070 105.840 ;
    RECT 0 105.910 0.070 105.980 ;
    RECT 0 106.050 0.070 106.120 ;
    RECT 0 106.190 0.070 106.260 ;
    RECT 0 106.330 0.070 106.400 ;
    RECT 0 106.470 0.070 106.540 ;
    RECT 0 106.610 0.070 106.680 ;
    RECT 0 106.750 0.070 106.820 ;
    RECT 0 106.890 0.070 106.960 ;
    RECT 0 107.030 0.070 107.100 ;
    RECT 0 107.170 0.070 107.240 ;
    RECT 0 107.310 0.070 107.380 ;
    RECT 0 107.450 0.070 107.520 ;
    RECT 0 107.590 0.070 107.660 ;
    RECT 0 107.730 0.070 107.800 ;
    RECT 0 107.870 0.070 107.940 ;
    RECT 0 108.010 0.070 108.080 ;
    RECT 0 108.150 0.070 108.220 ;
    RECT 0 108.290 0.070 108.360 ;
    RECT 0 108.430 0.070 108.500 ;
    RECT 0 108.570 0.070 108.640 ;
    RECT 0 108.710 0.070 108.780 ;
    RECT 0 108.850 0.070 108.920 ;
    RECT 0 108.990 0.070 109.060 ;
    RECT 0 109.130 0.070 109.200 ;
    RECT 0 109.270 0.070 109.340 ;
    RECT 0 109.410 0.070 109.480 ;
    RECT 0 109.550 0.070 109.620 ;
    RECT 0 109.690 0.070 109.760 ;
    RECT 0 109.830 0.070 109.900 ;
    RECT 0 109.970 0.070 110.040 ;
    RECT 0 110.110 0.070 110.180 ;
    RECT 0 110.250 0.070 110.320 ;
    RECT 0 110.390 0.070 110.460 ;
    RECT 0 110.530 0.070 110.600 ;
    RECT 0 110.670 0.070 110.740 ;
    RECT 0 110.810 0.070 110.880 ;
    RECT 0 110.950 0.070 111.020 ;
    RECT 0 111.090 0.070 111.160 ;
    RECT 0 111.230 0.070 111.300 ;
    RECT 0 111.370 0.070 111.440 ;
    RECT 0 111.510 0.070 111.580 ;
    RECT 0 111.650 0.070 111.720 ;
    RECT 0 111.790 0.070 111.860 ;
    RECT 0 111.930 0.070 112.000 ;
    RECT 0 112.070 0.070 112.140 ;
    RECT 0 112.210 0.070 112.280 ;
    RECT 0 112.350 0.070 112.420 ;
    RECT 0 112.490 0.070 112.560 ;
    RECT 0 112.630 0.070 112.700 ;
    RECT 0 112.770 0.070 112.840 ;
    RECT 0 112.910 0.070 112.980 ;
    RECT 0 113.050 0.070 113.120 ;
    RECT 0 113.190 0.070 113.260 ;
    RECT 0 113.330 0.070 113.400 ;
    RECT 0 113.470 0.070 113.540 ;
    RECT 0 113.610 0.070 113.680 ;
    RECT 0 113.750 0.070 113.820 ;
    RECT 0 113.890 0.070 113.960 ;
    RECT 0 114.030 0.070 114.100 ;
    RECT 0 114.170 0.070 114.240 ;
    RECT 0 114.310 0.070 114.380 ;
    RECT 0 114.450 0.070 114.520 ;
    RECT 0 114.590 0.070 114.660 ;
    RECT 0 114.730 0.070 114.800 ;
    RECT 0 114.870 0.070 114.940 ;
    RECT 0 115.010 0.070 115.080 ;
    RECT 0 115.150 0.070 115.220 ;
    RECT 0 115.290 0.070 115.360 ;
    RECT 0 115.430 0.070 115.500 ;
    RECT 0 115.570 0.070 115.640 ;
    RECT 0 115.710 0.070 115.780 ;
    RECT 0 115.850 0.070 115.920 ;
    RECT 0 115.990 0.070 116.060 ;
    RECT 0 116.130 0.070 116.200 ;
    RECT 0 116.270 0.070 116.340 ;
    RECT 0 116.410 0.070 116.480 ;
    RECT 0 116.550 0.070 116.620 ;
    RECT 0 116.690 0.070 116.760 ;
    RECT 0 116.830 0.070 116.900 ;
    RECT 0 116.970 0.070 117.040 ;
    RECT 0 117.110 0.070 117.180 ;
    RECT 0 117.250 0.070 117.320 ;
    RECT 0 117.390 0.070 117.460 ;
    RECT 0 117.530 0.070 117.600 ;
    RECT 0 117.670 0.070 117.740 ;
    RECT 0 117.810 0.070 117.880 ;
    RECT 0 117.950 0.070 118.020 ;
    RECT 0 118.090 0.070 118.160 ;
    RECT 0 118.230 0.070 118.300 ;
    RECT 0 118.370 0.070 118.440 ;
    RECT 0 118.510 0.070 118.580 ;
    RECT 0 118.650 0.070 118.720 ;
    RECT 0 118.790 0.070 118.860 ;
    RECT 0 118.930 0.070 119.000 ;
    RECT 0 119.070 0.070 119.140 ;
    RECT 0 119.210 0.070 119.280 ;
    RECT 0 119.350 0.070 119.420 ;
    RECT 0 119.490 0.070 119.560 ;
    RECT 0 119.630 0.070 119.700 ;
    RECT 0 119.770 0.070 119.840 ;
    RECT 0 119.910 0.070 119.980 ;
    RECT 0 120.050 0.070 120.120 ;
    RECT 0 120.190 0.070 120.260 ;
    RECT 0 120.330 0.070 120.400 ;
    RECT 0 120.470 0.070 120.540 ;
    RECT 0 120.610 0.070 120.680 ;
    RECT 0 120.750 0.070 120.820 ;
    RECT 0 120.890 0.070 120.960 ;
    RECT 0 121.030 0.070 121.100 ;
    RECT 0 121.170 0.070 121.240 ;
    RECT 0 121.310 0.070 121.380 ;
    RECT 0 121.450 0.070 121.520 ;
    RECT 0 121.590 0.070 121.660 ;
    RECT 0 121.730 0.070 121.800 ;
    RECT 0 121.870 0.070 121.940 ;
    RECT 0 122.010 0.070 122.080 ;
    RECT 0 122.150 0.070 122.220 ;
    RECT 0 122.290 0.070 122.360 ;
    RECT 0 122.430 0.070 122.500 ;
    RECT 0 122.570 0.070 122.640 ;
    RECT 0 122.710 0.070 122.780 ;
    RECT 0 122.850 0.070 122.920 ;
    RECT 0 122.990 0.070 123.060 ;
    RECT 0 123.130 0.070 123.200 ;
    RECT 0 123.270 0.070 123.340 ;
    RECT 0 123.410 0.070 123.480 ;
    RECT 0 123.550 0.070 123.620 ;
    RECT 0 123.690 0.070 123.760 ;
    RECT 0 123.830 0.070 123.900 ;
    RECT 0 123.970 0.070 124.040 ;
    RECT 0 124.110 0.070 124.180 ;
    RECT 0 124.250 0.070 124.320 ;
    RECT 0 124.390 0.070 124.460 ;
    RECT 0 124.530 0.070 124.600 ;
    RECT 0 124.670 0.070 124.740 ;
    RECT 0 124.810 0.070 124.880 ;
    RECT 0 124.950 0.070 125.020 ;
    RECT 0 125.090 0.070 125.160 ;
    RECT 0 125.230 0.070 125.300 ;
    RECT 0 125.370 0.070 125.440 ;
    RECT 0 125.510 0.070 125.580 ;
    RECT 0 125.650 0.070 125.720 ;
    RECT 0 125.790 0.070 125.860 ;
    RECT 0 125.930 0.070 126.000 ;
    RECT 0 126.070 0.070 126.140 ;
    RECT 0 126.210 0.070 126.280 ;
    RECT 0 126.350 0.070 126.420 ;
    RECT 0 126.490 0.070 126.560 ;
    RECT 0 126.630 0.070 126.700 ;
    RECT 0 126.770 0.070 126.840 ;
    RECT 0 126.910 0.070 126.980 ;
    RECT 0 127.050 0.070 127.120 ;
    RECT 0 127.190 0.070 127.260 ;
    RECT 0 127.330 0.070 127.400 ;
    RECT 0 127.470 0.070 127.540 ;
    RECT 0 127.610 0.070 127.680 ;
    RECT 0 127.750 0.070 127.820 ;
    RECT 0 127.890 0.070 127.960 ;
    RECT 0 128.030 0.070 128.100 ;
    RECT 0 128.170 0.070 128.240 ;
    RECT 0 128.310 0.070 128.380 ;
    RECT 0 128.450 0.070 128.520 ;
    RECT 0 128.590 0.070 128.660 ;
    RECT 0 128.730 0.070 128.800 ;
    RECT 0 128.870 0.070 128.940 ;
    RECT 0 129.010 0.070 129.080 ;
    RECT 0 129.150 0.070 129.220 ;
    RECT 0 129.290 0.070 129.360 ;
    RECT 0 129.430 0.070 129.500 ;
    RECT 0 129.570 0.070 140.000 ;
    RECT 0 140.070 0.070 140.140 ;
    RECT 0 140.210 0.070 140.280 ;
    RECT 0 140.350 0.070 140.420 ;
    RECT 0 140.490 0.070 140.560 ;
    RECT 0 140.630 0.070 140.700 ;
    RECT 0 140.770 0.070 140.840 ;
    RECT 0 140.910 0.070 151.340 ;
    RECT 0 151.410 0.070 151.480 ;
    RECT 0 151.550 0.070 151.620 ;
    RECT 0 151.690 0.070 154.000 ;
    LAYER metal4 ;
    RECT 0 0 151.810 1.400 ;
    RECT 0 152.600 151.810 154.000 ;
    RECT 0.000 1.400 1.260 152.600 ;
    RECT 1.540 1.400 2.380 152.600 ;
    RECT 2.660 1.400 3.500 152.600 ;
    RECT 3.780 1.400 4.620 152.600 ;
    RECT 4.900 1.400 5.740 152.600 ;
    RECT 6.020 1.400 6.860 152.600 ;
    RECT 7.140 1.400 7.980 152.600 ;
    RECT 8.260 1.400 9.100 152.600 ;
    RECT 9.380 1.400 10.220 152.600 ;
    RECT 10.500 1.400 11.340 152.600 ;
    RECT 11.620 1.400 12.460 152.600 ;
    RECT 12.740 1.400 13.580 152.600 ;
    RECT 13.860 1.400 14.700 152.600 ;
    RECT 14.980 1.400 15.820 152.600 ;
    RECT 16.100 1.400 16.940 152.600 ;
    RECT 17.220 1.400 18.060 152.600 ;
    RECT 18.340 1.400 19.180 152.600 ;
    RECT 19.460 1.400 20.300 152.600 ;
    RECT 20.580 1.400 21.420 152.600 ;
    RECT 21.700 1.400 22.540 152.600 ;
    RECT 22.820 1.400 23.660 152.600 ;
    RECT 23.940 1.400 24.780 152.600 ;
    RECT 25.060 1.400 25.900 152.600 ;
    RECT 26.180 1.400 27.020 152.600 ;
    RECT 27.300 1.400 28.140 152.600 ;
    RECT 28.420 1.400 29.260 152.600 ;
    RECT 29.540 1.400 30.380 152.600 ;
    RECT 30.660 1.400 31.500 152.600 ;
    RECT 31.780 1.400 32.620 152.600 ;
    RECT 32.900 1.400 33.740 152.600 ;
    RECT 34.020 1.400 34.860 152.600 ;
    RECT 35.140 1.400 35.980 152.600 ;
    RECT 36.260 1.400 37.100 152.600 ;
    RECT 37.380 1.400 38.220 152.600 ;
    RECT 38.500 1.400 39.340 152.600 ;
    RECT 39.620 1.400 40.460 152.600 ;
    RECT 40.740 1.400 41.580 152.600 ;
    RECT 41.860 1.400 42.700 152.600 ;
    RECT 42.980 1.400 43.820 152.600 ;
    RECT 44.100 1.400 44.940 152.600 ;
    RECT 45.220 1.400 46.060 152.600 ;
    RECT 46.340 1.400 47.180 152.600 ;
    RECT 47.460 1.400 48.300 152.600 ;
    RECT 48.580 1.400 49.420 152.600 ;
    RECT 49.700 1.400 50.540 152.600 ;
    RECT 50.820 1.400 51.660 152.600 ;
    RECT 51.940 1.400 52.780 152.600 ;
    RECT 53.060 1.400 53.900 152.600 ;
    RECT 54.180 1.400 55.020 152.600 ;
    RECT 55.300 1.400 56.140 152.600 ;
    RECT 56.420 1.400 57.260 152.600 ;
    RECT 57.540 1.400 58.380 152.600 ;
    RECT 58.660 1.400 59.500 152.600 ;
    RECT 59.780 1.400 60.620 152.600 ;
    RECT 60.900 1.400 61.740 152.600 ;
    RECT 62.020 1.400 62.860 152.600 ;
    RECT 63.140 1.400 63.980 152.600 ;
    RECT 64.260 1.400 65.100 152.600 ;
    RECT 65.380 1.400 66.220 152.600 ;
    RECT 66.500 1.400 67.340 152.600 ;
    RECT 67.620 1.400 68.460 152.600 ;
    RECT 68.740 1.400 69.580 152.600 ;
    RECT 69.860 1.400 70.700 152.600 ;
    RECT 70.980 1.400 71.820 152.600 ;
    RECT 72.100 1.400 72.940 152.600 ;
    RECT 73.220 1.400 74.060 152.600 ;
    RECT 74.340 1.400 75.180 152.600 ;
    RECT 75.460 1.400 76.300 152.600 ;
    RECT 76.580 1.400 77.420 152.600 ;
    RECT 77.700 1.400 78.540 152.600 ;
    RECT 78.820 1.400 79.660 152.600 ;
    RECT 79.940 1.400 80.780 152.600 ;
    RECT 81.060 1.400 81.900 152.600 ;
    RECT 82.180 1.400 83.020 152.600 ;
    RECT 83.300 1.400 84.140 152.600 ;
    RECT 84.420 1.400 85.260 152.600 ;
    RECT 85.540 1.400 86.380 152.600 ;
    RECT 86.660 1.400 87.500 152.600 ;
    RECT 87.780 1.400 88.620 152.600 ;
    RECT 88.900 1.400 89.740 152.600 ;
    RECT 90.020 1.400 90.860 152.600 ;
    RECT 91.140 1.400 91.980 152.600 ;
    RECT 92.260 1.400 93.100 152.600 ;
    RECT 93.380 1.400 94.220 152.600 ;
    RECT 94.500 1.400 95.340 152.600 ;
    RECT 95.620 1.400 96.460 152.600 ;
    RECT 96.740 1.400 97.580 152.600 ;
    RECT 97.860 1.400 98.700 152.600 ;
    RECT 98.980 1.400 99.820 152.600 ;
    RECT 100.100 1.400 100.940 152.600 ;
    RECT 101.220 1.400 102.060 152.600 ;
    RECT 102.340 1.400 103.180 152.600 ;
    RECT 103.460 1.400 104.300 152.600 ;
    RECT 104.580 1.400 105.420 152.600 ;
    RECT 105.700 1.400 106.540 152.600 ;
    RECT 106.820 1.400 107.660 152.600 ;
    RECT 107.940 1.400 108.780 152.600 ;
    RECT 109.060 1.400 109.900 152.600 ;
    RECT 110.180 1.400 111.020 152.600 ;
    RECT 111.300 1.400 112.140 152.600 ;
    RECT 112.420 1.400 113.260 152.600 ;
    RECT 113.540 1.400 114.380 152.600 ;
    RECT 114.660 1.400 115.500 152.600 ;
    RECT 115.780 1.400 116.620 152.600 ;
    RECT 116.900 1.400 117.740 152.600 ;
    RECT 118.020 1.400 118.860 152.600 ;
    RECT 119.140 1.400 119.980 152.600 ;
    RECT 120.260 1.400 121.100 152.600 ;
    RECT 121.380 1.400 122.220 152.600 ;
    RECT 122.500 1.400 123.340 152.600 ;
    RECT 123.620 1.400 124.460 152.600 ;
    RECT 124.740 1.400 125.580 152.600 ;
    RECT 125.860 1.400 126.700 152.600 ;
    RECT 126.980 1.400 127.820 152.600 ;
    RECT 128.100 1.400 128.940 152.600 ;
    RECT 129.220 1.400 130.060 152.600 ;
    RECT 130.340 1.400 131.180 152.600 ;
    RECT 131.460 1.400 132.300 152.600 ;
    RECT 132.580 1.400 133.420 152.600 ;
    RECT 133.700 1.400 134.540 152.600 ;
    RECT 134.820 1.400 135.660 152.600 ;
    RECT 135.940 1.400 136.780 152.600 ;
    RECT 137.060 1.400 137.900 152.600 ;
    RECT 138.180 1.400 139.020 152.600 ;
    RECT 139.300 1.400 140.140 152.600 ;
    RECT 140.420 1.400 141.260 152.600 ;
    RECT 141.540 1.400 142.380 152.600 ;
    RECT 142.660 1.400 143.500 152.600 ;
    RECT 143.780 1.400 144.620 152.600 ;
    RECT 144.900 1.400 145.740 152.600 ;
    RECT 146.020 1.400 146.860 152.600 ;
    RECT 147.140 1.400 147.980 152.600 ;
    RECT 148.260 1.400 149.100 152.600 ;
    RECT 149.380 1.400 150.220 152.600 ;
    RECT 150.500 1.400 151.810 152.600 ;
    LAYER OVERLAP ;
    RECT 0 0 151.810 154.000 ;
  END
END fakeram45_128x256

END LIBRARY
