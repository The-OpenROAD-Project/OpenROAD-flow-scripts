VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_512x8
  FOREIGN fakeram_512x8 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 1.140 BY 133.000 ;
  CLASS BLOCK ;
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.048 0.024 0.072 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.752 0.024 4.776 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.456 0.024 9.480 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.160 0.024 14.184 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.864 0.024 18.888 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.568 0.024 23.592 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 28.272 0.024 28.296 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 32.976 0.024 33.000 ;
    END
  END rd_out[7]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 37.680 0.024 37.704 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 42.384 0.024 42.408 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 47.088 0.024 47.112 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 51.792 0.024 51.816 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 56.496 0.024 56.520 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 61.200 0.024 61.224 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 65.904 0.024 65.928 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 70.608 0.024 70.632 ;
    END
  END wd_in[7]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 75.312 0.024 75.336 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 80.016 0.024 80.040 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 84.720 0.024 84.744 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 89.424 0.024 89.448 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 94.128 0.024 94.152 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 98.832 0.024 98.856 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 103.536 0.024 103.560 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 108.240 0.024 108.264 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 112.944 0.024 112.968 ;
    END
  END addr_in[8]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 117.648 0.024 117.672 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 122.352 0.024 122.376 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 127.056 0.024 127.080 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.048 0.000 1.092 0.096 ;
      RECT 0.048 0.768 1.092 0.864 ;
      RECT 0.048 1.536 1.092 1.632 ;
      RECT 0.048 2.304 1.092 2.400 ;
      RECT 0.048 3.072 1.092 3.168 ;
      RECT 0.048 3.840 1.092 3.936 ;
      RECT 0.048 4.608 1.092 4.704 ;
      RECT 0.048 5.376 1.092 5.472 ;
      RECT 0.048 6.144 1.092 6.240 ;
      RECT 0.048 6.912 1.092 7.008 ;
      RECT 0.048 7.680 1.092 7.776 ;
      RECT 0.048 8.448 1.092 8.544 ;
      RECT 0.048 9.216 1.092 9.312 ;
      RECT 0.048 9.984 1.092 10.080 ;
      RECT 0.048 10.752 1.092 10.848 ;
      RECT 0.048 11.520 1.092 11.616 ;
      RECT 0.048 12.288 1.092 12.384 ;
      RECT 0.048 13.056 1.092 13.152 ;
      RECT 0.048 13.824 1.092 13.920 ;
      RECT 0.048 14.592 1.092 14.688 ;
      RECT 0.048 15.360 1.092 15.456 ;
      RECT 0.048 16.128 1.092 16.224 ;
      RECT 0.048 16.896 1.092 16.992 ;
      RECT 0.048 17.664 1.092 17.760 ;
      RECT 0.048 18.432 1.092 18.528 ;
      RECT 0.048 19.200 1.092 19.296 ;
      RECT 0.048 19.968 1.092 20.064 ;
      RECT 0.048 20.736 1.092 20.832 ;
      RECT 0.048 21.504 1.092 21.600 ;
      RECT 0.048 22.272 1.092 22.368 ;
      RECT 0.048 23.040 1.092 23.136 ;
      RECT 0.048 23.808 1.092 23.904 ;
      RECT 0.048 24.576 1.092 24.672 ;
      RECT 0.048 25.344 1.092 25.440 ;
      RECT 0.048 26.112 1.092 26.208 ;
      RECT 0.048 26.880 1.092 26.976 ;
      RECT 0.048 27.648 1.092 27.744 ;
      RECT 0.048 28.416 1.092 28.512 ;
      RECT 0.048 29.184 1.092 29.280 ;
      RECT 0.048 29.952 1.092 30.048 ;
      RECT 0.048 30.720 1.092 30.816 ;
      RECT 0.048 31.488 1.092 31.584 ;
      RECT 0.048 32.256 1.092 32.352 ;
      RECT 0.048 33.024 1.092 33.120 ;
      RECT 0.048 33.792 1.092 33.888 ;
      RECT 0.048 34.560 1.092 34.656 ;
      RECT 0.048 35.328 1.092 35.424 ;
      RECT 0.048 36.096 1.092 36.192 ;
      RECT 0.048 36.864 1.092 36.960 ;
      RECT 0.048 37.632 1.092 37.728 ;
      RECT 0.048 38.400 1.092 38.496 ;
      RECT 0.048 39.168 1.092 39.264 ;
      RECT 0.048 39.936 1.092 40.032 ;
      RECT 0.048 40.704 1.092 40.800 ;
      RECT 0.048 41.472 1.092 41.568 ;
      RECT 0.048 42.240 1.092 42.336 ;
      RECT 0.048 43.008 1.092 43.104 ;
      RECT 0.048 43.776 1.092 43.872 ;
      RECT 0.048 44.544 1.092 44.640 ;
      RECT 0.048 45.312 1.092 45.408 ;
      RECT 0.048 46.080 1.092 46.176 ;
      RECT 0.048 46.848 1.092 46.944 ;
      RECT 0.048 47.616 1.092 47.712 ;
      RECT 0.048 48.384 1.092 48.480 ;
      RECT 0.048 49.152 1.092 49.248 ;
      RECT 0.048 49.920 1.092 50.016 ;
      RECT 0.048 50.688 1.092 50.784 ;
      RECT 0.048 51.456 1.092 51.552 ;
      RECT 0.048 52.224 1.092 52.320 ;
      RECT 0.048 52.992 1.092 53.088 ;
      RECT 0.048 53.760 1.092 53.856 ;
      RECT 0.048 54.528 1.092 54.624 ;
      RECT 0.048 55.296 1.092 55.392 ;
      RECT 0.048 56.064 1.092 56.160 ;
      RECT 0.048 56.832 1.092 56.928 ;
      RECT 0.048 57.600 1.092 57.696 ;
      RECT 0.048 58.368 1.092 58.464 ;
      RECT 0.048 59.136 1.092 59.232 ;
      RECT 0.048 59.904 1.092 60.000 ;
      RECT 0.048 60.672 1.092 60.768 ;
      RECT 0.048 61.440 1.092 61.536 ;
      RECT 0.048 62.208 1.092 62.304 ;
      RECT 0.048 62.976 1.092 63.072 ;
      RECT 0.048 63.744 1.092 63.840 ;
      RECT 0.048 64.512 1.092 64.608 ;
      RECT 0.048 65.280 1.092 65.376 ;
      RECT 0.048 66.048 1.092 66.144 ;
      RECT 0.048 66.816 1.092 66.912 ;
      RECT 0.048 67.584 1.092 67.680 ;
      RECT 0.048 68.352 1.092 68.448 ;
      RECT 0.048 69.120 1.092 69.216 ;
      RECT 0.048 69.888 1.092 69.984 ;
      RECT 0.048 70.656 1.092 70.752 ;
      RECT 0.048 71.424 1.092 71.520 ;
      RECT 0.048 72.192 1.092 72.288 ;
      RECT 0.048 72.960 1.092 73.056 ;
      RECT 0.048 73.728 1.092 73.824 ;
      RECT 0.048 74.496 1.092 74.592 ;
      RECT 0.048 75.264 1.092 75.360 ;
      RECT 0.048 76.032 1.092 76.128 ;
      RECT 0.048 76.800 1.092 76.896 ;
      RECT 0.048 77.568 1.092 77.664 ;
      RECT 0.048 78.336 1.092 78.432 ;
      RECT 0.048 79.104 1.092 79.200 ;
      RECT 0.048 79.872 1.092 79.968 ;
      RECT 0.048 80.640 1.092 80.736 ;
      RECT 0.048 81.408 1.092 81.504 ;
      RECT 0.048 82.176 1.092 82.272 ;
      RECT 0.048 82.944 1.092 83.040 ;
      RECT 0.048 83.712 1.092 83.808 ;
      RECT 0.048 84.480 1.092 84.576 ;
      RECT 0.048 85.248 1.092 85.344 ;
      RECT 0.048 86.016 1.092 86.112 ;
      RECT 0.048 86.784 1.092 86.880 ;
      RECT 0.048 87.552 1.092 87.648 ;
      RECT 0.048 88.320 1.092 88.416 ;
      RECT 0.048 89.088 1.092 89.184 ;
      RECT 0.048 89.856 1.092 89.952 ;
      RECT 0.048 90.624 1.092 90.720 ;
      RECT 0.048 91.392 1.092 91.488 ;
      RECT 0.048 92.160 1.092 92.256 ;
      RECT 0.048 92.928 1.092 93.024 ;
      RECT 0.048 93.696 1.092 93.792 ;
      RECT 0.048 94.464 1.092 94.560 ;
      RECT 0.048 95.232 1.092 95.328 ;
      RECT 0.048 96.000 1.092 96.096 ;
      RECT 0.048 96.768 1.092 96.864 ;
      RECT 0.048 97.536 1.092 97.632 ;
      RECT 0.048 98.304 1.092 98.400 ;
      RECT 0.048 99.072 1.092 99.168 ;
      RECT 0.048 99.840 1.092 99.936 ;
      RECT 0.048 100.608 1.092 100.704 ;
      RECT 0.048 101.376 1.092 101.472 ;
      RECT 0.048 102.144 1.092 102.240 ;
      RECT 0.048 102.912 1.092 103.008 ;
      RECT 0.048 103.680 1.092 103.776 ;
      RECT 0.048 104.448 1.092 104.544 ;
      RECT 0.048 105.216 1.092 105.312 ;
      RECT 0.048 105.984 1.092 106.080 ;
      RECT 0.048 106.752 1.092 106.848 ;
      RECT 0.048 107.520 1.092 107.616 ;
      RECT 0.048 108.288 1.092 108.384 ;
      RECT 0.048 109.056 1.092 109.152 ;
      RECT 0.048 109.824 1.092 109.920 ;
      RECT 0.048 110.592 1.092 110.688 ;
      RECT 0.048 111.360 1.092 111.456 ;
      RECT 0.048 112.128 1.092 112.224 ;
      RECT 0.048 112.896 1.092 112.992 ;
      RECT 0.048 113.664 1.092 113.760 ;
      RECT 0.048 114.432 1.092 114.528 ;
      RECT 0.048 115.200 1.092 115.296 ;
      RECT 0.048 115.968 1.092 116.064 ;
      RECT 0.048 116.736 1.092 116.832 ;
      RECT 0.048 117.504 1.092 117.600 ;
      RECT 0.048 118.272 1.092 118.368 ;
      RECT 0.048 119.040 1.092 119.136 ;
      RECT 0.048 119.808 1.092 119.904 ;
      RECT 0.048 120.576 1.092 120.672 ;
      RECT 0.048 121.344 1.092 121.440 ;
      RECT 0.048 122.112 1.092 122.208 ;
      RECT 0.048 122.880 1.092 122.976 ;
      RECT 0.048 123.648 1.092 123.744 ;
      RECT 0.048 124.416 1.092 124.512 ;
      RECT 0.048 125.184 1.092 125.280 ;
      RECT 0.048 125.952 1.092 126.048 ;
      RECT 0.048 126.720 1.092 126.816 ;
      RECT 0.048 127.488 1.092 127.584 ;
      RECT 0.048 128.256 1.092 128.352 ;
      RECT 0.048 129.024 1.092 129.120 ;
      RECT 0.048 129.792 1.092 129.888 ;
      RECT 0.048 130.560 1.092 130.656 ;
      RECT 0.048 131.328 1.092 131.424 ;
      RECT 0.048 132.096 1.092 132.192 ;
      RECT 0.048 132.864 1.092 132.960 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.048 0.384 1.092 0.480 ;
      RECT 0.048 1.152 1.092 1.248 ;
      RECT 0.048 1.920 1.092 2.016 ;
      RECT 0.048 2.688 1.092 2.784 ;
      RECT 0.048 3.456 1.092 3.552 ;
      RECT 0.048 4.224 1.092 4.320 ;
      RECT 0.048 4.992 1.092 5.088 ;
      RECT 0.048 5.760 1.092 5.856 ;
      RECT 0.048 6.528 1.092 6.624 ;
      RECT 0.048 7.296 1.092 7.392 ;
      RECT 0.048 8.064 1.092 8.160 ;
      RECT 0.048 8.832 1.092 8.928 ;
      RECT 0.048 9.600 1.092 9.696 ;
      RECT 0.048 10.368 1.092 10.464 ;
      RECT 0.048 11.136 1.092 11.232 ;
      RECT 0.048 11.904 1.092 12.000 ;
      RECT 0.048 12.672 1.092 12.768 ;
      RECT 0.048 13.440 1.092 13.536 ;
      RECT 0.048 14.208 1.092 14.304 ;
      RECT 0.048 14.976 1.092 15.072 ;
      RECT 0.048 15.744 1.092 15.840 ;
      RECT 0.048 16.512 1.092 16.608 ;
      RECT 0.048 17.280 1.092 17.376 ;
      RECT 0.048 18.048 1.092 18.144 ;
      RECT 0.048 18.816 1.092 18.912 ;
      RECT 0.048 19.584 1.092 19.680 ;
      RECT 0.048 20.352 1.092 20.448 ;
      RECT 0.048 21.120 1.092 21.216 ;
      RECT 0.048 21.888 1.092 21.984 ;
      RECT 0.048 22.656 1.092 22.752 ;
      RECT 0.048 23.424 1.092 23.520 ;
      RECT 0.048 24.192 1.092 24.288 ;
      RECT 0.048 24.960 1.092 25.056 ;
      RECT 0.048 25.728 1.092 25.824 ;
      RECT 0.048 26.496 1.092 26.592 ;
      RECT 0.048 27.264 1.092 27.360 ;
      RECT 0.048 28.032 1.092 28.128 ;
      RECT 0.048 28.800 1.092 28.896 ;
      RECT 0.048 29.568 1.092 29.664 ;
      RECT 0.048 30.336 1.092 30.432 ;
      RECT 0.048 31.104 1.092 31.200 ;
      RECT 0.048 31.872 1.092 31.968 ;
      RECT 0.048 32.640 1.092 32.736 ;
      RECT 0.048 33.408 1.092 33.504 ;
      RECT 0.048 34.176 1.092 34.272 ;
      RECT 0.048 34.944 1.092 35.040 ;
      RECT 0.048 35.712 1.092 35.808 ;
      RECT 0.048 36.480 1.092 36.576 ;
      RECT 0.048 37.248 1.092 37.344 ;
      RECT 0.048 38.016 1.092 38.112 ;
      RECT 0.048 38.784 1.092 38.880 ;
      RECT 0.048 39.552 1.092 39.648 ;
      RECT 0.048 40.320 1.092 40.416 ;
      RECT 0.048 41.088 1.092 41.184 ;
      RECT 0.048 41.856 1.092 41.952 ;
      RECT 0.048 42.624 1.092 42.720 ;
      RECT 0.048 43.392 1.092 43.488 ;
      RECT 0.048 44.160 1.092 44.256 ;
      RECT 0.048 44.928 1.092 45.024 ;
      RECT 0.048 45.696 1.092 45.792 ;
      RECT 0.048 46.464 1.092 46.560 ;
      RECT 0.048 47.232 1.092 47.328 ;
      RECT 0.048 48.000 1.092 48.096 ;
      RECT 0.048 48.768 1.092 48.864 ;
      RECT 0.048 49.536 1.092 49.632 ;
      RECT 0.048 50.304 1.092 50.400 ;
      RECT 0.048 51.072 1.092 51.168 ;
      RECT 0.048 51.840 1.092 51.936 ;
      RECT 0.048 52.608 1.092 52.704 ;
      RECT 0.048 53.376 1.092 53.472 ;
      RECT 0.048 54.144 1.092 54.240 ;
      RECT 0.048 54.912 1.092 55.008 ;
      RECT 0.048 55.680 1.092 55.776 ;
      RECT 0.048 56.448 1.092 56.544 ;
      RECT 0.048 57.216 1.092 57.312 ;
      RECT 0.048 57.984 1.092 58.080 ;
      RECT 0.048 58.752 1.092 58.848 ;
      RECT 0.048 59.520 1.092 59.616 ;
      RECT 0.048 60.288 1.092 60.384 ;
      RECT 0.048 61.056 1.092 61.152 ;
      RECT 0.048 61.824 1.092 61.920 ;
      RECT 0.048 62.592 1.092 62.688 ;
      RECT 0.048 63.360 1.092 63.456 ;
      RECT 0.048 64.128 1.092 64.224 ;
      RECT 0.048 64.896 1.092 64.992 ;
      RECT 0.048 65.664 1.092 65.760 ;
      RECT 0.048 66.432 1.092 66.528 ;
      RECT 0.048 67.200 1.092 67.296 ;
      RECT 0.048 67.968 1.092 68.064 ;
      RECT 0.048 68.736 1.092 68.832 ;
      RECT 0.048 69.504 1.092 69.600 ;
      RECT 0.048 70.272 1.092 70.368 ;
      RECT 0.048 71.040 1.092 71.136 ;
      RECT 0.048 71.808 1.092 71.904 ;
      RECT 0.048 72.576 1.092 72.672 ;
      RECT 0.048 73.344 1.092 73.440 ;
      RECT 0.048 74.112 1.092 74.208 ;
      RECT 0.048 74.880 1.092 74.976 ;
      RECT 0.048 75.648 1.092 75.744 ;
      RECT 0.048 76.416 1.092 76.512 ;
      RECT 0.048 77.184 1.092 77.280 ;
      RECT 0.048 77.952 1.092 78.048 ;
      RECT 0.048 78.720 1.092 78.816 ;
      RECT 0.048 79.488 1.092 79.584 ;
      RECT 0.048 80.256 1.092 80.352 ;
      RECT 0.048 81.024 1.092 81.120 ;
      RECT 0.048 81.792 1.092 81.888 ;
      RECT 0.048 82.560 1.092 82.656 ;
      RECT 0.048 83.328 1.092 83.424 ;
      RECT 0.048 84.096 1.092 84.192 ;
      RECT 0.048 84.864 1.092 84.960 ;
      RECT 0.048 85.632 1.092 85.728 ;
      RECT 0.048 86.400 1.092 86.496 ;
      RECT 0.048 87.168 1.092 87.264 ;
      RECT 0.048 87.936 1.092 88.032 ;
      RECT 0.048 88.704 1.092 88.800 ;
      RECT 0.048 89.472 1.092 89.568 ;
      RECT 0.048 90.240 1.092 90.336 ;
      RECT 0.048 91.008 1.092 91.104 ;
      RECT 0.048 91.776 1.092 91.872 ;
      RECT 0.048 92.544 1.092 92.640 ;
      RECT 0.048 93.312 1.092 93.408 ;
      RECT 0.048 94.080 1.092 94.176 ;
      RECT 0.048 94.848 1.092 94.944 ;
      RECT 0.048 95.616 1.092 95.712 ;
      RECT 0.048 96.384 1.092 96.480 ;
      RECT 0.048 97.152 1.092 97.248 ;
      RECT 0.048 97.920 1.092 98.016 ;
      RECT 0.048 98.688 1.092 98.784 ;
      RECT 0.048 99.456 1.092 99.552 ;
      RECT 0.048 100.224 1.092 100.320 ;
      RECT 0.048 100.992 1.092 101.088 ;
      RECT 0.048 101.760 1.092 101.856 ;
      RECT 0.048 102.528 1.092 102.624 ;
      RECT 0.048 103.296 1.092 103.392 ;
      RECT 0.048 104.064 1.092 104.160 ;
      RECT 0.048 104.832 1.092 104.928 ;
      RECT 0.048 105.600 1.092 105.696 ;
      RECT 0.048 106.368 1.092 106.464 ;
      RECT 0.048 107.136 1.092 107.232 ;
      RECT 0.048 107.904 1.092 108.000 ;
      RECT 0.048 108.672 1.092 108.768 ;
      RECT 0.048 109.440 1.092 109.536 ;
      RECT 0.048 110.208 1.092 110.304 ;
      RECT 0.048 110.976 1.092 111.072 ;
      RECT 0.048 111.744 1.092 111.840 ;
      RECT 0.048 112.512 1.092 112.608 ;
      RECT 0.048 113.280 1.092 113.376 ;
      RECT 0.048 114.048 1.092 114.144 ;
      RECT 0.048 114.816 1.092 114.912 ;
      RECT 0.048 115.584 1.092 115.680 ;
      RECT 0.048 116.352 1.092 116.448 ;
      RECT 0.048 117.120 1.092 117.216 ;
      RECT 0.048 117.888 1.092 117.984 ;
      RECT 0.048 118.656 1.092 118.752 ;
      RECT 0.048 119.424 1.092 119.520 ;
      RECT 0.048 120.192 1.092 120.288 ;
      RECT 0.048 120.960 1.092 121.056 ;
      RECT 0.048 121.728 1.092 121.824 ;
      RECT 0.048 122.496 1.092 122.592 ;
      RECT 0.048 123.264 1.092 123.360 ;
      RECT 0.048 124.032 1.092 124.128 ;
      RECT 0.048 124.800 1.092 124.896 ;
      RECT 0.048 125.568 1.092 125.664 ;
      RECT 0.048 126.336 1.092 126.432 ;
      RECT 0.048 127.104 1.092 127.200 ;
      RECT 0.048 127.872 1.092 127.968 ;
      RECT 0.048 128.640 1.092 128.736 ;
      RECT 0.048 129.408 1.092 129.504 ;
      RECT 0.048 130.176 1.092 130.272 ;
      RECT 0.048 130.944 1.092 131.040 ;
      RECT 0.048 131.712 1.092 131.808 ;
      RECT 0.048 132.480 1.092 132.576 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 1.140 133.000 ;
    LAYER M2 ;
    RECT 0 0 1.140 133.000 ;
    LAYER M3 ;
    RECT 0 0 1.140 133.000 ;
    LAYER M4 ;
    RECT 0.1 0 1.040 133.000 ;
  END
END fakeram_512x8

END LIBRARY
