module aes_cipher_top (clk,
    done,
    ld,
    rst,
    key,
    text_in,
    text_out);
 input clk;
 output done;
 input ld;
 input rst;
 input [127:0] key;
 input [127:0] text_in;
 output [127:0] text_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire clknet_leaf_0_clk;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire net754;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire net753;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire net752;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire net751;
 wire _01096_;
 wire _01097_;
 wire net750;
 wire _01099_;
 wire net749;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire net748;
 wire net747;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire net746;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire net745;
 wire _01115_;
 wire net744;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire net743;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire net742;
 wire _01127_;
 wire _01128_;
 wire net741;
 wire net740;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire net739;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire net738;
 wire _01140_;
 wire _01141_;
 wire net737;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire net736;
 wire _01148_;
 wire net735;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire net734;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire net733;
 wire _01162_;
 wire _01163_;
 wire net732;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire net731;
 wire net730;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire net729;
 wire _01190_;
 wire _01191_;
 wire net728;
 wire _01193_;
 wire _01194_;
 wire net727;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire net726;
 wire net725;
 wire _01202_;
 wire net724;
 wire _01204_;
 wire net723;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire net722;
 wire _01220_;
 wire _01221_;
 wire net721;
 wire net720;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire net719;
 wire _01228_;
 wire _01229_;
 wire net718;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire net717;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire net716;
 wire _01248_;
 wire net715;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire net714;
 wire _01259_;
 wire net713;
 wire net712;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire net711;
 wire _01276_;
 wire net710;
 wire _01278_;
 wire _01279_;
 wire net709;
 wire _01281_;
 wire net708;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire net707;
 wire net706;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire net705;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire net704;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire net703;
 wire _01310_;
 wire net702;
 wire net701;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire net700;
 wire net699;
 wire _01321_;
 wire _01322_;
 wire net698;
 wire net697;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire net696;
 wire _01336_;
 wire _01337_;
 wire net695;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire net694;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire net693;
 wire net692;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire net691;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire net690;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire net689;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire net688;
 wire net687;
 wire net686;
 wire _01491_;
 wire net685;
 wire net684;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire net683;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire net682;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire net681;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire net680;
 wire net679;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire net678;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire net677;
 wire net676;
 wire _01543_;
 wire net675;
 wire net674;
 wire net673;
 wire _01547_;
 wire net672;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire net671;
 wire _01555_;
 wire _01556_;
 wire net670;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire net669;
 wire _01567_;
 wire net668;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire net667;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire net666;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire net665;
 wire _01592_;
 wire net664;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire net663;
 wire _01602_;
 wire _01603_;
 wire net662;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire net661;
 wire net660;
 wire _01612_;
 wire net659;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire net658;
 wire _01624_;
 wire net657;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire net656;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire net655;
 wire _01644_;
 wire net654;
 wire net653;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire net652;
 wire net651;
 wire _01652_;
 wire _01653_;
 wire net650;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire net649;
 wire net648;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire net647;
 wire _01667_;
 wire _01668_;
 wire net646;
 wire _01670_;
 wire net645;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire net644;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire net643;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire net642;
 wire _01691_;
 wire net641;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire net640;
 wire _01701_;
 wire net639;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire net638;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire net637;
 wire _01715_;
 wire net636;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire net635;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire net634;
 wire _01727_;
 wire _01728_;
 wire net633;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire net632;
 wire net631;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire net630;
 wire _01756_;
 wire _01757_;
 wire net629;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire net628;
 wire net627;
 wire _01765_;
 wire net626;
 wire net625;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire net624;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire net623;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire net622;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire net621;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire net620;
 wire net619;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire net618;
 wire _01799_;
 wire net617;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire net616;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire net615;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire net614;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire net613;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire net612;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire net611;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire net610;
 wire _01894_;
 wire net609;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire net608;
 wire net607;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire net606;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire net605;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire net604;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire net603;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire net602;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire net601;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire net600;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire net599;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire net598;
 wire _01967_;
 wire net597;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire net596;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire net595;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire net594;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire net593;
 wire _02012_;
 wire _02013_;
 wire net592;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire net591;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire net590;
 wire _02109_;
 wire _02110_;
 wire net589;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire net588;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire net587;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire net586;
 wire net585;
 wire net584;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire net583;
 wire _02157_;
 wire net582;
 wire net581;
 wire _02160_;
 wire net580;
 wire _02162_;
 wire _02163_;
 wire net579;
 wire net578;
 wire net577;
 wire net576;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire net575;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire net574;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire net573;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire net572;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire net571;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire net570;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire net569;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire net568;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire net567;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire net566;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire net565;
 wire _02363_;
 wire net564;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire net563;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire net562;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire net561;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire net560;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire net559;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire net558;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire net557;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire net556;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire net555;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire net554;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire net553;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire net552;
 wire _02652_;
 wire net551;
 wire net550;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire net549;
 wire net548;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire net547;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire net546;
 wire _02701_;
 wire net545;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire net544;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire net543;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire net542;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire net541;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire net540;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire net539;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire net538;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire net537;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire net536;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire net535;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire net534;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire net533;
 wire net532;
 wire net531;
 wire _05056_;
 wire net530;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire net529;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire net528;
 wire _05072_;
 wire _05073_;
 wire net527;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire net526;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire net525;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire net524;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire net523;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire net522;
 wire _05131_;
 wire net521;
 wire net520;
 wire _05134_;
 wire _05135_;
 wire net519;
 wire net518;
 wire _05138_;
 wire net517;
 wire _05140_;
 wire net516;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire net515;
 wire net514;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire net513;
 wire _05165_;
 wire net512;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire net511;
 wire _05188_;
 wire net510;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire net509;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire net508;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire net507;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire net506;
 wire _05258_;
 wire _05259_;
 wire net505;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire net504;
 wire net503;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire net502;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire net501;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire net500;
 wire net499;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire net498;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire net497;
 wire _05362_;
 wire _05363_;
 wire net496;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire net495;
 wire _05407_;
 wire net494;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire net493;
 wire _05432_;
 wire net492;
 wire _05434_;
 wire _05435_;
 wire net491;
 wire net490;
 wire net489;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire net488;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire net487;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire net486;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire net485;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire net484;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire net483;
 wire _05490_;
 wire net482;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire net481;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire net480;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire net479;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire net478;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire net477;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire net476;
 wire _05527_;
 wire _05528_;
 wire net475;
 wire _05530_;
 wire net474;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire net473;
 wire _05537_;
 wire net472;
 wire net471;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire net470;
 wire _05547_;
 wire _05548_;
 wire net469;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire net468;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire net467;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire net466;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire net465;
 wire _05572_;
 wire net464;
 wire net463;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire net462;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire net461;
 wire net460;
 wire net459;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire net458;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire net457;
 wire _05615_;
 wire _05616_;
 wire net456;
 wire _05618_;
 wire _05619_;
 wire net455;
 wire _05621_;
 wire net454;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire net453;
 wire net452;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire net451;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire net450;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire net449;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire net1341;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire net1340;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire net1339;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire net448;
 wire _05734_;
 wire _05735_;
 wire net447;
 wire _05737_;
 wire net1338;
 wire net446;
 wire _05740_;
 wire _05741_;
 wire net445;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire net444;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire net443;
 wire net442;
 wire _05770_;
 wire net1337;
 wire _05772_;
 wire _05773_;
 wire net441;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire net440;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire net439;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire net438;
 wire _05796_;
 wire net437;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire net436;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire net435;
 wire _05807_;
 wire _05808_;
 wire net434;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire net1336;
 wire _05816_;
 wire _05817_;
 wire net433;
 wire _05819_;
 wire net432;
 wire _05821_;
 wire net431;
 wire net430;
 wire _05824_;
 wire _05825_;
 wire net1335;
 wire net429;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire net428;
 wire _05835_;
 wire net427;
 wire net1334;
 wire _05838_;
 wire _05839_;
 wire net426;
 wire _05841_;
 wire net425;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire net424;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire net423;
 wire _05856_;
 wire _05857_;
 wire net422;
 wire _05859_;
 wire _05860_;
 wire net421;
 wire net420;
 wire net419;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire net418;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire net417;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire net416;
 wire _05894_;
 wire net415;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire net414;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire net413;
 wire net412;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire net1333;
 wire _05915_;
 wire _05916_;
 wire net411;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire net410;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire net409;
 wire net408;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire net407;
 wire net406;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire net405;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire net404;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire net403;
 wire net402;
 wire net1332;
 wire _05970_;
 wire _05971_;
 wire net401;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire net1331;
 wire net400;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire net399;
 wire net398;
 wire net397;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire net396;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire net395;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire net394;
 wire net393;
 wire _06029_;
 wire _06030_;
 wire net392;
 wire net391;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire net390;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire net389;
 wire _06052_;
 wire net388;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire net387;
 wire _06061_;
 wire net386;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire net385;
 wire net1330;
 wire net384;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire net383;
 wire net382;
 wire _06075_;
 wire _06076_;
 wire net381;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire net380;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire net379;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire net1329;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire net378;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire net377;
 wire _06118_;
 wire net376;
 wire _06120_;
 wire _06121_;
 wire net375;
 wire _06123_;
 wire net374;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire net373;
 wire _06131_;
 wire net372;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire net371;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire net370;
 wire _06161_;
 wire net369;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire net368;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire net367;
 wire _06203_;
 wire net366;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire net365;
 wire net364;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire net363;
 wire _06226_;
 wire net362;
 wire _06228_;
 wire _06229_;
 wire net361;
 wire _06231_;
 wire net360;
 wire net1328;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire net359;
 wire _06239_;
 wire _06240_;
 wire net358;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire net357;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire net356;
 wire _06266_;
 wire net355;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire net354;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire net353;
 wire _06304_;
 wire net352;
 wire _06306_;
 wire net351;
 wire net350;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire net349;
 wire _06318_;
 wire _06319_;
 wire net1327;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire net348;
 wire _06333_;
 wire _06334_;
 wire net347;
 wire net346;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire net345;
 wire _06341_;
 wire _06342_;
 wire net344;
 wire net343;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire net342;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire net341;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire net340;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire net339;
 wire _06368_;
 wire net338;
 wire _06370_;
 wire net337;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire net336;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire net335;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire net1326;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire net334;
 wire net333;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire net332;
 wire _06411_;
 wire _06412_;
 wire net331;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire net330;
 wire net329;
 wire net328;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire net327;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire net326;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire net1325;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire net325;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire net1324;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire net324;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire net323;
 wire _06576_;
 wire net322;
 wire _06578_;
 wire net321;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire net320;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire net319;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire net318;
 wire _06605_;
 wire _06606_;
 wire net317;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire net316;
 wire _06612_;
 wire _06613_;
 wire net315;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire net314;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire net313;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire net312;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire net1323;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire net1322;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire net311;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire net1321;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire net310;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire net309;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire net308;
 wire _06735_;
 wire _06736_;
 wire net307;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire net306;
 wire net305;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire net304;
 wire net303;
 wire _06760_;
 wire net302;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire net301;
 wire net300;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire net299;
 wire net298;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire net1320;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire net297;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire net296;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire net295;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire net1319;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire net1318;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire net1317;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire net1316;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire net294;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire net1315;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire net1314;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire net293;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire net1313;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire net1312;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire net1311;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire net1310;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire net292;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire net1309;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire net291;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire net290;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire net1308;
 wire _07310_;
 wire net289;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire net1307;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire net288;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire net287;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire net1306;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire net286;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire net1305;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire net1304;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire net1303;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire net1302;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire net1301;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire net1300;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire net1299;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire net1298;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire net1297;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire net1296;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire net1295;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire net1294;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire net1293;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire net1292;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire net1291;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire net1290;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire net1289;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire net1288;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire net1287;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire net1286;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire net1285;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire net1284;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire net1283;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire net1282;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire net1281;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire net1280;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire net1279;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire net285;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire net284;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire net283;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire net282;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire net281;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire net1278;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire net280;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire net279;
 wire net278;
 wire net277;
 wire _09573_;
 wire _09574_;
 wire net276;
 wire net275;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire net274;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire net273;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire net272;
 wire _09599_;
 wire net271;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire net270;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire net269;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire net268;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire net267;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire net266;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire net265;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire net264;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire net263;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire net262;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire net261;
 wire _09674_;
 wire net260;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire net259;
 wire net258;
 wire _09681_;
 wire _09682_;
 wire net257;
 wire _09684_;
 wire net256;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire net255;
 wire _09691_;
 wire _09692_;
 wire net254;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire net253;
 wire _09700_;
 wire _09701_;
 wire net252;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire net251;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire net250;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire net249;
 wire net248;
 wire _09730_;
 wire _09731_;
 wire net247;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire net246;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire net245;
 wire _09772_;
 wire _09773_;
 wire net244;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire net243;
 wire net242;
 wire net241;
 wire net240;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire net239;
 wire _09797_;
 wire _09798_;
 wire net238;
 wire net237;
 wire _09801_;
 wire net236;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire net235;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire net234;
 wire _09819_;
 wire net233;
 wire _09821_;
 wire _09822_;
 wire net232;
 wire net231;
 wire _09825_;
 wire _09826_;
 wire net230;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire net229;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire net228;
 wire _09841_;
 wire net227;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire net226;
 wire net225;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire net224;
 wire net223;
 wire _09870_;
 wire _09871_;
 wire net222;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire net221;
 wire _09878_;
 wire net220;
 wire net219;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire net218;
 wire _09892_;
 wire _09893_;
 wire net217;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire net216;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire net215;
 wire _09925_;
 wire _09926_;
 wire net214;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire net213;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire net212;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire net211;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire net210;
 wire net209;
 wire net208;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire net207;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire net206;
 wire _09998_;
 wire net205;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire net1277;
 wire _10018_;
 wire net204;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire net203;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire net202;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire net201;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire net200;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire net199;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire net198;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire net1276;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire net197;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire net1275;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire net196;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire net195;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire net194;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire net193;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire net192;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire net191;
 wire net190;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire net189;
 wire _10207_;
 wire net188;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire net187;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire net186;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire net1274;
 wire net185;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire net184;
 wire net183;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire net1273;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire net182;
 wire _10244_;
 wire net181;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire net180;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire net179;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire net178;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire net177;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire net176;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire net175;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire net174;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire net173;
 wire net172;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire net171;
 wire net170;
 wire _10332_;
 wire _10333_;
 wire net169;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire net168;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire net167;
 wire _10345_;
 wire _10346_;
 wire net166;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire net165;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire net164;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire net163;
 wire _10372_;
 wire net162;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire net161;
 wire _10387_;
 wire net160;
 wire _10389_;
 wire _10390_;
 wire net159;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire net158;
 wire _10396_;
 wire net157;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire net156;
 wire _10410_;
 wire net155;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire net154;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire net153;
 wire net152;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire net151;
 wire net150;
 wire _10434_;
 wire _10435_;
 wire net149;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire net148;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire net147;
 wire _10451_;
 wire net146;
 wire _10453_;
 wire _10454_;
 wire net145;
 wire _10456_;
 wire net144;
 wire _10458_;
 wire _10459_;
 wire net143;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire net142;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire net141;
 wire _10470_;
 wire _10471_;
 wire net140;
 wire _10473_;
 wire net139;
 wire net138;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire net137;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire net136;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire net135;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire net134;
 wire _10504_;
 wire _10505_;
 wire net133;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire net132;
 wire net131;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire net130;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire net129;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire net128;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire net127;
 wire net126;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire net125;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire net124;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire net123;
 wire _10604_;
 wire _10605_;
 wire net122;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire net121;
 wire net120;
 wire _10618_;
 wire net119;
 wire net118;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire net117;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire net116;
 wire net115;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire net114;
 wire net113;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire net112;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire net111;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire net110;
 wire _10656_;
 wire net109;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire net108;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire net107;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire net106;
 wire _10671_;
 wire _10672_;
 wire net105;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire net104;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire net103;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire net102;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire net101;
 wire _10717_;
 wire net100;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire net99;
 wire net98;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire net97;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire net96;
 wire _10759_;
 wire net95;
 wire net94;
 wire _10762_;
 wire net93;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire net92;
 wire _10796_;
 wire _10797_;
 wire net91;
 wire _10799_;
 wire net90;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire net89;
 wire _10818_;
 wire _10819_;
 wire net88;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire net87;
 wire _10834_;
 wire _10835_;
 wire net86;
 wire net85;
 wire net84;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire net83;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire net82;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire net81;
 wire net80;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire net79;
 wire _10908_;
 wire _10909_;
 wire net78;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire net77;
 wire _10921_;
 wire net76;
 wire _10923_;
 wire net75;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire net74;
 wire _10932_;
 wire net73;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire net72;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire net71;
 wire net70;
 wire net69;
 wire _10950_;
 wire net68;
 wire _10952_;
 wire _10953_;
 wire net67;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire net66;
 wire _10961_;
 wire _10962_;
 wire net65;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire net64;
 wire _10971_;
 wire _10972_;
 wire net63;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire net62;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire net61;
 wire _11030_;
 wire net60;
 wire _11032_;
 wire _11033_;
 wire net59;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire net58;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire net57;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire net56;
 wire net55;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire net54;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire net53;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire net52;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire net51;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire net50;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire net49;
 wire net48;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire net1272;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire net47;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire net46;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire net45;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire net1271;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire net1270;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire net44;
 wire _11300_;
 wire _11301_;
 wire net1269;
 wire _11303_;
 wire _11304_;
 wire net43;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire net42;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire net41;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire net40;
 wire _11323_;
 wire net39;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire net38;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire net37;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire net36;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire net35;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire net1268;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire net34;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire net33;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire net32;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire net31;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire net30;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire net29;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire net1267;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire net1266;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire net1265;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire net1264;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire net1263;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire net1262;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire net1261;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire net28;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire net27;
 wire net1260;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire net26;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire net25;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire net1259;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire net24;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire net23;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire net22;
 wire net21;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire net20;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire net19;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire net18;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire net17;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire net16;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire net15;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire net14;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire net13;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire net12;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire net11;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire net10;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire net9;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire net8;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire net7;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire net6;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire net5;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire net4;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire net3;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire net2;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire net1;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire net1258;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire net1257;
 wire net1256;
 wire net1255;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire net1254;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire net1253;
 wire net1252;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire net1251;
 wire _14678_;
 wire net1250;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire net1249;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire net1248;
 wire _14694_;
 wire net1247;
 wire _14696_;
 wire net1246;
 wire net1245;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire net1244;
 wire _14708_;
 wire _14709_;
 wire net1243;
 wire net1242;
 wire _14712_;
 wire net1241;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire net1240;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire net1239;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire net1238;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire net1237;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire net1236;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire net1235;
 wire _14766_;
 wire net1234;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire net1233;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire net1232;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire net1231;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire net1230;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire net1229;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire net1228;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire net1227;
 wire net1226;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire net1225;
 wire net1224;
 wire _14850_;
 wire net1223;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire net1222;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire net1221;
 wire _14865_;
 wire net1220;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire net1219;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire net1218;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire net1217;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire net1216;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire net1215;
 wire net1214;
 wire _14943_;
 wire net1213;
 wire _14945_;
 wire _14946_;
 wire net1212;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire net1211;
 wire _14961_;
 wire net1210;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire net1209;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire net1208;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire net1207;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire net1206;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire net1205;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire _15104_;
 wire _15105_;
 wire _15106_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire _15123_;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire net1204;
 wire _15139_;
 wire net1203;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15168_;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire _15173_;
 wire _15174_;
 wire _15175_;
 wire _15176_;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15186_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire _15200_;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire net1202;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire net1201;
 wire _15270_;
 wire net1200;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire net1199;
 wire _15277_;
 wire _15278_;
 wire _15279_;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire net1198;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15353_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire net1197;
 wire net1196;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire _15403_;
 wire _15404_;
 wire net1195;
 wire _15406_;
 wire net1194;
 wire _15408_;
 wire _15409_;
 wire _15410_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire _15418_;
 wire _15419_;
 wire _15420_;
 wire _15421_;
 wire _15422_;
 wire _15423_;
 wire _15424_;
 wire _15425_;
 wire net1193;
 wire _15427_;
 wire _15428_;
 wire _15429_;
 wire net1192;
 wire _15431_;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire _15436_;
 wire _15437_;
 wire net1191;
 wire _15439_;
 wire _15440_;
 wire _15441_;
 wire _15442_;
 wire _15443_;
 wire _15444_;
 wire _15445_;
 wire net1190;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire _15460_;
 wire net1189;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire _15468_;
 wire _15469_;
 wire net1188;
 wire net1187;
 wire _15472_;
 wire _15473_;
 wire net1186;
 wire _15475_;
 wire _15476_;
 wire net1185;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire net1184;
 wire _15486_;
 wire net1183;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire net1182;
 wire _15492_;
 wire _15493_;
 wire net1181;
 wire _15495_;
 wire _15496_;
 wire net1180;
 wire _15498_;
 wire _15499_;
 wire net1179;
 wire _15501_;
 wire _15502_;
 wire _15503_;
 wire _15504_;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire _15508_;
 wire _15509_;
 wire _15510_;
 wire net1178;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire _15519_;
 wire _15520_;
 wire net1177;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire _15537_;
 wire _15538_;
 wire _15539_;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire _15543_;
 wire _15544_;
 wire net1176;
 wire _15546_;
 wire net1175;
 wire _15548_;
 wire _15549_;
 wire _15550_;
 wire net1174;
 wire _15552_;
 wire net1173;
 wire _15554_;
 wire _15555_;
 wire net1172;
 wire _15557_;
 wire net1171;
 wire _15559_;
 wire _15560_;
 wire _15561_;
 wire _15562_;
 wire _15563_;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire _15568_;
 wire _15569_;
 wire _15570_;
 wire _15571_;
 wire _15572_;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire _15576_;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire _15583_;
 wire _15584_;
 wire net1170;
 wire net1169;
 wire net1168;
 wire _15588_;
 wire _15589_;
 wire _15590_;
 wire _15591_;
 wire _15592_;
 wire _15593_;
 wire _15594_;
 wire _15595_;
 wire _15596_;
 wire _15597_;
 wire _15598_;
 wire _15599_;
 wire _15600_;
 wire net1167;
 wire _15602_;
 wire _15603_;
 wire _15604_;
 wire net1166;
 wire _15606_;
 wire _15607_;
 wire _15608_;
 wire _15609_;
 wire net1165;
 wire _15611_;
 wire _15612_;
 wire _15613_;
 wire _15614_;
 wire _15615_;
 wire net1164;
 wire _15617_;
 wire _15618_;
 wire net1163;
 wire _15620_;
 wire _15621_;
 wire net1162;
 wire _15623_;
 wire _15624_;
 wire _15625_;
 wire _15626_;
 wire _15627_;
 wire _15628_;
 wire _15629_;
 wire _15630_;
 wire _15631_;
 wire _15632_;
 wire _15633_;
 wire net1161;
 wire _15635_;
 wire net1160;
 wire _15637_;
 wire _15638_;
 wire _15639_;
 wire _15640_;
 wire _15641_;
 wire net1159;
 wire net1158;
 wire _15644_;
 wire _15645_;
 wire _15646_;
 wire _15647_;
 wire _15648_;
 wire _15649_;
 wire _15650_;
 wire _15651_;
 wire _15652_;
 wire _15653_;
 wire _15654_;
 wire _15655_;
 wire _15656_;
 wire _15657_;
 wire net1157;
 wire net1156;
 wire _15660_;
 wire _15661_;
 wire _15662_;
 wire _15663_;
 wire _15664_;
 wire _15665_;
 wire _15666_;
 wire _15667_;
 wire _15668_;
 wire _15669_;
 wire _15670_;
 wire _15671_;
 wire _15672_;
 wire _15673_;
 wire _15674_;
 wire _15675_;
 wire _15676_;
 wire _15677_;
 wire _15678_;
 wire _15679_;
 wire _15680_;
 wire _15681_;
 wire net1155;
 wire _15683_;
 wire _15684_;
 wire _15685_;
 wire _15686_;
 wire _15687_;
 wire net1154;
 wire _15689_;
 wire _15690_;
 wire _15691_;
 wire _15692_;
 wire _15693_;
 wire _15694_;
 wire _15695_;
 wire net1153;
 wire _15697_;
 wire _15698_;
 wire _15699_;
 wire net1152;
 wire _15701_;
 wire _15702_;
 wire _15703_;
 wire _15704_;
 wire net1151;
 wire _15706_;
 wire _15707_;
 wire _15708_;
 wire _15709_;
 wire _15710_;
 wire _15711_;
 wire _15712_;
 wire _15713_;
 wire net1150;
 wire net1149;
 wire _15716_;
 wire _15717_;
 wire _15718_;
 wire _15719_;
 wire _15720_;
 wire _15721_;
 wire _15722_;
 wire _15723_;
 wire _15724_;
 wire _15725_;
 wire _15726_;
 wire _15727_;
 wire _15728_;
 wire _15729_;
 wire _15730_;
 wire _15731_;
 wire _15732_;
 wire _15733_;
 wire _15734_;
 wire _15735_;
 wire _15736_;
 wire _15737_;
 wire _15738_;
 wire _15739_;
 wire _15740_;
 wire _15741_;
 wire _15742_;
 wire _15743_;
 wire _15744_;
 wire _15745_;
 wire _15746_;
 wire _15747_;
 wire _15748_;
 wire _15749_;
 wire _15750_;
 wire _15751_;
 wire _15752_;
 wire _15753_;
 wire _15754_;
 wire _15755_;
 wire _15756_;
 wire _15757_;
 wire _15758_;
 wire _15759_;
 wire _15760_;
 wire _15761_;
 wire _15762_;
 wire _15763_;
 wire _15764_;
 wire _15765_;
 wire _15766_;
 wire _15767_;
 wire _15768_;
 wire _15769_;
 wire _15770_;
 wire _15771_;
 wire _15772_;
 wire net1148;
 wire _15774_;
 wire net1147;
 wire _15776_;
 wire _15777_;
 wire _15778_;
 wire _15779_;
 wire _15780_;
 wire net1146;
 wire net1145;
 wire _15783_;
 wire _15784_;
 wire _15785_;
 wire net1144;
 wire _15787_;
 wire _15788_;
 wire _15789_;
 wire _15790_;
 wire _15791_;
 wire _15792_;
 wire _15793_;
 wire _15794_;
 wire _15795_;
 wire _15796_;
 wire _15797_;
 wire _15798_;
 wire _15799_;
 wire _15800_;
 wire _15801_;
 wire _15802_;
 wire _15803_;
 wire _15804_;
 wire _15805_;
 wire _15806_;
 wire _15807_;
 wire _15808_;
 wire _15809_;
 wire _15810_;
 wire _15811_;
 wire _15812_;
 wire _15813_;
 wire _15814_;
 wire _15815_;
 wire _15816_;
 wire _15817_;
 wire _15818_;
 wire _15819_;
 wire _15820_;
 wire _15821_;
 wire _15822_;
 wire _15823_;
 wire _15824_;
 wire _15825_;
 wire _15826_;
 wire _15827_;
 wire _15828_;
 wire _15829_;
 wire _15830_;
 wire _15831_;
 wire _15832_;
 wire _15833_;
 wire _15834_;
 wire _15835_;
 wire _15836_;
 wire _15837_;
 wire _15838_;
 wire _15839_;
 wire _15840_;
 wire _15841_;
 wire _15842_;
 wire _15843_;
 wire _15844_;
 wire _15845_;
 wire _15846_;
 wire _15847_;
 wire _15848_;
 wire _15849_;
 wire _15850_;
 wire _15851_;
 wire _15852_;
 wire _15853_;
 wire _15854_;
 wire _15855_;
 wire _15856_;
 wire _15857_;
 wire _15858_;
 wire _15859_;
 wire _15860_;
 wire _15861_;
 wire _15862_;
 wire _15863_;
 wire _15864_;
 wire _15865_;
 wire _15866_;
 wire _15867_;
 wire _15868_;
 wire _15869_;
 wire _15870_;
 wire _15871_;
 wire _15872_;
 wire _15873_;
 wire _15874_;
 wire _15875_;
 wire _15876_;
 wire _15877_;
 wire _15878_;
 wire _15879_;
 wire _15880_;
 wire _15881_;
 wire _15882_;
 wire _15883_;
 wire _15884_;
 wire _15885_;
 wire _15886_;
 wire _15887_;
 wire _15888_;
 wire _15889_;
 wire _15890_;
 wire _15891_;
 wire _15892_;
 wire _15893_;
 wire _15894_;
 wire _15895_;
 wire _15896_;
 wire _15897_;
 wire _15898_;
 wire _15899_;
 wire _15900_;
 wire _15901_;
 wire net1143;
 wire _15903_;
 wire _15904_;
 wire _15905_;
 wire _15906_;
 wire _15907_;
 wire _15908_;
 wire _15909_;
 wire _15910_;
 wire _15911_;
 wire _15912_;
 wire _15913_;
 wire _15914_;
 wire _15915_;
 wire _15916_;
 wire net1142;
 wire _15918_;
 wire _15919_;
 wire _15920_;
 wire _15921_;
 wire _15922_;
 wire _15923_;
 wire _15924_;
 wire _15925_;
 wire _15926_;
 wire _15927_;
 wire _15928_;
 wire _15929_;
 wire _15930_;
 wire _15931_;
 wire _15932_;
 wire _15933_;
 wire _15934_;
 wire _15935_;
 wire _15936_;
 wire _15937_;
 wire _15938_;
 wire _15939_;
 wire _15940_;
 wire _15941_;
 wire _15942_;
 wire _15943_;
 wire _15944_;
 wire _15945_;
 wire _15946_;
 wire _15947_;
 wire _15948_;
 wire _15949_;
 wire _15950_;
 wire _15951_;
 wire _15952_;
 wire _15953_;
 wire _15954_;
 wire _15955_;
 wire _15956_;
 wire _15957_;
 wire _15958_;
 wire _15959_;
 wire _15960_;
 wire _15961_;
 wire _15962_;
 wire _15963_;
 wire _15964_;
 wire _15965_;
 wire _15966_;
 wire _15967_;
 wire _15968_;
 wire _15969_;
 wire _15970_;
 wire _15971_;
 wire _15972_;
 wire _15973_;
 wire _15974_;
 wire _15975_;
 wire _15976_;
 wire _15977_;
 wire _15978_;
 wire _15979_;
 wire _15980_;
 wire net1141;
 wire _15982_;
 wire net1140;
 wire _15984_;
 wire _15985_;
 wire _15986_;
 wire _15987_;
 wire _15988_;
 wire _15989_;
 wire _15990_;
 wire _15991_;
 wire _15992_;
 wire _15993_;
 wire _15994_;
 wire _15995_;
 wire _15996_;
 wire _15997_;
 wire _15998_;
 wire _15999_;
 wire _16000_;
 wire _16001_;
 wire _16002_;
 wire _16003_;
 wire _16004_;
 wire _16005_;
 wire _16006_;
 wire _16007_;
 wire _16008_;
 wire _16009_;
 wire _16010_;
 wire _16011_;
 wire _16012_;
 wire _16013_;
 wire _16014_;
 wire _16015_;
 wire _16016_;
 wire _16017_;
 wire _16018_;
 wire _16019_;
 wire _16020_;
 wire _16021_;
 wire _16022_;
 wire _16023_;
 wire _16024_;
 wire _16025_;
 wire _16026_;
 wire _16027_;
 wire _16028_;
 wire _16029_;
 wire _16030_;
 wire _16031_;
 wire _16032_;
 wire _16033_;
 wire _16034_;
 wire _16035_;
 wire _16036_;
 wire _16037_;
 wire _16038_;
 wire _16039_;
 wire _16040_;
 wire _16041_;
 wire _16042_;
 wire _16043_;
 wire _16044_;
 wire _16045_;
 wire _16046_;
 wire _16047_;
 wire _16048_;
 wire _16049_;
 wire _16050_;
 wire net1139;
 wire _16052_;
 wire _16053_;
 wire _16054_;
 wire _16055_;
 wire _16056_;
 wire net1138;
 wire net1137;
 wire _16059_;
 wire _16060_;
 wire _16061_;
 wire _16062_;
 wire _16063_;
 wire _16064_;
 wire _16065_;
 wire _16066_;
 wire _16067_;
 wire _16068_;
 wire _16069_;
 wire _16070_;
 wire _16071_;
 wire _16072_;
 wire _16073_;
 wire _16074_;
 wire _16075_;
 wire _16076_;
 wire _16077_;
 wire _16078_;
 wire _16079_;
 wire _16080_;
 wire _16081_;
 wire _16082_;
 wire _16083_;
 wire _16084_;
 wire _16085_;
 wire _16086_;
 wire _16087_;
 wire _16088_;
 wire _16089_;
 wire _16090_;
 wire _16091_;
 wire _16092_;
 wire _16093_;
 wire _16094_;
 wire _16095_;
 wire _16096_;
 wire _16097_;
 wire _16098_;
 wire _16099_;
 wire _16100_;
 wire _16101_;
 wire _16102_;
 wire _16103_;
 wire _16104_;
 wire _16105_;
 wire _16106_;
 wire _16107_;
 wire _16108_;
 wire _16109_;
 wire _16110_;
 wire _16111_;
 wire _16112_;
 wire _16113_;
 wire _16114_;
 wire _16115_;
 wire _16116_;
 wire _16117_;
 wire _16118_;
 wire _16119_;
 wire _16120_;
 wire _16121_;
 wire _16122_;
 wire _16123_;
 wire _16124_;
 wire _16125_;
 wire _16126_;
 wire _16127_;
 wire net1136;
 wire _16129_;
 wire _16130_;
 wire _16131_;
 wire _16132_;
 wire _16133_;
 wire _16134_;
 wire _16135_;
 wire _16136_;
 wire _16137_;
 wire _16138_;
 wire _16139_;
 wire _16140_;
 wire _16141_;
 wire _16142_;
 wire _16143_;
 wire _16144_;
 wire _16145_;
 wire _16146_;
 wire _16147_;
 wire _16148_;
 wire _16149_;
 wire _16150_;
 wire _16151_;
 wire _16152_;
 wire _16153_;
 wire _16154_;
 wire _16155_;
 wire _16156_;
 wire _16157_;
 wire _16158_;
 wire _16159_;
 wire _16160_;
 wire _16161_;
 wire _16162_;
 wire _16163_;
 wire _16164_;
 wire _16165_;
 wire _16166_;
 wire _16167_;
 wire _16168_;
 wire _16169_;
 wire _16170_;
 wire _16171_;
 wire _16172_;
 wire _16173_;
 wire _16174_;
 wire _16175_;
 wire _16176_;
 wire _16177_;
 wire _16178_;
 wire _16179_;
 wire _16180_;
 wire _16181_;
 wire _16182_;
 wire _16183_;
 wire _16184_;
 wire _16185_;
 wire _16186_;
 wire _16187_;
 wire _16188_;
 wire _16189_;
 wire _16190_;
 wire _16191_;
 wire _16192_;
 wire _16193_;
 wire _16194_;
 wire _16195_;
 wire _16196_;
 wire _16197_;
 wire _16198_;
 wire _16199_;
 wire _16200_;
 wire _16201_;
 wire _16202_;
 wire _16203_;
 wire _16204_;
 wire _16205_;
 wire _16206_;
 wire _16207_;
 wire _16208_;
 wire _16209_;
 wire _16210_;
 wire _16211_;
 wire _16212_;
 wire _16213_;
 wire _16214_;
 wire _16215_;
 wire _16216_;
 wire _16217_;
 wire _16218_;
 wire _16219_;
 wire _16220_;
 wire _16221_;
 wire _16222_;
 wire _16223_;
 wire _16224_;
 wire _16225_;
 wire _16226_;
 wire _16227_;
 wire _16228_;
 wire _16229_;
 wire _16230_;
 wire _16231_;
 wire _16232_;
 wire _16233_;
 wire _16234_;
 wire _16235_;
 wire _16236_;
 wire _16237_;
 wire _16238_;
 wire _16239_;
 wire _16240_;
 wire _16241_;
 wire _16242_;
 wire _16243_;
 wire _16244_;
 wire _16245_;
 wire _16246_;
 wire _16247_;
 wire _16248_;
 wire _16249_;
 wire _16250_;
 wire _16251_;
 wire net1135;
 wire _16253_;
 wire _16254_;
 wire _16255_;
 wire _16256_;
 wire _16257_;
 wire _16258_;
 wire _16259_;
 wire _16260_;
 wire _16261_;
 wire _16262_;
 wire _16263_;
 wire net1134;
 wire _16265_;
 wire _16266_;
 wire _16267_;
 wire _16268_;
 wire _16269_;
 wire _16270_;
 wire _16271_;
 wire _16272_;
 wire _16273_;
 wire _16274_;
 wire _16275_;
 wire _16276_;
 wire _16277_;
 wire _16278_;
 wire _16279_;
 wire net1133;
 wire _16281_;
 wire _16282_;
 wire _16283_;
 wire _16284_;
 wire _16285_;
 wire _16286_;
 wire _16287_;
 wire _16288_;
 wire _16289_;
 wire _16290_;
 wire _16291_;
 wire _16292_;
 wire _16293_;
 wire _16294_;
 wire _16295_;
 wire _16296_;
 wire net1132;
 wire _16298_;
 wire _16299_;
 wire _16300_;
 wire _16301_;
 wire _16302_;
 wire _16303_;
 wire _16304_;
 wire net1131;
 wire _16306_;
 wire net1130;
 wire _16308_;
 wire _16309_;
 wire net1129;
 wire _16311_;
 wire _16312_;
 wire _16313_;
 wire _16314_;
 wire _16315_;
 wire _16316_;
 wire _16317_;
 wire _16318_;
 wire _16319_;
 wire net1128;
 wire _16321_;
 wire _16322_;
 wire _16323_;
 wire _16324_;
 wire _16325_;
 wire net1127;
 wire _16327_;
 wire net1126;
 wire _16329_;
 wire _16330_;
 wire net1125;
 wire _16332_;
 wire _16333_;
 wire _16334_;
 wire _16335_;
 wire _16336_;
 wire _16337_;
 wire _16338_;
 wire _16339_;
 wire _16340_;
 wire _16341_;
 wire _16342_;
 wire net1124;
 wire _16344_;
 wire _16345_;
 wire _16346_;
 wire _16347_;
 wire _16348_;
 wire _16349_;
 wire _16350_;
 wire _16351_;
 wire _16352_;
 wire _16353_;
 wire _16354_;
 wire net1123;
 wire _16356_;
 wire _16357_;
 wire net1122;
 wire net1121;
 wire _16360_;
 wire _16361_;
 wire _16362_;
 wire _16363_;
 wire _16364_;
 wire net1120;
 wire _16366_;
 wire net1119;
 wire _16368_;
 wire _16369_;
 wire _16370_;
 wire _16371_;
 wire _16372_;
 wire _16373_;
 wire _16374_;
 wire _16375_;
 wire _16376_;
 wire _16377_;
 wire _16378_;
 wire net1118;
 wire _16380_;
 wire _16381_;
 wire _16382_;
 wire _16383_;
 wire _16384_;
 wire _16385_;
 wire _16386_;
 wire _16387_;
 wire net1117;
 wire net1116;
 wire _16390_;
 wire _16391_;
 wire net1115;
 wire _16393_;
 wire _16394_;
 wire _16395_;
 wire net1114;
 wire _16397_;
 wire _16398_;
 wire net1113;
 wire _16400_;
 wire net1112;
 wire _16402_;
 wire _16403_;
 wire _16404_;
 wire _16405_;
 wire _16406_;
 wire _16407_;
 wire _16408_;
 wire _16409_;
 wire net1111;
 wire _16411_;
 wire net1110;
 wire _16413_;
 wire _16414_;
 wire _16415_;
 wire _16416_;
 wire _16417_;
 wire _16418_;
 wire _16419_;
 wire _16420_;
 wire _16421_;
 wire net1109;
 wire _16423_;
 wire _16424_;
 wire _16425_;
 wire _16426_;
 wire _16427_;
 wire _16428_;
 wire _16429_;
 wire _16430_;
 wire _16431_;
 wire _16432_;
 wire _16433_;
 wire _16434_;
 wire _16435_;
 wire _16436_;
 wire _16437_;
 wire net1108;
 wire _16439_;
 wire _16440_;
 wire net1107;
 wire net1106;
 wire _16443_;
 wire _16444_;
 wire _16445_;
 wire _16446_;
 wire _16447_;
 wire _16448_;
 wire _16449_;
 wire _16450_;
 wire _16451_;
 wire _16452_;
 wire net1105;
 wire _16454_;
 wire _16455_;
 wire _16456_;
 wire _16457_;
 wire _16458_;
 wire _16459_;
 wire _16460_;
 wire net1104;
 wire _16462_;
 wire _16463_;
 wire net1103;
 wire _16465_;
 wire _16466_;
 wire _16467_;
 wire net1102;
 wire _16469_;
 wire net1101;
 wire _16471_;
 wire _16472_;
 wire _16473_;
 wire _16474_;
 wire net1100;
 wire _16476_;
 wire _16477_;
 wire net1099;
 wire _16479_;
 wire _16480_;
 wire _16481_;
 wire _16482_;
 wire _16483_;
 wire _16484_;
 wire _16485_;
 wire _16486_;
 wire _16487_;
 wire _16488_;
 wire net1098;
 wire _16490_;
 wire _16491_;
 wire net1097;
 wire _16493_;
 wire _16494_;
 wire _16495_;
 wire net1096;
 wire _16497_;
 wire net1095;
 wire _16499_;
 wire _16500_;
 wire _16501_;
 wire net1094;
 wire _16503_;
 wire _16504_;
 wire _16505_;
 wire _16506_;
 wire _16507_;
 wire _16508_;
 wire _16509_;
 wire _16510_;
 wire _16511_;
 wire _16512_;
 wire _16513_;
 wire _16514_;
 wire _16515_;
 wire _16516_;
 wire _16517_;
 wire _16518_;
 wire _16519_;
 wire _16520_;
 wire _16521_;
 wire _16522_;
 wire _16523_;
 wire _16524_;
 wire _16525_;
 wire _16526_;
 wire _16527_;
 wire net1093;
 wire _16529_;
 wire _16530_;
 wire _16531_;
 wire _16532_;
 wire _16533_;
 wire _16534_;
 wire _16535_;
 wire _16536_;
 wire _16537_;
 wire _16538_;
 wire _16539_;
 wire _16540_;
 wire _16541_;
 wire _16542_;
 wire net1092;
 wire _16544_;
 wire _16545_;
 wire _16546_;
 wire _16547_;
 wire _16548_;
 wire _16549_;
 wire _16550_;
 wire _16551_;
 wire net1091;
 wire _16553_;
 wire _16554_;
 wire _16555_;
 wire _16556_;
 wire _16557_;
 wire _16558_;
 wire _16559_;
 wire _16560_;
 wire _16561_;
 wire net1090;
 wire _16563_;
 wire net1089;
 wire _16565_;
 wire _16566_;
 wire _16567_;
 wire _16568_;
 wire _16569_;
 wire _16570_;
 wire _16571_;
 wire net1088;
 wire _16573_;
 wire _16574_;
 wire _16575_;
 wire _16576_;
 wire _16577_;
 wire _16578_;
 wire _16579_;
 wire _16580_;
 wire _16581_;
 wire _16582_;
 wire _16583_;
 wire _16584_;
 wire _16585_;
 wire _16586_;
 wire _16587_;
 wire _16588_;
 wire _16589_;
 wire _16590_;
 wire _16591_;
 wire _16592_;
 wire _16593_;
 wire net1087;
 wire _16595_;
 wire _16596_;
 wire _16597_;
 wire _16598_;
 wire _16599_;
 wire _16600_;
 wire _16601_;
 wire _16602_;
 wire _16603_;
 wire _16604_;
 wire _16605_;
 wire _16606_;
 wire _16607_;
 wire net1086;
 wire _16609_;
 wire _16610_;
 wire _16611_;
 wire _16612_;
 wire _16613_;
 wire _16614_;
 wire _16615_;
 wire _16616_;
 wire _16617_;
 wire _16618_;
 wire _16619_;
 wire _16620_;
 wire _16621_;
 wire _16622_;
 wire _16623_;
 wire _16624_;
 wire _16625_;
 wire _16626_;
 wire _16627_;
 wire _16628_;
 wire _16629_;
 wire _16630_;
 wire _16631_;
 wire _16632_;
 wire _16633_;
 wire _16634_;
 wire _16635_;
 wire _16636_;
 wire _16637_;
 wire _16638_;
 wire net1085;
 wire _16640_;
 wire _16641_;
 wire _16642_;
 wire _16643_;
 wire _16644_;
 wire _16645_;
 wire _16646_;
 wire _16647_;
 wire net1084;
 wire _16649_;
 wire net1083;
 wire net1082;
 wire _16652_;
 wire _16653_;
 wire _16654_;
 wire _16655_;
 wire _16656_;
 wire _16657_;
 wire _16658_;
 wire _16659_;
 wire _16660_;
 wire _16661_;
 wire _16662_;
 wire _16663_;
 wire _16664_;
 wire _16665_;
 wire _16666_;
 wire _16667_;
 wire _16668_;
 wire _16669_;
 wire _16670_;
 wire _16671_;
 wire _16672_;
 wire _16673_;
 wire _16674_;
 wire _16675_;
 wire _16676_;
 wire _16677_;
 wire _16678_;
 wire _16679_;
 wire _16680_;
 wire _16681_;
 wire _16682_;
 wire _16683_;
 wire _16684_;
 wire _16685_;
 wire _16686_;
 wire _16687_;
 wire _16688_;
 wire _16689_;
 wire _16690_;
 wire _16691_;
 wire _16692_;
 wire _16693_;
 wire _16694_;
 wire _16695_;
 wire _16696_;
 wire _16697_;
 wire _16698_;
 wire _16699_;
 wire _16700_;
 wire _16701_;
 wire _16702_;
 wire _16703_;
 wire _16704_;
 wire _16705_;
 wire _16706_;
 wire _16707_;
 wire _16708_;
 wire _16709_;
 wire _16710_;
 wire _16711_;
 wire _16712_;
 wire _16713_;
 wire _16714_;
 wire _16715_;
 wire _16716_;
 wire _16717_;
 wire _16718_;
 wire _16719_;
 wire _16720_;
 wire _16721_;
 wire _16722_;
 wire _16723_;
 wire _16724_;
 wire _16725_;
 wire _16726_;
 wire _16727_;
 wire _16728_;
 wire _16729_;
 wire _16730_;
 wire _16731_;
 wire _16732_;
 wire _16733_;
 wire _16734_;
 wire _16735_;
 wire _16736_;
 wire _16737_;
 wire _16738_;
 wire _16739_;
 wire _16740_;
 wire _16741_;
 wire _16742_;
 wire _16743_;
 wire _16744_;
 wire _16745_;
 wire _16746_;
 wire _16747_;
 wire _16748_;
 wire _16749_;
 wire _16750_;
 wire _16751_;
 wire _16752_;
 wire _16753_;
 wire _16754_;
 wire _16755_;
 wire _16756_;
 wire _16757_;
 wire _16758_;
 wire _16759_;
 wire _16760_;
 wire _16761_;
 wire _16762_;
 wire _16763_;
 wire _16764_;
 wire _16765_;
 wire _16766_;
 wire _16767_;
 wire _16768_;
 wire _16769_;
 wire _16770_;
 wire _16771_;
 wire _16772_;
 wire _16773_;
 wire _16774_;
 wire _16775_;
 wire _16776_;
 wire _16777_;
 wire _16778_;
 wire _16779_;
 wire _16780_;
 wire _16781_;
 wire _16782_;
 wire _16783_;
 wire _16784_;
 wire _16785_;
 wire _16786_;
 wire _16787_;
 wire _16788_;
 wire _16789_;
 wire _16790_;
 wire _16791_;
 wire _16792_;
 wire _16793_;
 wire _16794_;
 wire _16795_;
 wire _16796_;
 wire _16797_;
 wire _16798_;
 wire _16799_;
 wire _16800_;
 wire _16801_;
 wire _16802_;
 wire _16803_;
 wire _16804_;
 wire _16805_;
 wire _16806_;
 wire _16807_;
 wire _16808_;
 wire _16809_;
 wire _16810_;
 wire _16811_;
 wire _16812_;
 wire _16813_;
 wire _16814_;
 wire _16815_;
 wire _16816_;
 wire _16817_;
 wire _16818_;
 wire _16819_;
 wire _16820_;
 wire _16821_;
 wire _16822_;
 wire _16823_;
 wire _16824_;
 wire _16825_;
 wire _16826_;
 wire _16827_;
 wire _16828_;
 wire _16829_;
 wire _16830_;
 wire _16831_;
 wire _16832_;
 wire _16833_;
 wire _16834_;
 wire _16835_;
 wire _16836_;
 wire _16837_;
 wire _16838_;
 wire _16839_;
 wire _16840_;
 wire _16841_;
 wire _16842_;
 wire _16843_;
 wire _16844_;
 wire _16845_;
 wire _16846_;
 wire _16847_;
 wire _16848_;
 wire _16849_;
 wire net1081;
 wire _16851_;
 wire _16852_;
 wire _16853_;
 wire net1080;
 wire _16855_;
 wire _16856_;
 wire _16857_;
 wire _16858_;
 wire _16859_;
 wire _16860_;
 wire _16861_;
 wire _16862_;
 wire _16863_;
 wire _16864_;
 wire _16865_;
 wire _16866_;
 wire _16867_;
 wire _16868_;
 wire _16869_;
 wire _16870_;
 wire _16871_;
 wire _16872_;
 wire _16873_;
 wire _16874_;
 wire _16875_;
 wire _16876_;
 wire _16877_;
 wire _16878_;
 wire _16879_;
 wire _16880_;
 wire _16881_;
 wire _16882_;
 wire _16883_;
 wire _16884_;
 wire _16885_;
 wire _16886_;
 wire _16887_;
 wire _16888_;
 wire _16889_;
 wire _16890_;
 wire _16891_;
 wire _16892_;
 wire _16893_;
 wire _16894_;
 wire _16895_;
 wire _16896_;
 wire _16897_;
 wire _16898_;
 wire _16899_;
 wire _16900_;
 wire _16901_;
 wire _16902_;
 wire _16903_;
 wire _16904_;
 wire _16905_;
 wire _16906_;
 wire _16907_;
 wire _16908_;
 wire _16909_;
 wire _16910_;
 wire _16911_;
 wire _16912_;
 wire _16913_;
 wire _16914_;
 wire _16915_;
 wire _16916_;
 wire _16917_;
 wire _16918_;
 wire _16919_;
 wire _16920_;
 wire _16921_;
 wire _16922_;
 wire _16923_;
 wire _16924_;
 wire _16925_;
 wire _16926_;
 wire _16927_;
 wire _16928_;
 wire _16929_;
 wire _16930_;
 wire _16931_;
 wire _16932_;
 wire _16933_;
 wire _16934_;
 wire _16935_;
 wire _16936_;
 wire _16937_;
 wire _16938_;
 wire _16939_;
 wire _16940_;
 wire _16941_;
 wire _16942_;
 wire _16943_;
 wire _16944_;
 wire _16945_;
 wire _16946_;
 wire _16947_;
 wire _16948_;
 wire _16949_;
 wire _16950_;
 wire _16951_;
 wire _16952_;
 wire _16953_;
 wire _16954_;
 wire _16955_;
 wire _16956_;
 wire _16957_;
 wire _16958_;
 wire _16959_;
 wire _16960_;
 wire _16961_;
 wire _16962_;
 wire _16963_;
 wire _16964_;
 wire _16965_;
 wire _16966_;
 wire _16967_;
 wire _16968_;
 wire _16969_;
 wire _16970_;
 wire _16971_;
 wire _16972_;
 wire _16973_;
 wire _16974_;
 wire _16975_;
 wire _16976_;
 wire _16977_;
 wire _16978_;
 wire _16979_;
 wire _16980_;
 wire _16981_;
 wire _16982_;
 wire _16983_;
 wire _16984_;
 wire _16985_;
 wire _16986_;
 wire _16987_;
 wire _16988_;
 wire _16989_;
 wire _16990_;
 wire _16991_;
 wire _16992_;
 wire _16993_;
 wire _16994_;
 wire _16995_;
 wire _16996_;
 wire _16997_;
 wire _16998_;
 wire _16999_;
 wire _17000_;
 wire _17001_;
 wire _17002_;
 wire _17003_;
 wire _17004_;
 wire _17005_;
 wire _17006_;
 wire _17007_;
 wire _17008_;
 wire _17009_;
 wire _17010_;
 wire _17011_;
 wire _17012_;
 wire _17013_;
 wire _17014_;
 wire _17015_;
 wire _17016_;
 wire _17017_;
 wire _17018_;
 wire _17019_;
 wire _17020_;
 wire _17021_;
 wire _17022_;
 wire _17023_;
 wire _17024_;
 wire _17025_;
 wire _17026_;
 wire _17027_;
 wire _17028_;
 wire _17029_;
 wire _17030_;
 wire _17031_;
 wire _17032_;
 wire _17033_;
 wire _17034_;
 wire _17035_;
 wire _17036_;
 wire _17037_;
 wire _17038_;
 wire _17039_;
 wire _17040_;
 wire _17041_;
 wire _17042_;
 wire _17043_;
 wire _17044_;
 wire _17045_;
 wire _17046_;
 wire _17047_;
 wire _17048_;
 wire _17049_;
 wire _17050_;
 wire _17051_;
 wire _17052_;
 wire _17053_;
 wire _17054_;
 wire net1079;
 wire _17056_;
 wire _17057_;
 wire _17058_;
 wire _17059_;
 wire _17060_;
 wire net1078;
 wire _17062_;
 wire _17063_;
 wire _17064_;
 wire _17065_;
 wire _17066_;
 wire _17067_;
 wire _17068_;
 wire _17069_;
 wire _17070_;
 wire _17071_;
 wire _17072_;
 wire _17073_;
 wire _17074_;
 wire _17075_;
 wire _17076_;
 wire _17077_;
 wire _17078_;
 wire _17079_;
 wire _17080_;
 wire _17081_;
 wire _17082_;
 wire _17083_;
 wire _17084_;
 wire _17085_;
 wire _17086_;
 wire _17087_;
 wire _17088_;
 wire _17089_;
 wire _17090_;
 wire _17091_;
 wire _17092_;
 wire _17093_;
 wire _17094_;
 wire _17095_;
 wire _17096_;
 wire _17097_;
 wire _17098_;
 wire _17099_;
 wire _17100_;
 wire _17101_;
 wire _17102_;
 wire _17103_;
 wire _17104_;
 wire _17105_;
 wire _17106_;
 wire _17107_;
 wire _17108_;
 wire _17109_;
 wire _17110_;
 wire _17111_;
 wire _17112_;
 wire _17113_;
 wire _17114_;
 wire _17115_;
 wire _17116_;
 wire _17117_;
 wire _17118_;
 wire _17119_;
 wire _17120_;
 wire _17121_;
 wire _17122_;
 wire _17123_;
 wire _17124_;
 wire _17125_;
 wire _17126_;
 wire _17127_;
 wire _17128_;
 wire _17129_;
 wire _17130_;
 wire _17131_;
 wire net1077;
 wire _17133_;
 wire _17134_;
 wire _17135_;
 wire _17136_;
 wire _17137_;
 wire _17138_;
 wire _17139_;
 wire _17140_;
 wire _17141_;
 wire _17142_;
 wire _17143_;
 wire _17144_;
 wire _17145_;
 wire _17146_;
 wire _17147_;
 wire _17148_;
 wire _17149_;
 wire net1076;
 wire _17151_;
 wire _17152_;
 wire _17153_;
 wire _17154_;
 wire _17155_;
 wire _17156_;
 wire _17157_;
 wire _17158_;
 wire _17159_;
 wire _17160_;
 wire _17161_;
 wire _17162_;
 wire _17163_;
 wire _17164_;
 wire _17165_;
 wire _17166_;
 wire _17167_;
 wire _17168_;
 wire _17169_;
 wire _17170_;
 wire _17171_;
 wire _17172_;
 wire _17173_;
 wire _17174_;
 wire net1075;
 wire _17176_;
 wire net1074;
 wire _17178_;
 wire _17179_;
 wire _17180_;
 wire _17181_;
 wire _17182_;
 wire _17183_;
 wire _17184_;
 wire _17185_;
 wire _17186_;
 wire _17187_;
 wire _17188_;
 wire _17189_;
 wire _17190_;
 wire _17191_;
 wire _17192_;
 wire _17193_;
 wire _17194_;
 wire _17195_;
 wire _17196_;
 wire _17197_;
 wire _17198_;
 wire _17199_;
 wire _17200_;
 wire _17201_;
 wire _17202_;
 wire _17203_;
 wire _17204_;
 wire _17205_;
 wire _17206_;
 wire _17207_;
 wire _17208_;
 wire _17209_;
 wire _17210_;
 wire _17211_;
 wire _17212_;
 wire _17213_;
 wire _17214_;
 wire _17215_;
 wire _17216_;
 wire _17217_;
 wire _17218_;
 wire _17219_;
 wire _17220_;
 wire _17221_;
 wire _17222_;
 wire _17223_;
 wire _17224_;
 wire _17225_;
 wire _17226_;
 wire _17227_;
 wire _17228_;
 wire _17229_;
 wire _17230_;
 wire _17231_;
 wire _17232_;
 wire _17233_;
 wire _17234_;
 wire _17235_;
 wire _17236_;
 wire _17237_;
 wire _17238_;
 wire _17239_;
 wire _17240_;
 wire _17241_;
 wire _17242_;
 wire _17243_;
 wire _17244_;
 wire _17245_;
 wire _17246_;
 wire _17247_;
 wire _17248_;
 wire _17249_;
 wire _17250_;
 wire _17251_;
 wire _17252_;
 wire _17253_;
 wire _17254_;
 wire _17255_;
 wire _17256_;
 wire _17257_;
 wire _17258_;
 wire _17259_;
 wire net1073;
 wire net1072;
 wire _17262_;
 wire _17263_;
 wire _17264_;
 wire _17265_;
 wire _17266_;
 wire _17267_;
 wire _17268_;
 wire _17269_;
 wire _17270_;
 wire _17271_;
 wire _17272_;
 wire _17273_;
 wire _17274_;
 wire _17275_;
 wire _17276_;
 wire _17277_;
 wire _17278_;
 wire _17279_;
 wire _17280_;
 wire _17281_;
 wire _17282_;
 wire _17283_;
 wire _17284_;
 wire _17285_;
 wire _17286_;
 wire _17287_;
 wire _17288_;
 wire _17289_;
 wire _17290_;
 wire _17291_;
 wire _17292_;
 wire _17293_;
 wire _17294_;
 wire _17295_;
 wire _17296_;
 wire _17297_;
 wire _17298_;
 wire _17299_;
 wire _17300_;
 wire _17301_;
 wire _17302_;
 wire _17303_;
 wire _17304_;
 wire net1071;
 wire _17306_;
 wire _17307_;
 wire _17308_;
 wire _17309_;
 wire _17310_;
 wire _17311_;
 wire _17312_;
 wire _17313_;
 wire _17314_;
 wire _17315_;
 wire _17316_;
 wire _17317_;
 wire _17318_;
 wire _17319_;
 wire _17320_;
 wire _17321_;
 wire _17322_;
 wire _17323_;
 wire _17324_;
 wire _17325_;
 wire _17326_;
 wire _17327_;
 wire _17328_;
 wire _17329_;
 wire _17330_;
 wire _17331_;
 wire _17332_;
 wire _17333_;
 wire _17334_;
 wire _17335_;
 wire _17336_;
 wire _17337_;
 wire _17338_;
 wire _17339_;
 wire _17340_;
 wire _17341_;
 wire _17342_;
 wire _17343_;
 wire _17344_;
 wire _17345_;
 wire _17346_;
 wire _17347_;
 wire _17348_;
 wire _17349_;
 wire _17350_;
 wire _17351_;
 wire _17352_;
 wire _17353_;
 wire net1070;
 wire _17355_;
 wire _17356_;
 wire _17357_;
 wire net1069;
 wire net1068;
 wire _17360_;
 wire _17361_;
 wire _17362_;
 wire _17363_;
 wire _17364_;
 wire _17365_;
 wire _17366_;
 wire _17367_;
 wire _17368_;
 wire _17369_;
 wire _17370_;
 wire _17371_;
 wire _17372_;
 wire _17373_;
 wire _17374_;
 wire _17375_;
 wire _17376_;
 wire _17377_;
 wire _17378_;
 wire _17379_;
 wire _17380_;
 wire _17381_;
 wire _17382_;
 wire _17383_;
 wire _17384_;
 wire _17385_;
 wire _17386_;
 wire _17387_;
 wire _17388_;
 wire net1067;
 wire _17390_;
 wire _17391_;
 wire _17392_;
 wire _17393_;
 wire _17394_;
 wire _17395_;
 wire _17396_;
 wire _17397_;
 wire _17398_;
 wire _17399_;
 wire _17400_;
 wire _17401_;
 wire _17402_;
 wire _17403_;
 wire _17404_;
 wire _17405_;
 wire _17406_;
 wire _17407_;
 wire _17408_;
 wire _17409_;
 wire _17410_;
 wire _17411_;
 wire _17412_;
 wire _17413_;
 wire _17414_;
 wire _17415_;
 wire _17416_;
 wire _17417_;
 wire _17418_;
 wire _17419_;
 wire _17420_;
 wire _17421_;
 wire _17422_;
 wire _17423_;
 wire _17424_;
 wire _17425_;
 wire _17426_;
 wire _17427_;
 wire _17428_;
 wire _17429_;
 wire _17430_;
 wire _17431_;
 wire _17432_;
 wire _17433_;
 wire _17434_;
 wire _17435_;
 wire _17436_;
 wire _17437_;
 wire _17438_;
 wire _17439_;
 wire _17440_;
 wire _17441_;
 wire _17442_;
 wire _17443_;
 wire _17444_;
 wire _17445_;
 wire _17446_;
 wire _17447_;
 wire _17448_;
 wire _17449_;
 wire _17450_;
 wire _17451_;
 wire _17452_;
 wire _17453_;
 wire net1066;
 wire net1065;
 wire _17456_;
 wire _17457_;
 wire _17458_;
 wire _17459_;
 wire _17460_;
 wire _17461_;
 wire _17462_;
 wire _17463_;
 wire _17464_;
 wire _17465_;
 wire _17466_;
 wire _17467_;
 wire _17468_;
 wire _17469_;
 wire _17470_;
 wire _17471_;
 wire _17472_;
 wire _17473_;
 wire _17474_;
 wire _17475_;
 wire _17476_;
 wire _17477_;
 wire _17478_;
 wire _17479_;
 wire _17480_;
 wire _17481_;
 wire _17482_;
 wire _17483_;
 wire _17484_;
 wire _17485_;
 wire _17486_;
 wire _17487_;
 wire net1064;
 wire _17489_;
 wire _17490_;
 wire _17491_;
 wire _17492_;
 wire _17493_;
 wire _17494_;
 wire _17495_;
 wire _17496_;
 wire _17497_;
 wire _17498_;
 wire _17499_;
 wire _17500_;
 wire _17501_;
 wire _17502_;
 wire _17503_;
 wire net1063;
 wire _17505_;
 wire _17506_;
 wire _17507_;
 wire _17508_;
 wire _17509_;
 wire _17510_;
 wire _17511_;
 wire _17512_;
 wire _17513_;
 wire _17514_;
 wire _17515_;
 wire _17516_;
 wire _17517_;
 wire _17518_;
 wire _17519_;
 wire _17520_;
 wire _17521_;
 wire _17522_;
 wire _17523_;
 wire _17524_;
 wire net1062;
 wire net1061;
 wire _17527_;
 wire _17528_;
 wire _17529_;
 wire _17530_;
 wire net1060;
 wire net1059;
 wire _17533_;
 wire _17534_;
 wire _17535_;
 wire _17536_;
 wire net1058;
 wire _17538_;
 wire _17539_;
 wire net1057;
 wire net1056;
 wire _17542_;
 wire _17543_;
 wire net1055;
 wire _17545_;
 wire _17546_;
 wire _17547_;
 wire _17548_;
 wire _17549_;
 wire _17550_;
 wire _17551_;
 wire net1054;
 wire _17553_;
 wire _17554_;
 wire _17555_;
 wire _17556_;
 wire _17557_;
 wire _17558_;
 wire _17559_;
 wire _17560_;
 wire _17561_;
 wire _17562_;
 wire _17563_;
 wire net1053;
 wire _17565_;
 wire _17566_;
 wire net1052;
 wire _17568_;
 wire _17569_;
 wire _17570_;
 wire _17571_;
 wire _17572_;
 wire _17573_;
 wire _17574_;
 wire _17575_;
 wire _17576_;
 wire _17577_;
 wire _17578_;
 wire _17579_;
 wire _17580_;
 wire _17581_;
 wire _17582_;
 wire net1051;
 wire net1050;
 wire net1049;
 wire _17586_;
 wire net1048;
 wire _17588_;
 wire _17589_;
 wire net1047;
 wire _17591_;
 wire _17592_;
 wire _17593_;
 wire net1046;
 wire net1045;
 wire _17596_;
 wire net1044;
 wire _17598_;
 wire _17599_;
 wire _17600_;
 wire _17601_;
 wire _17602_;
 wire _17603_;
 wire _17604_;
 wire _17605_;
 wire net1043;
 wire _17607_;
 wire _17608_;
 wire _17609_;
 wire _17610_;
 wire _17611_;
 wire _17612_;
 wire _17613_;
 wire _17614_;
 wire net1042;
 wire _17616_;
 wire _17617_;
 wire _17618_;
 wire _17619_;
 wire _17620_;
 wire _17621_;
 wire _17622_;
 wire _17623_;
 wire _17624_;
 wire net1041;
 wire _17626_;
 wire net1040;
 wire _17628_;
 wire _17629_;
 wire net1039;
 wire _17631_;
 wire _17632_;
 wire _17633_;
 wire _17634_;
 wire net1038;
 wire _17636_;
 wire _17637_;
 wire _17638_;
 wire _17639_;
 wire net1037;
 wire _17641_;
 wire net1036;
 wire net1035;
 wire _17644_;
 wire _17645_;
 wire _17646_;
 wire _17647_;
 wire _17648_;
 wire _17649_;
 wire _17650_;
 wire net1034;
 wire net1033;
 wire net1032;
 wire _17654_;
 wire _17655_;
 wire _17656_;
 wire _17657_;
 wire net1031;
 wire _17659_;
 wire _17660_;
 wire _17661_;
 wire _17662_;
 wire _17663_;
 wire net1030;
 wire _17665_;
 wire _17666_;
 wire _17667_;
 wire net1029;
 wire _17669_;
 wire _17670_;
 wire _17671_;
 wire _17672_;
 wire _17673_;
 wire _17674_;
 wire _17675_;
 wire _17676_;
 wire _17677_;
 wire _17678_;
 wire _17679_;
 wire _17680_;
 wire _17681_;
 wire _17682_;
 wire _17683_;
 wire _17684_;
 wire _17685_;
 wire net1028;
 wire _17687_;
 wire net1027;
 wire _17689_;
 wire _17690_;
 wire _17691_;
 wire _17692_;
 wire _17693_;
 wire _17694_;
 wire _17695_;
 wire net1026;
 wire _17697_;
 wire _17698_;
 wire net1025;
 wire _17700_;
 wire _17701_;
 wire net1024;
 wire _17703_;
 wire net1023;
 wire _17705_;
 wire _17706_;
 wire _17707_;
 wire net1022;
 wire _17709_;
 wire _17710_;
 wire _17711_;
 wire _17712_;
 wire _17713_;
 wire _17714_;
 wire _17715_;
 wire _17716_;
 wire _17717_;
 wire _17718_;
 wire net1021;
 wire _17720_;
 wire _17721_;
 wire _17722_;
 wire _17723_;
 wire net1020;
 wire _17725_;
 wire net1019;
 wire _17727_;
 wire _17728_;
 wire _17729_;
 wire _17730_;
 wire _17731_;
 wire _17732_;
 wire _17733_;
 wire _17734_;
 wire _17735_;
 wire net1018;
 wire _17737_;
 wire _17738_;
 wire _17739_;
 wire _17740_;
 wire _17741_;
 wire _17742_;
 wire _17743_;
 wire _17744_;
 wire _17745_;
 wire _17746_;
 wire _17747_;
 wire net1017;
 wire _17749_;
 wire _17750_;
 wire net1016;
 wire net1015;
 wire net1014;
 wire _17754_;
 wire _17755_;
 wire _17756_;
 wire _17757_;
 wire _17758_;
 wire _17759_;
 wire net1013;
 wire _17761_;
 wire _17762_;
 wire net1012;
 wire _17764_;
 wire _17765_;
 wire _17766_;
 wire _17767_;
 wire _17768_;
 wire _17769_;
 wire _17770_;
 wire _17771_;
 wire net1011;
 wire _17773_;
 wire _17774_;
 wire _17775_;
 wire _17776_;
 wire _17777_;
 wire net1010;
 wire _17779_;
 wire _17780_;
 wire _17781_;
 wire _17782_;
 wire _17783_;
 wire _17784_;
 wire _17785_;
 wire _17786_;
 wire _17787_;
 wire _17788_;
 wire net1009;
 wire _17790_;
 wire _17791_;
 wire _17792_;
 wire _17793_;
 wire _17794_;
 wire _17795_;
 wire _17796_;
 wire _17797_;
 wire net1008;
 wire _17799_;
 wire _17800_;
 wire _17801_;
 wire _17802_;
 wire _17803_;
 wire _17804_;
 wire _17805_;
 wire _17806_;
 wire _17807_;
 wire _17808_;
 wire _17809_;
 wire _17810_;
 wire _17811_;
 wire _17812_;
 wire _17813_;
 wire _17814_;
 wire _17815_;
 wire net1007;
 wire _17817_;
 wire _17818_;
 wire _17819_;
 wire _17820_;
 wire _17821_;
 wire _17822_;
 wire _17823_;
 wire _17824_;
 wire _17825_;
 wire _17826_;
 wire _17827_;
 wire _17828_;
 wire _17829_;
 wire _17830_;
 wire _17831_;
 wire _17832_;
 wire _17833_;
 wire _17834_;
 wire _17835_;
 wire _17836_;
 wire _17837_;
 wire _17838_;
 wire _17839_;
 wire net1006;
 wire _17841_;
 wire _17842_;
 wire _17843_;
 wire _17844_;
 wire _17845_;
 wire net1005;
 wire _17847_;
 wire _17848_;
 wire _17849_;
 wire _17850_;
 wire _17851_;
 wire _17852_;
 wire _17853_;
 wire _17854_;
 wire _17855_;
 wire _17856_;
 wire _17857_;
 wire _17858_;
 wire _17859_;
 wire _17860_;
 wire _17861_;
 wire _17862_;
 wire _17863_;
 wire _17864_;
 wire _17865_;
 wire _17866_;
 wire net1004;
 wire _17868_;
 wire _17869_;
 wire _17870_;
 wire _17871_;
 wire _17872_;
 wire _17873_;
 wire _17874_;
 wire _17875_;
 wire _17876_;
 wire _17877_;
 wire net1003;
 wire _17879_;
 wire _17880_;
 wire _17881_;
 wire _17882_;
 wire _17883_;
 wire _17884_;
 wire _17885_;
 wire _17886_;
 wire _17887_;
 wire _17888_;
 wire _17889_;
 wire _17890_;
 wire _17891_;
 wire _17892_;
 wire _17893_;
 wire _17894_;
 wire _17895_;
 wire _17896_;
 wire _17897_;
 wire _17898_;
 wire _17899_;
 wire _17900_;
 wire _17901_;
 wire _17902_;
 wire _17903_;
 wire _17904_;
 wire _17905_;
 wire _17906_;
 wire _17907_;
 wire _17908_;
 wire _17909_;
 wire _17910_;
 wire _17911_;
 wire _17912_;
 wire _17913_;
 wire _17914_;
 wire _17915_;
 wire _17916_;
 wire _17917_;
 wire _17918_;
 wire _17919_;
 wire _17920_;
 wire _17921_;
 wire net1002;
 wire _17923_;
 wire _17924_;
 wire _17925_;
 wire net1001;
 wire net1000;
 wire _17928_;
 wire net999;
 wire _17930_;
 wire _17931_;
 wire _17932_;
 wire _17933_;
 wire _17934_;
 wire net998;
 wire _17936_;
 wire _17937_;
 wire _17938_;
 wire net997;
 wire net996;
 wire _17941_;
 wire _17942_;
 wire _17943_;
 wire net995;
 wire _17945_;
 wire _17946_;
 wire _17947_;
 wire _17948_;
 wire _17949_;
 wire net994;
 wire _17951_;
 wire _17952_;
 wire _17953_;
 wire _17954_;
 wire _17955_;
 wire _17956_;
 wire _17957_;
 wire _17958_;
 wire _17959_;
 wire _17960_;
 wire _17961_;
 wire _17962_;
 wire _17963_;
 wire _17964_;
 wire _17965_;
 wire _17966_;
 wire _17967_;
 wire _17968_;
 wire net993;
 wire _17970_;
 wire _17971_;
 wire _17972_;
 wire _17973_;
 wire _17974_;
 wire _17975_;
 wire _17976_;
 wire _17977_;
 wire net992;
 wire net991;
 wire _17980_;
 wire net990;
 wire _17982_;
 wire _17983_;
 wire _17984_;
 wire _17985_;
 wire _17986_;
 wire _17987_;
 wire net989;
 wire net988;
 wire _17990_;
 wire _17991_;
 wire _17992_;
 wire _17993_;
 wire net987;
 wire _17995_;
 wire _17996_;
 wire _17997_;
 wire net986;
 wire _17999_;
 wire _18000_;
 wire net985;
 wire _18002_;
 wire _18003_;
 wire _18004_;
 wire _18005_;
 wire _18006_;
 wire _18007_;
 wire _18008_;
 wire _18009_;
 wire _18010_;
 wire net984;
 wire _18012_;
 wire _18013_;
 wire _18014_;
 wire net983;
 wire net982;
 wire _18017_;
 wire _18018_;
 wire _18019_;
 wire _18020_;
 wire _18021_;
 wire _18022_;
 wire net981;
 wire _18024_;
 wire _18025_;
 wire _18026_;
 wire _18027_;
 wire _18028_;
 wire net980;
 wire _18030_;
 wire _18031_;
 wire _18032_;
 wire _18033_;
 wire _18034_;
 wire net979;
 wire _18036_;
 wire _18037_;
 wire _18038_;
 wire _18039_;
 wire _18040_;
 wire net978;
 wire net977;
 wire net976;
 wire net975;
 wire _18045_;
 wire _18046_;
 wire _18047_;
 wire _18048_;
 wire _18049_;
 wire _18050_;
 wire net974;
 wire _18052_;
 wire net973;
 wire _18054_;
 wire net972;
 wire _18056_;
 wire _18057_;
 wire net971;
 wire _18059_;
 wire net970;
 wire _18061_;
 wire _18062_;
 wire _18063_;
 wire _18064_;
 wire _18065_;
 wire net969;
 wire _18067_;
 wire _18068_;
 wire _18069_;
 wire _18070_;
 wire _18071_;
 wire _18072_;
 wire _18073_;
 wire _18074_;
 wire net968;
 wire _18076_;
 wire _18077_;
 wire _18078_;
 wire _18079_;
 wire net967;
 wire _18081_;
 wire net966;
 wire _18083_;
 wire _18084_;
 wire _18085_;
 wire _18086_;
 wire _18087_;
 wire _18088_;
 wire _18089_;
 wire _18090_;
 wire net965;
 wire net964;
 wire _18093_;
 wire net963;
 wire _18095_;
 wire _18096_;
 wire net962;
 wire _18098_;
 wire _18099_;
 wire _18100_;
 wire _18101_;
 wire _18102_;
 wire _18103_;
 wire _18104_;
 wire _18105_;
 wire _18106_;
 wire _18107_;
 wire _18108_;
 wire net961;
 wire _18110_;
 wire _18111_;
 wire net960;
 wire _18113_;
 wire _18114_;
 wire _18115_;
 wire _18116_;
 wire net959;
 wire _18118_;
 wire _18119_;
 wire _18120_;
 wire _18121_;
 wire _18122_;
 wire _18123_;
 wire net958;
 wire _18125_;
 wire _18126_;
 wire _18127_;
 wire _18128_;
 wire _18129_;
 wire _18130_;
 wire _18131_;
 wire net957;
 wire _18133_;
 wire _18134_;
 wire _18135_;
 wire _18136_;
 wire _18137_;
 wire _18138_;
 wire _18139_;
 wire _18140_;
 wire net956;
 wire net955;
 wire _18143_;
 wire _18144_;
 wire net954;
 wire _18146_;
 wire _18147_;
 wire net953;
 wire _18149_;
 wire _18150_;
 wire _18151_;
 wire _18152_;
 wire _18153_;
 wire _18154_;
 wire _18155_;
 wire _18156_;
 wire _18157_;
 wire _18158_;
 wire net952;
 wire _18160_;
 wire _18161_;
 wire _18162_;
 wire _18163_;
 wire _18164_;
 wire _18165_;
 wire _18166_;
 wire _18167_;
 wire _18168_;
 wire _18169_;
 wire net951;
 wire _18171_;
 wire _18172_;
 wire _18173_;
 wire _18174_;
 wire _18175_;
 wire net950;
 wire _18177_;
 wire _18178_;
 wire net949;
 wire _18180_;
 wire _18181_;
 wire _18182_;
 wire _18183_;
 wire _18184_;
 wire _18185_;
 wire _18186_;
 wire _18187_;
 wire _18188_;
 wire _18189_;
 wire _18190_;
 wire _18191_;
 wire _18192_;
 wire _18193_;
 wire _18194_;
 wire _18195_;
 wire _18196_;
 wire _18197_;
 wire _18198_;
 wire _18199_;
 wire _18200_;
 wire _18201_;
 wire _18202_;
 wire _18203_;
 wire _18204_;
 wire _18205_;
 wire _18206_;
 wire _18207_;
 wire _18208_;
 wire _18209_;
 wire _18210_;
 wire _18211_;
 wire _18212_;
 wire _18213_;
 wire _18214_;
 wire _18215_;
 wire _18216_;
 wire _18217_;
 wire _18218_;
 wire _18219_;
 wire _18220_;
 wire _18221_;
 wire _18222_;
 wire _18223_;
 wire _18224_;
 wire _18225_;
 wire _18226_;
 wire _18227_;
 wire _18228_;
 wire _18229_;
 wire _18230_;
 wire _18231_;
 wire _18232_;
 wire _18233_;
 wire net948;
 wire _18235_;
 wire net947;
 wire _18237_;
 wire _18238_;
 wire _18239_;
 wire _18240_;
 wire _18241_;
 wire _18242_;
 wire _18243_;
 wire net946;
 wire net945;
 wire _18246_;
 wire _18247_;
 wire _18248_;
 wire _18249_;
 wire _18250_;
 wire net944;
 wire _18252_;
 wire _18253_;
 wire _18254_;
 wire _18255_;
 wire _18256_;
 wire _18257_;
 wire _18258_;
 wire _18259_;
 wire _18260_;
 wire _18261_;
 wire _18262_;
 wire _18263_;
 wire _18264_;
 wire _18265_;
 wire _18266_;
 wire net943;
 wire _18268_;
 wire _18269_;
 wire _18270_;
 wire _18271_;
 wire _18272_;
 wire _18273_;
 wire _18274_;
 wire _18275_;
 wire _18276_;
 wire _18277_;
 wire _18278_;
 wire _18279_;
 wire _18280_;
 wire _18281_;
 wire _18282_;
 wire _18283_;
 wire _18284_;
 wire _18285_;
 wire _18286_;
 wire _18287_;
 wire net942;
 wire _18289_;
 wire _18290_;
 wire _18291_;
 wire _18292_;
 wire _18293_;
 wire _18294_;
 wire _18295_;
 wire _18296_;
 wire _18297_;
 wire net941;
 wire _18299_;
 wire _18300_;
 wire net940;
 wire _18302_;
 wire _18303_;
 wire _18304_;
 wire _18305_;
 wire _18306_;
 wire _18307_;
 wire net939;
 wire _18309_;
 wire _18310_;
 wire _18311_;
 wire _18312_;
 wire _18313_;
 wire _18314_;
 wire net938;
 wire _18316_;
 wire net937;
 wire _18318_;
 wire net936;
 wire _18320_;
 wire clknet_1_1__leaf_clk;
 wire _18322_;
 wire clknet_1_0__leaf_clk;
 wire _18324_;
 wire _18325_;
 wire clknet_0_clk;
 wire _18327_;
 wire clknet_leaf_17_clk;
 wire _18329_;
 wire _18330_;
 wire clknet_leaf_16_clk;
 wire _18332_;
 wire _18333_;
 wire clknet_leaf_15_clk;
 wire _18335_;
 wire clknet_leaf_14_clk;
 wire _18337_;
 wire _18338_;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_11_clk;
 wire _18342_;
 wire _18343_;
 wire _18344_;
 wire _18345_;
 wire _18346_;
 wire _18347_;
 wire _18348_;
 wire _18349_;
 wire _18350_;
 wire _18351_;
 wire clknet_leaf_10_clk;
 wire _18353_;
 wire _18354_;
 wire clknet_leaf_9_clk;
 wire _18356_;
 wire _18357_;
 wire clknet_leaf_8_clk;
 wire _18359_;
 wire clknet_leaf_7_clk;
 wire _18361_;
 wire _18362_;
 wire clknet_leaf_6_clk;
 wire _18364_;
 wire clknet_leaf_5_clk;
 wire _18366_;
 wire clknet_leaf_4_clk;
 wire _18368_;
 wire _18369_;
 wire clknet_leaf_3_clk;
 wire _18371_;
 wire _18372_;
 wire _18373_;
 wire _18374_;
 wire _18375_;
 wire _18376_;
 wire _18377_;
 wire clknet_leaf_2_clk;
 wire _18379_;
 wire _18380_;
 wire _18381_;
 wire clknet_leaf_1_clk;
 wire _18383_;
 wire net935;
 wire net934;
 wire _18386_;
 wire _18387_;
 wire _18388_;
 wire net933;
 wire _18390_;
 wire _18391_;
 wire _18392_;
 wire _18393_;
 wire _18394_;
 wire _18395_;
 wire net932;
 wire _18397_;
 wire _18398_;
 wire _18399_;
 wire _18400_;
 wire _18401_;
 wire _18402_;
 wire net931;
 wire _18404_;
 wire _18405_;
 wire _18406_;
 wire _18407_;
 wire _18408_;
 wire _18409_;
 wire _18410_;
 wire _18411_;
 wire net930;
 wire _18413_;
 wire net929;
 wire _18415_;
 wire _18416_;
 wire _18417_;
 wire _18418_;
 wire _18419_;
 wire _18420_;
 wire _18421_;
 wire _18422_;
 wire net928;
 wire _18424_;
 wire _18425_;
 wire _18426_;
 wire _18427_;
 wire _18428_;
 wire net927;
 wire _18430_;
 wire _18431_;
 wire _18432_;
 wire _18433_;
 wire _18434_;
 wire _18435_;
 wire _18436_;
 wire _18437_;
 wire net926;
 wire _18439_;
 wire net925;
 wire _18441_;
 wire _18442_;
 wire _18443_;
 wire _18444_;
 wire _18445_;
 wire _18446_;
 wire _18447_;
 wire _18448_;
 wire _18449_;
 wire _18450_;
 wire _18451_;
 wire _18452_;
 wire _18453_;
 wire net924;
 wire _18455_;
 wire _18456_;
 wire net923;
 wire _18458_;
 wire _18459_;
 wire _18460_;
 wire _18461_;
 wire _18462_;
 wire _18463_;
 wire _18464_;
 wire net922;
 wire _18466_;
 wire _18467_;
 wire _18468_;
 wire _18469_;
 wire _18470_;
 wire _18471_;
 wire net921;
 wire _18473_;
 wire _18474_;
 wire _18475_;
 wire _18476_;
 wire _18477_;
 wire net920;
 wire _18479_;
 wire net919;
 wire _18481_;
 wire _18482_;
 wire _18483_;
 wire _18484_;
 wire _18485_;
 wire _18486_;
 wire _18487_;
 wire _18488_;
 wire _18489_;
 wire _18490_;
 wire net918;
 wire _18492_;
 wire _18493_;
 wire net917;
 wire _18495_;
 wire _18496_;
 wire _18497_;
 wire _18498_;
 wire _18499_;
 wire _18500_;
 wire _18501_;
 wire _18502_;
 wire _18503_;
 wire _18504_;
 wire _18505_;
 wire _18506_;
 wire _18507_;
 wire net916;
 wire net915;
 wire _18510_;
 wire _18511_;
 wire net914;
 wire net913;
 wire _18514_;
 wire _18515_;
 wire _18516_;
 wire _18517_;
 wire _18518_;
 wire net912;
 wire net911;
 wire _18521_;
 wire net910;
 wire _18523_;
 wire _18524_;
 wire _18525_;
 wire _18526_;
 wire _18527_;
 wire _18528_;
 wire net909;
 wire _18530_;
 wire _18531_;
 wire _18532_;
 wire _18533_;
 wire net908;
 wire _18535_;
 wire _18536_;
 wire _18537_;
 wire _18538_;
 wire _18539_;
 wire _18540_;
 wire net907;
 wire _18542_;
 wire _18543_;
 wire _18544_;
 wire _18545_;
 wire net906;
 wire _18547_;
 wire _18548_;
 wire _18549_;
 wire _18550_;
 wire _18551_;
 wire _18552_;
 wire _18553_;
 wire _18554_;
 wire _18555_;
 wire _18556_;
 wire net905;
 wire _18558_;
 wire _18559_;
 wire _18560_;
 wire _18561_;
 wire _18562_;
 wire _18563_;
 wire _18564_;
 wire _18565_;
 wire net904;
 wire _18567_;
 wire _18568_;
 wire _18569_;
 wire _18570_;
 wire _18571_;
 wire _18572_;
 wire _18573_;
 wire _18574_;
 wire _18575_;
 wire _18576_;
 wire _18577_;
 wire _18578_;
 wire _18579_;
 wire net903;
 wire _18581_;
 wire net902;
 wire _18583_;
 wire _18584_;
 wire _18585_;
 wire _18586_;
 wire _18587_;
 wire _18588_;
 wire _18589_;
 wire _18590_;
 wire _18591_;
 wire _18592_;
 wire _18593_;
 wire _18594_;
 wire _18595_;
 wire _18596_;
 wire _18597_;
 wire _18598_;
 wire _18599_;
 wire _18600_;
 wire _18601_;
 wire _18602_;
 wire _18603_;
 wire _18604_;
 wire _18605_;
 wire _18606_;
 wire _18607_;
 wire _18608_;
 wire net901;
 wire _18610_;
 wire _18611_;
 wire _18612_;
 wire _18613_;
 wire _18614_;
 wire _18615_;
 wire _18616_;
 wire _18617_;
 wire _18618_;
 wire _18619_;
 wire _18620_;
 wire _18621_;
 wire net900;
 wire _18623_;
 wire _18624_;
 wire _18625_;
 wire _18626_;
 wire _18627_;
 wire net899;
 wire _18629_;
 wire _18630_;
 wire _18631_;
 wire _18632_;
 wire _18633_;
 wire _18634_;
 wire _18635_;
 wire _18636_;
 wire _18637_;
 wire _18638_;
 wire _18639_;
 wire _18640_;
 wire _18641_;
 wire _18642_;
 wire _18643_;
 wire _18644_;
 wire _18645_;
 wire _18646_;
 wire _18647_;
 wire _18648_;
 wire _18649_;
 wire _18650_;
 wire _18651_;
 wire net898;
 wire _18653_;
 wire _18654_;
 wire _18655_;
 wire _18656_;
 wire _18657_;
 wire _18658_;
 wire _18659_;
 wire net897;
 wire _18661_;
 wire _18662_;
 wire _18663_;
 wire net896;
 wire net895;
 wire _18666_;
 wire net894;
 wire _18668_;
 wire _18669_;
 wire _18670_;
 wire _18671_;
 wire _18672_;
 wire _18673_;
 wire _18674_;
 wire _18675_;
 wire _18676_;
 wire _18677_;
 wire _18678_;
 wire _18679_;
 wire _18680_;
 wire _18681_;
 wire _18682_;
 wire _18683_;
 wire _18684_;
 wire _18685_;
 wire net893;
 wire _18687_;
 wire _18688_;
 wire _18689_;
 wire _18690_;
 wire _18691_;
 wire _18692_;
 wire _18693_;
 wire _18694_;
 wire _18695_;
 wire _18696_;
 wire _18697_;
 wire _18698_;
 wire _18699_;
 wire net892;
 wire net891;
 wire _18702_;
 wire _18703_;
 wire _18704_;
 wire _18705_;
 wire _18706_;
 wire _18707_;
 wire _18708_;
 wire net890;
 wire net889;
 wire _18711_;
 wire _18712_;
 wire _18713_;
 wire _18714_;
 wire _18715_;
 wire _18716_;
 wire _18717_;
 wire _18718_;
 wire _18719_;
 wire _18720_;
 wire _18721_;
 wire net888;
 wire _18723_;
 wire _18724_;
 wire _18725_;
 wire _18726_;
 wire _18727_;
 wire _18728_;
 wire _18729_;
 wire _18730_;
 wire _18731_;
 wire _18732_;
 wire _18733_;
 wire _18734_;
 wire _18735_;
 wire _18736_;
 wire _18737_;
 wire _18738_;
 wire _18739_;
 wire _18740_;
 wire _18741_;
 wire _18742_;
 wire _18743_;
 wire _18744_;
 wire _18745_;
 wire _18746_;
 wire _18747_;
 wire _18748_;
 wire net887;
 wire net886;
 wire _18751_;
 wire _18752_;
 wire _18753_;
 wire net885;
 wire net884;
 wire _18756_;
 wire _18757_;
 wire net883;
 wire _18759_;
 wire _18760_;
 wire _18761_;
 wire net882;
 wire _18763_;
 wire _18764_;
 wire _18765_;
 wire _18766_;
 wire _18767_;
 wire _18768_;
 wire _18769_;
 wire net881;
 wire _18771_;
 wire net880;
 wire _18773_;
 wire _18774_;
 wire _18775_;
 wire net879;
 wire _18777_;
 wire _18778_;
 wire _18779_;
 wire _18780_;
 wire _18781_;
 wire _18782_;
 wire _18783_;
 wire _18784_;
 wire _18785_;
 wire _18786_;
 wire _18787_;
 wire _18788_;
 wire _18789_;
 wire _18790_;
 wire _18791_;
 wire _18792_;
 wire net878;
 wire _18794_;
 wire _18795_;
 wire _18796_;
 wire _18797_;
 wire _18798_;
 wire _18799_;
 wire _18800_;
 wire _18801_;
 wire _18802_;
 wire net877;
 wire _18804_;
 wire _18805_;
 wire _18806_;
 wire _18807_;
 wire _18808_;
 wire _18809_;
 wire _18810_;
 wire _18811_;
 wire _18812_;
 wire _18813_;
 wire _18814_;
 wire _18815_;
 wire _18816_;
 wire _18817_;
 wire _18818_;
 wire _18819_;
 wire _18820_;
 wire _18821_;
 wire _18822_;
 wire _18823_;
 wire _18824_;
 wire _18825_;
 wire _18826_;
 wire _18827_;
 wire _18828_;
 wire _18829_;
 wire _18830_;
 wire _18831_;
 wire _18832_;
 wire _18833_;
 wire _18834_;
 wire _18835_;
 wire _18836_;
 wire _18837_;
 wire _18838_;
 wire _18839_;
 wire _18840_;
 wire _18841_;
 wire net876;
 wire _18843_;
 wire _18844_;
 wire _18845_;
 wire _18846_;
 wire _18847_;
 wire _18848_;
 wire _18849_;
 wire _18850_;
 wire _18851_;
 wire _18852_;
 wire _18853_;
 wire _18854_;
 wire net875;
 wire _18856_;
 wire _18857_;
 wire _18858_;
 wire _18859_;
 wire _18860_;
 wire _18861_;
 wire _18862_;
 wire _18863_;
 wire _18864_;
 wire _18865_;
 wire _18866_;
 wire _18867_;
 wire _18868_;
 wire _18869_;
 wire _18870_;
 wire net874;
 wire _18872_;
 wire _18873_;
 wire _18874_;
 wire _18875_;
 wire _18876_;
 wire _18877_;
 wire _18878_;
 wire _18879_;
 wire _18880_;
 wire _18881_;
 wire net873;
 wire _18883_;
 wire net872;
 wire _18885_;
 wire _18886_;
 wire _18887_;
 wire _18888_;
 wire _18889_;
 wire _18890_;
 wire net871;
 wire _18892_;
 wire _18893_;
 wire _18894_;
 wire _18895_;
 wire _18896_;
 wire _18897_;
 wire _18898_;
 wire _18899_;
 wire _18900_;
 wire _18901_;
 wire _18902_;
 wire _18903_;
 wire _18904_;
 wire _18905_;
 wire net870;
 wire _18907_;
 wire _18908_;
 wire _18909_;
 wire _18910_;
 wire _18911_;
 wire _18912_;
 wire _18913_;
 wire net869;
 wire _18915_;
 wire _18916_;
 wire _18917_;
 wire _18918_;
 wire net868;
 wire _18920_;
 wire _18921_;
 wire _18922_;
 wire _18923_;
 wire _18924_;
 wire _18925_;
 wire _18926_;
 wire _18927_;
 wire _18928_;
 wire _18929_;
 wire _18930_;
 wire _18931_;
 wire _18932_;
 wire _18933_;
 wire _18934_;
 wire _18935_;
 wire _18936_;
 wire _18937_;
 wire _18938_;
 wire _18939_;
 wire _18940_;
 wire _18941_;
 wire _18942_;
 wire _18943_;
 wire _18944_;
 wire _18945_;
 wire _18946_;
 wire _18947_;
 wire _18948_;
 wire _18949_;
 wire net867;
 wire _18951_;
 wire _18952_;
 wire _18953_;
 wire _18954_;
 wire _18955_;
 wire _18956_;
 wire _18957_;
 wire _18958_;
 wire _18959_;
 wire _18960_;
 wire _18961_;
 wire _18962_;
 wire _18963_;
 wire _18964_;
 wire _18965_;
 wire _18966_;
 wire _18967_;
 wire _18968_;
 wire _18969_;
 wire _18970_;
 wire _18971_;
 wire _18972_;
 wire net866;
 wire net865;
 wire _18975_;
 wire _18976_;
 wire _18977_;
 wire net864;
 wire net863;
 wire net862;
 wire _18981_;
 wire _18982_;
 wire _18983_;
 wire net861;
 wire net860;
 wire net859;
 wire _18987_;
 wire _18988_;
 wire _18989_;
 wire _18990_;
 wire _18991_;
 wire _18992_;
 wire net858;
 wire net857;
 wire _18995_;
 wire _18996_;
 wire _18997_;
 wire _18998_;
 wire _18999_;
 wire _19000_;
 wire _19001_;
 wire _19002_;
 wire _19003_;
 wire _19004_;
 wire net856;
 wire _19006_;
 wire _19007_;
 wire _19008_;
 wire net855;
 wire _19010_;
 wire _19011_;
 wire _19012_;
 wire _19013_;
 wire _19014_;
 wire _19015_;
 wire _19016_;
 wire _19017_;
 wire _19018_;
 wire _19019_;
 wire net854;
 wire _19021_;
 wire net853;
 wire _19023_;
 wire _19024_;
 wire _19025_;
 wire _19026_;
 wire net852;
 wire _19028_;
 wire _19029_;
 wire _19030_;
 wire _19031_;
 wire _19032_;
 wire _19033_;
 wire _19034_;
 wire _19035_;
 wire _19036_;
 wire net851;
 wire _19038_;
 wire net850;
 wire _19040_;
 wire _19041_;
 wire _19042_;
 wire net849;
 wire _19044_;
 wire _19045_;
 wire _19046_;
 wire _19047_;
 wire _19048_;
 wire _19049_;
 wire _19050_;
 wire net848;
 wire _19052_;
 wire _19053_;
 wire _19054_;
 wire _19055_;
 wire _19056_;
 wire _19057_;
 wire _19058_;
 wire _19059_;
 wire _19060_;
 wire _19061_;
 wire _19062_;
 wire _19063_;
 wire _19064_;
 wire _19065_;
 wire net847;
 wire _19067_;
 wire _19068_;
 wire _19069_;
 wire _19070_;
 wire _19071_;
 wire _19072_;
 wire _19073_;
 wire net846;
 wire _19075_;
 wire _19076_;
 wire net845;
 wire _19078_;
 wire _19079_;
 wire _19080_;
 wire _19081_;
 wire _19082_;
 wire _19083_;
 wire _19084_;
 wire _19085_;
 wire _19086_;
 wire _19087_;
 wire _19088_;
 wire net844;
 wire _19090_;
 wire _19091_;
 wire _19092_;
 wire _19093_;
 wire _19094_;
 wire _19095_;
 wire net843;
 wire _19097_;
 wire _19098_;
 wire _19099_;
 wire _19100_;
 wire _19101_;
 wire _19102_;
 wire _19103_;
 wire _19104_;
 wire _19105_;
 wire _19106_;
 wire _19107_;
 wire _19108_;
 wire _19109_;
 wire _19110_;
 wire _19111_;
 wire _19112_;
 wire _19113_;
 wire _19114_;
 wire _19115_;
 wire _19116_;
 wire _19117_;
 wire _19118_;
 wire _19119_;
 wire _19120_;
 wire _19121_;
 wire _19122_;
 wire _19123_;
 wire _19124_;
 wire _19125_;
 wire _19126_;
 wire _19127_;
 wire _19128_;
 wire _19129_;
 wire _19130_;
 wire _19131_;
 wire _19132_;
 wire _19133_;
 wire _19134_;
 wire _19135_;
 wire _19136_;
 wire _19137_;
 wire _19138_;
 wire _19139_;
 wire _19140_;
 wire _19141_;
 wire _19142_;
 wire _19143_;
 wire _19144_;
 wire _19145_;
 wire _19146_;
 wire _19147_;
 wire _19148_;
 wire _19149_;
 wire _19150_;
 wire _19151_;
 wire _19152_;
 wire _19153_;
 wire _19154_;
 wire _19155_;
 wire _19156_;
 wire _19157_;
 wire _19158_;
 wire _19159_;
 wire _19160_;
 wire _19161_;
 wire _19162_;
 wire _19163_;
 wire _19164_;
 wire _19165_;
 wire _19166_;
 wire _19167_;
 wire _19168_;
 wire _19169_;
 wire _19170_;
 wire _19171_;
 wire net842;
 wire _19173_;
 wire _19174_;
 wire _19175_;
 wire _19176_;
 wire _19177_;
 wire _19178_;
 wire net841;
 wire _19180_;
 wire _19181_;
 wire _19182_;
 wire _19183_;
 wire _19184_;
 wire _19185_;
 wire _19186_;
 wire _19187_;
 wire _19188_;
 wire _19189_;
 wire _19190_;
 wire _19191_;
 wire _19192_;
 wire _19193_;
 wire net840;
 wire _19195_;
 wire _19196_;
 wire _19197_;
 wire _19198_;
 wire _19199_;
 wire _19200_;
 wire _19201_;
 wire _19202_;
 wire _19203_;
 wire _19204_;
 wire _19205_;
 wire _19206_;
 wire _19207_;
 wire _19208_;
 wire _19209_;
 wire _19210_;
 wire _19211_;
 wire _19212_;
 wire _19213_;
 wire _19214_;
 wire _19215_;
 wire net839;
 wire _19217_;
 wire _19218_;
 wire _19219_;
 wire _19220_;
 wire _19221_;
 wire _19222_;
 wire _19223_;
 wire _19224_;
 wire _19225_;
 wire _19226_;
 wire _19227_;
 wire net838;
 wire _19229_;
 wire _19230_;
 wire _19231_;
 wire _19232_;
 wire _19233_;
 wire _19234_;
 wire net837;
 wire _19236_;
 wire _19237_;
 wire _19238_;
 wire _19239_;
 wire _19240_;
 wire net836;
 wire _19242_;
 wire _19243_;
 wire _19244_;
 wire _19245_;
 wire _19246_;
 wire _19247_;
 wire _19248_;
 wire _19249_;
 wire _19250_;
 wire _19251_;
 wire _19252_;
 wire _19253_;
 wire _19254_;
 wire _19255_;
 wire _19256_;
 wire _19257_;
 wire _19258_;
 wire _19259_;
 wire net835;
 wire net834;
 wire _19262_;
 wire _19263_;
 wire net833;
 wire _19265_;
 wire _19266_;
 wire _19267_;
 wire net832;
 wire _19269_;
 wire _19270_;
 wire net831;
 wire net830;
 wire _19273_;
 wire _19274_;
 wire _19275_;
 wire _19276_;
 wire _19277_;
 wire _19278_;
 wire _19279_;
 wire _19280_;
 wire _19281_;
 wire _19282_;
 wire _19283_;
 wire _19284_;
 wire _19285_;
 wire _19286_;
 wire _19287_;
 wire _19288_;
 wire _19289_;
 wire _19290_;
 wire _19291_;
 wire _19292_;
 wire _19293_;
 wire _19294_;
 wire _19295_;
 wire _19296_;
 wire _19297_;
 wire _19298_;
 wire _19299_;
 wire _19300_;
 wire _19301_;
 wire _19302_;
 wire _19303_;
 wire _19304_;
 wire _19305_;
 wire _19306_;
 wire _19307_;
 wire _19308_;
 wire _19309_;
 wire _19310_;
 wire _19311_;
 wire _19312_;
 wire _19313_;
 wire _19314_;
 wire _19315_;
 wire _19316_;
 wire _19317_;
 wire _19318_;
 wire _19319_;
 wire _19320_;
 wire _19321_;
 wire _19322_;
 wire _19323_;
 wire _19324_;
 wire _19325_;
 wire _19326_;
 wire _19327_;
 wire _19328_;
 wire _19329_;
 wire _19330_;
 wire _19331_;
 wire _19332_;
 wire _19333_;
 wire _19334_;
 wire _19335_;
 wire _19336_;
 wire _19337_;
 wire _19338_;
 wire _19339_;
 wire _19340_;
 wire _19341_;
 wire _19342_;
 wire _19343_;
 wire _19344_;
 wire _19345_;
 wire _19346_;
 wire _19347_;
 wire _19348_;
 wire _19349_;
 wire _19350_;
 wire _19351_;
 wire _19352_;
 wire _19353_;
 wire _19354_;
 wire _19355_;
 wire _19356_;
 wire _19357_;
 wire _19358_;
 wire _19359_;
 wire _19360_;
 wire _19361_;
 wire _19362_;
 wire _19363_;
 wire _19364_;
 wire _19365_;
 wire _19366_;
 wire _19367_;
 wire _19368_;
 wire _19369_;
 wire _19370_;
 wire _19371_;
 wire _19372_;
 wire _19373_;
 wire _19374_;
 wire _19375_;
 wire _19376_;
 wire _19377_;
 wire _19378_;
 wire _19379_;
 wire _19380_;
 wire _19381_;
 wire _19382_;
 wire _19383_;
 wire _19384_;
 wire _19385_;
 wire _19386_;
 wire _19387_;
 wire _19388_;
 wire _19389_;
 wire _19390_;
 wire _19391_;
 wire _19392_;
 wire _19393_;
 wire _19394_;
 wire _19395_;
 wire _19396_;
 wire _19397_;
 wire _19398_;
 wire _19399_;
 wire _19400_;
 wire _19401_;
 wire _19402_;
 wire _19403_;
 wire _19404_;
 wire _19405_;
 wire _19406_;
 wire _19407_;
 wire _19408_;
 wire _19409_;
 wire _19410_;
 wire _19411_;
 wire _19412_;
 wire _19413_;
 wire _19414_;
 wire _19415_;
 wire _19416_;
 wire _19417_;
 wire _19418_;
 wire _19419_;
 wire _19420_;
 wire _19421_;
 wire _19422_;
 wire _19423_;
 wire _19424_;
 wire _19425_;
 wire _19426_;
 wire _19427_;
 wire _19428_;
 wire _19429_;
 wire _19430_;
 wire _19431_;
 wire _19432_;
 wire _19433_;
 wire _19434_;
 wire _19435_;
 wire _19436_;
 wire _19437_;
 wire _19438_;
 wire _19439_;
 wire _19440_;
 wire _19441_;
 wire _19442_;
 wire _19443_;
 wire _19444_;
 wire _19445_;
 wire _19446_;
 wire _19447_;
 wire _19448_;
 wire _19449_;
 wire _19450_;
 wire _19451_;
 wire _19452_;
 wire _19453_;
 wire _19454_;
 wire _19455_;
 wire _19456_;
 wire _19457_;
 wire _19458_;
 wire _19459_;
 wire _19460_;
 wire _19461_;
 wire _19462_;
 wire _19463_;
 wire _19464_;
 wire _19465_;
 wire _19466_;
 wire _19467_;
 wire _19468_;
 wire _19469_;
 wire _19470_;
 wire _19471_;
 wire _19472_;
 wire _19473_;
 wire _19474_;
 wire _19475_;
 wire _19476_;
 wire _19477_;
 wire _19478_;
 wire _19479_;
 wire _19480_;
 wire _19481_;
 wire _19482_;
 wire _19483_;
 wire _19484_;
 wire _19485_;
 wire _19486_;
 wire _19487_;
 wire _19488_;
 wire _19489_;
 wire _19490_;
 wire _19491_;
 wire _19492_;
 wire _19493_;
 wire _19494_;
 wire _19495_;
 wire _19496_;
 wire _19497_;
 wire _19498_;
 wire _19499_;
 wire _19500_;
 wire _19501_;
 wire _19502_;
 wire _19503_;
 wire _19504_;
 wire _19505_;
 wire _19506_;
 wire _19507_;
 wire _19508_;
 wire _19509_;
 wire _19510_;
 wire _19511_;
 wire net829;
 wire _19513_;
 wire _19514_;
 wire _19515_;
 wire _19516_;
 wire _19517_;
 wire _19518_;
 wire _19519_;
 wire _19520_;
 wire _19521_;
 wire _19522_;
 wire _19523_;
 wire _19524_;
 wire _19525_;
 wire _19526_;
 wire _19527_;
 wire _19528_;
 wire _19529_;
 wire _19530_;
 wire _19531_;
 wire _19532_;
 wire _19533_;
 wire _19534_;
 wire _19535_;
 wire _19536_;
 wire _19537_;
 wire _19538_;
 wire _19539_;
 wire _19540_;
 wire _19541_;
 wire _19542_;
 wire _19543_;
 wire _19544_;
 wire _19545_;
 wire _19546_;
 wire _19547_;
 wire _19548_;
 wire _19549_;
 wire _19550_;
 wire _19551_;
 wire _19552_;
 wire _19553_;
 wire _19554_;
 wire _19555_;
 wire _19556_;
 wire _19557_;
 wire _19558_;
 wire _19559_;
 wire _19560_;
 wire _19561_;
 wire _19562_;
 wire _19563_;
 wire _19564_;
 wire _19565_;
 wire _19566_;
 wire _19567_;
 wire _19568_;
 wire _19569_;
 wire _19570_;
 wire _19571_;
 wire _19572_;
 wire _19573_;
 wire _19574_;
 wire _19575_;
 wire _19576_;
 wire _19577_;
 wire _19578_;
 wire _19579_;
 wire _19580_;
 wire _19581_;
 wire _19582_;
 wire net828;
 wire net827;
 wire _19585_;
 wire _19586_;
 wire _19587_;
 wire _19588_;
 wire _19589_;
 wire net826;
 wire _19591_;
 wire _19592_;
 wire _19593_;
 wire _19594_;
 wire _19595_;
 wire _19596_;
 wire _19597_;
 wire _19598_;
 wire _19599_;
 wire _19600_;
 wire _19601_;
 wire _19602_;
 wire _19603_;
 wire _19604_;
 wire _19605_;
 wire _19606_;
 wire _19607_;
 wire _19608_;
 wire _19609_;
 wire _19610_;
 wire _19611_;
 wire _19612_;
 wire _19613_;
 wire _19614_;
 wire _19615_;
 wire _19616_;
 wire _19617_;
 wire _19618_;
 wire _19619_;
 wire _19620_;
 wire _19621_;
 wire _19622_;
 wire _19623_;
 wire _19624_;
 wire _19625_;
 wire _19626_;
 wire _19627_;
 wire _19628_;
 wire _19629_;
 wire _19630_;
 wire _19631_;
 wire _19632_;
 wire _19633_;
 wire _19634_;
 wire _19635_;
 wire _19636_;
 wire _19637_;
 wire _19638_;
 wire _19639_;
 wire _19640_;
 wire _19641_;
 wire _19642_;
 wire _19643_;
 wire _19644_;
 wire _19645_;
 wire _19646_;
 wire _19647_;
 wire _19648_;
 wire _19649_;
 wire _19650_;
 wire _19651_;
 wire _19652_;
 wire _19653_;
 wire _19654_;
 wire _19655_;
 wire _19656_;
 wire _19657_;
 wire _19658_;
 wire _19659_;
 wire _19660_;
 wire _19661_;
 wire _19662_;
 wire _19663_;
 wire _19664_;
 wire _19665_;
 wire _19666_;
 wire _19667_;
 wire _19668_;
 wire _19669_;
 wire _19670_;
 wire _19671_;
 wire _19672_;
 wire _19673_;
 wire _19674_;
 wire _19675_;
 wire _19676_;
 wire _19677_;
 wire _19678_;
 wire _19679_;
 wire _19680_;
 wire _19681_;
 wire _19682_;
 wire net825;
 wire _19684_;
 wire _19685_;
 wire _19686_;
 wire _19687_;
 wire _19688_;
 wire _19689_;
 wire _19690_;
 wire _19691_;
 wire _19692_;
 wire _19693_;
 wire _19694_;
 wire _19695_;
 wire _19696_;
 wire _19697_;
 wire _19698_;
 wire _19699_;
 wire _19700_;
 wire _19701_;
 wire _19702_;
 wire _19703_;
 wire _19704_;
 wire _19705_;
 wire _19706_;
 wire _19707_;
 wire _19708_;
 wire _19709_;
 wire _19710_;
 wire _19711_;
 wire _19712_;
 wire _19713_;
 wire _19714_;
 wire _19715_;
 wire _19716_;
 wire _19717_;
 wire _19718_;
 wire net824;
 wire _19720_;
 wire _19721_;
 wire _19722_;
 wire _19723_;
 wire _19724_;
 wire _19725_;
 wire _19726_;
 wire _19727_;
 wire _19728_;
 wire _19729_;
 wire _19730_;
 wire _19731_;
 wire _19732_;
 wire _19733_;
 wire _19734_;
 wire _19735_;
 wire _19736_;
 wire _19737_;
 wire _19738_;
 wire _19739_;
 wire _19740_;
 wire _19741_;
 wire _19742_;
 wire _19743_;
 wire _19744_;
 wire _19745_;
 wire _19746_;
 wire _19747_;
 wire _19748_;
 wire _19749_;
 wire _19750_;
 wire _19751_;
 wire _19752_;
 wire _19753_;
 wire _19754_;
 wire _19755_;
 wire _19756_;
 wire _19757_;
 wire _19758_;
 wire _19759_;
 wire _19760_;
 wire _19761_;
 wire _19762_;
 wire _19763_;
 wire _19764_;
 wire _19765_;
 wire _19766_;
 wire _19767_;
 wire _19768_;
 wire _19769_;
 wire _19770_;
 wire _19771_;
 wire _19772_;
 wire _19773_;
 wire _19774_;
 wire _19775_;
 wire _19776_;
 wire _19777_;
 wire _19778_;
 wire _19779_;
 wire _19780_;
 wire _19781_;
 wire _19782_;
 wire _19783_;
 wire _19784_;
 wire _19785_;
 wire _19786_;
 wire _19787_;
 wire _19788_;
 wire _19789_;
 wire _19790_;
 wire _19791_;
 wire _19792_;
 wire _19793_;
 wire _19794_;
 wire _19795_;
 wire _19796_;
 wire _19797_;
 wire _19798_;
 wire _19799_;
 wire _19800_;
 wire _19801_;
 wire _19802_;
 wire _19803_;
 wire _19804_;
 wire _19805_;
 wire _19806_;
 wire _19807_;
 wire _19808_;
 wire _19809_;
 wire _19810_;
 wire _19811_;
 wire _19812_;
 wire _19813_;
 wire _19814_;
 wire _19815_;
 wire _19816_;
 wire _19817_;
 wire _19818_;
 wire _19819_;
 wire _19820_;
 wire _19821_;
 wire _19822_;
 wire _19823_;
 wire _19824_;
 wire _19825_;
 wire _19826_;
 wire _19827_;
 wire _19828_;
 wire _19829_;
 wire _19830_;
 wire _19831_;
 wire _19832_;
 wire _19833_;
 wire _19834_;
 wire _19835_;
 wire _19836_;
 wire _19837_;
 wire _19838_;
 wire _19839_;
 wire _19840_;
 wire _19841_;
 wire _19842_;
 wire _19843_;
 wire _19844_;
 wire _19845_;
 wire _19846_;
 wire _19847_;
 wire _19848_;
 wire _19849_;
 wire _19850_;
 wire _19851_;
 wire _19852_;
 wire _19853_;
 wire _19854_;
 wire _19855_;
 wire _19856_;
 wire _19857_;
 wire _19858_;
 wire _19859_;
 wire _19860_;
 wire _19861_;
 wire _19862_;
 wire _19863_;
 wire _19864_;
 wire _19865_;
 wire _19866_;
 wire _19867_;
 wire _19868_;
 wire _19869_;
 wire _19870_;
 wire _19871_;
 wire _19872_;
 wire _19873_;
 wire _19874_;
 wire _19875_;
 wire _19876_;
 wire _19877_;
 wire _19878_;
 wire _19879_;
 wire _19880_;
 wire _19881_;
 wire _19882_;
 wire _19883_;
 wire _19884_;
 wire _19885_;
 wire _19886_;
 wire _19887_;
 wire _19888_;
 wire _19889_;
 wire _19890_;
 wire _19891_;
 wire _19892_;
 wire _19893_;
 wire _19894_;
 wire _19895_;
 wire _19896_;
 wire _19897_;
 wire _19898_;
 wire _19899_;
 wire _19900_;
 wire _19901_;
 wire _19902_;
 wire _19903_;
 wire _19904_;
 wire _19905_;
 wire _19906_;
 wire _19907_;
 wire _19908_;
 wire _19909_;
 wire _19910_;
 wire _19911_;
 wire _19912_;
 wire _19913_;
 wire _19914_;
 wire _19915_;
 wire _19916_;
 wire _19917_;
 wire _19918_;
 wire _19919_;
 wire _19920_;
 wire _19921_;
 wire _19922_;
 wire _19923_;
 wire _19924_;
 wire _19925_;
 wire _19926_;
 wire _19927_;
 wire _19928_;
 wire _19929_;
 wire _19930_;
 wire _19931_;
 wire _19932_;
 wire _19933_;
 wire _19934_;
 wire _19935_;
 wire _19936_;
 wire _19937_;
 wire _19938_;
 wire _19939_;
 wire _19940_;
 wire _19941_;
 wire _19942_;
 wire _19943_;
 wire _19944_;
 wire _19945_;
 wire _19946_;
 wire _19947_;
 wire _19948_;
 wire _19949_;
 wire _19950_;
 wire _19951_;
 wire _19952_;
 wire _19953_;
 wire _19954_;
 wire _19955_;
 wire _19956_;
 wire _19957_;
 wire _19958_;
 wire _19959_;
 wire _19960_;
 wire _19961_;
 wire _19962_;
 wire _19963_;
 wire _19964_;
 wire _19965_;
 wire _19966_;
 wire _19967_;
 wire _19968_;
 wire _19969_;
 wire _19970_;
 wire _19971_;
 wire _19972_;
 wire _19973_;
 wire _19974_;
 wire _19975_;
 wire _19976_;
 wire _19977_;
 wire _19978_;
 wire _19979_;
 wire _19980_;
 wire _19981_;
 wire _19982_;
 wire _19983_;
 wire _19984_;
 wire _19985_;
 wire _19986_;
 wire _19987_;
 wire _19988_;
 wire _19989_;
 wire _19990_;
 wire _19991_;
 wire _19992_;
 wire _19993_;
 wire _19994_;
 wire _19995_;
 wire _19996_;
 wire _19997_;
 wire _19998_;
 wire _19999_;
 wire _20000_;
 wire _20001_;
 wire _20002_;
 wire _20003_;
 wire _20004_;
 wire _20005_;
 wire _20006_;
 wire _20007_;
 wire _20008_;
 wire _20009_;
 wire _20010_;
 wire _20011_;
 wire _20012_;
 wire _20013_;
 wire _20014_;
 wire _20015_;
 wire _20016_;
 wire _20017_;
 wire _20018_;
 wire _20019_;
 wire _20020_;
 wire _20021_;
 wire _20022_;
 wire _20023_;
 wire _20024_;
 wire _20025_;
 wire _20026_;
 wire _20027_;
 wire _20028_;
 wire _20029_;
 wire _20030_;
 wire _20031_;
 wire _20032_;
 wire _20033_;
 wire _20034_;
 wire _20035_;
 wire _20036_;
 wire _20037_;
 wire _20038_;
 wire _20039_;
 wire _20040_;
 wire _20041_;
 wire _20042_;
 wire _20043_;
 wire _20044_;
 wire _20045_;
 wire _20046_;
 wire _20047_;
 wire _20048_;
 wire _20049_;
 wire _20050_;
 wire _20051_;
 wire _20052_;
 wire _20053_;
 wire _20054_;
 wire _20055_;
 wire _20056_;
 wire _20057_;
 wire _20058_;
 wire _20059_;
 wire _20060_;
 wire _20061_;
 wire _20062_;
 wire _20063_;
 wire _20064_;
 wire _20065_;
 wire _20066_;
 wire _20067_;
 wire _20068_;
 wire _20069_;
 wire _20070_;
 wire _20071_;
 wire _20072_;
 wire _20073_;
 wire _20074_;
 wire _20075_;
 wire _20076_;
 wire _20077_;
 wire _20078_;
 wire _20079_;
 wire _20080_;
 wire _20081_;
 wire net823;
 wire _20083_;
 wire _20084_;
 wire _20085_;
 wire _20086_;
 wire _20087_;
 wire _20088_;
 wire _20089_;
 wire _20090_;
 wire _20091_;
 wire _20092_;
 wire _20093_;
 wire _20094_;
 wire _20095_;
 wire _20096_;
 wire _20097_;
 wire _20098_;
 wire _20099_;
 wire _20100_;
 wire _20101_;
 wire _20102_;
 wire _20103_;
 wire _20104_;
 wire _20105_;
 wire _20106_;
 wire _20107_;
 wire _20108_;
 wire _20109_;
 wire _20110_;
 wire _20111_;
 wire _20112_;
 wire _20113_;
 wire _20114_;
 wire _20115_;
 wire _20116_;
 wire _20117_;
 wire _20118_;
 wire _20119_;
 wire _20120_;
 wire _20121_;
 wire _20122_;
 wire _20123_;
 wire _20124_;
 wire _20125_;
 wire _20126_;
 wire _20127_;
 wire _20128_;
 wire _20129_;
 wire _20130_;
 wire _20131_;
 wire _20132_;
 wire _20133_;
 wire _20134_;
 wire _20135_;
 wire _20136_;
 wire _20137_;
 wire _20138_;
 wire _20139_;
 wire _20140_;
 wire _20141_;
 wire _20142_;
 wire _20143_;
 wire _20144_;
 wire _20145_;
 wire _20146_;
 wire _20147_;
 wire _20148_;
 wire _20149_;
 wire _20150_;
 wire _20151_;
 wire _20152_;
 wire _20153_;
 wire _20154_;
 wire _20155_;
 wire _20156_;
 wire _20157_;
 wire _20158_;
 wire _20159_;
 wire _20160_;
 wire _20161_;
 wire _20162_;
 wire _20163_;
 wire _20164_;
 wire _20165_;
 wire _20166_;
 wire _20167_;
 wire _20168_;
 wire _20169_;
 wire _20170_;
 wire _20171_;
 wire _20172_;
 wire _20173_;
 wire _20174_;
 wire _20175_;
 wire _20176_;
 wire _20177_;
 wire _20178_;
 wire _20179_;
 wire _20180_;
 wire _20181_;
 wire _20182_;
 wire _20183_;
 wire net822;
 wire _20185_;
 wire _20186_;
 wire _20187_;
 wire _20188_;
 wire _20189_;
 wire _20190_;
 wire _20191_;
 wire _20192_;
 wire _20193_;
 wire _20194_;
 wire _20195_;
 wire _20196_;
 wire _20197_;
 wire _20198_;
 wire _20199_;
 wire _20200_;
 wire _20201_;
 wire _20202_;
 wire _20203_;
 wire _20204_;
 wire _20205_;
 wire _20206_;
 wire _20207_;
 wire _20208_;
 wire _20209_;
 wire _20210_;
 wire _20211_;
 wire _20212_;
 wire _20213_;
 wire _20214_;
 wire _20215_;
 wire _20216_;
 wire _20217_;
 wire _20218_;
 wire _20219_;
 wire _20220_;
 wire _20221_;
 wire _20222_;
 wire _20223_;
 wire _20224_;
 wire _20225_;
 wire _20226_;
 wire _20227_;
 wire _20228_;
 wire _20229_;
 wire _20230_;
 wire _20231_;
 wire _20232_;
 wire _20233_;
 wire _20234_;
 wire _20235_;
 wire _20236_;
 wire _20237_;
 wire _20238_;
 wire _20239_;
 wire _20240_;
 wire _20241_;
 wire _20242_;
 wire _20243_;
 wire _20244_;
 wire _20245_;
 wire _20246_;
 wire _20247_;
 wire _20248_;
 wire _20249_;
 wire _20250_;
 wire _20251_;
 wire _20252_;
 wire _20253_;
 wire _20254_;
 wire _20255_;
 wire _20256_;
 wire _20257_;
 wire _20258_;
 wire _20259_;
 wire _20260_;
 wire _20261_;
 wire _20262_;
 wire _20263_;
 wire _20264_;
 wire _20265_;
 wire _20266_;
 wire _20267_;
 wire _20268_;
 wire _20269_;
 wire _20270_;
 wire _20271_;
 wire _20272_;
 wire _20273_;
 wire _20274_;
 wire _20275_;
 wire _20276_;
 wire _20277_;
 wire _20278_;
 wire _20279_;
 wire _20280_;
 wire _20281_;
 wire _20282_;
 wire _20283_;
 wire _20284_;
 wire _20285_;
 wire _20286_;
 wire _20287_;
 wire _20288_;
 wire _20289_;
 wire _20290_;
 wire _20291_;
 wire _20292_;
 wire _20293_;
 wire _20294_;
 wire _20295_;
 wire _20296_;
 wire _20297_;
 wire _20298_;
 wire _20299_;
 wire _20300_;
 wire _20301_;
 wire _20302_;
 wire _20303_;
 wire _20304_;
 wire _20305_;
 wire _20306_;
 wire _20307_;
 wire _20308_;
 wire _20309_;
 wire _20310_;
 wire _20311_;
 wire _20312_;
 wire _20313_;
 wire _20314_;
 wire _20315_;
 wire _20316_;
 wire _20317_;
 wire _20318_;
 wire _20319_;
 wire _20320_;
 wire _20321_;
 wire _20322_;
 wire _20323_;
 wire _20324_;
 wire _20325_;
 wire _20326_;
 wire _20327_;
 wire _20328_;
 wire _20329_;
 wire _20330_;
 wire _20331_;
 wire _20332_;
 wire _20333_;
 wire _20334_;
 wire _20335_;
 wire _20336_;
 wire _20337_;
 wire _20338_;
 wire _20339_;
 wire _20340_;
 wire _20341_;
 wire _20342_;
 wire _20343_;
 wire _20344_;
 wire _20345_;
 wire _20346_;
 wire _20347_;
 wire _20348_;
 wire _20349_;
 wire _20350_;
 wire _20351_;
 wire _20352_;
 wire _20353_;
 wire _20354_;
 wire _20355_;
 wire _20356_;
 wire _20357_;
 wire _20358_;
 wire _20359_;
 wire _20360_;
 wire _20361_;
 wire _20362_;
 wire _20363_;
 wire _20364_;
 wire _20365_;
 wire _20366_;
 wire _20367_;
 wire _20368_;
 wire _20369_;
 wire _20370_;
 wire _20371_;
 wire _20372_;
 wire _20373_;
 wire _20374_;
 wire _20375_;
 wire _20376_;
 wire _20377_;
 wire _20378_;
 wire _20379_;
 wire _20380_;
 wire _20381_;
 wire _20382_;
 wire _20383_;
 wire _20384_;
 wire _20385_;
 wire _20386_;
 wire _20387_;
 wire _20388_;
 wire _20389_;
 wire _20390_;
 wire _20391_;
 wire _20392_;
 wire _20393_;
 wire _20394_;
 wire _20395_;
 wire _20396_;
 wire _20397_;
 wire _20398_;
 wire _20399_;
 wire _20400_;
 wire _20401_;
 wire _20402_;
 wire _20403_;
 wire _20404_;
 wire _20405_;
 wire _20406_;
 wire _20407_;
 wire _20408_;
 wire _20409_;
 wire _20410_;
 wire _20411_;
 wire _20412_;
 wire _20413_;
 wire _20414_;
 wire _20415_;
 wire _20416_;
 wire _20417_;
 wire _20418_;
 wire _20419_;
 wire _20420_;
 wire _20421_;
 wire _20422_;
 wire _20423_;
 wire _20424_;
 wire _20425_;
 wire _20426_;
 wire _20427_;
 wire _20428_;
 wire _20429_;
 wire _20430_;
 wire _20431_;
 wire _20432_;
 wire _20433_;
 wire _20434_;
 wire _20435_;
 wire _20436_;
 wire _20437_;
 wire _20438_;
 wire _20439_;
 wire _20440_;
 wire _20441_;
 wire _20442_;
 wire _20443_;
 wire _20444_;
 wire _20445_;
 wire _20446_;
 wire _20447_;
 wire _20448_;
 wire _20449_;
 wire _20450_;
 wire _20451_;
 wire net821;
 wire net820;
 wire _20454_;
 wire _20455_;
 wire _20456_;
 wire _20457_;
 wire _20458_;
 wire _20459_;
 wire _20460_;
 wire _20461_;
 wire _20462_;
 wire _20463_;
 wire _20464_;
 wire _20465_;
 wire _20466_;
 wire _20467_;
 wire _20468_;
 wire _20469_;
 wire _20470_;
 wire _20471_;
 wire _20472_;
 wire _20473_;
 wire _20474_;
 wire _20475_;
 wire _20476_;
 wire _20477_;
 wire _20478_;
 wire _20479_;
 wire _20480_;
 wire _20481_;
 wire _20482_;
 wire _20483_;
 wire _20484_;
 wire _20485_;
 wire _20486_;
 wire _20487_;
 wire _20488_;
 wire _20489_;
 wire _20490_;
 wire _20491_;
 wire _20492_;
 wire _20493_;
 wire _20494_;
 wire _20495_;
 wire _20496_;
 wire _20497_;
 wire _20498_;
 wire _20499_;
 wire _20500_;
 wire _20501_;
 wire _20502_;
 wire _20503_;
 wire _20504_;
 wire _20505_;
 wire _20506_;
 wire _20507_;
 wire _20508_;
 wire _20509_;
 wire _20510_;
 wire _20511_;
 wire _20512_;
 wire _20513_;
 wire _20514_;
 wire _20515_;
 wire _20516_;
 wire _20517_;
 wire _20518_;
 wire _20519_;
 wire _20520_;
 wire _20521_;
 wire _20522_;
 wire _20523_;
 wire _20524_;
 wire _20525_;
 wire _20526_;
 wire _20527_;
 wire _20528_;
 wire _20529_;
 wire _20530_;
 wire _20531_;
 wire _20532_;
 wire _20533_;
 wire _20534_;
 wire _20535_;
 wire _20536_;
 wire _20537_;
 wire _20538_;
 wire _20539_;
 wire _20540_;
 wire _20541_;
 wire _20542_;
 wire _20543_;
 wire _20544_;
 wire _20545_;
 wire _20546_;
 wire _20547_;
 wire _20548_;
 wire _20549_;
 wire _20550_;
 wire _20551_;
 wire _20552_;
 wire _20553_;
 wire _20554_;
 wire _20555_;
 wire _20556_;
 wire _20557_;
 wire _20558_;
 wire _20559_;
 wire _20560_;
 wire _20561_;
 wire _20562_;
 wire _20563_;
 wire _20564_;
 wire _20565_;
 wire _20566_;
 wire _20567_;
 wire _20568_;
 wire _20569_;
 wire _20570_;
 wire _20571_;
 wire _20572_;
 wire _20573_;
 wire _20574_;
 wire _20575_;
 wire _20576_;
 wire _20577_;
 wire _20578_;
 wire _20579_;
 wire _20580_;
 wire _20581_;
 wire _20582_;
 wire _20583_;
 wire _20584_;
 wire _20585_;
 wire _20586_;
 wire _20587_;
 wire _20588_;
 wire _20589_;
 wire _20590_;
 wire _20591_;
 wire _20592_;
 wire _20593_;
 wire _20594_;
 wire _20595_;
 wire _20596_;
 wire _20597_;
 wire _20598_;
 wire _20599_;
 wire _20600_;
 wire _20601_;
 wire _20602_;
 wire _20603_;
 wire _20604_;
 wire _20605_;
 wire _20606_;
 wire _20607_;
 wire _20608_;
 wire _20609_;
 wire _20610_;
 wire _20611_;
 wire _20612_;
 wire _20613_;
 wire _20614_;
 wire _20615_;
 wire _20616_;
 wire _20617_;
 wire _20618_;
 wire _20619_;
 wire _20620_;
 wire _20621_;
 wire _20622_;
 wire _20623_;
 wire _20624_;
 wire _20625_;
 wire _20626_;
 wire _20627_;
 wire _20628_;
 wire _20629_;
 wire _20630_;
 wire _20631_;
 wire _20632_;
 wire _20633_;
 wire _20634_;
 wire _20635_;
 wire _20636_;
 wire _20637_;
 wire _20638_;
 wire _20639_;
 wire _20640_;
 wire _20641_;
 wire _20642_;
 wire _20643_;
 wire _20644_;
 wire _20645_;
 wire _20646_;
 wire _20647_;
 wire _20648_;
 wire _20649_;
 wire _20650_;
 wire _20651_;
 wire _20652_;
 wire _20653_;
 wire _20654_;
 wire _20655_;
 wire _20656_;
 wire _20657_;
 wire _20658_;
 wire _20659_;
 wire _20660_;
 wire _20661_;
 wire _20662_;
 wire _20663_;
 wire _20664_;
 wire _20665_;
 wire _20666_;
 wire _20667_;
 wire _20668_;
 wire _20669_;
 wire _20670_;
 wire _20671_;
 wire _20672_;
 wire _20673_;
 wire _20674_;
 wire _20675_;
 wire _20676_;
 wire _20677_;
 wire _20678_;
 wire _20679_;
 wire _20680_;
 wire _20681_;
 wire _20682_;
 wire _20683_;
 wire _20684_;
 wire _20685_;
 wire _20686_;
 wire _20687_;
 wire _20688_;
 wire _20689_;
 wire _20690_;
 wire _20691_;
 wire _20692_;
 wire _20693_;
 wire _20694_;
 wire _20695_;
 wire _20696_;
 wire _20697_;
 wire _20698_;
 wire _20699_;
 wire _20700_;
 wire _20701_;
 wire _20702_;
 wire _20703_;
 wire _20704_;
 wire _20705_;
 wire _20706_;
 wire _20707_;
 wire _20708_;
 wire _20709_;
 wire _20710_;
 wire _20711_;
 wire _20712_;
 wire _20713_;
 wire _20714_;
 wire _20715_;
 wire _20716_;
 wire _20717_;
 wire _20718_;
 wire _20719_;
 wire _20720_;
 wire _20721_;
 wire _20722_;
 wire _20723_;
 wire _20724_;
 wire _20725_;
 wire _20726_;
 wire _20727_;
 wire _20728_;
 wire _20729_;
 wire _20730_;
 wire _20731_;
 wire _20732_;
 wire _20733_;
 wire _20734_;
 wire _20735_;
 wire _20736_;
 wire _20737_;
 wire _20738_;
 wire _20739_;
 wire _20740_;
 wire _20741_;
 wire _20742_;
 wire _20743_;
 wire _20744_;
 wire _20745_;
 wire _20746_;
 wire _20747_;
 wire _20748_;
 wire _20749_;
 wire _20750_;
 wire _20751_;
 wire _20752_;
 wire _20753_;
 wire _20754_;
 wire _20755_;
 wire _20756_;
 wire _20757_;
 wire _20758_;
 wire _20759_;
 wire _20760_;
 wire _20761_;
 wire _20762_;
 wire _20763_;
 wire _20764_;
 wire _20765_;
 wire _20766_;
 wire _20767_;
 wire _20768_;
 wire _20769_;
 wire _20770_;
 wire _20771_;
 wire _20772_;
 wire _20773_;
 wire _20774_;
 wire _20775_;
 wire _20776_;
 wire _20777_;
 wire _20778_;
 wire _20779_;
 wire _20780_;
 wire _20781_;
 wire _20782_;
 wire _20783_;
 wire _20784_;
 wire _20785_;
 wire _20786_;
 wire _20787_;
 wire _20788_;
 wire _20789_;
 wire _20790_;
 wire _20791_;
 wire _20792_;
 wire _20793_;
 wire _20794_;
 wire _20795_;
 wire _20796_;
 wire _20797_;
 wire _20798_;
 wire _20799_;
 wire _20800_;
 wire _20801_;
 wire _20802_;
 wire _20803_;
 wire _20804_;
 wire _20805_;
 wire _20806_;
 wire _20807_;
 wire _20808_;
 wire _20809_;
 wire _20810_;
 wire _20811_;
 wire _20812_;
 wire _20813_;
 wire _20814_;
 wire _20815_;
 wire _20816_;
 wire _20817_;
 wire _20818_;
 wire _20819_;
 wire _20820_;
 wire _20821_;
 wire _20822_;
 wire _20823_;
 wire _20824_;
 wire _20825_;
 wire _20826_;
 wire _20827_;
 wire _20828_;
 wire _20829_;
 wire _20830_;
 wire _20831_;
 wire _20832_;
 wire _20833_;
 wire _20834_;
 wire _20835_;
 wire _20836_;
 wire _20837_;
 wire _20838_;
 wire _20839_;
 wire _20840_;
 wire _20841_;
 wire _20842_;
 wire _20843_;
 wire _20844_;
 wire _20845_;
 wire _20846_;
 wire _20847_;
 wire _20848_;
 wire _20849_;
 wire _20850_;
 wire _20851_;
 wire _20852_;
 wire _20853_;
 wire _20854_;
 wire _20855_;
 wire _20856_;
 wire _20857_;
 wire _20858_;
 wire _20859_;
 wire _20860_;
 wire _20861_;
 wire _20862_;
 wire _20863_;
 wire _20864_;
 wire _20865_;
 wire _20866_;
 wire _20867_;
 wire _20868_;
 wire _20869_;
 wire _20870_;
 wire _20871_;
 wire _20872_;
 wire _20873_;
 wire _20874_;
 wire _20875_;
 wire _20876_;
 wire _20877_;
 wire _20878_;
 wire _20879_;
 wire _20880_;
 wire _20881_;
 wire _20882_;
 wire _20883_;
 wire _20884_;
 wire _20885_;
 wire _20886_;
 wire _20887_;
 wire _20888_;
 wire _20889_;
 wire _20890_;
 wire _20891_;
 wire _20892_;
 wire _20893_;
 wire _20894_;
 wire _20895_;
 wire _20896_;
 wire _20897_;
 wire _20898_;
 wire _20899_;
 wire _20900_;
 wire _20901_;
 wire _20902_;
 wire _20903_;
 wire _20904_;
 wire _20905_;
 wire _20906_;
 wire _20907_;
 wire _20908_;
 wire _20909_;
 wire _20910_;
 wire _20911_;
 wire _20912_;
 wire _20913_;
 wire _20914_;
 wire _20915_;
 wire _20916_;
 wire _20917_;
 wire _20918_;
 wire _20919_;
 wire _20920_;
 wire _20921_;
 wire _20922_;
 wire _20923_;
 wire _20924_;
 wire _20925_;
 wire _20926_;
 wire _20927_;
 wire _20928_;
 wire _20929_;
 wire _20930_;
 wire _20931_;
 wire _20932_;
 wire _20933_;
 wire _20934_;
 wire _20935_;
 wire _20936_;
 wire _20937_;
 wire _20938_;
 wire _20939_;
 wire _20940_;
 wire _20941_;
 wire _20942_;
 wire _20943_;
 wire _20944_;
 wire _20945_;
 wire _20946_;
 wire _20947_;
 wire _20948_;
 wire _20949_;
 wire _20950_;
 wire _20951_;
 wire _20952_;
 wire _20953_;
 wire _20954_;
 wire _20955_;
 wire _20956_;
 wire _20957_;
 wire _20958_;
 wire _20959_;
 wire _20960_;
 wire _20961_;
 wire _20962_;
 wire _20963_;
 wire _20964_;
 wire _20965_;
 wire _20966_;
 wire _20967_;
 wire _20968_;
 wire _20969_;
 wire _20970_;
 wire _20971_;
 wire _20972_;
 wire _20973_;
 wire _20974_;
 wire _20975_;
 wire _20976_;
 wire _20977_;
 wire _20978_;
 wire _20979_;
 wire _20980_;
 wire _20981_;
 wire _20982_;
 wire _20983_;
 wire _20984_;
 wire _20985_;
 wire _20986_;
 wire _20987_;
 wire _20988_;
 wire _20989_;
 wire _20990_;
 wire _20991_;
 wire _20992_;
 wire _20993_;
 wire _20994_;
 wire _20995_;
 wire _20996_;
 wire _20997_;
 wire _20998_;
 wire _20999_;
 wire _21000_;
 wire _21001_;
 wire _21002_;
 wire _21003_;
 wire _21004_;
 wire _21005_;
 wire _21006_;
 wire _21007_;
 wire _21008_;
 wire _21009_;
 wire _21010_;
 wire _21011_;
 wire _21012_;
 wire _21013_;
 wire _21014_;
 wire _21015_;
 wire _21016_;
 wire _21017_;
 wire _21018_;
 wire _21019_;
 wire _21020_;
 wire _21021_;
 wire _21022_;
 wire _21023_;
 wire _21024_;
 wire _21025_;
 wire _21026_;
 wire _21027_;
 wire _21028_;
 wire _21029_;
 wire _21030_;
 wire _21031_;
 wire _21032_;
 wire _21033_;
 wire _21034_;
 wire _21035_;
 wire _21036_;
 wire _21037_;
 wire _21038_;
 wire _21039_;
 wire _21040_;
 wire _21041_;
 wire _21042_;
 wire _21043_;
 wire _21044_;
 wire _21045_;
 wire _21046_;
 wire _21047_;
 wire _21048_;
 wire _21049_;
 wire _21050_;
 wire _21051_;
 wire _21052_;
 wire _21053_;
 wire _21054_;
 wire _21055_;
 wire _21056_;
 wire _21057_;
 wire _21058_;
 wire _21059_;
 wire _21060_;
 wire _21061_;
 wire _21062_;
 wire _21063_;
 wire _21064_;
 wire _21065_;
 wire _21066_;
 wire _21067_;
 wire _21068_;
 wire _21069_;
 wire _21070_;
 wire _21071_;
 wire _21072_;
 wire _21073_;
 wire _21074_;
 wire _21075_;
 wire _21076_;
 wire _21077_;
 wire _21078_;
 wire _21079_;
 wire _21080_;
 wire _21081_;
 wire _21082_;
 wire _21083_;
 wire _21084_;
 wire _21085_;
 wire _21086_;
 wire _21087_;
 wire _21088_;
 wire _21089_;
 wire _21090_;
 wire _21091_;
 wire _21092_;
 wire _21093_;
 wire _21094_;
 wire _21095_;
 wire _21096_;
 wire _21097_;
 wire _21098_;
 wire _21099_;
 wire _21100_;
 wire _21101_;
 wire _21102_;
 wire _21103_;
 wire _21104_;
 wire _21105_;
 wire _21106_;
 wire _21107_;
 wire _21108_;
 wire _21109_;
 wire _21110_;
 wire _21111_;
 wire _21112_;
 wire _21113_;
 wire _21114_;
 wire _21115_;
 wire _21116_;
 wire _21117_;
 wire _21118_;
 wire _21119_;
 wire _21120_;
 wire _21121_;
 wire _21122_;
 wire _21123_;
 wire _21124_;
 wire _21125_;
 wire _21126_;
 wire _21127_;
 wire _21128_;
 wire _21129_;
 wire _21130_;
 wire _21131_;
 wire _21132_;
 wire _21133_;
 wire _21134_;
 wire net819;
 wire _21136_;
 wire net818;
 wire _21138_;
 wire _21139_;
 wire _21140_;
 wire _21141_;
 wire _21142_;
 wire _21143_;
 wire _21144_;
 wire _21145_;
 wire _21146_;
 wire _21147_;
 wire _21148_;
 wire _21149_;
 wire _21150_;
 wire _21151_;
 wire _21152_;
 wire _21153_;
 wire _21154_;
 wire _21155_;
 wire _21156_;
 wire _21157_;
 wire _21158_;
 wire _21159_;
 wire _21160_;
 wire _21161_;
 wire _21162_;
 wire _21163_;
 wire _21164_;
 wire _21165_;
 wire _21166_;
 wire _21167_;
 wire _21168_;
 wire _21169_;
 wire _21170_;
 wire _21171_;
 wire _21172_;
 wire _21173_;
 wire _21174_;
 wire _21175_;
 wire _21176_;
 wire _21177_;
 wire _21178_;
 wire _21179_;
 wire _21180_;
 wire _21181_;
 wire _21182_;
 wire _21183_;
 wire _21184_;
 wire _21185_;
 wire _21186_;
 wire _21187_;
 wire _21188_;
 wire _21189_;
 wire _21190_;
 wire _21191_;
 wire _21192_;
 wire _21193_;
 wire _21194_;
 wire _21195_;
 wire _21196_;
 wire _21197_;
 wire _21198_;
 wire _21199_;
 wire _21200_;
 wire _21201_;
 wire _21202_;
 wire _21203_;
 wire _21204_;
 wire _21205_;
 wire _21206_;
 wire _21207_;
 wire _21208_;
 wire _21209_;
 wire _21210_;
 wire _21211_;
 wire _21212_;
 wire _21213_;
 wire _21214_;
 wire _21215_;
 wire _21216_;
 wire _21217_;
 wire _21218_;
 wire _21219_;
 wire _21220_;
 wire _21221_;
 wire _21222_;
 wire _21223_;
 wire _21224_;
 wire _21225_;
 wire _21226_;
 wire _21227_;
 wire _21228_;
 wire _21229_;
 wire _21230_;
 wire _21231_;
 wire _21232_;
 wire _21233_;
 wire _21234_;
 wire _21235_;
 wire _21236_;
 wire _21237_;
 wire _21238_;
 wire _21239_;
 wire _21240_;
 wire _21241_;
 wire _21242_;
 wire _21243_;
 wire _21244_;
 wire _21245_;
 wire _21246_;
 wire _21247_;
 wire _21248_;
 wire _21249_;
 wire _21250_;
 wire _21251_;
 wire _21252_;
 wire _21253_;
 wire _21254_;
 wire _21255_;
 wire _21256_;
 wire _21257_;
 wire _21258_;
 wire _21259_;
 wire _21260_;
 wire _21261_;
 wire _21262_;
 wire _21263_;
 wire _21264_;
 wire _21265_;
 wire _21266_;
 wire _21267_;
 wire _21268_;
 wire _21269_;
 wire _21270_;
 wire _21271_;
 wire _21272_;
 wire _21273_;
 wire _21274_;
 wire _21275_;
 wire _21276_;
 wire _21277_;
 wire _21278_;
 wire _21279_;
 wire _21280_;
 wire _21281_;
 wire _21282_;
 wire _21283_;
 wire _21284_;
 wire _21285_;
 wire _21286_;
 wire _21287_;
 wire _21288_;
 wire _21289_;
 wire _21290_;
 wire _21291_;
 wire _21292_;
 wire _21293_;
 wire _21294_;
 wire _21295_;
 wire _21296_;
 wire _21297_;
 wire _21298_;
 wire _21299_;
 wire _21300_;
 wire _21301_;
 wire _21302_;
 wire _21303_;
 wire _21304_;
 wire _21305_;
 wire _21306_;
 wire _21307_;
 wire _21308_;
 wire _21309_;
 wire _21310_;
 wire _21311_;
 wire _21312_;
 wire _21313_;
 wire _21314_;
 wire _21315_;
 wire _21316_;
 wire _21317_;
 wire _21318_;
 wire _21319_;
 wire _21320_;
 wire _21321_;
 wire _21322_;
 wire _21323_;
 wire _21324_;
 wire _21325_;
 wire _21326_;
 wire _21327_;
 wire _21328_;
 wire _21329_;
 wire _21330_;
 wire _21331_;
 wire _21332_;
 wire _21333_;
 wire _21334_;
 wire _21335_;
 wire _21336_;
 wire _21337_;
 wire _21338_;
 wire _21339_;
 wire _21340_;
 wire _21341_;
 wire _21342_;
 wire _21343_;
 wire _21344_;
 wire _21345_;
 wire _21346_;
 wire _21347_;
 wire _21348_;
 wire _21349_;
 wire _21350_;
 wire _21351_;
 wire _21352_;
 wire _21353_;
 wire _21354_;
 wire _21355_;
 wire _21356_;
 wire _21357_;
 wire _21358_;
 wire _21359_;
 wire _21360_;
 wire _21361_;
 wire _21362_;
 wire _21363_;
 wire _21364_;
 wire _21365_;
 wire _21366_;
 wire _21367_;
 wire _21368_;
 wire _21369_;
 wire _21370_;
 wire _21371_;
 wire _21372_;
 wire _21373_;
 wire _21374_;
 wire _21375_;
 wire _21376_;
 wire _21377_;
 wire _21378_;
 wire _21379_;
 wire _21380_;
 wire _21381_;
 wire _21382_;
 wire _21383_;
 wire _21384_;
 wire _21385_;
 wire _21386_;
 wire _21387_;
 wire _21388_;
 wire _21389_;
 wire _21390_;
 wire _21391_;
 wire _21392_;
 wire _21393_;
 wire _21394_;
 wire _21395_;
 wire _21396_;
 wire _21397_;
 wire _21398_;
 wire _21399_;
 wire _21400_;
 wire _21401_;
 wire _21402_;
 wire _21403_;
 wire _21404_;
 wire _21405_;
 wire _21406_;
 wire _21407_;
 wire _21408_;
 wire _21409_;
 wire _21410_;
 wire _21411_;
 wire _21412_;
 wire _21413_;
 wire _21414_;
 wire _21415_;
 wire _21416_;
 wire _21417_;
 wire _21418_;
 wire _21419_;
 wire _21420_;
 wire _21421_;
 wire _21422_;
 wire _21423_;
 wire _21424_;
 wire _21425_;
 wire _21426_;
 wire net817;
 wire _21428_;
 wire _21429_;
 wire _21430_;
 wire _21431_;
 wire _21432_;
 wire _21433_;
 wire _21434_;
 wire _21435_;
 wire _21436_;
 wire _21437_;
 wire _21438_;
 wire _21439_;
 wire _21440_;
 wire _21441_;
 wire _21442_;
 wire _21443_;
 wire _21444_;
 wire _21445_;
 wire _21446_;
 wire _21447_;
 wire _21448_;
 wire _21449_;
 wire _21450_;
 wire _21451_;
 wire _21452_;
 wire _21453_;
 wire _21454_;
 wire _21455_;
 wire _21456_;
 wire _21457_;
 wire _21458_;
 wire _21459_;
 wire _21460_;
 wire _21461_;
 wire _21462_;
 wire net816;
 wire _21464_;
 wire _21465_;
 wire _21466_;
 wire _21467_;
 wire _21468_;
 wire _21469_;
 wire _21470_;
 wire _21471_;
 wire _21472_;
 wire _21473_;
 wire _21474_;
 wire _21475_;
 wire _21476_;
 wire _21477_;
 wire net815;
 wire _21479_;
 wire _21480_;
 wire _21481_;
 wire net814;
 wire _21483_;
 wire _21484_;
 wire _21485_;
 wire _21486_;
 wire _21487_;
 wire _21488_;
 wire _21489_;
 wire _21490_;
 wire _21491_;
 wire _21492_;
 wire _21493_;
 wire net813;
 wire _21495_;
 wire _21496_;
 wire _21497_;
 wire _21498_;
 wire _21499_;
 wire _21500_;
 wire _21501_;
 wire _21502_;
 wire _21503_;
 wire _21504_;
 wire _21505_;
 wire _21506_;
 wire _21507_;
 wire _21508_;
 wire _21509_;
 wire _21510_;
 wire _21511_;
 wire _21512_;
 wire _21513_;
 wire _21514_;
 wire _21515_;
 wire _21516_;
 wire _21517_;
 wire _21518_;
 wire _21519_;
 wire _21520_;
 wire _21521_;
 wire _21522_;
 wire _21523_;
 wire _21524_;
 wire _21525_;
 wire _21526_;
 wire _21527_;
 wire _21528_;
 wire _21529_;
 wire _21530_;
 wire _21531_;
 wire _21532_;
 wire _21533_;
 wire _21534_;
 wire _21535_;
 wire _21536_;
 wire _21537_;
 wire _21538_;
 wire _21539_;
 wire _21540_;
 wire _21541_;
 wire _21542_;
 wire _21543_;
 wire _21544_;
 wire _21545_;
 wire _21546_;
 wire _21547_;
 wire _21548_;
 wire _21549_;
 wire _21550_;
 wire net812;
 wire _21552_;
 wire _21553_;
 wire _21554_;
 wire _21555_;
 wire _21556_;
 wire _21557_;
 wire _21558_;
 wire _21559_;
 wire _21560_;
 wire _21561_;
 wire _21562_;
 wire _21563_;
 wire _21564_;
 wire _21565_;
 wire _21566_;
 wire _21567_;
 wire _21568_;
 wire _21569_;
 wire _21570_;
 wire _21571_;
 wire _21572_;
 wire _21573_;
 wire _21574_;
 wire _21575_;
 wire net811;
 wire _21577_;
 wire _21578_;
 wire _21579_;
 wire _21580_;
 wire _21581_;
 wire _21582_;
 wire _21583_;
 wire _21584_;
 wire _21585_;
 wire _21586_;
 wire _21587_;
 wire _21588_;
 wire _21589_;
 wire _21590_;
 wire _21591_;
 wire _21592_;
 wire _21593_;
 wire _21594_;
 wire _21595_;
 wire _21596_;
 wire _21597_;
 wire _21598_;
 wire _21599_;
 wire _21600_;
 wire _21601_;
 wire _21602_;
 wire _21603_;
 wire _21604_;
 wire _21605_;
 wire _21606_;
 wire _21607_;
 wire _21608_;
 wire _21609_;
 wire _21610_;
 wire _21611_;
 wire _21612_;
 wire _21613_;
 wire _21614_;
 wire _21615_;
 wire _21616_;
 wire _21617_;
 wire _21618_;
 wire _21619_;
 wire _21620_;
 wire _21621_;
 wire _21622_;
 wire _21623_;
 wire _21624_;
 wire _21625_;
 wire _21626_;
 wire _21627_;
 wire _21628_;
 wire _21629_;
 wire _21630_;
 wire _21631_;
 wire _21632_;
 wire _21633_;
 wire _21634_;
 wire _21635_;
 wire _21636_;
 wire _21637_;
 wire _21638_;
 wire _21639_;
 wire _21640_;
 wire _21641_;
 wire _21642_;
 wire _21643_;
 wire _21644_;
 wire _21645_;
 wire _21646_;
 wire _21647_;
 wire _21648_;
 wire _21649_;
 wire _21650_;
 wire _21651_;
 wire _21652_;
 wire _21653_;
 wire _21654_;
 wire _21655_;
 wire _21656_;
 wire _21657_;
 wire _21658_;
 wire _21659_;
 wire _21660_;
 wire _21661_;
 wire _21662_;
 wire _21663_;
 wire _21664_;
 wire _21665_;
 wire _21666_;
 wire _21667_;
 wire _21668_;
 wire _21669_;
 wire _21670_;
 wire _21671_;
 wire _21672_;
 wire _21673_;
 wire _21674_;
 wire _21675_;
 wire _21676_;
 wire _21677_;
 wire _21678_;
 wire _21679_;
 wire _21680_;
 wire _21681_;
 wire _21682_;
 wire _21683_;
 wire _21684_;
 wire _21685_;
 wire _21686_;
 wire _21687_;
 wire _21688_;
 wire _21689_;
 wire net810;
 wire _21691_;
 wire _21692_;
 wire _21693_;
 wire _21694_;
 wire _21695_;
 wire _21696_;
 wire _21697_;
 wire _21698_;
 wire _21699_;
 wire _21700_;
 wire _21701_;
 wire _21702_;
 wire _21703_;
 wire _21704_;
 wire net809;
 wire _21706_;
 wire _21707_;
 wire net808;
 wire _21709_;
 wire _21710_;
 wire _21711_;
 wire _21712_;
 wire _21713_;
 wire _21714_;
 wire _21715_;
 wire _21716_;
 wire _21717_;
 wire net807;
 wire _21719_;
 wire _21720_;
 wire _21721_;
 wire _21722_;
 wire _21723_;
 wire _21724_;
 wire _21725_;
 wire _21726_;
 wire _21727_;
 wire _21728_;
 wire _21729_;
 wire _21730_;
 wire _21731_;
 wire _21732_;
 wire _21733_;
 wire _21734_;
 wire _21735_;
 wire _21736_;
 wire _21737_;
 wire _21738_;
 wire _21739_;
 wire _21740_;
 wire _21741_;
 wire _21742_;
 wire _21743_;
 wire _21744_;
 wire _21745_;
 wire net806;
 wire _21747_;
 wire _21748_;
 wire _21749_;
 wire _21750_;
 wire _21751_;
 wire _21752_;
 wire _21753_;
 wire _21754_;
 wire _21755_;
 wire _21756_;
 wire _21757_;
 wire _21758_;
 wire _21759_;
 wire _21760_;
 wire _21761_;
 wire _21762_;
 wire _21763_;
 wire _21764_;
 wire _21765_;
 wire _21766_;
 wire _21767_;
 wire _21768_;
 wire _21769_;
 wire _21770_;
 wire _21771_;
 wire _21772_;
 wire _21773_;
 wire _21774_;
 wire net805;
 wire _21776_;
 wire _21777_;
 wire _21778_;
 wire _21779_;
 wire _21780_;
 wire _21781_;
 wire _21782_;
 wire _21783_;
 wire _21784_;
 wire _21785_;
 wire _21786_;
 wire _21787_;
 wire _21788_;
 wire _21789_;
 wire _21790_;
 wire _21791_;
 wire _21792_;
 wire _21793_;
 wire _21794_;
 wire _21795_;
 wire net804;
 wire _21797_;
 wire _21798_;
 wire _21799_;
 wire _21800_;
 wire _21801_;
 wire _21802_;
 wire _21803_;
 wire _21804_;
 wire _21805_;
 wire _21806_;
 wire _21807_;
 wire _21808_;
 wire _21809_;
 wire _21810_;
 wire _21811_;
 wire _21812_;
 wire _21813_;
 wire _21814_;
 wire _21815_;
 wire _21816_;
 wire _21817_;
 wire _21818_;
 wire _21819_;
 wire _21820_;
 wire _21821_;
 wire _21822_;
 wire _21823_;
 wire _21824_;
 wire _21825_;
 wire _21826_;
 wire _21827_;
 wire _21828_;
 wire _21829_;
 wire _21830_;
 wire _21831_;
 wire _21832_;
 wire _21833_;
 wire _21834_;
 wire _21835_;
 wire _21836_;
 wire _21837_;
 wire _21838_;
 wire _21839_;
 wire _21840_;
 wire _21841_;
 wire _21842_;
 wire _21843_;
 wire _21844_;
 wire _21845_;
 wire _21846_;
 wire _21847_;
 wire _21848_;
 wire _21849_;
 wire _21850_;
 wire _21851_;
 wire _21852_;
 wire _21853_;
 wire _21854_;
 wire _21855_;
 wire _21856_;
 wire _21857_;
 wire _21858_;
 wire _21859_;
 wire _21860_;
 wire _21861_;
 wire _21862_;
 wire _21863_;
 wire _21864_;
 wire _21865_;
 wire net803;
 wire _21867_;
 wire _21868_;
 wire _21869_;
 wire net802;
 wire net801;
 wire _21872_;
 wire _21873_;
 wire net800;
 wire net799;
 wire _21876_;
 wire _21877_;
 wire _21878_;
 wire _21879_;
 wire net798;
 wire _21881_;
 wire net797;
 wire _21883_;
 wire _21884_;
 wire _21885_;
 wire _21886_;
 wire _21887_;
 wire _21888_;
 wire _21889_;
 wire _21890_;
 wire _21891_;
 wire _21892_;
 wire _21893_;
 wire _21894_;
 wire _21895_;
 wire net796;
 wire _21897_;
 wire _21898_;
 wire _21899_;
 wire _21900_;
 wire _21901_;
 wire net795;
 wire net794;
 wire _21904_;
 wire net793;
 wire net792;
 wire _21907_;
 wire _21908_;
 wire _21909_;
 wire _21910_;
 wire _21911_;
 wire _21912_;
 wire _21913_;
 wire _21914_;
 wire _21915_;
 wire _21916_;
 wire _21917_;
 wire _21918_;
 wire _21919_;
 wire _21920_;
 wire net791;
 wire _21922_;
 wire net790;
 wire _21924_;
 wire _21925_;
 wire _21926_;
 wire _21927_;
 wire net789;
 wire _21929_;
 wire net788;
 wire _21931_;
 wire _21932_;
 wire net787;
 wire _21934_;
 wire net786;
 wire _21936_;
 wire _21937_;
 wire _21938_;
 wire net785;
 wire _21940_;
 wire net784;
 wire _21942_;
 wire _21943_;
 wire _21944_;
 wire _21945_;
 wire net783;
 wire net782;
 wire net781;
 wire net780;
 wire _21950_;
 wire _21951_;
 wire _21952_;
 wire _21953_;
 wire _21954_;
 wire _21955_;
 wire _21956_;
 wire _21957_;
 wire _21958_;
 wire net779;
 wire _21960_;
 wire _21961_;
 wire _21962_;
 wire _21963_;
 wire _21964_;
 wire net778;
 wire _21966_;
 wire _21967_;
 wire net777;
 wire _21969_;
 wire net776;
 wire _21971_;
 wire _21972_;
 wire _21973_;
 wire _21974_;
 wire _21975_;
 wire _21976_;
 wire net775;
 wire _21978_;
 wire _21979_;
 wire _21980_;
 wire _21981_;
 wire _21982_;
 wire _21983_;
 wire net774;
 wire _21985_;
 wire net773;
 wire _21987_;
 wire _21988_;
 wire _21989_;
 wire _21990_;
 wire _21991_;
 wire _21992_;
 wire net772;
 wire _21994_;
 wire _21995_;
 wire _21996_;
 wire _21997_;
 wire net771;
 wire _21999_;
 wire _22000_;
 wire _22001_;
 wire _22002_;
 wire _22003_;
 wire _22004_;
 wire _22005_;
 wire _22006_;
 wire _22007_;
 wire _22008_;
 wire net770;
 wire _22010_;
 wire _22011_;
 wire _22012_;
 wire _22013_;
 wire _22014_;
 wire _22015_;
 wire _22016_;
 wire _22017_;
 wire _22018_;
 wire _22019_;
 wire net769;
 wire net768;
 wire _22022_;
 wire _22023_;
 wire _22024_;
 wire _22025_;
 wire _22026_;
 wire _22027_;
 wire _22028_;
 wire net767;
 wire net766;
 wire _22031_;
 wire _22032_;
 wire _22033_;
 wire _22034_;
 wire _22035_;
 wire net765;
 wire _22037_;
 wire _22038_;
 wire _22039_;
 wire _22040_;
 wire _22041_;
 wire _22042_;
 wire _22043_;
 wire _22044_;
 wire _22045_;
 wire _22046_;
 wire net764;
 wire _22048_;
 wire _22049_;
 wire net763;
 wire _22051_;
 wire _22052_;
 wire _22053_;
 wire _22054_;
 wire _22055_;
 wire _22056_;
 wire _22057_;
 wire net762;
 wire _22059_;
 wire _22060_;
 wire _22061_;
 wire _22062_;
 wire _22063_;
 wire _22064_;
 wire net761;
 wire net760;
 wire _22067_;
 wire _22068_;
 wire _22069_;
 wire _22070_;
 wire net759;
 wire net758;
 wire _22073_;
 wire _22074_;
 wire _22075_;
 wire _22076_;
 wire _22077_;
 wire net757;
 wire _22079_;
 wire _22080_;
 wire _22081_;
 wire _22082_;
 wire _22083_;
 wire _22084_;
 wire _22085_;
 wire _22086_;
 wire _22087_;
 wire _22088_;
 wire _22089_;
 wire _22090_;
 wire _22091_;
 wire _22092_;
 wire net756;
 wire _22094_;
 wire _22095_;
 wire _22096_;
 wire net755;
 wire _22098_;
 wire _22099_;
 wire _22100_;
 wire _22101_;
 wire _22102_;
 wire _22103_;
 wire _22104_;
 wire _22105_;
 wire _22106_;
 wire _22107_;
 wire \u0.r0.rcnt[0] ;
 wire \u0.r0.rcnt[1] ;
 wire \u0.r0.rcnt[2] ;
 wire \u0.r0.rcnt_next[0] ;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3164;
 wire net3165;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3965;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3973;
 wire net3974;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3983;
 wire net3984;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net3990;
 wire net3991;
 wire net3992;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net3999;
 wire net4000;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4004;
 wire net4005;
 wire net4006;
 wire net4007;
 wire net4008;
 wire net4009;
 wire net4010;
 wire net4011;
 wire net4012;
 wire net4013;
 wire net4014;
 wire net4015;
 wire net4016;
 wire net4017;
 wire net4018;
 wire net4019;
 wire net4020;
 wire net4021;
 wire net4022;
 wire net4023;
 wire net4024;
 wire net4025;
 wire net4026;
 wire net4027;
 wire net4028;
 wire net4029;
 wire net4030;
 wire net4031;
 wire net4032;
 wire net4033;
 wire net4034;
 wire net4035;
 wire net4036;
 wire net4037;
 wire net4038;
 wire net4039;
 wire net4040;
 wire net4041;
 wire net4042;
 wire net4043;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net4050;
 wire net4051;
 wire net4052;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4058;
 wire net4059;
 wire net4060;
 wire net4061;
 wire net4062;
 wire net4063;
 wire net4064;
 wire net4065;
 wire net4066;
 wire net4067;
 wire net4068;
 wire net4069;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net4075;
 wire net4076;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4083;
 wire net4084;
 wire net4085;
 wire net4086;
 wire net4087;
 wire net4088;
 wire net4089;
 wire net4090;
 wire net4091;
 wire net4092;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net4096;
 wire net4097;
 wire net4098;
 wire net4099;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4103;
 wire net4104;
 wire net4105;
 wire net4106;
 wire net4107;
 wire net4108;
 wire net4109;
 wire net4110;
 wire net4111;
 wire net4112;
 wire net4113;
 wire net4114;
 wire net4115;
 wire net4116;
 wire net4117;
 wire net4118;
 wire net4119;
 wire net4120;
 wire net4121;
 wire net4122;
 wire net4123;
 wire net4124;
 wire net4125;
 wire net4126;
 wire net4127;
 wire net4128;
 wire net4129;
 wire net4130;
 wire net4131;
 wire net4132;
 wire net4133;
 wire net4134;
 wire net4135;
 wire net4136;
 wire net4137;
 wire net4138;
 wire net4139;
 wire net4140;
 wire net4141;
 wire net4142;
 wire net4143;
 wire net4144;
 wire net4145;
 wire net4146;
 wire net4147;
 wire net4148;
 wire net4149;
 wire net4150;
 wire net4151;
 wire net4152;
 wire net4153;
 wire net4154;
 wire net4155;
 wire net4156;
 wire net4157;
 wire net4158;
 wire net4159;
 wire net4160;
 wire net4161;
 wire net4162;
 wire net4163;
 wire net4164;
 wire net4165;
 wire net4166;
 wire net4167;
 wire net4168;
 wire net4169;
 wire net4170;
 wire net4171;
 wire net4172;
 wire net4173;
 wire net4174;
 wire net4175;
 wire net4176;
 wire net4177;
 wire net4178;
 wire net4179;
 wire net4180;
 wire net4181;
 wire net4182;
 wire net4183;
 wire net4184;
 wire net4185;
 wire net4186;
 wire net4187;
 wire net4188;
 wire net4189;
 wire net4190;
 wire net4191;
 wire net4192;
 wire net4193;
 wire net4194;
 wire net4195;
 wire net4196;
 wire net4197;
 wire net4198;
 wire net4199;
 wire net4200;
 wire net4201;
 wire net4202;
 wire net4203;
 wire net4204;
 wire net4205;
 wire net4206;
 wire net4207;
 wire net4208;
 wire net4209;
 wire net4210;
 wire net4211;
 wire net4212;
 wire net4213;
 wire net4214;
 wire net4215;
 wire net4216;
 wire net4217;
 wire net4218;
 wire net4219;
 wire net4220;
 wire net4221;
 wire net4222;
 wire net4223;
 wire net4224;
 wire net4225;
 wire net4226;
 wire net4227;
 wire net4228;
 wire net4229;
 wire net4230;
 wire net4231;
 wire net4232;
 wire net4233;
 wire net4234;

 AND2x2_ASAP7_75t_R _22108_ (.A(_00786_),
    .B(_00787_),
    .Y(_22107_));
 INVx1_ASAP7_75t_R _22109_ (.A(_00917_),
    .Y(_22105_));
 INVx1_ASAP7_75t_R _98_128 (.A(clknet_leaf_14_clk),
    .Y(net533));
 INVx1_ASAP7_75t_R _98_127 (.A(clknet_leaf_14_clk),
    .Y(net532));
 NAND2x2_ASAP7_75t_R _22112_ (.A(net403),
    .B(net1),
    .Y(_05716_));
 INVx1_ASAP7_75t_R _98_126 (.A(clknet_leaf_14_clk),
    .Y(net531));
 INVx1_ASAP7_75t_R _98_125 (.A(clknet_leaf_15_clk),
    .Y(net530));
 INVx5_ASAP7_75t_R _22115_ (.A(_00424_),
    .Y(_05749_));
 NAND2x2_ASAP7_75t_R _22116_ (.A(_00423_),
    .B(_05749_),
    .Y(_05760_));
 INVx1_ASAP7_75t_R _98_124 (.A(clknet_leaf_15_clk),
    .Y(net529));
 AND2x4_ASAP7_75t_R _22118_ (.A(_00421_),
    .B(_00422_),
    .Y(_05782_));
 INVx3_ASAP7_75t_R _22119_ (.A(_05782_),
    .Y(_05793_));
 NOR2x2_ASAP7_75t_R _22120_ (.A(_05760_),
    .B(_05793_),
    .Y(_05804_));
 INVx1_ASAP7_75t_R _98_123 (.A(clknet_leaf_15_clk),
    .Y(net528));
 INVx1_ASAP7_75t_R _98_122 (.A(clknet_leaf_15_clk),
    .Y(net527));
 INVx1_ASAP7_75t_R _98_121 (.A(clknet_leaf_0_clk),
    .Y(net526));
 INVx2_ASAP7_75t_R _22124_ (.A(net3395),
    .Y(_05848_));
 NAND2x2_ASAP7_75t_R _22125_ (.A(net3402),
    .B(_05848_),
    .Y(_05859_));
 NAND2x2_ASAP7_75t_R _22126_ (.A(_00423_),
    .B(_00424_),
    .Y(_05870_));
 NOR2x2_ASAP7_75t_R _22127_ (.A(_05870_),
    .B(_05793_),
    .Y(_05881_));
 CKINVDCx6p67_ASAP7_75t_R _22128_ (.A(_05881_),
    .Y(_05892_));
 NAND2x2_ASAP7_75t_R _22129_ (.A(net3399),
    .B(net3395),
    .Y(_05903_));
 INVx1_ASAP7_75t_R _98_120 (.A(clknet_leaf_15_clk),
    .Y(net525));
 CKINVDCx9p33_ASAP7_75t_R _22131_ (.A(_00428_),
    .Y(_05925_));
 NAND2x2_ASAP7_75t_R _22132_ (.A(_00427_),
    .B(_05925_),
    .Y(_05936_));
 NOR2x2_ASAP7_75t_R _22133_ (.A(_05903_),
    .B(_05936_),
    .Y(_05947_));
 CKINVDCx10_ASAP7_75t_R _22134_ (.A(_05947_),
    .Y(_05958_));
 INVx1_ASAP7_75t_R _98_119 (.A(clknet_leaf_16_clk),
    .Y(net524));
 INVx1_ASAP7_75t_R _98_118 (.A(clknet_leaf_1_clk),
    .Y(net523));
 NOR2x2_ASAP7_75t_R _22137_ (.A(net1614),
    .B(net1654),
    .Y(_05991_));
 INVx2_ASAP7_75t_R _22138_ (.A(_05991_),
    .Y(_06002_));
 AO21x1_ASAP7_75t_R _22139_ (.A1(_05958_),
    .A2(_06002_),
    .B(_05892_),
    .Y(_06013_));
 OA21x2_ASAP7_75t_R _22140_ (.A1(net2858),
    .A2(_05892_),
    .B(_06013_),
    .Y(_06024_));
 INVx2_ASAP7_75t_R _22141_ (.A(_06024_),
    .Y(_06035_));
 NOR2x2_ASAP7_75t_R _22142_ (.A(net3399),
    .B(net3395),
    .Y(_06046_));
 CKINVDCx9p33_ASAP7_75t_R _22143_ (.A(_06046_),
    .Y(_06057_));
 INVx1_ASAP7_75t_R _98_117 (.A(clknet_leaf_2_clk),
    .Y(net522));
 NOR2x2_ASAP7_75t_R _22145_ (.A(net1614),
    .B(_06057_),
    .Y(_06079_));
 INVx3_ASAP7_75t_R _22146_ (.A(_06079_),
    .Y(_06090_));
 INVx1_ASAP7_75t_R _98_116 (.A(clknet_leaf_16_clk),
    .Y(net521));
 AND2x6_ASAP7_75t_R _22148_ (.A(net1614),
    .B(net2133),
    .Y(_06112_));
 NAND2x2_ASAP7_75t_R _22149_ (.A(_06046_),
    .B(_06112_),
    .Y(_06123_));
 INVx1_ASAP7_75t_R _22150_ (.A(_05936_),
    .Y(_06134_));
 NAND2x2_ASAP7_75t_R _22151_ (.A(_06046_),
    .B(_06134_),
    .Y(_06145_));
 AO21x1_ASAP7_75t_R _22152_ (.A1(_06123_),
    .A2(_06145_),
    .B(_05892_),
    .Y(_06156_));
 OA21x2_ASAP7_75t_R _22153_ (.A1(_05892_),
    .A2(_06090_),
    .B(_06156_),
    .Y(_06167_));
 INVx1_ASAP7_75t_R _22154_ (.A(_06167_),
    .Y(_06178_));
 INVx4_ASAP7_75t_R _22155_ (.A(net3399),
    .Y(_06189_));
 NAND2x2_ASAP7_75t_R _22156_ (.A(net3395),
    .B(_06189_),
    .Y(_06200_));
 NOR2x2_ASAP7_75t_R _22157_ (.A(net1615),
    .B(net1935),
    .Y(_06211_));
 CKINVDCx6p67_ASAP7_75t_R _22158_ (.A(_06211_),
    .Y(_06222_));
 INVx1_ASAP7_75t_R _98_115 (.A(clknet_leaf_6_clk),
    .Y(net520));
 NOR2x1_ASAP7_75t_R _22160_ (.A(_06222_),
    .B(_05892_),
    .Y(_06244_));
 NOR2x2_ASAP7_75t_R _22161_ (.A(net1012),
    .B(net1936),
    .Y(_06255_));
 INVx6_ASAP7_75t_R _22162_ (.A(_06200_),
    .Y(_06266_));
 NAND2x2_ASAP7_75t_R _22163_ (.A(_06112_),
    .B(_06266_),
    .Y(_06277_));
 NOR2x2_ASAP7_75t_R _22164_ (.A(_06277_),
    .B(_05892_),
    .Y(_06288_));
 AO21x1_ASAP7_75t_R _22165_ (.A1(_06255_),
    .A2(_05881_),
    .B(_06288_),
    .Y(_06299_));
 OR5x1_ASAP7_75t_R _22166_ (.A(_05804_),
    .B(_06035_),
    .C(_06178_),
    .D(_06244_),
    .E(_06299_),
    .Y(_06309_));
 INVx1_ASAP7_75t_R _98_114 (.A(clknet_leaf_6_clk),
    .Y(net519));
 INVx2_ASAP7_75t_R _22168_ (.A(_00421_),
    .Y(_06331_));
 CKINVDCx6p67_ASAP7_75t_R _22169_ (.A(_00422_),
    .Y(_06342_));
 INVx2_ASAP7_75t_R _22170_ (.A(_00423_),
    .Y(_06353_));
 AND3x1_ASAP7_75t_R _22171_ (.A(_06353_),
    .B(_00421_),
    .C(_00422_),
    .Y(_06364_));
 OR4x2_ASAP7_75t_R _22172_ (.A(_06309_),
    .B(_06331_),
    .C(_06342_),
    .D(_06364_),
    .Y(_06375_));
 INVx1_ASAP7_75t_R _98_113 (.A(clknet_leaf_14_clk),
    .Y(net518));
 INVx6_ASAP7_75t_R _22174_ (.A(_00427_),
    .Y(_06397_));
 NAND2x2_ASAP7_75t_R _22175_ (.A(net2130),
    .B(_06397_),
    .Y(_06408_));
 NOR2x2_ASAP7_75t_R _22176_ (.A(net1658),
    .B(_06408_),
    .Y(_06419_));
 INVx5_ASAP7_75t_R _22177_ (.A(_06419_),
    .Y(_06430_));
 NOR2x2_ASAP7_75t_R _22178_ (.A(net3387),
    .B(_00422_),
    .Y(_06441_));
 INVx4_ASAP7_75t_R _22179_ (.A(_06441_),
    .Y(_06452_));
 NOR2x2_ASAP7_75t_R _22180_ (.A(net3389),
    .B(_06452_),
    .Y(_06463_));
 INVx6_ASAP7_75t_R _22181_ (.A(_06463_),
    .Y(_06474_));
 NOR2x1_ASAP7_75t_R _22182_ (.A(_06430_),
    .B(_06474_),
    .Y(_06485_));
 INVx1_ASAP7_75t_R _98_112 (.A(clknet_leaf_11_clk),
    .Y(net517));
 NOR2x2_ASAP7_75t_R _22184_ (.A(net3390),
    .B(_06474_),
    .Y(_06507_));
 NOR2x2_ASAP7_75t_R _22185_ (.A(net2134),
    .B(net1937),
    .Y(_06518_));
 AND2x2_ASAP7_75t_R _22186_ (.A(_06463_),
    .B(_06518_),
    .Y(_06529_));
 NOR2x2_ASAP7_75t_R _22187_ (.A(_06408_),
    .B(_06057_),
    .Y(_06540_));
 AND2x2_ASAP7_75t_R _22188_ (.A(_06463_),
    .B(_06540_),
    .Y(_06551_));
 INVx1_ASAP7_75t_R _98_111 (.A(clknet_leaf_11_clk),
    .Y(net516));
 NOR2x2_ASAP7_75t_R _22190_ (.A(net2321),
    .B(_06474_),
    .Y(_06573_));
 OR4x1_ASAP7_75t_R _22191_ (.A(_06507_),
    .B(_06529_),
    .C(_06551_),
    .D(_06573_),
    .Y(_06584_));
 NOR2x2_ASAP7_75t_R _22192_ (.A(_05760_),
    .B(_06452_),
    .Y(_06595_));
 INVx6_ASAP7_75t_R _22193_ (.A(_06595_),
    .Y(_06606_));
 NOR2x1_ASAP7_75t_R _22194_ (.A(net1940),
    .B(_06606_),
    .Y(_06617_));
 NOR2x2_ASAP7_75t_R _22195_ (.A(_05936_),
    .B(net2858),
    .Y(_06628_));
 INVx1_ASAP7_75t_R _98_110 (.A(clknet_leaf_4_clk),
    .Y(net515));
 INVx1_ASAP7_75t_R _98_109 (.A(clknet_leaf_4_clk),
    .Y(net514));
 NOR2x2_ASAP7_75t_R _22198_ (.A(_06430_),
    .B(_06606_),
    .Y(_06661_));
 AO21x1_ASAP7_75t_R _22199_ (.A1(_06628_),
    .A2(_06595_),
    .B(_06661_),
    .Y(_06672_));
 INVx1_ASAP7_75t_R _98_108 (.A(clknet_leaf_7_clk),
    .Y(net513));
 NOR2x1_ASAP7_75t_R _22201_ (.A(net2321),
    .B(_06606_),
    .Y(_06694_));
 AO21x1_ASAP7_75t_R _22202_ (.A1(_06595_),
    .A2(_06540_),
    .B(_06694_),
    .Y(_06705_));
 OR5x1_ASAP7_75t_R _22203_ (.A(_06485_),
    .B(_06584_),
    .C(_06617_),
    .D(_06672_),
    .E(_06705_),
    .Y(_06716_));
 CKINVDCx5p33_ASAP7_75t_R _22204_ (.A(net2858),
    .Y(_06727_));
 NAND2x2_ASAP7_75t_R _22205_ (.A(net1616),
    .B(_06727_),
    .Y(_06738_));
 NAND2x2_ASAP7_75t_R _22206_ (.A(_00424_),
    .B(_06353_),
    .Y(_06749_));
 NOR2x2_ASAP7_75t_R _22207_ (.A(_06749_),
    .B(_06452_),
    .Y(_06760_));
 INVx4_ASAP7_75t_R _22208_ (.A(_06760_),
    .Y(_06771_));
 NOR2x1_ASAP7_75t_R _22209_ (.A(_06738_),
    .B(_06771_),
    .Y(_06782_));
 INVx1_ASAP7_75t_R _98_107 (.A(clknet_leaf_5_clk),
    .Y(net512));
 NOR2x2_ASAP7_75t_R _22211_ (.A(_00423_),
    .B(_00424_),
    .Y(_06804_));
 AND2x6_ASAP7_75t_R _22212_ (.A(_06441_),
    .B(_06804_),
    .Y(_06815_));
 CKINVDCx6p67_ASAP7_75t_R _22213_ (.A(_06815_),
    .Y(_06826_));
 INVx1_ASAP7_75t_R _98_106 (.A(clknet_leaf_6_clk),
    .Y(net511));
 NOR2x1_ASAP7_75t_R _22215_ (.A(net3393),
    .B(_06826_),
    .Y(_06848_));
 INVx1_ASAP7_75t_R _98_105 (.A(clknet_leaf_6_clk),
    .Y(net510));
 AND2x2_ASAP7_75t_R _22217_ (.A(_06815_),
    .B(_06255_),
    .Y(_06870_));
 AND2x2_ASAP7_75t_R _22218_ (.A(_06815_),
    .B(_06540_),
    .Y(_06881_));
 NOR2x1_ASAP7_75t_R _22219_ (.A(_06222_),
    .B(_06826_),
    .Y(_06892_));
 OR4x1_ASAP7_75t_R _22220_ (.A(_06848_),
    .B(_06870_),
    .C(_06881_),
    .D(_06892_),
    .Y(_06903_));
 CKINVDCx6p67_ASAP7_75t_R _22221_ (.A(net1658),
    .Y(_06914_));
 NAND2x2_ASAP7_75t_R _22222_ (.A(_06112_),
    .B(_06914_),
    .Y(_06925_));
 INVx2_ASAP7_75t_R _22223_ (.A(_06925_),
    .Y(_06936_));
 NOR2x2_ASAP7_75t_R _22224_ (.A(net1618),
    .B(net2134),
    .Y(_06946_));
 INVx5_ASAP7_75t_R _22225_ (.A(_06946_),
    .Y(_06957_));
 NOR2x2_ASAP7_75t_R _22226_ (.A(net1655),
    .B(_06957_),
    .Y(_06968_));
 INVx1_ASAP7_75t_R _98_104 (.A(clknet_leaf_7_clk),
    .Y(net509));
 INVx1_ASAP7_75t_R _98_103 (.A(clknet_leaf_11_clk),
    .Y(net508));
 OA21x2_ASAP7_75t_R _22229_ (.A1(_06936_),
    .A2(_06968_),
    .B(_06760_),
    .Y(_07001_));
 INVx1_ASAP7_75t_R _98_102 (.A(clknet_leaf_11_clk),
    .Y(net507));
 AND3x1_ASAP7_75t_R _22231_ (.A(_06760_),
    .B(_05936_),
    .C(_06266_),
    .Y(_07023_));
 INVx1_ASAP7_75t_R _22232_ (.A(_07023_),
    .Y(_07034_));
 INVx1_ASAP7_75t_R _98_101 (.A(clknet_leaf_6_clk),
    .Y(net506));
 AND3x1_ASAP7_75t_R _22234_ (.A(_06760_),
    .B(_05925_),
    .C(net2586),
    .Y(_07056_));
 INVx1_ASAP7_75t_R _22235_ (.A(_07056_),
    .Y(_07067_));
 NAND2x1_ASAP7_75t_R _22236_ (.A(_07034_),
    .B(_07067_),
    .Y(_07078_));
 INVx2_ASAP7_75t_R _22237_ (.A(_06112_),
    .Y(_07089_));
 NOR2x2_ASAP7_75t_R _22238_ (.A(net2859),
    .B(_07089_),
    .Y(_07100_));
 CKINVDCx6p67_ASAP7_75t_R _22239_ (.A(_07100_),
    .Y(_07111_));
 INVx1_ASAP7_75t_R _98_100 (.A(clknet_leaf_8_clk),
    .Y(net505));
 NOR2x1_ASAP7_75t_R _22241_ (.A(_06826_),
    .B(_07111_),
    .Y(_07133_));
 NOR2x1_ASAP7_75t_R _22242_ (.A(_06002_),
    .B(_06826_),
    .Y(_07144_));
 INVx1_ASAP7_75t_R _98_99 (.A(clknet_leaf_1_clk),
    .Y(net504));
 NOR2x1_ASAP7_75t_R _22244_ (.A(_05958_),
    .B(_06826_),
    .Y(_07166_));
 OR3x1_ASAP7_75t_R _22245_ (.A(_07133_),
    .B(_07144_),
    .C(_07166_),
    .Y(_07177_));
 OR5x1_ASAP7_75t_R _22246_ (.A(_06782_),
    .B(_06903_),
    .C(_07001_),
    .D(_07078_),
    .E(_07177_),
    .Y(_07188_));
 NOR2x1_ASAP7_75t_R _22247_ (.A(_06716_),
    .B(_07188_),
    .Y(_07199_));
 CKINVDCx9p33_ASAP7_75t_R _22248_ (.A(_06255_),
    .Y(_07210_));
 INVx1_ASAP7_75t_R _98 (.A(clknet_leaf_16_clk),
    .Y(net503));
 INVx1_ASAP7_75t_R _48_97 (.A(clknet_leaf_7_clk),
    .Y(net502));
 AO21x1_ASAP7_75t_R _22251_ (.A1(_07210_),
    .A2(_06222_),
    .B(_05892_),
    .Y(_07243_));
 NOR2x2_ASAP7_75t_R _22252_ (.A(net2858),
    .B(_06957_),
    .Y(_07254_));
 INVx8_ASAP7_75t_R _22253_ (.A(_07254_),
    .Y(_07265_));
 INVx1_ASAP7_75t_R _48_96 (.A(clknet_leaf_14_clk),
    .Y(net501));
 NOR2x2_ASAP7_75t_R _22255_ (.A(_06408_),
    .B(net2858),
    .Y(_07287_));
 CKINVDCx10_ASAP7_75t_R _22256_ (.A(_07287_),
    .Y(_07298_));
 INVx1_ASAP7_75t_R _48_95 (.A(clknet_leaf_14_clk),
    .Y(net500));
 INVx1_ASAP7_75t_R _48_94 (.A(clknet_leaf_13_clk),
    .Y(net499));
 AO21x1_ASAP7_75t_R _22259_ (.A1(_07265_),
    .A2(_07298_),
    .B(_05892_),
    .Y(_07331_));
 CKINVDCx6p67_ASAP7_75t_R _22260_ (.A(_06540_),
    .Y(_07342_));
 INVx1_ASAP7_75t_R _48_93 (.A(clknet_leaf_2_clk),
    .Y(net498));
 AO21x1_ASAP7_75t_R _22262_ (.A1(_07342_),
    .A2(net1047),
    .B(_05892_),
    .Y(_07364_));
 NOR2x1_ASAP7_75t_R _22263_ (.A(_06002_),
    .B(_05892_),
    .Y(_07375_));
 INVx1_ASAP7_75t_R _22264_ (.A(_07375_),
    .Y(_07386_));
 NAND2x1_ASAP7_75t_R _22265_ (.A(_06628_),
    .B(_05881_),
    .Y(_07396_));
 AND5x1_ASAP7_75t_R _22266_ (.A(_07243_),
    .B(_07331_),
    .C(_07364_),
    .D(_07386_),
    .E(_07396_),
    .Y(_07407_));
 NOR2x2_ASAP7_75t_R _22267_ (.A(_06749_),
    .B(_05793_),
    .Y(_07418_));
 AND3x1_ASAP7_75t_R _22268_ (.A(_07418_),
    .B(_06957_),
    .C(_06914_),
    .Y(_07429_));
 INVx1_ASAP7_75t_R _22269_ (.A(_07429_),
    .Y(_07440_));
 AND3x1_ASAP7_75t_R _22270_ (.A(_07418_),
    .B(_06266_),
    .C(_07089_),
    .Y(_07451_));
 INVx1_ASAP7_75t_R _22271_ (.A(_07451_),
    .Y(_07462_));
 INVx1_ASAP7_75t_R _48_92 (.A(clknet_leaf_15_clk),
    .Y(net497));
 INVx8_ASAP7_75t_R _22273_ (.A(_07418_),
    .Y(_07484_));
 INVx1_ASAP7_75t_R _48_91 (.A(clknet_leaf_15_clk),
    .Y(net496));
 AO21x1_ASAP7_75t_R _22275_ (.A1(_06090_),
    .A2(net2055),
    .B(_07484_),
    .Y(_07506_));
 CKINVDCx8_ASAP7_75t_R _22276_ (.A(_06628_),
    .Y(_07517_));
 INVx1_ASAP7_75t_R _48_90 (.A(clknet_leaf_1_clk),
    .Y(net495));
 AO21x1_ASAP7_75t_R _22278_ (.A1(_07517_),
    .A2(_07298_),
    .B(_07484_),
    .Y(_07539_));
 AND4x1_ASAP7_75t_R _22279_ (.A(_07440_),
    .B(_07462_),
    .C(_07506_),
    .D(_07539_),
    .Y(_07550_));
 NOR2x2_ASAP7_75t_R _22280_ (.A(net1936),
    .B(_06957_),
    .Y(_07561_));
 INVx4_ASAP7_75t_R _22281_ (.A(_07561_),
    .Y(_07572_));
 INVx5_ASAP7_75t_R _22282_ (.A(_05804_),
    .Y(_07583_));
 INVx1_ASAP7_75t_R _48_89 (.A(clknet_leaf_1_clk),
    .Y(net494));
 AO21x1_ASAP7_75t_R _22284_ (.A1(_07572_),
    .A2(_06277_),
    .B(_07583_),
    .Y(_07605_));
 AO21x1_ASAP7_75t_R _22285_ (.A1(_07517_),
    .A2(_07298_),
    .B(_07583_),
    .Y(_07616_));
 INVx1_ASAP7_75t_R _48_88 (.A(clknet_leaf_1_clk),
    .Y(net493));
 NAND2x1_ASAP7_75t_R _22287_ (.A(_06419_),
    .B(_05804_),
    .Y(_07638_));
 NAND2x1_ASAP7_75t_R _22288_ (.A(_06968_),
    .B(_05804_),
    .Y(_07649_));
 AND4x1_ASAP7_75t_R _22289_ (.A(_07605_),
    .B(_07616_),
    .C(_07638_),
    .D(_07649_),
    .Y(_07660_));
 NAND2x2_ASAP7_75t_R _22290_ (.A(_05925_),
    .B(_06914_),
    .Y(_07671_));
 NAND2x2_ASAP7_75t_R _22291_ (.A(_06804_),
    .B(_05782_),
    .Y(_07682_));
 INVx1_ASAP7_75t_R _48_87 (.A(clknet_leaf_1_clk),
    .Y(net492));
 AO21x1_ASAP7_75t_R _22293_ (.A1(_06430_),
    .A2(_07671_),
    .B(_07682_),
    .Y(_07704_));
 AO21x1_ASAP7_75t_R _22294_ (.A1(_06145_),
    .A2(_06123_),
    .B(_07682_),
    .Y(_07715_));
 AND2x6_ASAP7_75t_R _22295_ (.A(_06946_),
    .B(_06046_),
    .Y(_07726_));
 CKINVDCx8_ASAP7_75t_R _22296_ (.A(_07726_),
    .Y(_07737_));
 INVx1_ASAP7_75t_R _48_86 (.A(clknet_leaf_2_clk),
    .Y(net491));
 NOR2x1_ASAP7_75t_R _22298_ (.A(_07682_),
    .B(_07737_),
    .Y(_07759_));
 INVx1_ASAP7_75t_R _22299_ (.A(_07759_),
    .Y(_07770_));
 INVx3_ASAP7_75t_R _22300_ (.A(_07682_),
    .Y(_07781_));
 INVx1_ASAP7_75t_R _22301_ (.A(_06277_),
    .Y(_07792_));
 NAND2x1_ASAP7_75t_R _22302_ (.A(_07781_),
    .B(_07792_),
    .Y(_07803_));
 INVx1_ASAP7_75t_R _48_85 (.A(clknet_leaf_2_clk),
    .Y(net490));
 NAND2x1_ASAP7_75t_R _22304_ (.A(net2582),
    .B(_07781_),
    .Y(_07824_));
 AND5x1_ASAP7_75t_R _22305_ (.A(_07704_),
    .B(_07715_),
    .C(_07770_),
    .D(_07803_),
    .E(_07824_),
    .Y(_07835_));
 AND4x1_ASAP7_75t_R _22306_ (.A(_07407_),
    .B(_07550_),
    .C(_07660_),
    .D(_07835_),
    .Y(_07846_));
 NAND2x2_ASAP7_75t_R _22307_ (.A(net3387),
    .B(_06342_),
    .Y(_07857_));
 NOR2x2_ASAP7_75t_R _22308_ (.A(_07857_),
    .B(_05760_),
    .Y(_07868_));
 INVx4_ASAP7_75t_R _22309_ (.A(_07868_),
    .Y(_07879_));
 INVx1_ASAP7_75t_R _48_84 (.A(clknet_leaf_3_clk),
    .Y(net489));
 AO21x1_ASAP7_75t_R _22311_ (.A1(_07265_),
    .A2(_07298_),
    .B(_07879_),
    .Y(_07901_));
 INVx1_ASAP7_75t_R _48_83 (.A(clknet_leaf_6_clk),
    .Y(net488));
 AO21x1_ASAP7_75t_R _22313_ (.A1(net3398),
    .A2(_06925_),
    .B(_07879_),
    .Y(_07923_));
 AND2x2_ASAP7_75t_R _22314_ (.A(_07726_),
    .B(_07868_),
    .Y(_07934_));
 INVx1_ASAP7_75t_R _22315_ (.A(_07934_),
    .Y(_07945_));
 AND2x2_ASAP7_75t_R _22316_ (.A(_06968_),
    .B(_07868_),
    .Y(_07956_));
 INVx1_ASAP7_75t_R _22317_ (.A(_07956_),
    .Y(_07967_));
 NAND2x1_ASAP7_75t_R _22318_ (.A(_06518_),
    .B(_07868_),
    .Y(_07978_));
 AND5x1_ASAP7_75t_R _22319_ (.A(_07901_),
    .B(_07923_),
    .C(_07945_),
    .D(_07967_),
    .E(_07978_),
    .Y(_07989_));
 NOR2x2_ASAP7_75t_R _22320_ (.A(net3388),
    .B(_07857_),
    .Y(_08000_));
 INVx6_ASAP7_75t_R _22321_ (.A(_08000_),
    .Y(_08011_));
 INVx1_ASAP7_75t_R _48_82 (.A(clknet_leaf_6_clk),
    .Y(net487));
 NOR2x1_ASAP7_75t_R _22323_ (.A(_06946_),
    .B(_06057_),
    .Y(_08033_));
 INVx1_ASAP7_75t_R _48_81 (.A(clknet_leaf_8_clk),
    .Y(net486));
 OA21x2_ASAP7_75t_R _22325_ (.A1(_08033_),
    .A2(_06518_),
    .B(_08000_),
    .Y(_08055_));
 INVx1_ASAP7_75t_R _22326_ (.A(_08055_),
    .Y(_08066_));
 AO21x1_ASAP7_75t_R _22327_ (.A1(net3392),
    .A2(_06925_),
    .B(_08011_),
    .Y(_08077_));
 OA211x2_ASAP7_75t_R _22328_ (.A1(_07111_),
    .A2(_08011_),
    .B(_08066_),
    .C(_08077_),
    .Y(_08088_));
 NOR2x2_ASAP7_75t_R _22329_ (.A(_00423_),
    .B(_05749_),
    .Y(_08099_));
 INVx1_ASAP7_75t_R _22330_ (.A(_07857_),
    .Y(_08110_));
 NAND2x2_ASAP7_75t_R _22331_ (.A(_08099_),
    .B(_08110_),
    .Y(_08121_));
 INVx1_ASAP7_75t_R _48_80 (.A(clknet_leaf_11_clk),
    .Y(net485));
 AO21x1_ASAP7_75t_R _22333_ (.A1(_07572_),
    .A2(net3393),
    .B(_08121_),
    .Y(_08143_));
 NOR2x1_ASAP7_75t_R _22334_ (.A(_08121_),
    .B(_07210_),
    .Y(_08154_));
 INVx1_ASAP7_75t_R _22335_ (.A(_08154_),
    .Y(_08165_));
 NOR2x1_ASAP7_75t_R _22336_ (.A(_08121_),
    .B(_07342_),
    .Y(_08176_));
 INVx1_ASAP7_75t_R _22337_ (.A(_08176_),
    .Y(_08186_));
 AO21x1_ASAP7_75t_R _22338_ (.A1(_07671_),
    .A2(net2858),
    .B(_08121_),
    .Y(_08197_));
 AND4x1_ASAP7_75t_R _22339_ (.A(_08143_),
    .B(_08165_),
    .C(_08186_),
    .D(_08197_),
    .Y(_08208_));
 INVx1_ASAP7_75t_R _22340_ (.A(_06804_),
    .Y(_08219_));
 NOR2x2_ASAP7_75t_R _22341_ (.A(_07857_),
    .B(_08219_),
    .Y(_08230_));
 AND2x2_ASAP7_75t_R _22342_ (.A(_07561_),
    .B(_08230_),
    .Y(_08241_));
 INVx3_ASAP7_75t_R _22343_ (.A(net2322),
    .Y(_08252_));
 OA21x2_ASAP7_75t_R _22344_ (.A1(_08252_),
    .A2(_06540_),
    .B(_08230_),
    .Y(_08263_));
 NOR2x1_ASAP7_75t_R _22345_ (.A(_08241_),
    .B(_08263_),
    .Y(_08274_));
 INVx4_ASAP7_75t_R _22346_ (.A(_08230_),
    .Y(_08285_));
 AO21x1_ASAP7_75t_R _22347_ (.A1(_07265_),
    .A2(_07517_),
    .B(_08285_),
    .Y(_08296_));
 INVx4_ASAP7_75t_R _22348_ (.A(_06408_),
    .Y(_08307_));
 OR3x1_ASAP7_75t_R _22349_ (.A(_08285_),
    .B(_08307_),
    .C(net1656),
    .Y(_08318_));
 AND3x1_ASAP7_75t_R _22350_ (.A(_08274_),
    .B(_08296_),
    .C(_08318_),
    .Y(_08329_));
 AND4x1_ASAP7_75t_R _22351_ (.A(_07989_),
    .B(_08088_),
    .C(_08208_),
    .D(_08329_),
    .Y(_08340_));
 INVx1_ASAP7_75t_R _48_79 (.A(clknet_leaf_11_clk),
    .Y(net484));
 AND4x2_ASAP7_75t_R _22353_ (.A(_06331_),
    .B(_00422_),
    .C(_00423_),
    .D(_00424_),
    .Y(_08362_));
 INVx1_ASAP7_75t_R _48_78 (.A(clknet_leaf_4_clk),
    .Y(net483));
 INVx1_ASAP7_75t_R _48_77 (.A(clknet_leaf_4_clk),
    .Y(net482));
 OA211x2_ASAP7_75t_R _22356_ (.A1(net1146),
    .A2(_05925_),
    .B(_08362_),
    .C(_06727_),
    .Y(_08395_));
 OR3x4_ASAP7_75t_R _22357_ (.A(_05760_),
    .B(_00421_),
    .C(_06342_),
    .Y(_08406_));
 INVx2_ASAP7_75t_R _22358_ (.A(_08406_),
    .Y(_08417_));
 OA31x2_ASAP7_75t_R _22359_ (.A1(_06419_),
    .A2(_05947_),
    .A3(_06079_),
    .B1(_08417_),
    .Y(_08428_));
 AND3x1_ASAP7_75t_R _22360_ (.A(_08362_),
    .B(_07089_),
    .C(net2586),
    .Y(_08439_));
 OA21x2_ASAP7_75t_R _22361_ (.A1(_06936_),
    .A2(_06419_),
    .B(_08362_),
    .Y(_08450_));
 OR3x4_ASAP7_75t_R _22362_ (.A(_05870_),
    .B(_00421_),
    .C(_06342_),
    .Y(_08461_));
 INVx1_ASAP7_75t_R _48_76 (.A(clknet_leaf_7_clk),
    .Y(net481));
 NOR2x1_ASAP7_75t_R _22364_ (.A(_07210_),
    .B(_08461_),
    .Y(_08483_));
 AO21x1_ASAP7_75t_R _22365_ (.A1(_07561_),
    .A2(_08362_),
    .B(_08483_),
    .Y(_08494_));
 OR5x1_ASAP7_75t_R _22366_ (.A(_08395_),
    .B(_08428_),
    .C(_08439_),
    .D(_08450_),
    .E(_08494_),
    .Y(_08505_));
 AND3x4_ASAP7_75t_R _22367_ (.A(_08099_),
    .B(_06331_),
    .C(_00422_),
    .Y(_08516_));
 INVx1_ASAP7_75t_R _48_75 (.A(clknet_leaf_5_clk),
    .Y(net480));
 NAND2x1_ASAP7_75t_R _22369_ (.A(_07210_),
    .B(_07737_),
    .Y(_08537_));
 AND3x1_ASAP7_75t_R _22370_ (.A(_08516_),
    .B(net1146),
    .C(_06046_),
    .Y(_08548_));
 AO21x1_ASAP7_75t_R _22371_ (.A1(_08516_),
    .A2(_08537_),
    .B(_08548_),
    .Y(_08559_));
 AND3x4_ASAP7_75t_R _22372_ (.A(_06804_),
    .B(_06331_),
    .C(_00422_),
    .Y(_08570_));
 INVx1_ASAP7_75t_R _48_74 (.A(clknet_leaf_6_clk),
    .Y(net479));
 AND3x1_ASAP7_75t_R _22374_ (.A(_08570_),
    .B(_05936_),
    .C(_06914_),
    .Y(_08592_));
 NOR2x2_ASAP7_75t_R _22375_ (.A(net2858),
    .B(_08307_),
    .Y(_08603_));
 INVx1_ASAP7_75t_R _22376_ (.A(_08603_),
    .Y(_08614_));
 CKINVDCx5p33_ASAP7_75t_R _22377_ (.A(_08570_),
    .Y(_08625_));
 INVx1_ASAP7_75t_R _48_73 (.A(clknet_leaf_6_clk),
    .Y(net478));
 NOR2x1_ASAP7_75t_R _22379_ (.A(_08614_),
    .B(_08625_),
    .Y(_08647_));
 NOR2x1_ASAP7_75t_R _22380_ (.A(net2055),
    .B(_08625_),
    .Y(_08658_));
 OR3x4_ASAP7_75t_R _22381_ (.A(_06749_),
    .B(_00421_),
    .C(_06342_),
    .Y(_08669_));
 INVx1_ASAP7_75t_R _48_72 (.A(clknet_leaf_7_clk),
    .Y(net477));
 NOR2x1_ASAP7_75t_R _22383_ (.A(_07111_),
    .B(_08669_),
    .Y(_08691_));
 OR5x1_ASAP7_75t_R _22384_ (.A(_08559_),
    .B(_08592_),
    .C(_08647_),
    .D(_08658_),
    .E(_08691_),
    .Y(_08702_));
 NOR2x1_ASAP7_75t_R _22385_ (.A(_08505_),
    .B(_08702_),
    .Y(_08713_));
 AND4x2_ASAP7_75t_R _22386_ (.A(_07199_),
    .B(_07846_),
    .C(_08340_),
    .D(_08713_),
    .Y(_08724_));
 INVx1_ASAP7_75t_R _48_71 (.A(clknet_leaf_11_clk),
    .Y(net476));
 XOR2x1_ASAP7_75t_R _22388_ (.A(_00409_),
    .Y(_08746_),
    .B(net3512));
 INVx3_ASAP7_75t_R _22389_ (.A(_00484_),
    .Y(_08757_));
 XOR2x1_ASAP7_75t_R _22390_ (.A(_08746_),
    .Y(_08768_),
    .B(_08757_));
 INVx6_ASAP7_75t_R _22391_ (.A(_00500_),
    .Y(_08779_));
 XOR2x1_ASAP7_75t_R _22392_ (.A(_08768_),
    .Y(_08790_),
    .B(_08779_));
 AOI21x1_ASAP7_75t_R _22393_ (.A1(net2609),
    .A2(_08724_),
    .B(_08790_),
    .Y(_08801_));
 AND3x1_ASAP7_75t_R _22394_ (.A(_08724_),
    .B(_06375_),
    .C(_08790_),
    .Y(_08812_));
 INVx13_ASAP7_75t_R _22395_ (.A(net401),
    .Y(_08823_));
 INVx1_ASAP7_75t_R _48_70 (.A(clknet_leaf_11_clk),
    .Y(net475));
 OAI21x1_ASAP7_75t_R _22397_ (.A1(_08801_),
    .A2(_08812_),
    .B(net400),
    .Y(_08845_));
 NAND2x1_ASAP7_75t_R _22398_ (.A(_05716_),
    .B(_08845_),
    .Y(_00353_));
 INVx1_ASAP7_75t_R _48_69 (.A(clknet_leaf_6_clk),
    .Y(net474));
 INVx1_ASAP7_75t_R _48_68 (.A(clknet_leaf_6_clk),
    .Y(net473));
 INVx1_ASAP7_75t_R _22401_ (.A(net4017),
    .Y(_08887_));
 AO21x1_ASAP7_75t_R _22402_ (.A1(_06430_),
    .A2(_06925_),
    .B(_08625_),
    .Y(_08898_));
 AO21x1_ASAP7_75t_R _22403_ (.A1(_07210_),
    .A2(_07572_),
    .B(_08625_),
    .Y(_08909_));
 NAND2x1_ASAP7_75t_R _22404_ (.A(_06540_),
    .B(_08570_),
    .Y(_08920_));
 NAND2x1_ASAP7_75t_R _22405_ (.A(_07287_),
    .B(_08570_),
    .Y(_08931_));
 NAND2x1_ASAP7_75t_R _22406_ (.A(_08252_),
    .B(_08570_),
    .Y(_08942_));
 AND5x1_ASAP7_75t_R _22407_ (.A(_08898_),
    .B(_08909_),
    .C(_08920_),
    .D(_08931_),
    .E(_08942_),
    .Y(_08953_));
 OA211x2_ASAP7_75t_R _22408_ (.A1(net1146),
    .A2(_05925_),
    .B(_08516_),
    .C(_06266_),
    .Y(_08964_));
 INVx1_ASAP7_75t_R _22409_ (.A(_08964_),
    .Y(_08975_));
 NAND2x2_ASAP7_75t_R _22410_ (.A(_05947_),
    .B(_08516_),
    .Y(_08986_));
 OA21x2_ASAP7_75t_R _22411_ (.A1(_06419_),
    .A2(_06968_),
    .B(_08516_),
    .Y(_08997_));
 INVx1_ASAP7_75t_R _22412_ (.A(_08997_),
    .Y(_09008_));
 NAND2x1_ASAP7_75t_R _22413_ (.A(_06628_),
    .B(_08516_),
    .Y(_09019_));
 AND4x1_ASAP7_75t_R _22414_ (.A(_08975_),
    .B(_08986_),
    .C(_09008_),
    .D(_09019_),
    .Y(_09030_));
 NAND2x1_ASAP7_75t_R _22415_ (.A(_08953_),
    .B(_09030_),
    .Y(_09041_));
 NOR2x2_ASAP7_75t_R _22416_ (.A(_06408_),
    .B(net1939),
    .Y(_09052_));
 INVx1_ASAP7_75t_R _48_67 (.A(clknet_leaf_1_clk),
    .Y(net472));
 AO21x1_ASAP7_75t_R _22418_ (.A1(_09052_),
    .A2(_08362_),
    .B(_08483_),
    .Y(_09074_));
 OA21x2_ASAP7_75t_R _22419_ (.A1(_06419_),
    .A2(_08603_),
    .B(_08362_),
    .Y(_09085_));
 NOR2x1_ASAP7_75t_R _22420_ (.A(_07737_),
    .B(_08461_),
    .Y(_09096_));
 OR3x1_ASAP7_75t_R _22421_ (.A(_09074_),
    .B(_09085_),
    .C(_09096_),
    .Y(_09107_));
 INVx1_ASAP7_75t_R _48_66 (.A(clknet_leaf_15_clk),
    .Y(net471));
 AO21x1_ASAP7_75t_R _22423_ (.A1(_07210_),
    .A2(net3403),
    .B(_08406_),
    .Y(_09128_));
 AO21x1_ASAP7_75t_R _22424_ (.A1(_06738_),
    .A2(_06430_),
    .B(_08406_),
    .Y(_09138_));
 NOR2x1_ASAP7_75t_R _22425_ (.A(_06057_),
    .B(_08406_),
    .Y(_09149_));
 INVx1_ASAP7_75t_R _22426_ (.A(_09149_),
    .Y(_09159_));
 NAND3x1_ASAP7_75t_R _22427_ (.A(_09128_),
    .B(_09138_),
    .C(_09159_),
    .Y(_09170_));
 OR3x2_ASAP7_75t_R _22428_ (.A(_09041_),
    .B(_09107_),
    .C(_09170_),
    .Y(_09179_));
 AND2x2_ASAP7_75t_R _22429_ (.A(_06760_),
    .B(net2349),
    .Y(_09190_));
 OA21x2_ASAP7_75t_R _22430_ (.A1(_07726_),
    .A2(_06540_),
    .B(_06815_),
    .Y(_09201_));
 AO21x1_ASAP7_75t_R _22431_ (.A1(_07561_),
    .A2(_06815_),
    .B(_09201_),
    .Y(_09211_));
 NAND2x2_ASAP7_75t_R _22432_ (.A(net1620),
    .B(_06266_),
    .Y(_09221_));
 NOR2x2_ASAP7_75t_R _22433_ (.A(_09221_),
    .B(_06771_),
    .Y(_09232_));
 AO21x1_ASAP7_75t_R _22434_ (.A1(_09052_),
    .A2(_06760_),
    .B(_09232_),
    .Y(_09243_));
 AO21x1_ASAP7_75t_R _22435_ (.A1(_07737_),
    .A2(net3390),
    .B(_06771_),
    .Y(_09253_));
 INVx1_ASAP7_75t_R _22436_ (.A(_09253_),
    .Y(_09263_));
 NOR2x2_ASAP7_75t_R _22437_ (.A(_06738_),
    .B(_06826_),
    .Y(_09274_));
 AO21x1_ASAP7_75t_R _22438_ (.A1(_06815_),
    .A2(net2349),
    .B(_09274_),
    .Y(_09285_));
 OR5x1_ASAP7_75t_R _22439_ (.A(_09190_),
    .B(_09211_),
    .C(_09243_),
    .D(_09263_),
    .E(_09285_),
    .Y(_09295_));
 AND2x2_ASAP7_75t_R _22440_ (.A(_07254_),
    .B(_06463_),
    .Y(_09306_));
 AO21x1_ASAP7_75t_R _22441_ (.A1(_06628_),
    .A2(_06463_),
    .B(_09306_),
    .Y(_09317_));
 INVx1_ASAP7_75t_R _48_65 (.A(clknet_leaf_8_clk),
    .Y(net470));
 AND2x2_ASAP7_75t_R _22443_ (.A(_07561_),
    .B(_06463_),
    .Y(_09337_));
 AO21x1_ASAP7_75t_R _22444_ (.A1(_07737_),
    .A2(_07342_),
    .B(_06474_),
    .Y(_09348_));
 INVx1_ASAP7_75t_R _22445_ (.A(_09348_),
    .Y(_09359_));
 AND2x2_ASAP7_75t_R _22446_ (.A(_06408_),
    .B(_05936_),
    .Y(_09369_));
 AND3x1_ASAP7_75t_R _22447_ (.A(_09369_),
    .B(_06463_),
    .C(_06914_),
    .Y(_09380_));
 OR5x1_ASAP7_75t_R _22448_ (.A(_06507_),
    .B(_09317_),
    .C(_09337_),
    .D(_09359_),
    .E(_09380_),
    .Y(_09391_));
 NOR2x2_ASAP7_75t_R _22449_ (.A(net1653),
    .B(_06606_),
    .Y(_09401_));
 AND2x2_ASAP7_75t_R _22450_ (.A(_06595_),
    .B(_07287_),
    .Y(_09412_));
 INVx1_ASAP7_75t_R _22451_ (.A(_09412_),
    .Y(_09422_));
 AND2x2_ASAP7_75t_R _22452_ (.A(_07254_),
    .B(_06595_),
    .Y(_09433_));
 INVx1_ASAP7_75t_R _22453_ (.A(_09433_),
    .Y(_09443_));
 NAND2x1_ASAP7_75t_R _22454_ (.A(_09422_),
    .B(_09443_),
    .Y(_09454_));
 AO221x1_ASAP7_75t_R _22455_ (.A1(_05925_),
    .A2(_09401_),
    .B1(_06628_),
    .B2(_06595_),
    .C(_09454_),
    .Y(_09464_));
 AND2x2_ASAP7_75t_R _22456_ (.A(_07726_),
    .B(_06595_),
    .Y(_09474_));
 AND2x2_ASAP7_75t_R _22457_ (.A(_06595_),
    .B(_09052_),
    .Y(_09485_));
 NOR2x1_ASAP7_75t_R _22458_ (.A(net2055),
    .B(_06606_),
    .Y(_09495_));
 OR3x1_ASAP7_75t_R _22459_ (.A(_09474_),
    .B(_09485_),
    .C(_09495_),
    .Y(_09505_));
 OR4x2_ASAP7_75t_R _22460_ (.A(_09295_),
    .B(_09391_),
    .C(_09464_),
    .D(_09505_),
    .Y(_09516_));
 NOR2x2_ASAP7_75t_R _22461_ (.A(_09179_),
    .B(_09516_),
    .Y(_09526_));
 AO21x1_ASAP7_75t_R _22462_ (.A1(_07210_),
    .A2(_06277_),
    .B(_07682_),
    .Y(_09537_));
 NOR2x1_ASAP7_75t_R _22463_ (.A(_07682_),
    .B(_07342_),
    .Y(_09547_));
 INVx1_ASAP7_75t_R _22464_ (.A(_09547_),
    .Y(_09557_));
 NOR2x1_ASAP7_75t_R _22465_ (.A(_07682_),
    .B(_07572_),
    .Y(_09567_));
 INVx1_ASAP7_75t_R _22466_ (.A(_09567_),
    .Y(_09577_));
 AND4x1_ASAP7_75t_R _22467_ (.A(_09537_),
    .B(_07715_),
    .C(_09557_),
    .D(_09577_),
    .Y(_09588_));
 OR3x1_ASAP7_75t_R _22468_ (.A(_07484_),
    .B(_06946_),
    .C(net2858),
    .Y(_09599_));
 OR3x1_ASAP7_75t_R _22469_ (.A(_07484_),
    .B(_06134_),
    .C(net1655),
    .Y(_09610_));
 AO21x1_ASAP7_75t_R _22470_ (.A1(_07265_),
    .A2(_07517_),
    .B(_07682_),
    .Y(_09621_));
 AND5x1_ASAP7_75t_R _22471_ (.A(_07704_),
    .B(_09588_),
    .C(_09599_),
    .D(_09610_),
    .E(_09621_),
    .Y(_09632_));
 INVx1_ASAP7_75t_R _22472_ (.A(_06244_),
    .Y(_09643_));
 AO21x1_ASAP7_75t_R _22473_ (.A1(_07111_),
    .A2(_07298_),
    .B(_07583_),
    .Y(_09654_));
 AO21x1_ASAP7_75t_R _22474_ (.A1(_06925_),
    .A2(_05958_),
    .B(_07583_),
    .Y(_09665_));
 NAND2x1_ASAP7_75t_R _22475_ (.A(_06211_),
    .B(_05804_),
    .Y(_09676_));
 NAND2x1_ASAP7_75t_R _22476_ (.A(_06540_),
    .B(_05804_),
    .Y(_09687_));
 AND4x1_ASAP7_75t_R _22477_ (.A(_09654_),
    .B(_09665_),
    .C(_09676_),
    .D(_09687_),
    .Y(_09698_));
 OA211x2_ASAP7_75t_R _22478_ (.A1(net1617),
    .A2(net2131),
    .B(_05881_),
    .C(_06727_),
    .Y(_09709_));
 INVx1_ASAP7_75t_R _22479_ (.A(_09709_),
    .Y(_09720_));
 AND5x1_ASAP7_75t_R _22480_ (.A(_09643_),
    .B(_09698_),
    .C(_07386_),
    .D(_06167_),
    .E(_09720_),
    .Y(_09731_));
 NAND2x1_ASAP7_75t_R _22481_ (.A(_09632_),
    .B(_09731_),
    .Y(_09742_));
 AND2x2_ASAP7_75t_R _22482_ (.A(_05947_),
    .B(_08000_),
    .Y(_09753_));
 NAND2x1_ASAP7_75t_R _22483_ (.A(_08000_),
    .B(_06540_),
    .Y(_09764_));
 NOR2x1_ASAP7_75t_R _22484_ (.A(_06145_),
    .B(_08011_),
    .Y(_09775_));
 INVx1_ASAP7_75t_R _22485_ (.A(_09775_),
    .Y(_09786_));
 NAND2x1_ASAP7_75t_R _22486_ (.A(_09764_),
    .B(_09786_),
    .Y(_09797_));
 NOR2x1_ASAP7_75t_R _22487_ (.A(net1938),
    .B(_08011_),
    .Y(_09808_));
 AND3x1_ASAP7_75t_R _22488_ (.A(_08000_),
    .B(_06957_),
    .C(_06727_),
    .Y(_09819_));
 NAND2x1_ASAP7_75t_R _22489_ (.A(_08000_),
    .B(_06968_),
    .Y(_09830_));
 INVx1_ASAP7_75t_R _22490_ (.A(_09830_),
    .Y(_09841_));
 OR5x1_ASAP7_75t_R _22491_ (.A(_09753_),
    .B(_09797_),
    .C(_09808_),
    .D(_09819_),
    .E(_09841_),
    .Y(_09852_));
 INVx4_ASAP7_75t_R _22492_ (.A(_08121_),
    .Y(_09863_));
 AO21x1_ASAP7_75t_R _22493_ (.A1(_09863_),
    .A2(_06211_),
    .B(_08176_),
    .Y(_09874_));
 NOR2x1_ASAP7_75t_R _22494_ (.A(_08121_),
    .B(_07298_),
    .Y(_09885_));
 AO21x1_ASAP7_75t_R _22495_ (.A1(_09863_),
    .A2(_07100_),
    .B(_09885_),
    .Y(_09896_));
 NOR2x1_ASAP7_75t_R _22496_ (.A(net1657),
    .B(_08121_),
    .Y(_09907_));
 INVx1_ASAP7_75t_R _22497_ (.A(_09907_),
    .Y(_09918_));
 NOR2x1_ASAP7_75t_R _22498_ (.A(_06112_),
    .B(_09918_),
    .Y(_09929_));
 OR3x1_ASAP7_75t_R _22499_ (.A(_09874_),
    .B(_09896_),
    .C(_09929_),
    .Y(_09940_));
 INVx1_ASAP7_75t_R _22500_ (.A(_06123_),
    .Y(_09951_));
 AO21x1_ASAP7_75t_R _22501_ (.A1(_09951_),
    .A2(_07868_),
    .B(_07934_),
    .Y(_09962_));
 AND2x2_ASAP7_75t_R _22502_ (.A(_09052_),
    .B(_07868_),
    .Y(_09973_));
 OA21x2_ASAP7_75t_R _22503_ (.A1(_07792_),
    .A2(_06255_),
    .B(_07868_),
    .Y(_09984_));
 OA21x2_ASAP7_75t_R _22504_ (.A1(_06936_),
    .A2(_07254_),
    .B(_07868_),
    .Y(_09995_));
 OR4x1_ASAP7_75t_R _22505_ (.A(_09962_),
    .B(_09973_),
    .C(_09984_),
    .D(_09995_),
    .Y(_10006_));
 INVx1_ASAP7_75t_R _48_64 (.A(clknet_leaf_14_clk),
    .Y(net469));
 NOR2x1_ASAP7_75t_R _22507_ (.A(net3398),
    .B(_08285_),
    .Y(_10028_));
 AO21x1_ASAP7_75t_R _22508_ (.A1(_06968_),
    .A2(_08230_),
    .B(_10028_),
    .Y(_10039_));
 AO21x1_ASAP7_75t_R _22509_ (.A1(_07100_),
    .A2(_08230_),
    .B(_10039_),
    .Y(_10050_));
 NOR2x1_ASAP7_75t_R _22510_ (.A(_06057_),
    .B(_08285_),
    .Y(_10061_));
 AND2x2_ASAP7_75t_R _22511_ (.A(_08230_),
    .B(_09052_),
    .Y(_10072_));
 AO221x1_ASAP7_75t_R _22512_ (.A1(_06255_),
    .A2(_08230_),
    .B1(_07089_),
    .B2(_10061_),
    .C(_10072_),
    .Y(_10083_));
 OR5x1_ASAP7_75t_R _22513_ (.A(_09852_),
    .B(_09940_),
    .C(_10006_),
    .D(_10050_),
    .E(_10083_),
    .Y(_10094_));
 NOR2x1_ASAP7_75t_R _22514_ (.A(_09742_),
    .B(_10094_),
    .Y(_10105_));
 NAND2x2_ASAP7_75t_R _22515_ (.A(_09526_),
    .B(_10105_),
    .Y(_10116_));
 INVx4_ASAP7_75t_R _22516_ (.A(_06375_),
    .Y(_10127_));
 INVx1_ASAP7_75t_R _48_63 (.A(clknet_leaf_13_clk),
    .Y(net468));
 INVx1_ASAP7_75t_R _48_62 (.A(clknet_leaf_13_clk),
    .Y(net467));
 XOR2x1_ASAP7_75t_R _22519_ (.A(_00410_),
    .Y(_10160_),
    .B(net2196));
 INVx4_ASAP7_75t_R _22520_ (.A(_00483_),
    .Y(_10171_));
 XOR2x1_ASAP7_75t_R _22521_ (.A(_10160_),
    .Y(_10182_),
    .B(_10171_));
 XOR2x1_ASAP7_75t_R _22522_ (.A(_10182_),
    .Y(_10193_),
    .B(_00499_));
 NOR3x1_ASAP7_75t_R _22523_ (.A(_10116_),
    .B(_10127_),
    .C(_10193_),
    .Y(_10204_));
 OA21x2_ASAP7_75t_R _22524_ (.A1(_10116_),
    .A2(_10127_),
    .B(_10193_),
    .Y(_10215_));
 INVx1_ASAP7_75t_R _48_61 (.A(clknet_leaf_1_clk),
    .Y(net466));
 INVx1_ASAP7_75t_R _48_60 (.A(clknet_leaf_1_clk),
    .Y(net465));
 OAI21x1_ASAP7_75t_R _22527_ (.A1(_10204_),
    .A2(_10215_),
    .B(net400),
    .Y(_10248_));
 OAI21x1_ASAP7_75t_R _22528_ (.A1(net400),
    .A2(_08887_),
    .B(_10248_),
    .Y(_00364_));
 INVx1_ASAP7_75t_R _22529_ (.A(_08592_),
    .Y(_10269_));
 OR3x1_ASAP7_75t_R _22530_ (.A(_08461_),
    .B(_06419_),
    .C(_06079_),
    .Y(_10280_));
 NAND2x1_ASAP7_75t_R _22531_ (.A(_05991_),
    .B(_08417_),
    .Y(_10291_));
 AO21x1_ASAP7_75t_R _22532_ (.A1(net3391),
    .A2(net1047),
    .B(_08406_),
    .Y(_10302_));
 AO21x1_ASAP7_75t_R _22533_ (.A1(_07572_),
    .A2(_09221_),
    .B(_08406_),
    .Y(_10313_));
 AND4x1_ASAP7_75t_R _22534_ (.A(_10280_),
    .B(_10291_),
    .C(_10302_),
    .D(_10313_),
    .Y(_10324_));
 AO21x1_ASAP7_75t_R _22535_ (.A1(_07265_),
    .A2(_07298_),
    .B(_08669_),
    .Y(_10335_));
 AO21x1_ASAP7_75t_R _22536_ (.A1(_07342_),
    .A2(net2321),
    .B(_08669_),
    .Y(_10346_));
 NAND2x1_ASAP7_75t_R _22537_ (.A(_09052_),
    .B(_08516_),
    .Y(_10357_));
 AND4x1_ASAP7_75t_R _22538_ (.A(_10335_),
    .B(_10346_),
    .C(_09019_),
    .D(_10357_),
    .Y(_10368_));
 AO21x1_ASAP7_75t_R _22539_ (.A1(net2055),
    .A2(_07342_),
    .B(_08625_),
    .Y(_10379_));
 NAND2x1_ASAP7_75t_R _22540_ (.A(_09052_),
    .B(_08570_),
    .Y(_10390_));
 OA211x2_ASAP7_75t_R _22541_ (.A1(_09221_),
    .A2(_08625_),
    .B(_10379_),
    .C(_10390_),
    .Y(_10401_));
 AO21x1_ASAP7_75t_R _22542_ (.A1(_07298_),
    .A2(_06738_),
    .B(_08625_),
    .Y(_10412_));
 AND5x1_ASAP7_75t_R _22543_ (.A(_10269_),
    .B(_10324_),
    .C(_10368_),
    .D(_10401_),
    .E(_10412_),
    .Y(_10423_));
 INVx1_ASAP7_75t_R _22544_ (.A(_06892_),
    .Y(_10434_));
 AND3x1_ASAP7_75t_R _22545_ (.A(_06760_),
    .B(_06408_),
    .C(_06046_),
    .Y(_10445_));
 INVx1_ASAP7_75t_R _22546_ (.A(_10445_),
    .Y(_10456_));
 AO21x1_ASAP7_75t_R _22547_ (.A1(_07265_),
    .A2(_07298_),
    .B(_06771_),
    .Y(_10467_));
 CKINVDCx5p33_ASAP7_75t_R _22548_ (.A(_09052_),
    .Y(_10478_));
 AO21x1_ASAP7_75t_R _22549_ (.A1(_07210_),
    .A2(_10478_),
    .B(_06771_),
    .Y(_10489_));
 AND3x1_ASAP7_75t_R _22550_ (.A(_10456_),
    .B(_10467_),
    .C(_10489_),
    .Y(_10500_));
 INVx1_ASAP7_75t_R _22551_ (.A(_09274_),
    .Y(_10511_));
 AO21x1_ASAP7_75t_R _22552_ (.A1(_07737_),
    .A2(net1047),
    .B(_06826_),
    .Y(_10522_));
 INVx4_ASAP7_75t_R _22553_ (.A(_06968_),
    .Y(_10533_));
 AO21x1_ASAP7_75t_R _22554_ (.A1(_10533_),
    .A2(_06925_),
    .B(_06826_),
    .Y(_10544_));
 AND5x1_ASAP7_75t_R _22555_ (.A(_10434_),
    .B(_10500_),
    .C(_10511_),
    .D(_10522_),
    .E(_10544_),
    .Y(_10555_));
 AO21x1_ASAP7_75t_R _22556_ (.A1(_06463_),
    .A2(net2582),
    .B(_09317_),
    .Y(_10566_));
 NOR2x1_ASAP7_75t_R _22557_ (.A(_06474_),
    .B(_07111_),
    .Y(_10577_));
 NOR2x1_ASAP7_75t_R _22558_ (.A(net3400),
    .B(_05936_),
    .Y(_10588_));
 OA21x2_ASAP7_75t_R _22559_ (.A1(_06211_),
    .A2(_10588_),
    .B(_06463_),
    .Y(_10599_));
 AO21x1_ASAP7_75t_R _22560_ (.A1(_06968_),
    .A2(_06463_),
    .B(_06485_),
    .Y(_10610_));
 OR4x1_ASAP7_75t_R _22561_ (.A(_10566_),
    .B(_10577_),
    .C(_10599_),
    .D(_10610_),
    .Y(_10621_));
 AO21x1_ASAP7_75t_R _22562_ (.A1(_06968_),
    .A2(_06595_),
    .B(_06661_),
    .Y(_10632_));
 NOR2x1_ASAP7_75t_R _22563_ (.A(net3392),
    .B(_06606_),
    .Y(_10643_));
 OR3x1_ASAP7_75t_R _22564_ (.A(_10632_),
    .B(_09454_),
    .C(_10643_),
    .Y(_10654_));
 AND2x2_ASAP7_75t_R _22565_ (.A(_06595_),
    .B(_06079_),
    .Y(_10665_));
 AND2x2_ASAP7_75t_R _22566_ (.A(_06595_),
    .B(_06255_),
    .Y(_10676_));
 OR4x1_ASAP7_75t_R _22567_ (.A(_10665_),
    .B(_10676_),
    .C(_09485_),
    .D(_09495_),
    .Y(_10687_));
 NOR3x1_ASAP7_75t_R _22568_ (.A(_10621_),
    .B(_10654_),
    .C(_10687_),
    .Y(_10698_));
 AND3x2_ASAP7_75t_R _22569_ (.A(_10423_),
    .B(_10555_),
    .C(_10698_),
    .Y(_10709_));
 NOR2x1_ASAP7_75t_R _22570_ (.A(_08011_),
    .B(_07737_),
    .Y(_10720_));
 INVx1_ASAP7_75t_R _22571_ (.A(_10720_),
    .Y(_10731_));
 NOR2x1_ASAP7_75t_R _22572_ (.A(_08011_),
    .B(_10478_),
    .Y(_10742_));
 INVx1_ASAP7_75t_R _22573_ (.A(_10742_),
    .Y(_10753_));
 NOR2x1_ASAP7_75t_R _22574_ (.A(_08011_),
    .B(_07517_),
    .Y(_10764_));
 INVx1_ASAP7_75t_R _22575_ (.A(_10764_),
    .Y(_10775_));
 AND2x2_ASAP7_75t_R _22576_ (.A(_06419_),
    .B(_08000_),
    .Y(_10786_));
 INVx1_ASAP7_75t_R _22577_ (.A(_10786_),
    .Y(_10797_));
 AND5x1_ASAP7_75t_R _22578_ (.A(_09764_),
    .B(_10731_),
    .C(_10753_),
    .D(_10775_),
    .E(_10797_),
    .Y(_10808_));
 NAND2x1_ASAP7_75t_R _22579_ (.A(_06628_),
    .B(_07868_),
    .Y(_10819_));
 INVx1_ASAP7_75t_R _22580_ (.A(_09973_),
    .Y(_10830_));
 AO21x1_ASAP7_75t_R _22581_ (.A1(_07737_),
    .A2(net1047),
    .B(_07879_),
    .Y(_10841_));
 AND5x1_ASAP7_75t_R _22582_ (.A(_07967_),
    .B(_10808_),
    .C(_10819_),
    .D(_10830_),
    .E(_10841_),
    .Y(_10852_));
 AO21x1_ASAP7_75t_R _22583_ (.A1(_07298_),
    .A2(_10533_),
    .B(_07583_),
    .Y(_10863_));
 NAND2x1_ASAP7_75t_R _22584_ (.A(_06727_),
    .B(_07418_),
    .Y(_10874_));
 OR3x1_ASAP7_75t_R _22585_ (.A(_07484_),
    .B(_08307_),
    .C(net1654),
    .Y(_10885_));
 NAND2x1_ASAP7_75t_R _22586_ (.A(_07726_),
    .B(_07418_),
    .Y(_10896_));
 AO21x1_ASAP7_75t_R _22587_ (.A1(_10478_),
    .A2(_09221_),
    .B(_07484_),
    .Y(_10906_));
 AND4x1_ASAP7_75t_R _22588_ (.A(_10874_),
    .B(_10885_),
    .C(_10896_),
    .D(_10906_),
    .Y(_10917_));
 NOR2x2_ASAP7_75t_R _22589_ (.A(_06057_),
    .B(_08307_),
    .Y(_10928_));
 OA21x2_ASAP7_75t_R _22590_ (.A1(_10928_),
    .A2(_09052_),
    .B(_05881_),
    .Y(_10939_));
 INVx1_ASAP7_75t_R _22591_ (.A(_10939_),
    .Y(_10950_));
 AO21x1_ASAP7_75t_R _22592_ (.A1(_06430_),
    .A2(net3398),
    .B(_05892_),
    .Y(_10961_));
 AND3x1_ASAP7_75t_R _22593_ (.A(_10950_),
    .B(_07331_),
    .C(_10961_),
    .Y(_10972_));
 AO21x1_ASAP7_75t_R _22594_ (.A1(_07210_),
    .A2(_06277_),
    .B(_07583_),
    .Y(_10983_));
 AO21x1_ASAP7_75t_R _22595_ (.A1(_06123_),
    .A2(net1047),
    .B(_07583_),
    .Y(_10994_));
 NAND2x1_ASAP7_75t_R _22596_ (.A(_07561_),
    .B(_05804_),
    .Y(_11005_));
 AND3x1_ASAP7_75t_R _22597_ (.A(_10983_),
    .B(_10994_),
    .C(_11005_),
    .Y(_11016_));
 AO21x1_ASAP7_75t_R _22598_ (.A1(_07737_),
    .A2(_06145_),
    .B(_07682_),
    .Y(_11027_));
 AO21x1_ASAP7_75t_R _22599_ (.A1(_07517_),
    .A2(_07298_),
    .B(_07682_),
    .Y(_11038_));
 AO21x1_ASAP7_75t_R _22600_ (.A1(_05958_),
    .A2(_06925_),
    .B(_07682_),
    .Y(_11049_));
 AND4x1_ASAP7_75t_R _22601_ (.A(_11027_),
    .B(_11038_),
    .C(_11049_),
    .D(_07803_),
    .Y(_11060_));
 AND5x1_ASAP7_75t_R _22602_ (.A(_10863_),
    .B(_10917_),
    .C(_10972_),
    .D(_11016_),
    .E(_11060_),
    .Y(_11071_));
 NOR2x1_ASAP7_75t_R _22603_ (.A(_08121_),
    .B(_07265_),
    .Y(_11082_));
 INVx1_ASAP7_75t_R _22604_ (.A(_11082_),
    .Y(_11093_));
 AO21x1_ASAP7_75t_R _22605_ (.A1(_07210_),
    .A2(net3393),
    .B(_08285_),
    .Y(_11104_));
 NAND2x1_ASAP7_75t_R _22606_ (.A(_08230_),
    .B(_08252_),
    .Y(_11115_));
 NAND2x1_ASAP7_75t_R _22607_ (.A(_08230_),
    .B(_06968_),
    .Y(_11126_));
 AND4x1_ASAP7_75t_R _22608_ (.A(_08296_),
    .B(_11104_),
    .C(_11115_),
    .D(_11126_),
    .Y(_11137_));
 NAND2x1_ASAP7_75t_R _22609_ (.A(_06628_),
    .B(_09863_),
    .Y(_11148_));
 NAND2x1_ASAP7_75t_R _22610_ (.A(_05947_),
    .B(_09863_),
    .Y(_11159_));
 NAND2x1_ASAP7_75t_R _22611_ (.A(_08252_),
    .B(_09863_),
    .Y(_11170_));
 AND3x1_ASAP7_75t_R _22612_ (.A(_08143_),
    .B(_08186_),
    .C(_11170_),
    .Y(_11181_));
 AND5x1_ASAP7_75t_R _22613_ (.A(_11093_),
    .B(_11137_),
    .C(_11148_),
    .D(_11159_),
    .E(_11181_),
    .Y(_11192_));
 AND3x1_ASAP7_75t_R _22614_ (.A(_10852_),
    .B(_11071_),
    .C(_11192_),
    .Y(_11203_));
 NAND2x2_ASAP7_75t_R _22615_ (.A(_10709_),
    .B(_11203_),
    .Y(_11214_));
 INVx1_ASAP7_75t_R _48_59 (.A(clknet_leaf_15_clk),
    .Y(net464));
 XOR2x1_ASAP7_75t_R _22617_ (.A(_00385_),
    .Y(_11236_),
    .B(net3530));
 XNOR2x2_ASAP7_75t_R _22618_ (.A(_00482_),
    .B(_00524_),
    .Y(_11247_));
 XNOR2x1_ASAP7_75t_R _22619_ (.B(_11247_),
    .Y(_11258_),
    .A(_11236_));
 XOR2x1_ASAP7_75t_R _22620_ (.A(_11214_),
    .Y(_11269_),
    .B(_11258_));
 INVx1_ASAP7_75t_R _48_58 (.A(clknet_leaf_12_clk),
    .Y(net463));
 INVx1_ASAP7_75t_R _48_57 (.A(clknet_leaf_1_clk),
    .Y(net462));
 INVx1_ASAP7_75t_R _48_56 (.A(clknet_leaf_11_clk),
    .Y(net461));
 AND2x2_ASAP7_75t_R _22624_ (.A(net403),
    .B(net4164),
    .Y(_11313_));
 AO21x1_ASAP7_75t_R _22625_ (.A1(_11269_),
    .A2(net400),
    .B(_11313_),
    .Y(_00375_));
 NAND2x1_ASAP7_75t_R _22626_ (.A(_07100_),
    .B(_08362_),
    .Y(_11334_));
 AO21x1_ASAP7_75t_R _22627_ (.A1(net3392),
    .A2(_06925_),
    .B(_08461_),
    .Y(_11345_));
 AO21x1_ASAP7_75t_R _22628_ (.A1(_07342_),
    .A2(net1047),
    .B(_08461_),
    .Y(_11356_));
 NOR2x1_ASAP7_75t_R _22629_ (.A(_06222_),
    .B(_08461_),
    .Y(_11367_));
 INVx1_ASAP7_75t_R _22630_ (.A(_11367_),
    .Y(_11378_));
 NAND2x1_ASAP7_75t_R _22631_ (.A(_06968_),
    .B(_08362_),
    .Y(_11389_));
 AND5x1_ASAP7_75t_R _22632_ (.A(_11334_),
    .B(_11345_),
    .C(_11356_),
    .D(_11378_),
    .E(_11389_),
    .Y(_11400_));
 AO21x1_ASAP7_75t_R _22633_ (.A1(_07210_),
    .A2(_10478_),
    .B(_08406_),
    .Y(_11411_));
 AO21x1_ASAP7_75t_R _22634_ (.A1(_07517_),
    .A2(_07265_),
    .B(_08406_),
    .Y(_11422_));
 AND4x1_ASAP7_75t_R _22635_ (.A(_11411_),
    .B(_11422_),
    .C(_09159_),
    .D(_10291_),
    .Y(_11433_));
 AO21x1_ASAP7_75t_R _22636_ (.A1(_07111_),
    .A2(_07265_),
    .B(_08669_),
    .Y(_11444_));
 AO21x1_ASAP7_75t_R _22637_ (.A1(_07737_),
    .A2(_10478_),
    .B(_08669_),
    .Y(_11454_));
 AND3x1_ASAP7_75t_R _22638_ (.A(_09008_),
    .B(_11444_),
    .C(_11454_),
    .Y(_11465_));
 INVx1_ASAP7_75t_R _48_55 (.A(clknet_leaf_1_clk),
    .Y(net460));
 OA211x2_ASAP7_75t_R _22640_ (.A1(_06397_),
    .A2(net2132),
    .B(_08570_),
    .C(_06727_),
    .Y(_11487_));
 INVx1_ASAP7_75t_R _22641_ (.A(_11487_),
    .Y(_11498_));
 OR3x1_ASAP7_75t_R _22642_ (.A(_08625_),
    .B(_06112_),
    .C(_06057_),
    .Y(_11509_));
 AO21x1_ASAP7_75t_R _22643_ (.A1(_10533_),
    .A2(net3392),
    .B(_08625_),
    .Y(_11520_));
 AO21x1_ASAP7_75t_R _22644_ (.A1(net3403),
    .A2(_07572_),
    .B(_08625_),
    .Y(_11531_));
 AND4x1_ASAP7_75t_R _22645_ (.A(_11498_),
    .B(_11509_),
    .C(_11520_),
    .D(_11531_),
    .Y(_11542_));
 AND4x2_ASAP7_75t_R _22646_ (.A(_11400_),
    .B(_11433_),
    .C(_11465_),
    .D(_11542_),
    .Y(_11553_));
 OA21x2_ASAP7_75t_R _22647_ (.A1(_06419_),
    .A2(_05947_),
    .B(_06760_),
    .Y(_11564_));
 OR3x1_ASAP7_75t_R _22648_ (.A(_11564_),
    .B(_06782_),
    .C(_09190_),
    .Y(_11575_));
 AND2x2_ASAP7_75t_R _22649_ (.A(_07561_),
    .B(_06760_),
    .Y(_11586_));
 OA21x2_ASAP7_75t_R _22650_ (.A1(_09951_),
    .A2(_06079_),
    .B(_06760_),
    .Y(_11597_));
 OR4x2_ASAP7_75t_R _22651_ (.A(_11575_),
    .B(_11586_),
    .C(_09232_),
    .D(_11597_),
    .Y(_11608_));
 OR3x1_ASAP7_75t_R _22652_ (.A(_06870_),
    .B(_06881_),
    .C(_06892_),
    .Y(_11619_));
 NOR2x1_ASAP7_75t_R _22653_ (.A(_06925_),
    .B(_06826_),
    .Y(_11630_));
 AND2x2_ASAP7_75t_R _22654_ (.A(_06815_),
    .B(_07254_),
    .Y(_11641_));
 OR5x2_ASAP7_75t_R _22655_ (.A(_11619_),
    .B(_07144_),
    .C(_07133_),
    .D(_11630_),
    .E(_11641_),
    .Y(_11652_));
 NOR2x2_ASAP7_75t_R _22656_ (.A(_11608_),
    .B(_11652_),
    .Y(_11663_));
 NOR2x1_ASAP7_75t_R _22657_ (.A(_09221_),
    .B(_06474_),
    .Y(_11674_));
 OR5x2_ASAP7_75t_R _22658_ (.A(_06507_),
    .B(_09359_),
    .C(_06573_),
    .D(_11674_),
    .E(_09337_),
    .Y(_11685_));
 NOR2x1_ASAP7_75t_R _22659_ (.A(net1653),
    .B(_06474_),
    .Y(_11696_));
 OA21x2_ASAP7_75t_R _22660_ (.A1(_11696_),
    .A2(_09401_),
    .B(net1146),
    .Y(_11707_));
 AO221x2_ASAP7_75t_R _22661_ (.A1(_06968_),
    .A2(_06463_),
    .B1(_00424_),
    .B2(_11707_),
    .C(_10577_),
    .Y(_11718_));
 AND2x2_ASAP7_75t_R _22662_ (.A(_07561_),
    .B(_06595_),
    .Y(_11729_));
 NOR2x1_ASAP7_75t_R _22663_ (.A(_06606_),
    .B(_07111_),
    .Y(_11740_));
 OR5x2_ASAP7_75t_R _22664_ (.A(_11729_),
    .B(_11740_),
    .C(_09433_),
    .D(_10665_),
    .E(_10643_),
    .Y(_11751_));
 NOR3x2_ASAP7_75t_R _22665_ (.B(_11718_),
    .C(_11751_),
    .Y(_11762_),
    .A(_11685_));
 NAND3x2_ASAP7_75t_R _22666_ (.B(_11663_),
    .C(_11762_),
    .Y(_11773_),
    .A(_11553_));
 NOR2x1_ASAP7_75t_R _22667_ (.A(_06123_),
    .B(_07682_),
    .Y(_11784_));
 INVx1_ASAP7_75t_R _22668_ (.A(_11784_),
    .Y(_11795_));
 OA211x2_ASAP7_75t_R _22669_ (.A1(_06397_),
    .A2(net2131),
    .B(_05804_),
    .C(_06914_),
    .Y(_11806_));
 INVx1_ASAP7_75t_R _22670_ (.A(_11806_),
    .Y(_11817_));
 AO21x1_ASAP7_75t_R _22671_ (.A1(_07111_),
    .A2(_07517_),
    .B(_07583_),
    .Y(_11828_));
 NAND2x1_ASAP7_75t_R _22672_ (.A(_09951_),
    .B(_05804_),
    .Y(_11839_));
 AND4x1_ASAP7_75t_R _22673_ (.A(_11817_),
    .B(_07605_),
    .C(_11828_),
    .D(_11839_),
    .Y(_11850_));
 AO21x1_ASAP7_75t_R _22674_ (.A1(_07517_),
    .A2(_07298_),
    .B(_05892_),
    .Y(_11861_));
 AO21x1_ASAP7_75t_R _22675_ (.A1(net3392),
    .A2(_10533_),
    .B(_05892_),
    .Y(_11872_));
 AO21x1_ASAP7_75t_R _22676_ (.A1(_07342_),
    .A2(_06123_),
    .B(_05892_),
    .Y(_11883_));
 NAND2x1_ASAP7_75t_R _22677_ (.A(_07561_),
    .B(_05881_),
    .Y(_11894_));
 AND4x1_ASAP7_75t_R _22678_ (.A(_11861_),
    .B(_11872_),
    .C(_11883_),
    .D(_11894_),
    .Y(_11904_));
 AO21x1_ASAP7_75t_R _22679_ (.A1(_07265_),
    .A2(_07517_),
    .B(_07484_),
    .Y(_11915_));
 NOR2x1_ASAP7_75t_R _22680_ (.A(_06145_),
    .B(_07484_),
    .Y(_11926_));
 INVx1_ASAP7_75t_R _22681_ (.A(_11926_),
    .Y(_11937_));
 OA211x2_ASAP7_75t_R _22682_ (.A1(_07484_),
    .A2(net3392),
    .B(_11915_),
    .C(_11937_),
    .Y(_11948_));
 AO21x1_ASAP7_75t_R _22683_ (.A1(_07111_),
    .A2(_07265_),
    .B(_07682_),
    .Y(_11959_));
 AND5x1_ASAP7_75t_R _22684_ (.A(_11795_),
    .B(_11850_),
    .C(_11904_),
    .D(_11948_),
    .E(_11959_),
    .Y(_11970_));
 INVx1_ASAP7_75t_R _22685_ (.A(_09929_),
    .Y(_11981_));
 AND2x2_ASAP7_75t_R _22686_ (.A(_09863_),
    .B(_06518_),
    .Y(_11992_));
 INVx1_ASAP7_75t_R _22687_ (.A(_11992_),
    .Y(_12003_));
 NAND2x1_ASAP7_75t_R _22688_ (.A(_06079_),
    .B(_09863_),
    .Y(_12014_));
 AND5x1_ASAP7_75t_R _22689_ (.A(_11981_),
    .B(_11148_),
    .C(_12003_),
    .D(_11170_),
    .E(_12014_),
    .Y(_12025_));
 OA211x2_ASAP7_75t_R _22690_ (.A1(_06397_),
    .A2(net2135),
    .B(_08000_),
    .C(_06914_),
    .Y(_12036_));
 NOR2x1_ASAP7_75t_R _22691_ (.A(_09819_),
    .B(_12036_),
    .Y(_12047_));
 AO21x1_ASAP7_75t_R _22692_ (.A1(_07342_),
    .A2(net2055),
    .B(_08011_),
    .Y(_12058_));
 OA211x2_ASAP7_75t_R _22693_ (.A1(_07210_),
    .A2(_08011_),
    .B(_12047_),
    .C(_12058_),
    .Y(_12069_));
 NOR2x1_ASAP7_75t_R _22694_ (.A(_06057_),
    .B(_07879_),
    .Y(_12080_));
 NOR2x1_ASAP7_75t_R _22695_ (.A(_12080_),
    .B(_09984_),
    .Y(_12091_));
 NOR2x1_ASAP7_75t_R _22696_ (.A(_06222_),
    .B(_07879_),
    .Y(_12102_));
 INVx1_ASAP7_75t_R _22697_ (.A(_12102_),
    .Y(_12113_));
 AO21x1_ASAP7_75t_R _22698_ (.A1(_07265_),
    .A2(_07517_),
    .B(_07879_),
    .Y(_12124_));
 AND4x1_ASAP7_75t_R _22699_ (.A(_12091_),
    .B(_07967_),
    .C(_12113_),
    .D(_12124_),
    .Y(_12135_));
 AO21x1_ASAP7_75t_R _22700_ (.A1(_07517_),
    .A2(_07298_),
    .B(_08285_),
    .Y(_12146_));
 AO21x1_ASAP7_75t_R _22701_ (.A1(_10478_),
    .A2(net3394),
    .B(_08285_),
    .Y(_12157_));
 AND4x1_ASAP7_75t_R _22702_ (.A(_12146_),
    .B(_12157_),
    .C(_11115_),
    .D(_11126_),
    .Y(_12168_));
 AND4x1_ASAP7_75t_R _22703_ (.A(_12025_),
    .B(_12069_),
    .C(_12135_),
    .D(_12168_),
    .Y(_12179_));
 AND2x2_ASAP7_75t_R _22704_ (.A(_11970_),
    .B(_12179_),
    .Y(_12190_));
 INVx1_ASAP7_75t_R _22705_ (.A(_12190_),
    .Y(_12201_));
 NOR2x2_ASAP7_75t_R _22706_ (.A(_11773_),
    .B(_12201_),
    .Y(_12212_));
 INVx1_ASAP7_75t_R _48_54 (.A(clknet_leaf_1_clk),
    .Y(net459));
 XNOR2x2_ASAP7_75t_R _22708_ (.A(_00481_),
    .B(_00523_),
    .Y(_12234_));
 INVx1_ASAP7_75t_R _48_53 (.A(clknet_leaf_2_clk),
    .Y(net458));
 XOR2x1_ASAP7_75t_R _22710_ (.A(_00386_),
    .Y(_12256_),
    .B(net3534));
 XOR2x1_ASAP7_75t_R _22711_ (.A(_12234_),
    .Y(_12267_),
    .B(_12256_));
 XOR2x1_ASAP7_75t_R _22712_ (.A(_12212_),
    .Y(_12278_),
    .B(_12267_));
 AND2x2_ASAP7_75t_R _22713_ (.A(net404),
    .B(net4130),
    .Y(_12289_));
 AO21x1_ASAP7_75t_R _22714_ (.A1(_12278_),
    .A2(net399),
    .B(_12289_),
    .Y(_00378_));
 NAND2x2_ASAP7_75t_R _22715_ (.A(net1619),
    .B(_06914_),
    .Y(_12310_));
 OR3x1_ASAP7_75t_R _22716_ (.A(_12310_),
    .B(_07857_),
    .C(_05760_),
    .Y(_12321_));
 INVx1_ASAP7_75t_R _22717_ (.A(_09885_),
    .Y(_12332_));
 AND4x1_ASAP7_75t_R _22718_ (.A(_11378_),
    .B(_12321_),
    .C(_12332_),
    .D(_08186_),
    .Y(_12343_));
 AO21x1_ASAP7_75t_R _22719_ (.A1(_08669_),
    .A2(_06771_),
    .B(_07265_),
    .Y(_12354_));
 AND4x1_ASAP7_75t_R _22720_ (.A(_12343_),
    .B(_08942_),
    .C(_09830_),
    .D(_12354_),
    .Y(_12365_));
 NAND2x1_ASAP7_75t_R _22721_ (.A(_10928_),
    .B(_05881_),
    .Y(_12376_));
 NAND2x1_ASAP7_75t_R _22722_ (.A(_05881_),
    .B(_07100_),
    .Y(_12387_));
 AND4x1_ASAP7_75t_R _22723_ (.A(_10390_),
    .B(_12387_),
    .C(_10819_),
    .D(_11839_),
    .Y(_12398_));
 NOR2x1_ASAP7_75t_R _22724_ (.A(_07298_),
    .B(_08406_),
    .Y(_12408_));
 INVx1_ASAP7_75t_R _22725_ (.A(_12408_),
    .Y(_12419_));
 AO21x1_ASAP7_75t_R _22726_ (.A1(net1047),
    .A2(net2055),
    .B(_08121_),
    .Y(_12430_));
 NAND2x1_ASAP7_75t_R _22727_ (.A(_08603_),
    .B(_07781_),
    .Y(_12441_));
 AND5x1_ASAP7_75t_R _22728_ (.A(_12376_),
    .B(_12398_),
    .C(_12419_),
    .D(_12430_),
    .E(_12441_),
    .Y(_12452_));
 NAND2x1_ASAP7_75t_R _22729_ (.A(_12365_),
    .B(_12452_),
    .Y(_12463_));
 OR4x1_ASAP7_75t_R _22730_ (.A(_07111_),
    .B(_06353_),
    .C(_05749_),
    .D(_06452_),
    .Y(_12474_));
 INVx1_ASAP7_75t_R _22731_ (.A(_10665_),
    .Y(_12485_));
 AND4x1_ASAP7_75t_R _22732_ (.A(_12474_),
    .B(_07901_),
    .C(_07067_),
    .D(_12485_),
    .Y(_12496_));
 OA211x2_ASAP7_75t_R _22733_ (.A1(_07210_),
    .A2(_07583_),
    .B(_06013_),
    .C(_12113_),
    .Y(_12507_));
 NOR2x1_ASAP7_75t_R _22734_ (.A(_07682_),
    .B(_06090_),
    .Y(_12518_));
 INVx1_ASAP7_75t_R _22735_ (.A(_12518_),
    .Y(_12529_));
 OA21x2_ASAP7_75t_R _22736_ (.A1(net3403),
    .A2(_07484_),
    .B(_12529_),
    .Y(_12540_));
 OA211x2_ASAP7_75t_R _22737_ (.A1(_06826_),
    .A2(_06057_),
    .B(_12507_),
    .C(_12540_),
    .Y(_12551_));
 NAND2x1_ASAP7_75t_R _22738_ (.A(_12496_),
    .B(_12551_),
    .Y(_12562_));
 AO22x1_ASAP7_75t_R _22739_ (.A1(_06727_),
    .A2(_08000_),
    .B1(_08417_),
    .B2(_06266_),
    .Y(_12573_));
 AO21x1_ASAP7_75t_R _22740_ (.A1(_06463_),
    .A2(_07287_),
    .B(_06288_),
    .Y(_12584_));
 NAND2x1_ASAP7_75t_R _22741_ (.A(_06419_),
    .B(_08516_),
    .Y(_12595_));
 NAND2x1_ASAP7_75t_R _22742_ (.A(_08986_),
    .B(_12595_),
    .Y(_12606_));
 OR3x1_ASAP7_75t_R _22743_ (.A(_12584_),
    .B(_11992_),
    .C(_12606_),
    .Y(_12617_));
 AO21x1_ASAP7_75t_R _22744_ (.A1(_08307_),
    .A2(_12573_),
    .B(_12617_),
    .Y(_12628_));
 AO32x1_ASAP7_75t_R _22745_ (.A1(_06112_),
    .A2(_06727_),
    .A3(_08000_),
    .B1(_06760_),
    .B2(_06968_),
    .Y(_12639_));
 AND2x2_ASAP7_75t_R _22746_ (.A(_08417_),
    .B(_10928_),
    .Y(_12650_));
 AND2x2_ASAP7_75t_R _22747_ (.A(_05804_),
    .B(_08603_),
    .Y(_12661_));
 NOR2x1_ASAP7_75t_R _22748_ (.A(_07572_),
    .B(_07484_),
    .Y(_12672_));
 AO21x1_ASAP7_75t_R _22749_ (.A1(_08417_),
    .A2(_06968_),
    .B(_12672_),
    .Y(_12683_));
 OR4x1_ASAP7_75t_R _22750_ (.A(_12639_),
    .B(_12650_),
    .C(_12661_),
    .D(_12683_),
    .Y(_12694_));
 AO32x1_ASAP7_75t_R _22751_ (.A1(_06957_),
    .A2(_07418_),
    .A3(_06727_),
    .B1(_06266_),
    .B2(_08000_),
    .Y(_12705_));
 OR3x1_ASAP7_75t_R _22752_ (.A(_08559_),
    .B(_08439_),
    .C(_12705_),
    .Y(_12716_));
 OR3x1_ASAP7_75t_R _22753_ (.A(_12628_),
    .B(_12694_),
    .C(_12716_),
    .Y(_12727_));
 OR3x1_ASAP7_75t_R _22754_ (.A(_12463_),
    .B(_12562_),
    .C(_12727_),
    .Y(_12738_));
 INVx1_ASAP7_75t_R _22755_ (.A(_09687_),
    .Y(_12749_));
 OR4x1_ASAP7_75t_R _22756_ (.A(_09085_),
    .B(_07429_),
    .C(_09232_),
    .D(_07133_),
    .Y(_12760_));
 AND3x1_ASAP7_75t_R _22757_ (.A(_08417_),
    .B(_06266_),
    .C(_06946_),
    .Y(_12771_));
 AND3x1_ASAP7_75t_R _22758_ (.A(_05804_),
    .B(_05925_),
    .C(_05991_),
    .Y(_12782_));
 OR5x1_ASAP7_75t_R _22759_ (.A(_12749_),
    .B(_12760_),
    .C(_12771_),
    .D(_10599_),
    .E(_12782_),
    .Y(_12793_));
 AND2x2_ASAP7_75t_R _22760_ (.A(_07254_),
    .B(_08230_),
    .Y(_12804_));
 AO21x1_ASAP7_75t_R _22761_ (.A1(_08230_),
    .A2(net2349),
    .B(_12804_),
    .Y(_12815_));
 AO21x1_ASAP7_75t_R _22762_ (.A1(_06123_),
    .A2(_06145_),
    .B(_07484_),
    .Y(_12826_));
 INVx1_ASAP7_75t_R _22763_ (.A(_12826_),
    .Y(_12837_));
 OAI22x1_ASAP7_75t_R _22764_ (.A1(_08285_),
    .A2(_06738_),
    .B1(_06090_),
    .B2(_07484_),
    .Y(_12848_));
 OR3x1_ASAP7_75t_R _22765_ (.A(_12815_),
    .B(_12837_),
    .C(_12848_),
    .Y(_12859_));
 INVx1_ASAP7_75t_R _22766_ (.A(_08898_),
    .Y(_12869_));
 OA21x2_ASAP7_75t_R _22767_ (.A1(_12869_),
    .A2(_06617_),
    .B(_06397_),
    .Y(_12880_));
 INVx1_ASAP7_75t_R _22768_ (.A(_11104_),
    .Y(_12891_));
 AO21x1_ASAP7_75t_R _22769_ (.A1(_09052_),
    .A2(_08230_),
    .B(_12891_),
    .Y(_12902_));
 AND2x2_ASAP7_75t_R _22770_ (.A(_06760_),
    .B(_06628_),
    .Y(_12913_));
 OR4x1_ASAP7_75t_R _22771_ (.A(_12913_),
    .B(_06870_),
    .C(_09412_),
    .D(_06661_),
    .Y(_12924_));
 OR5x1_ASAP7_75t_R _22772_ (.A(_10061_),
    .B(_12859_),
    .C(_12880_),
    .D(_12902_),
    .E(_12924_),
    .Y(_12935_));
 AO32x1_ASAP7_75t_R _22773_ (.A1(_08307_),
    .A2(net2586),
    .A3(_07868_),
    .B1(_06628_),
    .B2(_08570_),
    .Y(_12946_));
 AO32x1_ASAP7_75t_R _22774_ (.A1(_00422_),
    .A2(_06255_),
    .A3(_06804_),
    .B1(_08230_),
    .B2(_06936_),
    .Y(_12957_));
 AO21x1_ASAP7_75t_R _22775_ (.A1(_09907_),
    .A2(_09369_),
    .B(_11564_),
    .Y(_12968_));
 OR5x1_ASAP7_75t_R _22776_ (.A(_10676_),
    .B(_12946_),
    .C(_11707_),
    .D(_12957_),
    .E(_12968_),
    .Y(_12979_));
 OR3x1_ASAP7_75t_R _22777_ (.A(_12793_),
    .B(_12935_),
    .C(_12979_),
    .Y(_12990_));
 NOR2x2_ASAP7_75t_R _22778_ (.A(_12738_),
    .B(_12990_),
    .Y(_13001_));
 INVx1_ASAP7_75t_R _48_52 (.A(clknet_leaf_2_clk),
    .Y(net457));
 XOR2x2_ASAP7_75t_R _22780_ (.A(_00480_),
    .B(_00522_),
    .Y(_13023_));
 INVx1_ASAP7_75t_R _48_51 (.A(clknet_leaf_7_clk),
    .Y(net456));
 INVx1_ASAP7_75t_R _48_50 (.A(clknet_leaf_6_clk),
    .Y(net455));
 XOR2x1_ASAP7_75t_R _22783_ (.A(_00387_),
    .Y(_13056_),
    .B(_00448_));
 XNOR2x1_ASAP7_75t_R _22784_ (.B(_13056_),
    .Y(_13067_),
    .A(_13023_));
 XOR2x1_ASAP7_75t_R _22785_ (.A(_13001_),
    .Y(_13078_),
    .B(_13067_));
 AND2x2_ASAP7_75t_R _22786_ (.A(net405),
    .B(net73),
    .Y(_13089_));
 AO21x1_ASAP7_75t_R _22787_ (.A1(_13078_),
    .A2(net399),
    .B(_13089_),
    .Y(_00379_));
 INVx1_ASAP7_75t_R _48_49 (.A(clknet_leaf_8_clk),
    .Y(net454));
 INVx1_ASAP7_75t_R _48 (.A(clknet_leaf_11_clk),
    .Y(net453));
 XNOR2x1_ASAP7_75t_R _22790_ (.B(_00479_),
    .Y(_13132_),
    .A(_00447_));
 XNOR2x2_ASAP7_75t_R _22791_ (.A(_00498_),
    .B(_00521_),
    .Y(_13143_));
 XNOR2x1_ASAP7_75t_R _22792_ (.B(_13143_),
    .Y(_13154_),
    .A(_13132_));
 OR5x1_ASAP7_75t_R _22793_ (.A(_08263_),
    .B(_12815_),
    .C(_08241_),
    .D(_10028_),
    .E(_12891_),
    .Y(_13165_));
 NAND2x1_ASAP7_75t_R _22794_ (.A(_06957_),
    .B(_06727_),
    .Y(_13176_));
 AO21x1_ASAP7_75t_R _22795_ (.A1(_06222_),
    .A2(net3403),
    .B(_07879_),
    .Y(_13187_));
 OA211x2_ASAP7_75t_R _22796_ (.A1(_07879_),
    .A2(_13176_),
    .B(_13187_),
    .C(_07967_),
    .Y(_13197_));
 NOR2x1_ASAP7_75t_R _22797_ (.A(_08011_),
    .B(_07265_),
    .Y(_13208_));
 INVx1_ASAP7_75t_R _22798_ (.A(_13208_),
    .Y(_13219_));
 AND4x1_ASAP7_75t_R _22799_ (.A(_08066_),
    .B(_10775_),
    .C(_10797_),
    .D(_13219_),
    .Y(_13230_));
 NAND2x1_ASAP7_75t_R _22800_ (.A(_13197_),
    .B(_13230_),
    .Y(_13241_));
 OA21x2_ASAP7_75t_R _22801_ (.A1(_08252_),
    .A2(_07726_),
    .B(_09863_),
    .Y(_13252_));
 OR4x1_ASAP7_75t_R _22802_ (.A(_09929_),
    .B(_13252_),
    .C(_09885_),
    .D(_11992_),
    .Y(_13263_));
 OR3x1_ASAP7_75t_R _22803_ (.A(_13165_),
    .B(_13241_),
    .C(_13263_),
    .Y(_13274_));
 AO21x1_ASAP7_75t_R _22804_ (.A1(_06090_),
    .A2(net2055),
    .B(_05892_),
    .Y(_13285_));
 INVx1_ASAP7_75t_R _22805_ (.A(_06288_),
    .Y(_13296_));
 AND5x1_ASAP7_75t_R _22806_ (.A(_09643_),
    .B(_09720_),
    .C(_13285_),
    .D(_06013_),
    .E(_13296_),
    .Y(_13307_));
 AO21x1_ASAP7_75t_R _22807_ (.A1(_06222_),
    .A2(_09221_),
    .B(_07484_),
    .Y(_13318_));
 AO21x1_ASAP7_75t_R _22808_ (.A1(_07342_),
    .A2(_06123_),
    .B(_07484_),
    .Y(_13329_));
 AND4x1_ASAP7_75t_R _22809_ (.A(_09599_),
    .B(_10885_),
    .C(_13318_),
    .D(_13329_),
    .Y(_13340_));
 NAND2x1_ASAP7_75t_R _22810_ (.A(_06419_),
    .B(_07781_),
    .Y(_13351_));
 AND3x1_ASAP7_75t_R _22811_ (.A(_07715_),
    .B(_12529_),
    .C(_09577_),
    .Y(_13362_));
 AND3x1_ASAP7_75t_R _22812_ (.A(_13340_),
    .B(_13351_),
    .C(_13362_),
    .Y(_13373_));
 AND3x1_ASAP7_75t_R _22813_ (.A(_05804_),
    .B(_08603_),
    .C(net1012),
    .Y(_13384_));
 INVx1_ASAP7_75t_R _22814_ (.A(_13384_),
    .Y(_13395_));
 AO21x1_ASAP7_75t_R _22815_ (.A1(_06222_),
    .A2(_06277_),
    .B(_07583_),
    .Y(_13406_));
 AO21x1_ASAP7_75t_R _22816_ (.A1(_07342_),
    .A2(net1047),
    .B(_07583_),
    .Y(_13417_));
 AND4x1_ASAP7_75t_R _22817_ (.A(_13395_),
    .B(_07649_),
    .C(_13406_),
    .D(_13417_),
    .Y(_13428_));
 AND3x1_ASAP7_75t_R _22818_ (.A(_13307_),
    .B(_13373_),
    .C(_13428_),
    .Y(_13439_));
 INVx1_ASAP7_75t_R _22819_ (.A(_13439_),
    .Y(_13450_));
 NOR2x2_ASAP7_75t_R _22820_ (.A(_13274_),
    .B(_13450_),
    .Y(_13461_));
 OA211x2_ASAP7_75t_R _22821_ (.A1(_06397_),
    .A2(net2131),
    .B(_08570_),
    .C(_06266_),
    .Y(_13472_));
 INVx1_ASAP7_75t_R _22822_ (.A(_13472_),
    .Y(_13483_));
 NAND2x1_ASAP7_75t_R _22823_ (.A(_07254_),
    .B(_08570_),
    .Y(_13494_));
 OR3x1_ASAP7_75t_R _22824_ (.A(_08625_),
    .B(_06397_),
    .C(_06057_),
    .Y(_13505_));
 AND5x2_ASAP7_75t_R _22825_ (.A(_10269_),
    .B(_13483_),
    .C(_13494_),
    .D(_13505_),
    .E(_08920_),
    .Y(_13516_));
 AO21x1_ASAP7_75t_R _22826_ (.A1(_06738_),
    .A2(_06925_),
    .B(_08406_),
    .Y(_13527_));
 AO21x1_ASAP7_75t_R _22827_ (.A1(_07210_),
    .A2(_06222_),
    .B(_08461_),
    .Y(_13537_));
 AO21x1_ASAP7_75t_R _22828_ (.A1(net2055),
    .A2(_07737_),
    .B(_08461_),
    .Y(_13548_));
 AND5x2_ASAP7_75t_R _22829_ (.A(_11389_),
    .B(_11411_),
    .C(_13527_),
    .D(_13537_),
    .E(_13548_),
    .Y(_13559_));
 NOR2x1_ASAP7_75t_R _22830_ (.A(_06925_),
    .B(_08669_),
    .Y(_13570_));
 INVx1_ASAP7_75t_R _22831_ (.A(_13570_),
    .Y(_13581_));
 OR3x1_ASAP7_75t_R _22832_ (.A(_08669_),
    .B(net3401),
    .C(net1146),
    .Y(_13592_));
 NAND2x1_ASAP7_75t_R _22833_ (.A(net2582),
    .B(_08516_),
    .Y(_13603_));
 AND5x2_ASAP7_75t_R _22834_ (.A(_13581_),
    .B(_13592_),
    .C(_08986_),
    .D(_12595_),
    .E(_13603_),
    .Y(_13614_));
 NAND3x2_ASAP7_75t_R _22835_ (.B(_13559_),
    .C(_13614_),
    .Y(_13625_),
    .A(_13516_));
 NOR2x1_ASAP7_75t_R _22836_ (.A(_09221_),
    .B(_06606_),
    .Y(_13636_));
 OR4x1_ASAP7_75t_R _22837_ (.A(_11729_),
    .B(_09412_),
    .C(_13636_),
    .D(_09401_),
    .Y(_13647_));
 AND3x1_ASAP7_75t_R _22838_ (.A(_06463_),
    .B(net2133),
    .C(_06266_),
    .Y(_13658_));
 OA21x2_ASAP7_75t_R _22839_ (.A1(_06628_),
    .A2(net2582),
    .B(_06463_),
    .Y(_13669_));
 OR5x2_ASAP7_75t_R _22840_ (.A(_06573_),
    .B(_13647_),
    .C(_11696_),
    .D(_13658_),
    .E(_13669_),
    .Y(_13680_));
 AND3x1_ASAP7_75t_R _22841_ (.A(_06815_),
    .B(net2133),
    .C(net2586),
    .Y(_13691_));
 AO21x1_ASAP7_75t_R _22842_ (.A1(_09052_),
    .A2(_06815_),
    .B(_13691_),
    .Y(_13702_));
 OR3x1_ASAP7_75t_R _22843_ (.A(_07166_),
    .B(_11641_),
    .C(_09274_),
    .Y(_13713_));
 NOR2x1_ASAP7_75t_R _22844_ (.A(_12310_),
    .B(_06771_),
    .Y(_13724_));
 AO21x1_ASAP7_75t_R _22845_ (.A1(_06760_),
    .A2(_07100_),
    .B(_13724_),
    .Y(_13735_));
 AO21x1_ASAP7_75t_R _22846_ (.A1(_06760_),
    .A2(_06540_),
    .B(_11586_),
    .Y(_13746_));
 OR4x2_ASAP7_75t_R _22847_ (.A(_13702_),
    .B(_13713_),
    .C(_13735_),
    .D(_13746_),
    .Y(_13757_));
 NOR3x2_ASAP7_75t_R _22848_ (.B(_13680_),
    .C(_13757_),
    .Y(_13768_),
    .A(_13625_));
 NAND2x2_ASAP7_75t_R _22849_ (.A(_13461_),
    .B(_13768_),
    .Y(_13779_));
 NOR2x2_ASAP7_75t_R _22850_ (.A(_13779_),
    .B(_10127_),
    .Y(_13790_));
 NAND2x1_ASAP7_75t_R _22851_ (.A(_13154_),
    .B(_13790_),
    .Y(_13801_));
 INVx1_ASAP7_75t_R _22852_ (.A(_13779_),
    .Y(_13812_));
 AO21x1_ASAP7_75t_R _22853_ (.A1(_13812_),
    .A2(net2609),
    .B(_13154_),
    .Y(_13822_));
 NAND2x1_ASAP7_75t_R _22854_ (.A(_13801_),
    .B(_13822_),
    .Y(_13833_));
 INVx1_ASAP7_75t_R net399_47 (.A(clknet_leaf_11_clk),
    .Y(net452));
 NAND2x2_ASAP7_75t_R _22856_ (.A(net403),
    .B(net4044),
    .Y(_13855_));
 OAI21x1_ASAP7_75t_R _22857_ (.A1(net404),
    .A2(_13833_),
    .B(_13855_),
    .Y(_00380_));
 INVx1_ASAP7_75t_R _22858_ (.A(net4056),
    .Y(_13875_));
 NOR2x1_ASAP7_75t_R _22859_ (.A(_07210_),
    .B(_07583_),
    .Y(_13886_));
 AO21x1_ASAP7_75t_R _22860_ (.A1(_05804_),
    .A2(_07726_),
    .B(_12749_),
    .Y(_13897_));
 NOR2x1_ASAP7_75t_R _22861_ (.A(_13886_),
    .B(_13897_),
    .Y(_13907_));
 OA211x2_ASAP7_75t_R _22862_ (.A1(net2858),
    .A2(_07583_),
    .B(_13907_),
    .C(_11817_),
    .Y(_13918_));
 NOR2x1_ASAP7_75t_R _22863_ (.A(_10939_),
    .B(_06035_),
    .Y(_13928_));
 AO21x1_ASAP7_75t_R _22864_ (.A1(_07265_),
    .A2(_07298_),
    .B(_07484_),
    .Y(_13939_));
 INVx1_ASAP7_75t_R _22865_ (.A(_13939_),
    .Y(_13949_));
 AO21x1_ASAP7_75t_R _22866_ (.A1(_07418_),
    .A2(_05947_),
    .B(_13949_),
    .Y(_13960_));
 NOR2x1_ASAP7_75t_R _22867_ (.A(_06222_),
    .B(_07484_),
    .Y(_13970_));
 OR3x1_ASAP7_75t_R _22868_ (.A(_13960_),
    .B(_13970_),
    .C(_12837_),
    .Y(_13981_));
 INVx1_ASAP7_75t_R _22869_ (.A(_13981_),
    .Y(_13992_));
 NOR2x1_ASAP7_75t_R _22870_ (.A(_07682_),
    .B(_07671_),
    .Y(_14003_));
 INVx1_ASAP7_75t_R _22871_ (.A(_14003_),
    .Y(_14013_));
 AND4x1_ASAP7_75t_R _22872_ (.A(_07770_),
    .B(_09577_),
    .C(_11795_),
    .D(_14013_),
    .Y(_14024_));
 AND4x2_ASAP7_75t_R _22873_ (.A(_13918_),
    .B(_13928_),
    .C(_13992_),
    .D(_14024_),
    .Y(_14034_));
 AND3x1_ASAP7_75t_R _22874_ (.A(_12124_),
    .B(_07923_),
    .C(_07967_),
    .Y(_14044_));
 AO21x1_ASAP7_75t_R _22875_ (.A1(_07517_),
    .A2(_07298_),
    .B(_08011_),
    .Y(_14055_));
 AO21x1_ASAP7_75t_R _22876_ (.A1(_10478_),
    .A2(net3403),
    .B(_08011_),
    .Y(_14066_));
 AND5x2_ASAP7_75t_R _22877_ (.A(_09786_),
    .B(_12091_),
    .C(_14044_),
    .D(_14055_),
    .E(_14066_),
    .Y(_14076_));
 NOR2x1_ASAP7_75t_R _22878_ (.A(_06430_),
    .B(_08285_),
    .Y(_14087_));
 AO21x1_ASAP7_75t_R _22879_ (.A1(_08230_),
    .A2(_06936_),
    .B(_14087_),
    .Y(_14097_));
 AND3x1_ASAP7_75t_R _22880_ (.A(_08230_),
    .B(_07089_),
    .C(net2586),
    .Y(_14107_));
 OR4x1_ASAP7_75t_R _22881_ (.A(_14097_),
    .B(_12804_),
    .C(_10072_),
    .D(_14107_),
    .Y(_14118_));
 OA211x2_ASAP7_75t_R _22882_ (.A1(_08121_),
    .A2(net2055),
    .B(_08143_),
    .C(_08165_),
    .Y(_14128_));
 OA211x2_ASAP7_75t_R _22883_ (.A1(net1146),
    .A2(_05925_),
    .B(_09863_),
    .C(_06914_),
    .Y(_14139_));
 INVx1_ASAP7_75t_R _22884_ (.A(_14139_),
    .Y(_14149_));
 OA211x2_ASAP7_75t_R _22885_ (.A1(_08121_),
    .A2(_07111_),
    .B(_14149_),
    .C(_11148_),
    .Y(_14160_));
 NAND2x1_ASAP7_75t_R _22886_ (.A(_14128_),
    .B(_14160_),
    .Y(_14170_));
 NOR2x2_ASAP7_75t_R _22887_ (.A(_14118_),
    .B(_14170_),
    .Y(_14181_));
 NAND3x2_ASAP7_75t_R _22888_ (.B(_14076_),
    .C(_14181_),
    .Y(_14191_),
    .A(_14034_));
 AO21x1_ASAP7_75t_R _22889_ (.A1(net2055),
    .A2(net1047),
    .B(_08461_),
    .Y(_14202_));
 AO21x1_ASAP7_75t_R _22890_ (.A1(_06277_),
    .A2(_10478_),
    .B(_08461_),
    .Y(_14212_));
 OA211x2_ASAP7_75t_R _22891_ (.A1(_08461_),
    .A2(_07737_),
    .B(_14202_),
    .C(_14212_),
    .Y(_14222_));
 AO21x1_ASAP7_75t_R _22892_ (.A1(_10533_),
    .A2(_06925_),
    .B(_08461_),
    .Y(_14232_));
 OA211x2_ASAP7_75t_R _22893_ (.A1(_08461_),
    .A2(_07298_),
    .B(_14232_),
    .C(_11334_),
    .Y(_14243_));
 INVx1_ASAP7_75t_R _22894_ (.A(_12650_),
    .Y(_14253_));
 AO21x1_ASAP7_75t_R _22895_ (.A1(_06002_),
    .A2(_06925_),
    .B(_08406_),
    .Y(_14264_));
 AND5x2_ASAP7_75t_R _22896_ (.A(_09128_),
    .B(_14222_),
    .C(_14243_),
    .D(_14253_),
    .E(_14264_),
    .Y(_14274_));
 NAND2x1_ASAP7_75t_R _22897_ (.A(_06079_),
    .B(_08516_),
    .Y(_14285_));
 AND4x1_ASAP7_75t_R _22898_ (.A(_08975_),
    .B(_13581_),
    .C(_14285_),
    .D(_11444_),
    .Y(_14295_));
 NAND2x1_ASAP7_75t_R _22899_ (.A(_06266_),
    .B(_08570_),
    .Y(_14305_));
 AO21x1_ASAP7_75t_R _22900_ (.A1(_10533_),
    .A2(_12310_),
    .B(_08625_),
    .Y(_14316_));
 AO21x1_ASAP7_75t_R _22901_ (.A1(_07517_),
    .A2(_07298_),
    .B(_08625_),
    .Y(_14326_));
 AND4x1_ASAP7_75t_R _22902_ (.A(_13505_),
    .B(_14305_),
    .C(_14316_),
    .D(_14326_),
    .Y(_14337_));
 AND2x2_ASAP7_75t_R _22903_ (.A(_14295_),
    .B(_14337_),
    .Y(_14339_));
 OR4x1_ASAP7_75t_R _22904_ (.A(_10445_),
    .B(_06782_),
    .C(_11586_),
    .D(_13724_),
    .Y(_14340_));
 INVx1_ASAP7_75t_R _22905_ (.A(_14340_),
    .Y(_14341_));
 OA211x2_ASAP7_75t_R _22906_ (.A1(_06397_),
    .A2(_05925_),
    .B(_06815_),
    .C(_06727_),
    .Y(_14342_));
 INVx1_ASAP7_75t_R _22907_ (.A(_14342_),
    .Y(_14343_));
 AO21x1_ASAP7_75t_R _22908_ (.A1(net3403),
    .A2(net1047),
    .B(_06826_),
    .Y(_14344_));
 AND3x1_ASAP7_75t_R _22909_ (.A(_14341_),
    .B(_14343_),
    .C(_14344_),
    .Y(_14345_));
 AO21x1_ASAP7_75t_R _22910_ (.A1(_09052_),
    .A2(_06463_),
    .B(_11674_),
    .Y(_14346_));
 NOR2x1_ASAP7_75t_R _22911_ (.A(net3398),
    .B(_06474_),
    .Y(_14347_));
 OR4x1_ASAP7_75t_R _22912_ (.A(_14346_),
    .B(_06507_),
    .C(_09306_),
    .D(_14347_),
    .Y(_14348_));
 INVx1_ASAP7_75t_R _22913_ (.A(_14348_),
    .Y(_14349_));
 NOR2x1_ASAP7_75t_R _22914_ (.A(_05925_),
    .B(net1941),
    .Y(_14350_));
 AO221x1_ASAP7_75t_R _22915_ (.A1(_07100_),
    .A2(_06595_),
    .B1(_09369_),
    .B2(_09401_),
    .C(_09412_),
    .Y(_14351_));
 AOI211x1_ASAP7_75t_R _22916_ (.A1(_06595_),
    .A2(_14350_),
    .B(_14351_),
    .C(_06694_),
    .Y(_14352_));
 AND3x2_ASAP7_75t_R _22917_ (.A(_14345_),
    .B(_14349_),
    .C(_14352_),
    .Y(_14353_));
 NAND3x2_ASAP7_75t_R _22918_ (.B(_14339_),
    .C(_14353_),
    .Y(_14354_),
    .A(_14274_));
 NOR2x2_ASAP7_75t_R _22919_ (.A(_14191_),
    .B(_14354_),
    .Y(_14355_));
 INVx1_ASAP7_75t_R net399_46 (.A(clknet_leaf_4_clk),
    .Y(net451));
 XOR2x1_ASAP7_75t_R _22921_ (.A(_00411_),
    .Y(_14357_),
    .B(_00446_));
 INVx5_ASAP7_75t_R _22922_ (.A(_00478_),
    .Y(_14358_));
 XOR2x1_ASAP7_75t_R _22923_ (.A(_14357_),
    .Y(_14359_),
    .B(_14358_));
 CKINVDCx5p33_ASAP7_75t_R _22924_ (.A(_00497_),
    .Y(_14360_));
 XOR2x1_ASAP7_75t_R _22925_ (.A(_14359_),
    .Y(_14361_),
    .B(_14360_));
 AOI21x1_ASAP7_75t_R _22926_ (.A1(net2609),
    .A2(_14355_),
    .B(_14361_),
    .Y(_14362_));
 AND3x1_ASAP7_75t_R _22927_ (.A(_14355_),
    .B(net2609),
    .C(_14361_),
    .Y(_14363_));
 OAI21x1_ASAP7_75t_R _22928_ (.A1(_14362_),
    .A2(_14363_),
    .B(net399),
    .Y(_14364_));
 OAI21x1_ASAP7_75t_R _22929_ (.A1(net399),
    .A2(_13875_),
    .B(_14364_),
    .Y(_00381_));
 INVx1_ASAP7_75t_R _22930_ (.A(_12913_),
    .Y(_14375_));
 AO21x1_ASAP7_75t_R _22931_ (.A1(_06430_),
    .A2(_12310_),
    .B(_06771_),
    .Y(_14382_));
 AND5x1_ASAP7_75t_R _22932_ (.A(_07034_),
    .B(_14375_),
    .C(_09253_),
    .D(_10467_),
    .E(_14382_),
    .Y(_14388_));
 INVx1_ASAP7_75t_R _22933_ (.A(_14388_),
    .Y(_14395_));
 OR3x1_ASAP7_75t_R _22934_ (.A(_09359_),
    .B(_06573_),
    .C(_11674_),
    .Y(_14401_));
 NOR2x1_ASAP7_75t_R _22935_ (.A(_06925_),
    .B(_06474_),
    .Y(_14407_));
 OR3x1_ASAP7_75t_R _22936_ (.A(_14401_),
    .B(_10566_),
    .C(_14407_),
    .Y(_14414_));
 OA211x2_ASAP7_75t_R _22937_ (.A1(net1146),
    .A2(net2133),
    .B(_06815_),
    .C(_06914_),
    .Y(_14420_));
 OR4x1_ASAP7_75t_R _22938_ (.A(_14420_),
    .B(_06870_),
    .C(_09274_),
    .D(_13691_),
    .Y(_14427_));
 AND3x1_ASAP7_75t_R _22939_ (.A(_06595_),
    .B(net1146),
    .C(net2586),
    .Y(_14433_));
 OR5x1_ASAP7_75t_R _22940_ (.A(_06661_),
    .B(_14433_),
    .C(_11729_),
    .D(_09412_),
    .E(_09474_),
    .Y(_14440_));
 OR4x1_ASAP7_75t_R _22941_ (.A(_14395_),
    .B(_14414_),
    .C(_14427_),
    .D(_14440_),
    .Y(_14446_));
 AO21x1_ASAP7_75t_R _22942_ (.A1(_07342_),
    .A2(_06222_),
    .B(_08625_),
    .Y(_14453_));
 AO21x1_ASAP7_75t_R _22943_ (.A1(_07265_),
    .A2(_07298_),
    .B(_08406_),
    .Y(_14459_));
 AO21x1_ASAP7_75t_R _22944_ (.A1(_10533_),
    .A2(net3392),
    .B(_08406_),
    .Y(_14466_));
 AO21x1_ASAP7_75t_R _22945_ (.A1(net2055),
    .A2(_07737_),
    .B(_08406_),
    .Y(_14472_));
 AND4x1_ASAP7_75t_R _22946_ (.A(_11411_),
    .B(_14459_),
    .C(_14466_),
    .D(_14472_),
    .Y(_14478_));
 AO21x1_ASAP7_75t_R _22947_ (.A1(_07210_),
    .A2(net3403),
    .B(_08461_),
    .Y(_14485_));
 OA211x2_ASAP7_75t_R _22948_ (.A1(_07517_),
    .A2(_08461_),
    .B(_14485_),
    .C(_14232_),
    .Y(_14491_));
 AOI221x1_ASAP7_75t_R _22949_ (.A1(_06397_),
    .A2(_05925_),
    .B1(net1935),
    .B2(_06057_),
    .C(_08669_),
    .Y(_14498_));
 NOR2x1_ASAP7_75t_R _22950_ (.A(_13570_),
    .B(_14498_),
    .Y(_14504_));
 AO21x1_ASAP7_75t_R _22951_ (.A1(_12310_),
    .A2(_08614_),
    .B(_08625_),
    .Y(_14511_));
 AND5x1_ASAP7_75t_R _22952_ (.A(_14453_),
    .B(_14478_),
    .C(_14491_),
    .D(_14504_),
    .E(_14511_),
    .Y(_14517_));
 INVx1_ASAP7_75t_R _22953_ (.A(_14517_),
    .Y(_14524_));
 NOR2x1_ASAP7_75t_R _22954_ (.A(_14446_),
    .B(_14524_),
    .Y(_14530_));
 INVx2_ASAP7_75t_R _22955_ (.A(_14530_),
    .Y(_14536_));
 INVx1_ASAP7_75t_R _22956_ (.A(_09753_),
    .Y(_14542_));
 AO21x1_ASAP7_75t_R _22957_ (.A1(_07572_),
    .A2(_10478_),
    .B(_08011_),
    .Y(_14550_));
 AND5x1_ASAP7_75t_R _22958_ (.A(_14542_),
    .B(_14550_),
    .C(_10731_),
    .D(_13219_),
    .E(_09786_),
    .Y(_14558_));
 AO21x1_ASAP7_75t_R _22959_ (.A1(_07517_),
    .A2(_07298_),
    .B(_07879_),
    .Y(_14564_));
 AO21x1_ASAP7_75t_R _22960_ (.A1(_07210_),
    .A2(_10478_),
    .B(_07879_),
    .Y(_14569_));
 AO21x1_ASAP7_75t_R _22961_ (.A1(_10533_),
    .A2(net3392),
    .B(_07879_),
    .Y(_14571_));
 AND4x1_ASAP7_75t_R _22962_ (.A(_14564_),
    .B(_14569_),
    .C(_14571_),
    .D(_07945_),
    .Y(_14572_));
 NOR2x1_ASAP7_75t_R _22963_ (.A(_14107_),
    .B(_12902_),
    .Y(_14573_));
 AND4x1_ASAP7_75t_R _22964_ (.A(_11093_),
    .B(_08165_),
    .C(_09918_),
    .D(_12014_),
    .Y(_14574_));
 AOI21x1_ASAP7_75t_R _22965_ (.A1(_08230_),
    .A2(_08603_),
    .B(_10039_),
    .Y(_14575_));
 AND5x1_ASAP7_75t_R _22966_ (.A(_14558_),
    .B(_14572_),
    .C(_14573_),
    .D(_14574_),
    .E(_14575_),
    .Y(_14576_));
 AO21x1_ASAP7_75t_R _22967_ (.A1(_07111_),
    .A2(_07265_),
    .B(_05892_),
    .Y(_14577_));
 OA211x2_ASAP7_75t_R _22968_ (.A1(_05892_),
    .A2(_07342_),
    .B(_14577_),
    .C(_06156_),
    .Y(_14578_));
 AND3x1_ASAP7_75t_R _22969_ (.A(_13395_),
    .B(_07638_),
    .C(_09665_),
    .Y(_14579_));
 NAND2x1_ASAP7_75t_R _22970_ (.A(_07726_),
    .B(_05804_),
    .Y(_14580_));
 AND4x1_ASAP7_75t_R _22971_ (.A(_10983_),
    .B(_09676_),
    .C(_10994_),
    .D(_14580_),
    .Y(_14581_));
 AND3x1_ASAP7_75t_R _22972_ (.A(_14578_),
    .B(_14579_),
    .C(_14581_),
    .Y(_14582_));
 AND4x1_ASAP7_75t_R _22973_ (.A(_07440_),
    .B(_07462_),
    .C(_11937_),
    .D(_13939_),
    .Y(_14583_));
 NAND2x1_ASAP7_75t_R _22974_ (.A(_06211_),
    .B(_07781_),
    .Y(_14584_));
 AND5x1_ASAP7_75t_R _22975_ (.A(_11795_),
    .B(_09621_),
    .C(_14013_),
    .D(_09557_),
    .E(_14584_),
    .Y(_14585_));
 AND3x1_ASAP7_75t_R _22976_ (.A(_14582_),
    .B(_14583_),
    .C(_14585_),
    .Y(_14586_));
 AND2x2_ASAP7_75t_R _22977_ (.A(_14576_),
    .B(_14586_),
    .Y(_14587_));
 INVx2_ASAP7_75t_R _22978_ (.A(_14587_),
    .Y(_14588_));
 NOR2x2_ASAP7_75t_R _22979_ (.A(_14536_),
    .B(_14588_),
    .Y(_14589_));
 XNOR2x2_ASAP7_75t_R _22980_ (.A(_00477_),
    .B(_00520_),
    .Y(_14590_));
 INVx1_ASAP7_75t_R net399_45 (.A(clknet_leaf_7_clk),
    .Y(net450));
 XOR2x1_ASAP7_75t_R _22982_ (.A(_00388_),
    .Y(_14592_),
    .B(_00445_));
 XOR2x1_ASAP7_75t_R _22983_ (.A(_14590_),
    .Y(_14593_),
    .B(_14592_));
 XOR2x1_ASAP7_75t_R _22984_ (.A(_14589_),
    .Y(_14594_),
    .B(_14593_));
 AND2x2_ASAP7_75t_R _22985_ (.A(net404),
    .B(net106),
    .Y(_14595_));
 AO21x1_ASAP7_75t_R _22986_ (.A1(_14594_),
    .A2(net399),
    .B(_14595_),
    .Y(_00382_));
 INVx3_ASAP7_75t_R _22987_ (.A(net4074),
    .Y(_14596_));
 INVx1_ASAP7_75t_R net399_44 (.A(clknet_leaf_7_clk),
    .Y(net449));
 INVx1_ASAP7_75t_R net399_43 (.A(clknet_leaf_8_clk),
    .Y(net448));
 INVx1_ASAP7_75t_R net399_42 (.A(clknet_leaf_8_clk),
    .Y(net447));
 XOR2x1_ASAP7_75t_R _22991_ (.A(_00412_),
    .Y(_14600_),
    .B(net3552));
 INVx5_ASAP7_75t_R _22992_ (.A(_00476_),
    .Y(_14601_));
 XOR2x1_ASAP7_75t_R _22993_ (.A(_14600_),
    .Y(_14602_),
    .B(_14601_));
 INVx4_ASAP7_75t_R _22994_ (.A(_00496_),
    .Y(_14603_));
 XOR2x1_ASAP7_75t_R _22995_ (.A(_14602_),
    .Y(_14604_),
    .B(_14603_));
 NOR2x2_ASAP7_75t_R _22996_ (.A(_00449_),
    .B(net3526),
    .Y(_14605_));
 INVx5_ASAP7_75t_R _22997_ (.A(net1983),
    .Y(_14606_));
 NAND2x2_ASAP7_75t_R _22998_ (.A(_00445_),
    .B(_00446_),
    .Y(_14607_));
 NAND2x2_ASAP7_75t_R _22999_ (.A(_00447_),
    .B(_00448_),
    .Y(_14608_));
 NOR2x2_ASAP7_75t_R _23000_ (.A(_14607_),
    .B(_14608_),
    .Y(_14609_));
 INVx6_ASAP7_75t_R _23001_ (.A(_14609_),
    .Y(_14610_));
 NOR2x1_ASAP7_75t_R _23002_ (.A(_14606_),
    .B(_14610_),
    .Y(_14611_));
 INVx1_ASAP7_75t_R _23003_ (.A(_14611_),
    .Y(_14612_));
 INVx2_ASAP7_75t_R _23004_ (.A(net3529),
    .Y(_14613_));
 NOR2x2_ASAP7_75t_R _23005_ (.A(_00449_),
    .B(_14613_),
    .Y(_14614_));
 NAND2x2_ASAP7_75t_R _23006_ (.A(net2199),
    .B(net3516),
    .Y(_14615_));
 INVx1_ASAP7_75t_R _23007_ (.A(_14615_),
    .Y(_14616_));
 NAND2x2_ASAP7_75t_R _23008_ (.A(_14614_),
    .B(_14616_),
    .Y(_14617_));
 INVx3_ASAP7_75t_R _23009_ (.A(_14617_),
    .Y(_14618_));
 NAND2x1_ASAP7_75t_R _23010_ (.A(_14609_),
    .B(_14618_),
    .Y(_14619_));
 INVx13_ASAP7_75t_R _23011_ (.A(net2197),
    .Y(_14620_));
 NOR2x2_ASAP7_75t_R _23012_ (.A(net3513),
    .B(_14620_),
    .Y(_14621_));
 NAND2x2_ASAP7_75t_R _23013_ (.A(_14614_),
    .B(_14621_),
    .Y(_14622_));
 INVx2_ASAP7_75t_R _23014_ (.A(_14622_),
    .Y(_14623_));
 NAND2x1_ASAP7_75t_R _23015_ (.A(_14609_),
    .B(_14623_),
    .Y(_14624_));
 NAND2x2_ASAP7_75t_R _23016_ (.A(_14620_),
    .B(_14614_),
    .Y(_14625_));
 INVx2_ASAP7_75t_R _23017_ (.A(_14625_),
    .Y(_14626_));
 NAND2x1_ASAP7_75t_R _23018_ (.A(_14609_),
    .B(_14626_),
    .Y(_14627_));
 AND4x1_ASAP7_75t_R _23019_ (.A(_14612_),
    .B(_14619_),
    .C(_14624_),
    .D(_14627_),
    .Y(_14628_));
 INVx4_ASAP7_75t_R _23020_ (.A(_00449_),
    .Y(_14629_));
 NOR2x2_ASAP7_75t_R _23021_ (.A(net3526),
    .B(_14629_),
    .Y(_14630_));
 INVx6_ASAP7_75t_R _23022_ (.A(_14630_),
    .Y(_14631_));
 INVx1_ASAP7_75t_R net399_41 (.A(clknet_leaf_6_clk),
    .Y(net446));
 NAND2x2_ASAP7_75t_R _23024_ (.A(net3532),
    .B(net3526),
    .Y(_14633_));
 INVx2_ASAP7_75t_R _23025_ (.A(_14621_),
    .Y(_14634_));
 NOR2x2_ASAP7_75t_R _23026_ (.A(_14633_),
    .B(_14634_),
    .Y(_14635_));
 CKINVDCx8_ASAP7_75t_R _23027_ (.A(_14635_),
    .Y(_14636_));
 INVx8_ASAP7_75t_R _23028_ (.A(_14633_),
    .Y(_14637_));
 NAND2x2_ASAP7_75t_R _23029_ (.A(_14620_),
    .B(_14637_),
    .Y(_14638_));
 AO21x1_ASAP7_75t_R _23030_ (.A1(_14636_),
    .A2(_14638_),
    .B(_14610_),
    .Y(_14639_));
 OA21x2_ASAP7_75t_R _23031_ (.A1(_14631_),
    .A2(_14610_),
    .B(_14639_),
    .Y(_14640_));
 AND2x2_ASAP7_75t_R _23032_ (.A(_14628_),
    .B(_14640_),
    .Y(_14641_));
 AND5x2_ASAP7_75t_R _23033_ (.A(_00445_),
    .B(_14641_),
    .C(_00446_),
    .D(_00447_),
    .E(_00448_),
    .Y(_14642_));
 INVx3_ASAP7_75t_R _23034_ (.A(_00447_),
    .Y(_14643_));
 NAND2x2_ASAP7_75t_R _23035_ (.A(_00448_),
    .B(_14643_),
    .Y(_14644_));
 INVx2_ASAP7_75t_R _23036_ (.A(_00445_),
    .Y(_14645_));
 NAND2x2_ASAP7_75t_R _23037_ (.A(_00446_),
    .B(_14645_),
    .Y(_14646_));
 NOR2x2_ASAP7_75t_R _23038_ (.A(_14644_),
    .B(_14646_),
    .Y(_14647_));
 NOR2x2_ASAP7_75t_R _23039_ (.A(net1769),
    .B(_14631_),
    .Y(_14648_));
 NAND2x1_ASAP7_75t_R _23040_ (.A(_14647_),
    .B(_14648_),
    .Y(_14649_));
 NAND2x2_ASAP7_75t_R _23041_ (.A(net3516),
    .B(_14620_),
    .Y(_14650_));
 NOR2x2_ASAP7_75t_R _23042_ (.A(_14633_),
    .B(_14650_),
    .Y(_14651_));
 INVx8_ASAP7_75t_R _23043_ (.A(_14651_),
    .Y(_14652_));
 NOR2x2_ASAP7_75t_R _23044_ (.A(net1770),
    .B(net3505),
    .Y(_14653_));
 CKINVDCx11_ASAP7_75t_R _23045_ (.A(_14653_),
    .Y(_14654_));
 NOR2x2_ASAP7_75t_R _23046_ (.A(_00447_),
    .B(_00448_),
    .Y(_14655_));
 INVx1_ASAP7_75t_R _23047_ (.A(_14646_),
    .Y(_14656_));
 NAND2x2_ASAP7_75t_R _23048_ (.A(_14655_),
    .B(_14656_),
    .Y(_14657_));
 AO21x1_ASAP7_75t_R _23049_ (.A1(_14652_),
    .A2(_14654_),
    .B(_14657_),
    .Y(_14658_));
 NOR2x2_ASAP7_75t_R _23050_ (.A(net2199),
    .B(net3515),
    .Y(_14659_));
 NAND2x2_ASAP7_75t_R _23051_ (.A(_14659_),
    .B(_14637_),
    .Y(_14660_));
 INVx4_ASAP7_75t_R _23052_ (.A(_14660_),
    .Y(_14661_));
 INVx4_ASAP7_75t_R _23053_ (.A(_14657_),
    .Y(_14662_));
 NAND2x1_ASAP7_75t_R _23054_ (.A(_14661_),
    .B(_14662_),
    .Y(_14663_));
 AND2x2_ASAP7_75t_R _23055_ (.A(_14658_),
    .B(_14663_),
    .Y(_14664_));
 INVx1_ASAP7_75t_R net399_40 (.A(clknet_leaf_11_clk),
    .Y(net445));
 INVx1_ASAP7_75t_R net399_39 (.A(clknet_leaf_11_clk),
    .Y(net444));
 NAND2x2_ASAP7_75t_R _23058_ (.A(net1985),
    .B(_14650_),
    .Y(_14667_));
 INVx3_ASAP7_75t_R _23059_ (.A(_14647_),
    .Y(_14668_));
 AO21x1_ASAP7_75t_R _23060_ (.A1(net1819),
    .A2(_14667_),
    .B(_14668_),
    .Y(_14669_));
 NOR2x2_ASAP7_75t_R _23061_ (.A(_14615_),
    .B(_14606_),
    .Y(_14670_));
 NAND2x1_ASAP7_75t_R _23062_ (.A(_14670_),
    .B(_14662_),
    .Y(_14671_));
 CKINVDCx10_ASAP7_75t_R _23063_ (.A(net3513),
    .Y(_14672_));
 NOR2x2_ASAP7_75t_R _23064_ (.A(net2200),
    .B(_14672_),
    .Y(_14673_));
 NOR2x2_ASAP7_75t_R _23065_ (.A(_14673_),
    .B(_14631_),
    .Y(_14674_));
 NAND2x1_ASAP7_75t_R _23066_ (.A(_14674_),
    .B(_14662_),
    .Y(_14675_));
 AND5x1_ASAP7_75t_R _23067_ (.A(_14649_),
    .B(_14664_),
    .C(_14669_),
    .D(_14671_),
    .E(_14675_),
    .Y(_14676_));
 INVx1_ASAP7_75t_R net399_38 (.A(clknet_leaf_11_clk),
    .Y(net443));
 NOR2x2_ASAP7_75t_R _23069_ (.A(_14608_),
    .B(_14646_),
    .Y(_14678_));
 INVx1_ASAP7_75t_R net399_37 (.A(clknet_leaf_6_clk),
    .Y(net442));
 OA211x2_ASAP7_75t_R _23071_ (.A1(net2201),
    .A2(_14672_),
    .B(_14678_),
    .C(net2721),
    .Y(_14680_));
 INVx1_ASAP7_75t_R _23072_ (.A(_14680_),
    .Y(_14681_));
 INVx3_ASAP7_75t_R _23073_ (.A(_00448_),
    .Y(_14682_));
 NAND2x2_ASAP7_75t_R _23074_ (.A(_00447_),
    .B(_14682_),
    .Y(_14683_));
 NOR2x2_ASAP7_75t_R _23075_ (.A(_14646_),
    .B(_14683_),
    .Y(_14684_));
 NAND2x1_ASAP7_75t_R _23076_ (.A(net1987),
    .B(_14684_),
    .Y(_14685_));
 INVx4_ASAP7_75t_R _23077_ (.A(_14684_),
    .Y(_14686_));
 INVx1_ASAP7_75t_R net399_36 (.A(clknet_leaf_6_clk),
    .Y(net441));
 AO21x1_ASAP7_75t_R _23079_ (.A1(_14636_),
    .A2(_14652_),
    .B(_14686_),
    .Y(_14688_));
 OA21x2_ASAP7_75t_R _23080_ (.A1(net2201),
    .A2(_14685_),
    .B(_14688_),
    .Y(_14689_));
 AND3x1_ASAP7_75t_R _23081_ (.A(_14678_),
    .B(net1988),
    .C(_14615_),
    .Y(_14690_));
 INVx1_ASAP7_75t_R _23082_ (.A(_14690_),
    .Y(_14691_));
 NAND2x2_ASAP7_75t_R _23083_ (.A(_14659_),
    .B(_14614_),
    .Y(_14692_));
 INVx1_ASAP7_75t_R net399_35 (.A(clknet_leaf_1_clk),
    .Y(net440));
 INVx6_ASAP7_75t_R _23085_ (.A(_14678_),
    .Y(_14694_));
 INVx1_ASAP7_75t_R net399_34 (.A(clknet_leaf_15_clk),
    .Y(net439));
 AO21x1_ASAP7_75t_R _23087_ (.A1(net1820),
    .A2(net3510),
    .B(_14694_),
    .Y(_14696_));
 INVx1_ASAP7_75t_R net399_33 (.A(clknet_leaf_7_clk),
    .Y(net438));
 INVx1_ASAP7_75t_R net399_32 (.A(clknet_leaf_15_clk),
    .Y(net437));
 AO21x1_ASAP7_75t_R _23090_ (.A1(_14652_),
    .A2(_14654_),
    .B(_14694_),
    .Y(_14699_));
 AND5x1_ASAP7_75t_R _23091_ (.A(_14681_),
    .B(_14689_),
    .C(_14691_),
    .D(_14696_),
    .E(_14699_),
    .Y(_14700_));
 NAND2x1_ASAP7_75t_R _23092_ (.A(_14676_),
    .B(_14700_),
    .Y(_14701_));
 NOR2x2_ASAP7_75t_R _23093_ (.A(_00445_),
    .B(_00446_),
    .Y(_14702_));
 INVx4_ASAP7_75t_R _23094_ (.A(_14702_),
    .Y(_14703_));
 NOR2x2_ASAP7_75t_R _23095_ (.A(_14644_),
    .B(_14703_),
    .Y(_14704_));
 AND3x1_ASAP7_75t_R _23096_ (.A(_14704_),
    .B(_00451_),
    .C(_14630_),
    .Y(_14705_));
 INVx1_ASAP7_75t_R _23097_ (.A(_14705_),
    .Y(_14706_));
 INVx1_ASAP7_75t_R net399_31 (.A(clknet_leaf_14_clk),
    .Y(net436));
 AND3x1_ASAP7_75t_R _23099_ (.A(_14704_),
    .B(_14614_),
    .C(_14634_),
    .Y(_14708_));
 INVx1_ASAP7_75t_R _23100_ (.A(_14708_),
    .Y(_14709_));
 INVx1_ASAP7_75t_R net399_30 (.A(clknet_leaf_14_clk),
    .Y(net435));
 INVx1_ASAP7_75t_R net399_29 (.A(clknet_leaf_2_clk),
    .Y(net434));
 INVx4_ASAP7_75t_R _23103_ (.A(_14704_),
    .Y(_14712_));
 INVx1_ASAP7_75t_R net399_28 (.A(clknet_leaf_1_clk),
    .Y(net433));
 AO21x1_ASAP7_75t_R _23105_ (.A1(_14654_),
    .A2(net3522),
    .B(_14712_),
    .Y(_14714_));
 NAND2x2_ASAP7_75t_R _23106_ (.A(_14659_),
    .B(net1983),
    .Y(_14715_));
 NAND2x2_ASAP7_75t_R _23107_ (.A(_14605_),
    .B(_14621_),
    .Y(_14716_));
 INVx1_ASAP7_75t_R net399_27 (.A(clknet_leaf_15_clk),
    .Y(net432));
 AO21x1_ASAP7_75t_R _23109_ (.A1(net1873),
    .A2(_14716_),
    .B(_14712_),
    .Y(_14718_));
 AND4x1_ASAP7_75t_R _23110_ (.A(_14706_),
    .B(_14709_),
    .C(_14714_),
    .D(_14718_),
    .Y(_14719_));
 NOR2x2_ASAP7_75t_R _23111_ (.A(_14608_),
    .B(_14703_),
    .Y(_14720_));
 OA211x2_ASAP7_75t_R _23112_ (.A1(net2197),
    .A2(net3513),
    .B(_14720_),
    .C(net1989),
    .Y(_14721_));
 INVx1_ASAP7_75t_R _23113_ (.A(_14721_),
    .Y(_14722_));
 INVx1_ASAP7_75t_R net399_26 (.A(clknet_leaf_1_clk),
    .Y(net431));
 NAND2x1_ASAP7_75t_R _23115_ (.A(_14651_),
    .B(_14720_),
    .Y(_14724_));
 INVx4_ASAP7_75t_R _23116_ (.A(_14720_),
    .Y(_14725_));
 AO21x1_ASAP7_75t_R _23117_ (.A1(net1818),
    .A2(_14692_),
    .B(_14725_),
    .Y(_14726_));
 AND3x1_ASAP7_75t_R _23118_ (.A(_14722_),
    .B(_14724_),
    .C(_14726_),
    .Y(_14727_));
 NAND2x2_ASAP7_75t_R _23119_ (.A(net3528),
    .B(_14629_),
    .Y(_14728_));
 NOR2x2_ASAP7_75t_R _23120_ (.A(_14683_),
    .B(_14703_),
    .Y(_14729_));
 CKINVDCx6p67_ASAP7_75t_R _23121_ (.A(_14729_),
    .Y(_14730_));
 INVx1_ASAP7_75t_R net399_25 (.A(clknet_leaf_0_clk),
    .Y(net430));
 NOR2x2_ASAP7_75t_R _23123_ (.A(_14650_),
    .B(_14606_),
    .Y(_14732_));
 CKINVDCx11_ASAP7_75t_R _23124_ (.A(_14732_),
    .Y(_14733_));
 AO21x1_ASAP7_75t_R _23125_ (.A1(_14733_),
    .A2(_14716_),
    .B(_14730_),
    .Y(_14734_));
 NAND2x2_ASAP7_75t_R _23126_ (.A(_14630_),
    .B(_14621_),
    .Y(_14735_));
 INVx1_ASAP7_75t_R net399_24 (.A(clknet_leaf_1_clk),
    .Y(net429));
 AO21x1_ASAP7_75t_R _23128_ (.A1(net1830),
    .A2(_14652_),
    .B(_14730_),
    .Y(_14737_));
 OA211x2_ASAP7_75t_R _23129_ (.A1(_14728_),
    .A2(_14730_),
    .B(_14734_),
    .C(_14737_),
    .Y(_14738_));
 AND2x6_ASAP7_75t_R _23130_ (.A(_14702_),
    .B(_14655_),
    .Y(_14739_));
 INVx6_ASAP7_75t_R _23131_ (.A(_14739_),
    .Y(_14740_));
 AO21x1_ASAP7_75t_R _23132_ (.A1(net3521),
    .A2(_14652_),
    .B(_14740_),
    .Y(_14741_));
 INVx1_ASAP7_75t_R _23133_ (.A(_14741_),
    .Y(_14742_));
 INVx1_ASAP7_75t_R net399_23 (.A(clknet_leaf_1_clk),
    .Y(net428));
 CKINVDCx6p67_ASAP7_75t_R _23135_ (.A(_14648_),
    .Y(_14744_));
 NOR2x1_ASAP7_75t_R _23136_ (.A(_14740_),
    .B(_14744_),
    .Y(_14745_));
 NOR2x1_ASAP7_75t_R _23137_ (.A(_14740_),
    .B(_14636_),
    .Y(_14746_));
 OR3x1_ASAP7_75t_R _23138_ (.A(_14742_),
    .B(_14745_),
    .C(_14746_),
    .Y(_14747_));
 NOR2x2_ASAP7_75t_R _23139_ (.A(net1818),
    .B(_14740_),
    .Y(_14748_));
 AO21x1_ASAP7_75t_R _23140_ (.A1(_14618_),
    .A2(_14739_),
    .B(_14748_),
    .Y(_14749_));
 AND2x2_ASAP7_75t_R _23141_ (.A(_14739_),
    .B(_14732_),
    .Y(_14750_));
 NOR2x1_ASAP7_75t_R _23142_ (.A(net3506),
    .B(_14740_),
    .Y(_14751_));
 OR3x1_ASAP7_75t_R _23143_ (.A(_14749_),
    .B(_14750_),
    .C(_14751_),
    .Y(_14752_));
 NOR2x1_ASAP7_75t_R _23144_ (.A(_14747_),
    .B(_14752_),
    .Y(_14753_));
 AND4x1_ASAP7_75t_R _23145_ (.A(_14719_),
    .B(_14727_),
    .C(_14738_),
    .D(_14753_),
    .Y(_14754_));
 INVx1_ASAP7_75t_R _23146_ (.A(_14754_),
    .Y(_14755_));
 NOR2x1_ASAP7_75t_R _23147_ (.A(_14701_),
    .B(_14755_),
    .Y(_14756_));
 NAND2x2_ASAP7_75t_R _23148_ (.A(_14650_),
    .B(_14637_),
    .Y(_14757_));
 INVx4_ASAP7_75t_R _23149_ (.A(_00446_),
    .Y(_14758_));
 NAND2x2_ASAP7_75t_R _23150_ (.A(_00445_),
    .B(_14758_),
    .Y(_14759_));
 OR3x1_ASAP7_75t_R _23151_ (.A(_14757_),
    .B(_14683_),
    .C(_14759_),
    .Y(_14760_));
 NOR2x2_ASAP7_75t_R _23152_ (.A(_14683_),
    .B(_14759_),
    .Y(_14761_));
 INVx3_ASAP7_75t_R _23153_ (.A(_14715_),
    .Y(_14762_));
 NAND2x1_ASAP7_75t_R _23154_ (.A(_14761_),
    .B(_14762_),
    .Y(_14763_));
 NAND2x2_ASAP7_75t_R _23155_ (.A(_14659_),
    .B(_14630_),
    .Y(_14764_));
 INVx1_ASAP7_75t_R net399_22 (.A(clknet_leaf_1_clk),
    .Y(net427));
 NAND2x2_ASAP7_75t_R _23157_ (.A(_14673_),
    .B(_14630_),
    .Y(_14766_));
 INVx1_ASAP7_75t_R net399_21 (.A(clknet_leaf_2_clk),
    .Y(net426));
 CKINVDCx5p33_ASAP7_75t_R _23159_ (.A(_14761_),
    .Y(_14768_));
 AO21x1_ASAP7_75t_R _23160_ (.A1(_14764_),
    .A2(net3535),
    .B(_14768_),
    .Y(_14769_));
 AO21x1_ASAP7_75t_R _23161_ (.A1(net3510),
    .A2(net3524),
    .B(_14768_),
    .Y(_14770_));
 AND4x1_ASAP7_75t_R _23162_ (.A(_14760_),
    .B(_14763_),
    .C(_14769_),
    .D(_14770_),
    .Y(_14771_));
 INVx1_ASAP7_75t_R net399_20 (.A(clknet_leaf_4_clk),
    .Y(net425));
 AO21x1_ASAP7_75t_R _23164_ (.A1(_14620_),
    .A2(_14672_),
    .B(_14606_),
    .Y(_14773_));
 NAND2x2_ASAP7_75t_R _23165_ (.A(_14672_),
    .B(net3525),
    .Y(_14774_));
 NOR2x2_ASAP7_75t_R _23166_ (.A(_14608_),
    .B(_14759_),
    .Y(_14775_));
 CKINVDCx5p33_ASAP7_75t_R _23167_ (.A(_14775_),
    .Y(_14776_));
 INVx1_ASAP7_75t_R net399_19 (.A(clknet_leaf_7_clk),
    .Y(net424));
 AO21x1_ASAP7_75t_R _23169_ (.A1(_14773_),
    .A2(_14774_),
    .B(_14776_),
    .Y(_14778_));
 NAND2x1_ASAP7_75t_R _23170_ (.A(_14775_),
    .B(_14648_),
    .Y(_14779_));
 AO21x1_ASAP7_75t_R _23171_ (.A1(_14636_),
    .A2(_14654_),
    .B(_14776_),
    .Y(_14780_));
 AND3x1_ASAP7_75t_R _23172_ (.A(_14778_),
    .B(_14779_),
    .C(_14780_),
    .Y(_14781_));
 NOR2x2_ASAP7_75t_R _23173_ (.A(_14644_),
    .B(_14759_),
    .Y(_14782_));
 CKINVDCx5p33_ASAP7_75t_R _23174_ (.A(_14782_),
    .Y(_14783_));
 NOR2x1_ASAP7_75t_R _23175_ (.A(_14633_),
    .B(_14783_),
    .Y(_14784_));
 INVx1_ASAP7_75t_R net399_18 (.A(clknet_leaf_6_clk),
    .Y(net423));
 AOI22x1_ASAP7_75t_R _23177_ (.A1(_14784_),
    .A2(_14672_),
    .B1(net2722),
    .B2(_14782_),
    .Y(_14786_));
 AND2x2_ASAP7_75t_R _23178_ (.A(_14732_),
    .B(_14782_),
    .Y(_14787_));
 INVx1_ASAP7_75t_R _23179_ (.A(_14787_),
    .Y(_14788_));
 AO21x1_ASAP7_75t_R _23180_ (.A1(net3518),
    .A2(_14774_),
    .B(_14783_),
    .Y(_14789_));
 AND3x1_ASAP7_75t_R _23181_ (.A(_14786_),
    .B(_14788_),
    .C(_14789_),
    .Y(_14790_));
 NOR2x1_ASAP7_75t_R _23182_ (.A(_00446_),
    .B(_14645_),
    .Y(_14791_));
 AND2x6_ASAP7_75t_R _23183_ (.A(_14791_),
    .B(_14655_),
    .Y(_14792_));
 INVx5_ASAP7_75t_R _23184_ (.A(_14792_),
    .Y(_14793_));
 INVx1_ASAP7_75t_R net399_17 (.A(clknet_leaf_6_clk),
    .Y(net422));
 AO21x1_ASAP7_75t_R _23186_ (.A1(net3539),
    .A2(_14764_),
    .B(_14793_),
    .Y(_14795_));
 OA21x2_ASAP7_75t_R _23187_ (.A1(_14757_),
    .A2(_14793_),
    .B(_14795_),
    .Y(_14796_));
 INVx4_ASAP7_75t_R _23188_ (.A(_14692_),
    .Y(_14797_));
 INVx1_ASAP7_75t_R net399_16 (.A(clknet_leaf_11_clk),
    .Y(net421));
 NAND2x1_ASAP7_75t_R _23190_ (.A(_14797_),
    .B(_14792_),
    .Y(_14799_));
 AO21x1_ASAP7_75t_R _23191_ (.A1(_14733_),
    .A2(_14716_),
    .B(_14793_),
    .Y(_14800_));
 AND3x1_ASAP7_75t_R _23192_ (.A(_14796_),
    .B(_14799_),
    .C(_14800_),
    .Y(_14801_));
 AND4x1_ASAP7_75t_R _23193_ (.A(_14771_),
    .B(_14781_),
    .C(_14790_),
    .D(_14801_),
    .Y(_14802_));
 INVx1_ASAP7_75t_R _23194_ (.A(_14802_),
    .Y(_14803_));
 CKINVDCx8_ASAP7_75t_R _23195_ (.A(_14670_),
    .Y(_14804_));
 NAND2x2_ASAP7_75t_R _23196_ (.A(_14620_),
    .B(net1984),
    .Y(_14805_));
 NOR2x2_ASAP7_75t_R _23197_ (.A(_14607_),
    .B(_14644_),
    .Y(_14806_));
 CKINVDCx5p33_ASAP7_75t_R _23198_ (.A(_14806_),
    .Y(_14807_));
 AO21x1_ASAP7_75t_R _23199_ (.A1(_14804_),
    .A2(_14805_),
    .B(_14807_),
    .Y(_14808_));
 NAND2x2_ASAP7_75t_R _23200_ (.A(net2199),
    .B(_14637_),
    .Y(_14809_));
 AO21x1_ASAP7_75t_R _23201_ (.A1(_14652_),
    .A2(_14809_),
    .B(_14807_),
    .Y(_14810_));
 AO21x1_ASAP7_75t_R _23202_ (.A1(net1817),
    .A2(_14625_),
    .B(_14807_),
    .Y(_14811_));
 AO21x1_ASAP7_75t_R _23203_ (.A1(net3539),
    .A2(net3537),
    .B(_14807_),
    .Y(_14812_));
 AND4x1_ASAP7_75t_R _23204_ (.A(_14808_),
    .B(_14810_),
    .C(_14811_),
    .D(_14812_),
    .Y(_14813_));
 NAND2x2_ASAP7_75t_R _23205_ (.A(_14672_),
    .B(_14637_),
    .Y(_14814_));
 AND3x4_ASAP7_75t_R _23206_ (.A(_14655_),
    .B(_00445_),
    .C(_00446_),
    .Y(_14815_));
 CKINVDCx6p67_ASAP7_75t_R _23207_ (.A(_14815_),
    .Y(_14816_));
 INVx1_ASAP7_75t_R net399_15 (.A(clknet_leaf_11_clk),
    .Y(net420));
 AO21x1_ASAP7_75t_R _23209_ (.A1(_14652_),
    .A2(_14814_),
    .B(_14816_),
    .Y(_14818_));
 INVx4_ASAP7_75t_R _23210_ (.A(_14766_),
    .Y(_14819_));
 NAND2x1_ASAP7_75t_R _23211_ (.A(_14819_),
    .B(_14815_),
    .Y(_14820_));
 AO21x1_ASAP7_75t_R _23212_ (.A1(_14804_),
    .A2(_14716_),
    .B(_14816_),
    .Y(_14821_));
 NOR2x1_ASAP7_75t_R _23213_ (.A(_14715_),
    .B(_14816_),
    .Y(_14822_));
 INVx1_ASAP7_75t_R _23214_ (.A(_14822_),
    .Y(_14823_));
 NAND2x1_ASAP7_75t_R _23215_ (.A(_14618_),
    .B(_14815_),
    .Y(_14824_));
 AND3x1_ASAP7_75t_R _23216_ (.A(_14821_),
    .B(_14823_),
    .C(_14824_),
    .Y(_14825_));
 AND4x1_ASAP7_75t_R _23217_ (.A(_14813_),
    .B(_14818_),
    .C(_14820_),
    .D(_14825_),
    .Y(_14826_));
 AO21x1_ASAP7_75t_R _23218_ (.A1(net3537),
    .A2(_14764_),
    .B(_14610_),
    .Y(_14827_));
 NOR2x1_ASAP7_75t_R _23219_ (.A(_14638_),
    .B(_14610_),
    .Y(_14828_));
 INVx1_ASAP7_75t_R _23220_ (.A(_14828_),
    .Y(_14829_));
 OA211x2_ASAP7_75t_R _23221_ (.A1(net3539),
    .A2(_14610_),
    .B(_14827_),
    .C(_14829_),
    .Y(_14830_));
 INVx1_ASAP7_75t_R net399_14 (.A(clknet_leaf_5_clk),
    .Y(net419));
 INVx1_ASAP7_75t_R net399_13 (.A(clknet_leaf_7_clk),
    .Y(net418));
 AO21x1_ASAP7_75t_R _23224_ (.A1(_14733_),
    .A2(net2179),
    .B(_14610_),
    .Y(_14833_));
 NOR2x2_ASAP7_75t_R _23225_ (.A(_14607_),
    .B(_14683_),
    .Y(_14834_));
 CKINVDCx6p67_ASAP7_75t_R _23226_ (.A(_14834_),
    .Y(_14835_));
 AO21x1_ASAP7_75t_R _23227_ (.A1(_14652_),
    .A2(_14660_),
    .B(_14835_),
    .Y(_14836_));
 AO21x1_ASAP7_75t_R _23228_ (.A1(_14692_),
    .A2(net3518),
    .B(_14835_),
    .Y(_14837_));
 AO21x1_ASAP7_75t_R _23229_ (.A1(net3539),
    .A2(_14766_),
    .B(_14835_),
    .Y(_14838_));
 AND3x1_ASAP7_75t_R _23230_ (.A(_14836_),
    .B(_14837_),
    .C(_14838_),
    .Y(_14839_));
 AND5x1_ASAP7_75t_R _23231_ (.A(_14627_),
    .B(_14830_),
    .C(_14624_),
    .D(_14833_),
    .E(_14839_),
    .Y(_14840_));
 NAND2x1_ASAP7_75t_R _23232_ (.A(_14826_),
    .B(_14840_),
    .Y(_14841_));
 NOR2x1_ASAP7_75t_R _23233_ (.A(_14803_),
    .B(_14841_),
    .Y(_14842_));
 NAND2x1_ASAP7_75t_R _23234_ (.A(_14756_),
    .B(_14842_),
    .Y(_14843_));
 NOR2x2_ASAP7_75t_R _23235_ (.A(_14642_),
    .B(_14843_),
    .Y(_14844_));
 NOR2x1_ASAP7_75t_R _23236_ (.A(_14604_),
    .B(_14844_),
    .Y(_14845_));
 AND2x2_ASAP7_75t_R _23237_ (.A(_14844_),
    .B(_14604_),
    .Y(_14846_));
 OAI21x1_ASAP7_75t_R _23238_ (.A1(_14845_),
    .A2(_14846_),
    .B(net399),
    .Y(_14847_));
 OAI21x1_ASAP7_75t_R _23239_ (.A1(net399),
    .A2(_14596_),
    .B(_14847_),
    .Y(_00383_));
 INVx1_ASAP7_75t_R net399_12 (.A(clknet_leaf_2_clk),
    .Y(net417));
 INVx1_ASAP7_75t_R net399_11 (.A(clknet_leaf_4_clk),
    .Y(net416));
 AO21x1_ASAP7_75t_R _23242_ (.A1(_14733_),
    .A2(_14625_),
    .B(_14835_),
    .Y(_14850_));
 INVx1_ASAP7_75t_R net399_10 (.A(clknet_leaf_6_clk),
    .Y(net415));
 AO21x1_ASAP7_75t_R _23244_ (.A1(_14744_),
    .A2(net3536),
    .B(_14835_),
    .Y(_14852_));
 OR3x1_ASAP7_75t_R _23245_ (.A(_14809_),
    .B(_14683_),
    .C(_14607_),
    .Y(_14853_));
 AND3x1_ASAP7_75t_R _23246_ (.A(_14850_),
    .B(_14852_),
    .C(_14853_),
    .Y(_14854_));
 OR3x1_ASAP7_75t_R _23247_ (.A(_14610_),
    .B(_14659_),
    .C(_14631_),
    .Y(_14855_));
 AND5x1_ASAP7_75t_R _23248_ (.A(_14612_),
    .B(_14854_),
    .C(_14829_),
    .D(_14627_),
    .E(_14855_),
    .Y(_14856_));
 OR3x1_ASAP7_75t_R _23249_ (.A(_14807_),
    .B(_14659_),
    .C(_14631_),
    .Y(_14857_));
 INVx1_ASAP7_75t_R net399_9 (.A(clknet_leaf_6_clk),
    .Y(net414));
 AO21x1_ASAP7_75t_R _23251_ (.A1(net1817),
    .A2(net3519),
    .B(_14816_),
    .Y(_14859_));
 NAND2x2_ASAP7_75t_R _23252_ (.A(net2200),
    .B(net1985),
    .Y(_14860_));
 AO21x1_ASAP7_75t_R _23253_ (.A1(_14733_),
    .A2(_14860_),
    .B(_14816_),
    .Y(_14861_));
 NAND2x1_ASAP7_75t_R _23254_ (.A(_14797_),
    .B(_14815_),
    .Y(_14862_));
 AND3x1_ASAP7_75t_R _23255_ (.A(_14859_),
    .B(_14861_),
    .C(_14862_),
    .Y(_14863_));
 INVx1_ASAP7_75t_R net399_8 (.A(clknet_leaf_1_clk),
    .Y(net413));
 AO21x1_ASAP7_75t_R _23257_ (.A1(_14764_),
    .A2(net3539),
    .B(_14816_),
    .Y(_14865_));
 INVx1_ASAP7_75t_R net399_7 (.A(clknet_leaf_7_clk),
    .Y(net412));
 AO21x1_ASAP7_75t_R _23259_ (.A1(_14654_),
    .A2(_14638_),
    .B(_14807_),
    .Y(_14867_));
 AND5x1_ASAP7_75t_R _23260_ (.A(_14857_),
    .B(_14863_),
    .C(_14818_),
    .D(_14865_),
    .E(_14867_),
    .Y(_14868_));
 NAND2x1_ASAP7_75t_R _23261_ (.A(_14856_),
    .B(_14868_),
    .Y(_14869_));
 NOR2x2_ASAP7_75t_R _23262_ (.A(_14728_),
    .B(_14650_),
    .Y(_14870_));
 AND2x2_ASAP7_75t_R _23263_ (.A(_14870_),
    .B(_14761_),
    .Y(_14871_));
 INVx1_ASAP7_75t_R _23264_ (.A(_14763_),
    .Y(_14872_));
 AO21x1_ASAP7_75t_R _23265_ (.A1(_14761_),
    .A2(_14670_),
    .B(_14872_),
    .Y(_14873_));
 INVx1_ASAP7_75t_R net399_6 (.A(clknet_leaf_11_clk),
    .Y(net411));
 NOR2x1_ASAP7_75t_R _23267_ (.A(_14622_),
    .B(_14768_),
    .Y(_14875_));
 AO21x1_ASAP7_75t_R _23268_ (.A1(_14761_),
    .A2(_14618_),
    .B(_14875_),
    .Y(_14876_));
 NOR2x1_ASAP7_75t_R _23269_ (.A(_14764_),
    .B(_14768_),
    .Y(_14877_));
 NOR2x1_ASAP7_75t_R _23270_ (.A(_14654_),
    .B(_14768_),
    .Y(_14878_));
 OR5x1_ASAP7_75t_R _23271_ (.A(_14871_),
    .B(_14873_),
    .C(_14876_),
    .D(_14877_),
    .E(_14878_),
    .Y(_14879_));
 AO21x1_ASAP7_75t_R _23272_ (.A1(_14735_),
    .A2(net3535),
    .B(_14776_),
    .Y(_14880_));
 NAND2x1_ASAP7_75t_R _23273_ (.A(_14779_),
    .B(_14880_),
    .Y(_14881_));
 NAND2x1_ASAP7_75t_R _23274_ (.A(_14775_),
    .B(_14661_),
    .Y(_14882_));
 NOR2x1_ASAP7_75t_R _23275_ (.A(_14776_),
    .B(_14636_),
    .Y(_14883_));
 INVx1_ASAP7_75t_R _23276_ (.A(_14883_),
    .Y(_14884_));
 NAND2x1_ASAP7_75t_R _23277_ (.A(_14882_),
    .B(_14884_),
    .Y(_14885_));
 NOR2x1_ASAP7_75t_R _23278_ (.A(_14716_),
    .B(_14776_),
    .Y(_14886_));
 AO21x1_ASAP7_75t_R _23279_ (.A1(_14732_),
    .A2(_14775_),
    .B(_14886_),
    .Y(_14887_));
 NAND2x1_ASAP7_75t_R _23280_ (.A(_14775_),
    .B(_14623_),
    .Y(_14888_));
 AO21x1_ASAP7_75t_R _23281_ (.A1(net3518),
    .A2(net3506),
    .B(_14776_),
    .Y(_14889_));
 NAND2x1_ASAP7_75t_R _23282_ (.A(_14888_),
    .B(_14889_),
    .Y(_14890_));
 OR4x1_ASAP7_75t_R _23283_ (.A(_14881_),
    .B(_14885_),
    .C(_14887_),
    .D(_14890_),
    .Y(_14891_));
 AO21x1_ASAP7_75t_R _23284_ (.A1(_14626_),
    .A2(_14782_),
    .B(_14787_),
    .Y(_14892_));
 NOR2x1_ASAP7_75t_R _23285_ (.A(net3535),
    .B(_14783_),
    .Y(_14893_));
 AO21x1_ASAP7_75t_R _23286_ (.A1(_14648_),
    .A2(_14782_),
    .B(_14893_),
    .Y(_14894_));
 AND3x1_ASAP7_75t_R _23287_ (.A(_14782_),
    .B(_14615_),
    .C(_14637_),
    .Y(_14895_));
 OR3x1_ASAP7_75t_R _23288_ (.A(_14892_),
    .B(_14894_),
    .C(_14895_),
    .Y(_14896_));
 NOR2x1_ASAP7_75t_R _23289_ (.A(_14814_),
    .B(_14793_),
    .Y(_14897_));
 AO21x1_ASAP7_75t_R _23290_ (.A1(_14648_),
    .A2(_14792_),
    .B(_14897_),
    .Y(_14898_));
 OA211x2_ASAP7_75t_R _23291_ (.A1(_14620_),
    .A2(_14672_),
    .B(_14792_),
    .C(net1985),
    .Y(_14899_));
 NOR2x1_ASAP7_75t_R _23292_ (.A(_14622_),
    .B(_14793_),
    .Y(_14900_));
 AO21x1_ASAP7_75t_R _23293_ (.A1(_14870_),
    .A2(_14792_),
    .B(_14900_),
    .Y(_14901_));
 OR3x1_ASAP7_75t_R _23294_ (.A(_14898_),
    .B(_14899_),
    .C(_14901_),
    .Y(_14902_));
 OR4x2_ASAP7_75t_R _23295_ (.A(_14879_),
    .B(_14891_),
    .C(_14896_),
    .D(_14902_),
    .Y(_14903_));
 NOR2x2_ASAP7_75t_R _23296_ (.A(_14869_),
    .B(_14903_),
    .Y(_14904_));
 INVx6_ASAP7_75t_R _23297_ (.A(_14642_),
    .Y(_14905_));
 OA21x2_ASAP7_75t_R _23298_ (.A1(_14674_),
    .A2(_14651_),
    .B(_14678_),
    .Y(_14906_));
 INVx1_ASAP7_75t_R _23299_ (.A(_14906_),
    .Y(_14907_));
 AO21x1_ASAP7_75t_R _23300_ (.A1(_14744_),
    .A2(_14735_),
    .B(_14686_),
    .Y(_14908_));
 NAND2x2_ASAP7_75t_R _23301_ (.A(net2197),
    .B(_14629_),
    .Y(_14909_));
 NOR2x2_ASAP7_75t_R _23302_ (.A(_14613_),
    .B(_14909_),
    .Y(_14910_));
 NAND2x1_ASAP7_75t_R _23303_ (.A(_14910_),
    .B(_14684_),
    .Y(_14911_));
 NAND2x1_ASAP7_75t_R _23304_ (.A(_14651_),
    .B(_14684_),
    .Y(_14912_));
 AND4x1_ASAP7_75t_R _23305_ (.A(_14908_),
    .B(_14911_),
    .C(_14685_),
    .D(_14912_),
    .Y(_14913_));
 INVx1_ASAP7_75t_R net399_5 (.A(clknet_leaf_7_clk),
    .Y(net410));
 AO21x1_ASAP7_75t_R _23307_ (.A1(_14733_),
    .A2(_14716_),
    .B(_14657_),
    .Y(_14915_));
 NAND2x1_ASAP7_75t_R _23308_ (.A(_14819_),
    .B(_14662_),
    .Y(_14916_));
 AO21x1_ASAP7_75t_R _23309_ (.A1(net1819),
    .A2(net3510),
    .B(_14657_),
    .Y(_14917_));
 AND4x1_ASAP7_75t_R _23310_ (.A(_14915_),
    .B(_14658_),
    .C(_14916_),
    .D(_14917_),
    .Y(_14918_));
 INVx5_ASAP7_75t_R _23311_ (.A(_14910_),
    .Y(_14919_));
 AO21x1_ASAP7_75t_R _23312_ (.A1(_14919_),
    .A2(net3510),
    .B(_14668_),
    .Y(_14920_));
 AO21x1_ASAP7_75t_R _23313_ (.A1(_14652_),
    .A2(net3521),
    .B(_14668_),
    .Y(_14921_));
 INVx4_ASAP7_75t_R _23314_ (.A(_14735_),
    .Y(_14922_));
 NAND2x1_ASAP7_75t_R _23315_ (.A(_14647_),
    .B(_14922_),
    .Y(_14923_));
 NAND2x1_ASAP7_75t_R _23316_ (.A(_14647_),
    .B(net3523),
    .Y(_14924_));
 AND4x1_ASAP7_75t_R _23317_ (.A(_14920_),
    .B(_14921_),
    .C(_14923_),
    .D(_14924_),
    .Y(_14925_));
 CKINVDCx6p67_ASAP7_75t_R _23318_ (.A(_14870_),
    .Y(_14926_));
 INVx1_ASAP7_75t_R net399_4 (.A(clknet_leaf_7_clk),
    .Y(net409));
 NAND2x1_ASAP7_75t_R _23320_ (.A(_14678_),
    .B(_14623_),
    .Y(_14928_));
 NAND2x1_ASAP7_75t_R _23321_ (.A(_14678_),
    .B(_14762_),
    .Y(_14929_));
 OA211x2_ASAP7_75t_R _23322_ (.A1(_14926_),
    .A2(_14694_),
    .B(_14928_),
    .C(_14929_),
    .Y(_14930_));
 AND5x1_ASAP7_75t_R _23323_ (.A(_14907_),
    .B(_14913_),
    .C(_14918_),
    .D(_14925_),
    .E(_14930_),
    .Y(_14931_));
 NAND2x1_ASAP7_75t_R _23324_ (.A(_14720_),
    .B(_14797_),
    .Y(_14932_));
 INVx1_ASAP7_75t_R net399_3 (.A(clknet_leaf_0_clk),
    .Y(net408));
 AO21x1_ASAP7_75t_R _23326_ (.A1(_14654_),
    .A2(net3521),
    .B(_14725_),
    .Y(_14934_));
 AO21x1_ASAP7_75t_R _23327_ (.A1(_14735_),
    .A2(_14764_),
    .B(_14725_),
    .Y(_14935_));
 OR3x1_ASAP7_75t_R _23328_ (.A(_14805_),
    .B(_14608_),
    .C(_14703_),
    .Y(_14936_));
 NAND2x1_ASAP7_75t_R _23329_ (.A(_14670_),
    .B(_14720_),
    .Y(_14937_));
 AND5x1_ASAP7_75t_R _23330_ (.A(_14932_),
    .B(_14934_),
    .C(_14935_),
    .D(_14936_),
    .E(_14937_),
    .Y(_14938_));
 OR3x1_ASAP7_75t_R _23331_ (.A(_14730_),
    .B(_14631_),
    .C(_14616_),
    .Y(_14939_));
 NAND2x1_ASAP7_75t_R _23332_ (.A(_14870_),
    .B(_14729_),
    .Y(_14940_));
 INVx1_ASAP7_75t_R net399_2 (.A(clknet_leaf_15_clk),
    .Y(net407));
 INVx1_ASAP7_75t_R _43355__1 (.A(clknet_leaf_8_clk),
    .Y(net406));
 AO21x1_ASAP7_75t_R _23335_ (.A1(_14636_),
    .A2(_14660_),
    .B(_14730_),
    .Y(_14943_));
 BUFx16f_ASAP7_75t_R load_slew405 (.A(net129),
    .Y(net405));
 AO21x1_ASAP7_75t_R _23337_ (.A1(_14804_),
    .A2(net1873),
    .B(_14730_),
    .Y(_14945_));
 AND4x1_ASAP7_75t_R _23338_ (.A(_14939_),
    .B(_14940_),
    .C(_14943_),
    .D(_14945_),
    .Y(_14946_));
 BUFx16f_ASAP7_75t_R load_slew404 (.A(net405),
    .Y(net404));
 AO21x1_ASAP7_75t_R _23340_ (.A1(_14804_),
    .A2(net1873),
    .B(_14712_),
    .Y(_14948_));
 AO21x1_ASAP7_75t_R _23341_ (.A1(_14926_),
    .A2(_14919_),
    .B(_14712_),
    .Y(_14949_));
 NAND2x1_ASAP7_75t_R _23342_ (.A(_14704_),
    .B(_14819_),
    .Y(_14950_));
 AND3x1_ASAP7_75t_R _23343_ (.A(_14948_),
    .B(_14949_),
    .C(_14950_),
    .Y(_14951_));
 AO21x2_ASAP7_75t_R _23344_ (.A1(_14744_),
    .A2(_14735_),
    .B(_14740_),
    .Y(_14952_));
 NAND2x1_ASAP7_75t_R _23345_ (.A(_14739_),
    .B(_14797_),
    .Y(_14953_));
 NAND2x1_ASAP7_75t_R _23346_ (.A(_14739_),
    .B(_14819_),
    .Y(_14954_));
 AO21x1_ASAP7_75t_R _23347_ (.A1(_14733_),
    .A2(net1873),
    .B(_14740_),
    .Y(_14955_));
 AND4x1_ASAP7_75t_R _23348_ (.A(_14952_),
    .B(_14953_),
    .C(_14954_),
    .D(_14955_),
    .Y(_14956_));
 AND4x1_ASAP7_75t_R _23349_ (.A(_14938_),
    .B(_14946_),
    .C(_14951_),
    .D(_14956_),
    .Y(_14957_));
 AND2x2_ASAP7_75t_R _23350_ (.A(_14931_),
    .B(_14957_),
    .Y(_14958_));
 AND3x4_ASAP7_75t_R _23351_ (.A(_14904_),
    .B(_14905_),
    .C(_14958_),
    .Y(_14959_));
 BUFx16f_ASAP7_75t_R load_slew403 (.A(net404),
    .Y(net403));
 XNOR2x1_ASAP7_75t_R _23353_ (.B(_00475_),
    .Y(_14961_),
    .A(net3543));
 BUFx16f_ASAP7_75t_R load_slew402 (.A(net405),
    .Y(net402));
 XNOR2x2_ASAP7_75t_R _23355_ (.A(_00495_),
    .B(_00519_),
    .Y(_14963_));
 XNOR2x1_ASAP7_75t_R _23356_ (.B(_14963_),
    .Y(_14964_),
    .A(_14961_));
 XOR2x1_ASAP7_75t_R _23357_ (.A(_14959_),
    .Y(_14965_),
    .B(_14964_));
 AND2x2_ASAP7_75t_R _23358_ (.A(net402),
    .B(net128),
    .Y(_14966_));
 AO21x1_ASAP7_75t_R _23359_ (.A1(_14965_),
    .A2(net399),
    .B(_14966_),
    .Y(_00384_));
 NAND2x1_ASAP7_75t_R _23360_ (.A(_14782_),
    .B(_14922_),
    .Y(_14967_));
 NOR2x1_ASAP7_75t_R _23361_ (.A(_14919_),
    .B(_14793_),
    .Y(_14968_));
 INVx1_ASAP7_75t_R _23362_ (.A(_14968_),
    .Y(_14969_));
 INVx2_ASAP7_75t_R _23363_ (.A(_14716_),
    .Y(_14970_));
 NAND2x1_ASAP7_75t_R _23364_ (.A(_14970_),
    .B(_14792_),
    .Y(_14971_));
 NAND2x1_ASAP7_75t_R _23365_ (.A(_14661_),
    .B(_14792_),
    .Y(_14972_));
 AND4x1_ASAP7_75t_R _23366_ (.A(_14795_),
    .B(_14969_),
    .C(_14971_),
    .D(_14972_),
    .Y(_14973_));
 AO21x1_ASAP7_75t_R _23367_ (.A1(net3510),
    .A2(net2178),
    .B(_14783_),
    .Y(_14974_));
 NAND2x1_ASAP7_75t_R _23368_ (.A(_14782_),
    .B(_14970_),
    .Y(_14975_));
 AND3x1_ASAP7_75t_R _23369_ (.A(_14974_),
    .B(_14975_),
    .C(_14788_),
    .Y(_14976_));
 BUFx16f_ASAP7_75t_R wire401 (.A(net405),
    .Y(net401));
 NOR2x1_ASAP7_75t_R _23371_ (.A(_14764_),
    .B(_14783_),
    .Y(_14978_));
 INVx1_ASAP7_75t_R _23372_ (.A(_14978_),
    .Y(_14979_));
 NAND2x1_ASAP7_75t_R _23373_ (.A(_14782_),
    .B(_14635_),
    .Y(_14980_));
 AND5x2_ASAP7_75t_R _23374_ (.A(_14967_),
    .B(_14973_),
    .C(_14976_),
    .D(_14979_),
    .E(_14980_),
    .Y(_14981_));
 AO21x1_ASAP7_75t_R _23375_ (.A1(_14654_),
    .A2(_14636_),
    .B(_14816_),
    .Y(_14982_));
 AO21x1_ASAP7_75t_R _23376_ (.A1(net1830),
    .A2(net2136),
    .B(_14816_),
    .Y(_14983_));
 AO21x1_ASAP7_75t_R _23377_ (.A1(_14715_),
    .A2(net2179),
    .B(_14816_),
    .Y(_14984_));
 AND4x1_ASAP7_75t_R _23378_ (.A(_14982_),
    .B(_14983_),
    .C(_14984_),
    .D(_14824_),
    .Y(_14985_));
 AO21x1_ASAP7_75t_R _23379_ (.A1(_14636_),
    .A2(_14652_),
    .B(_14610_),
    .Y(_14986_));
 AO21x1_ASAP7_75t_R _23380_ (.A1(_14926_),
    .A2(_14667_),
    .B(_14610_),
    .Y(_14987_));
 AND3x1_ASAP7_75t_R _23381_ (.A(_14986_),
    .B(_14827_),
    .C(_14987_),
    .Y(_14988_));
 AO21x1_ASAP7_75t_R _23382_ (.A1(_14804_),
    .A2(_14716_),
    .B(_14835_),
    .Y(_14989_));
 BUFx16f_ASAP7_75t_R wire400 (.A(_08823_),
    .Y(net400));
 AO21x1_ASAP7_75t_R _23384_ (.A1(net2136),
    .A2(net1943),
    .B(_14835_),
    .Y(_14991_));
 AO21x1_ASAP7_75t_R _23385_ (.A1(_14919_),
    .A2(net3510),
    .B(_14835_),
    .Y(_14992_));
 AND3x1_ASAP7_75t_R _23386_ (.A(_14989_),
    .B(_14991_),
    .C(_14992_),
    .Y(_14993_));
 AO21x1_ASAP7_75t_R _23387_ (.A1(_14926_),
    .A2(_14919_),
    .B(_14807_),
    .Y(_14994_));
 AO21x1_ASAP7_75t_R _23388_ (.A1(_14631_),
    .A2(_14757_),
    .B(_14807_),
    .Y(_14995_));
 OA211x2_ASAP7_75t_R _23389_ (.A1(_14715_),
    .A2(_14807_),
    .B(_14994_),
    .C(_14995_),
    .Y(_14996_));
 AND4x2_ASAP7_75t_R _23390_ (.A(_14985_),
    .B(_14988_),
    .C(_14993_),
    .D(_14996_),
    .Y(_14997_));
 NAND2x1_ASAP7_75t_R _23391_ (.A(_14651_),
    .B(_14775_),
    .Y(_14998_));
 AO21x1_ASAP7_75t_R _23392_ (.A1(net1874),
    .A2(net2179),
    .B(_14768_),
    .Y(_14999_));
 INVx1_ASAP7_75t_R _23393_ (.A(_14871_),
    .Y(_15000_));
 NAND2x1_ASAP7_75t_R _23394_ (.A(_14761_),
    .B(_14661_),
    .Y(_15001_));
 NAND2x2_ASAP7_75t_R _23395_ (.A(_14761_),
    .B(_14922_),
    .Y(_15002_));
 AND4x1_ASAP7_75t_R _23396_ (.A(_14999_),
    .B(_15000_),
    .C(_15001_),
    .D(_15002_),
    .Y(_15003_));
 NAND2x1_ASAP7_75t_R _23397_ (.A(_14775_),
    .B(_14922_),
    .Y(_15004_));
 NAND2x1_ASAP7_75t_R _23398_ (.A(_14775_),
    .B(_14870_),
    .Y(_15005_));
 BUFx16f_ASAP7_75t_R load_slew399 (.A(_08823_),
    .Y(net399));
 AO21x1_ASAP7_75t_R _23400_ (.A1(_14733_),
    .A2(net1874),
    .B(_14776_),
    .Y(_15007_));
 AND5x2_ASAP7_75t_R _23401_ (.A(_14998_),
    .B(_15003_),
    .C(_15004_),
    .D(_15005_),
    .E(_15007_),
    .Y(_15008_));
 NAND3x2_ASAP7_75t_R _23402_ (.B(_14997_),
    .C(_15008_),
    .Y(_15009_),
    .A(_14981_));
 AO21x1_ASAP7_75t_R _23403_ (.A1(_14744_),
    .A2(net1830),
    .B(_14657_),
    .Y(_15010_));
 AO21x1_ASAP7_75t_R _23404_ (.A1(_14926_),
    .A2(_14919_),
    .B(_14657_),
    .Y(_15011_));
 AO21x1_ASAP7_75t_R _23405_ (.A1(_14733_),
    .A2(_14804_),
    .B(_14657_),
    .Y(_15012_));
 AND5x1_ASAP7_75t_R _23406_ (.A(_14664_),
    .B(_15010_),
    .C(_14916_),
    .D(_15011_),
    .E(_15012_),
    .Y(_15013_));
 AO21x1_ASAP7_75t_R _23407_ (.A1(_14757_),
    .A2(_14631_),
    .B(_14694_),
    .Y(_15014_));
 OR3x1_ASAP7_75t_R _23408_ (.A(_14638_),
    .B(_14646_),
    .C(_14683_),
    .Y(_15015_));
 AO21x1_ASAP7_75t_R _23409_ (.A1(_14919_),
    .A2(net3510),
    .B(_14686_),
    .Y(_15016_));
 OR3x1_ASAP7_75t_R _23410_ (.A(_14860_),
    .B(_14646_),
    .C(_14683_),
    .Y(_15017_));
 AO21x1_ASAP7_75t_R _23411_ (.A1(_14728_),
    .A2(_14860_),
    .B(_14694_),
    .Y(_15018_));
 AND5x1_ASAP7_75t_R _23412_ (.A(_15014_),
    .B(_15015_),
    .C(_15016_),
    .D(_15017_),
    .E(_15018_),
    .Y(_15019_));
 NAND2x1_ASAP7_75t_R _23413_ (.A(_14647_),
    .B(_14870_),
    .Y(_15020_));
 AO21x1_ASAP7_75t_R _23414_ (.A1(_14733_),
    .A2(net2179),
    .B(_14668_),
    .Y(_15021_));
 NOR2x1_ASAP7_75t_R _23415_ (.A(_14764_),
    .B(_14668_),
    .Y(_15022_));
 INVx1_ASAP7_75t_R _23416_ (.A(_15022_),
    .Y(_15023_));
 NAND2x1_ASAP7_75t_R _23417_ (.A(_14647_),
    .B(_14819_),
    .Y(_15024_));
 AND5x1_ASAP7_75t_R _23418_ (.A(_15020_),
    .B(_15021_),
    .C(_14923_),
    .D(_15023_),
    .E(_15024_),
    .Y(_15025_));
 AND3x2_ASAP7_75t_R _23419_ (.A(_15013_),
    .B(_15019_),
    .C(_15025_),
    .Y(_15026_));
 NAND2x1_ASAP7_75t_R _23420_ (.A(_14630_),
    .B(_14720_),
    .Y(_15027_));
 AO21x1_ASAP7_75t_R _23421_ (.A1(_14926_),
    .A2(net3524),
    .B(_14730_),
    .Y(_15028_));
 OR3x1_ASAP7_75t_R _23422_ (.A(_14805_),
    .B(_14683_),
    .C(_14703_),
    .Y(_15029_));
 OA211x2_ASAP7_75t_R _23423_ (.A1(_14804_),
    .A2(_14730_),
    .B(_15028_),
    .C(_15029_),
    .Y(_15030_));
 AO21x1_ASAP7_75t_R _23424_ (.A1(net1943),
    .A2(_14652_),
    .B(_14730_),
    .Y(_15031_));
 NAND2x1_ASAP7_75t_R _23425_ (.A(_14729_),
    .B(net3523),
    .Y(_15032_));
 NOR2x1_ASAP7_75t_R _23426_ (.A(_14766_),
    .B(_14730_),
    .Y(_15033_));
 INVx1_ASAP7_75t_R _23427_ (.A(_15033_),
    .Y(_15034_));
 INVx2_ASAP7_75t_R _23428_ (.A(_14764_),
    .Y(_15035_));
 NAND2x1_ASAP7_75t_R _23429_ (.A(_14729_),
    .B(_15035_),
    .Y(_15036_));
 AND4x1_ASAP7_75t_R _23430_ (.A(_15031_),
    .B(_15032_),
    .C(_15034_),
    .D(_15036_),
    .Y(_15037_));
 AO21x1_ASAP7_75t_R _23431_ (.A1(_14652_),
    .A2(net1943),
    .B(_14725_),
    .Y(_15038_));
 NAND2x1_ASAP7_75t_R _23432_ (.A(_14629_),
    .B(_14621_),
    .Y(_15039_));
 AO21x1_ASAP7_75t_R _23433_ (.A1(_14625_),
    .A2(_15039_),
    .B(_14725_),
    .Y(_15040_));
 AND5x2_ASAP7_75t_R _23434_ (.A(_15027_),
    .B(_15030_),
    .C(_15037_),
    .D(_15038_),
    .E(_15040_),
    .Y(_15041_));
 NAND2x1_ASAP7_75t_R _23435_ (.A(_14672_),
    .B(net1987),
    .Y(_15042_));
 AO21x1_ASAP7_75t_R _23436_ (.A1(net3506),
    .A2(_15042_),
    .B(_14740_),
    .Y(_15043_));
 AO21x1_ASAP7_75t_R _23437_ (.A1(_14654_),
    .A2(net1943),
    .B(_14740_),
    .Y(_15044_));
 AND3x1_ASAP7_75t_R _23438_ (.A(_14952_),
    .B(_15043_),
    .C(_15044_),
    .Y(_15045_));
 BUFx16f_ASAP7_75t_R max_length398 (.A(net399),
    .Y(net398));
 AO21x1_ASAP7_75t_R _23440_ (.A1(net3509),
    .A2(net2136),
    .B(_14712_),
    .Y(_15047_));
 AO21x1_ASAP7_75t_R _23441_ (.A1(_14926_),
    .A2(net1819),
    .B(_14712_),
    .Y(_15048_));
 OA211x2_ASAP7_75t_R _23442_ (.A1(_00451_),
    .A2(_14672_),
    .B(_14704_),
    .C(net1989),
    .Y(_15049_));
 INVx1_ASAP7_75t_R _23443_ (.A(_15049_),
    .Y(_15050_));
 AND4x2_ASAP7_75t_R _23444_ (.A(_15045_),
    .B(_15047_),
    .C(_15048_),
    .D(_15050_),
    .Y(_15051_));
 NAND3x2_ASAP7_75t_R _23445_ (.B(_15041_),
    .C(_15051_),
    .Y(_15052_),
    .A(_15026_));
 NOR2x2_ASAP7_75t_R _23446_ (.A(_15009_),
    .B(_15052_),
    .Y(_15053_));
 XOR2x2_ASAP7_75t_R _23447_ (.A(_00474_),
    .B(_00518_),
    .Y(_15054_));
 BUFx16f_ASAP7_75t_R load_slew397 (.A(_00528_),
    .Y(net397));
 XOR2x1_ASAP7_75t_R _23449_ (.A(_00389_),
    .Y(_15056_),
    .B(_00442_));
 XNOR2x1_ASAP7_75t_R _23450_ (.B(_15056_),
    .Y(_15057_),
    .A(_15054_));
 XOR2x1_ASAP7_75t_R _23451_ (.A(_15053_),
    .Y(_15058_),
    .B(_15057_));
 AND2x2_ASAP7_75t_R _23452_ (.A(net402),
    .B(net12),
    .Y(_15059_));
 AO21x1_ASAP7_75t_R _23453_ (.A1(_15058_),
    .A2(net399),
    .B(_15059_),
    .Y(_00354_));
 AO21x1_ASAP7_75t_R _23454_ (.A1(_14733_),
    .A2(_14804_),
    .B(_14776_),
    .Y(_15060_));
 AO21x1_ASAP7_75t_R _23455_ (.A1(_14654_),
    .A2(_14638_),
    .B(_14776_),
    .Y(_15061_));
 AND5x1_ASAP7_75t_R _23456_ (.A(_14779_),
    .B(_15060_),
    .C(_15061_),
    .D(_14880_),
    .E(_14888_),
    .Y(_15062_));
 AO21x1_ASAP7_75t_R _23457_ (.A1(_14606_),
    .A2(_14909_),
    .B(_14768_),
    .Y(_15063_));
 NOR2x1_ASAP7_75t_R _23458_ (.A(net3508),
    .B(_14768_),
    .Y(_15064_));
 INVx1_ASAP7_75t_R _23459_ (.A(_15064_),
    .Y(_15065_));
 INVx1_ASAP7_75t_R _23460_ (.A(_14877_),
    .Y(_15066_));
 AND5x1_ASAP7_75t_R _23461_ (.A(_15063_),
    .B(_15065_),
    .C(_15066_),
    .D(_15001_),
    .E(_15002_),
    .Y(_15067_));
 INVx1_ASAP7_75t_R _23462_ (.A(_14895_),
    .Y(_15068_));
 AO21x1_ASAP7_75t_R _23463_ (.A1(net3510),
    .A2(net3524),
    .B(_14783_),
    .Y(_15069_));
 AO21x1_ASAP7_75t_R _23464_ (.A1(net2179),
    .A2(_14805_),
    .B(_14783_),
    .Y(_15070_));
 AND4x1_ASAP7_75t_R _23465_ (.A(_15068_),
    .B(_14967_),
    .C(_15069_),
    .D(_15070_),
    .Y(_15071_));
 AO21x1_ASAP7_75t_R _23466_ (.A1(net1830),
    .A2(net2136),
    .B(_14793_),
    .Y(_15072_));
 AO21x1_ASAP7_75t_R _23467_ (.A1(_14926_),
    .A2(net2178),
    .B(_14793_),
    .Y(_15073_));
 AND4x1_ASAP7_75t_R _23468_ (.A(_15072_),
    .B(_15073_),
    .C(_14971_),
    .D(_14972_),
    .Y(_15074_));
 AND4x2_ASAP7_75t_R _23469_ (.A(_15062_),
    .B(_15067_),
    .C(_15071_),
    .D(_15074_),
    .Y(_15075_));
 NOR2x1_ASAP7_75t_R _23470_ (.A(_14804_),
    .B(_14816_),
    .Y(_15076_));
 INVx1_ASAP7_75t_R _23471_ (.A(_15076_),
    .Y(_15077_));
 AO21x1_ASAP7_75t_R _23472_ (.A1(_14744_),
    .A2(net1830),
    .B(_14835_),
    .Y(_15078_));
 AND3x1_ASAP7_75t_R _23473_ (.A(_14834_),
    .B(_14634_),
    .C(_14637_),
    .Y(_15079_));
 INVx1_ASAP7_75t_R _23474_ (.A(_15079_),
    .Y(_15080_));
 NAND2x1_ASAP7_75t_R _23475_ (.A(_14834_),
    .B(_14670_),
    .Y(_15081_));
 AND4x1_ASAP7_75t_R _23476_ (.A(_15078_),
    .B(_15080_),
    .C(_15081_),
    .D(_14837_),
    .Y(_15082_));
 OR3x1_ASAP7_75t_R _23477_ (.A(_14814_),
    .B(_14607_),
    .C(_14608_),
    .Y(_15083_));
 NAND2x1_ASAP7_75t_R _23478_ (.A(_14609_),
    .B(_14797_),
    .Y(_15084_));
 AO21x1_ASAP7_75t_R _23479_ (.A1(_14733_),
    .A2(_14804_),
    .B(_14610_),
    .Y(_15085_));
 AO21x1_ASAP7_75t_R _23480_ (.A1(net1830),
    .A2(net2136),
    .B(_14610_),
    .Y(_15086_));
 AND4x1_ASAP7_75t_R _23481_ (.A(_15083_),
    .B(_15084_),
    .C(_15085_),
    .D(_15086_),
    .Y(_15087_));
 AO21x1_ASAP7_75t_R _23482_ (.A1(net3509),
    .A2(net1830),
    .B(_14807_),
    .Y(_15088_));
 NAND2x1_ASAP7_75t_R _23483_ (.A(_14806_),
    .B(_14635_),
    .Y(_15089_));
 NAND2x1_ASAP7_75t_R _23484_ (.A(_14806_),
    .B(_14970_),
    .Y(_15090_));
 AND3x1_ASAP7_75t_R _23485_ (.A(_15088_),
    .B(_15089_),
    .C(_15090_),
    .Y(_15091_));
 AO21x1_ASAP7_75t_R _23486_ (.A1(net3509),
    .A2(_14744_),
    .B(_14816_),
    .Y(_15092_));
 AND5x2_ASAP7_75t_R _23487_ (.A(_15077_),
    .B(_15082_),
    .C(_15087_),
    .D(_15091_),
    .E(_15092_),
    .Y(_15093_));
 NAND2x2_ASAP7_75t_R _23488_ (.A(_15075_),
    .B(_15093_),
    .Y(_15094_));
 AO21x1_ASAP7_75t_R _23489_ (.A1(_14744_),
    .A2(_14757_),
    .B(_14694_),
    .Y(_15095_));
 NOR2x1_ASAP7_75t_R _23490_ (.A(net3506),
    .B(_14694_),
    .Y(_15096_));
 INVx1_ASAP7_75t_R _23491_ (.A(_15096_),
    .Y(_15097_));
 AO21x1_ASAP7_75t_R _23492_ (.A1(_14733_),
    .A2(net2179),
    .B(_14694_),
    .Y(_15098_));
 AND3x1_ASAP7_75t_R _23493_ (.A(_15095_),
    .B(_15097_),
    .C(_15098_),
    .Y(_15099_));
 OA211x2_ASAP7_75t_R _23494_ (.A1(_14620_),
    .A2(net3517),
    .B(_14662_),
    .C(net2721),
    .Y(_15100_));
 INVx1_ASAP7_75t_R _23495_ (.A(_15100_),
    .Y(_15101_));
 OA211x2_ASAP7_75t_R _23496_ (.A1(_14636_),
    .A2(_14657_),
    .B(_15101_),
    .C(_14663_),
    .Y(_15102_));
 AO21x1_ASAP7_75t_R _23497_ (.A1(_14926_),
    .A2(net1819),
    .B(_14686_),
    .Y(_15103_));
 AO21x1_ASAP7_75t_R _23498_ (.A1(net3509),
    .A2(net1830),
    .B(_14686_),
    .Y(_15104_));
 AND4x1_ASAP7_75t_R _23499_ (.A(_15015_),
    .B(_14685_),
    .C(_15103_),
    .D(_15104_),
    .Y(_15105_));
 AO21x1_ASAP7_75t_R _23500_ (.A1(_14926_),
    .A2(net1875),
    .B(_14668_),
    .Y(_15106_));
 AND4x1_ASAP7_75t_R _23501_ (.A(_15106_),
    .B(_14921_),
    .C(_14649_),
    .D(_15023_),
    .Y(_15107_));
 AO21x1_ASAP7_75t_R _23502_ (.A1(net2178),
    .A2(net3510),
    .B(_14657_),
    .Y(_15108_));
 NOR2x1_ASAP7_75t_R _23503_ (.A(_14716_),
    .B(_14657_),
    .Y(_15109_));
 INVx1_ASAP7_75t_R _23504_ (.A(_15109_),
    .Y(_15110_));
 OA211x2_ASAP7_75t_R _23505_ (.A1(_14805_),
    .A2(_14657_),
    .B(_15108_),
    .C(_15110_),
    .Y(_15111_));
 AND5x1_ASAP7_75t_R _23506_ (.A(_15099_),
    .B(_15102_),
    .C(_15105_),
    .D(_15107_),
    .E(_15111_),
    .Y(_15112_));
 NOR3x1_ASAP7_75t_R _23507_ (.A(_14750_),
    .B(_14751_),
    .C(_14748_),
    .Y(_15113_));
 INVx1_ASAP7_75t_R _23508_ (.A(_14745_),
    .Y(_15114_));
 NAND2x1_ASAP7_75t_R _23509_ (.A(_14653_),
    .B(_14739_),
    .Y(_15115_));
 NOR2x1_ASAP7_75t_R _23510_ (.A(_14764_),
    .B(_14740_),
    .Y(_15116_));
 INVx1_ASAP7_75t_R _23511_ (.A(_15116_),
    .Y(_15117_));
 AND5x1_ASAP7_75t_R _23512_ (.A(_15113_),
    .B(_15114_),
    .C(_14741_),
    .D(_15115_),
    .E(_15117_),
    .Y(_15118_));
 NOR2x2_ASAP7_75t_R _23513_ (.A(_14692_),
    .B(_14730_),
    .Y(_15119_));
 INVx1_ASAP7_75t_R _23514_ (.A(_15119_),
    .Y(_15120_));
 NAND2x1_ASAP7_75t_R _23515_ (.A(_14729_),
    .B(_14648_),
    .Y(_15121_));
 AND5x1_ASAP7_75t_R _23516_ (.A(_15032_),
    .B(_15029_),
    .C(_15120_),
    .D(_15036_),
    .E(_15121_),
    .Y(_15122_));
 NAND2x1_ASAP7_75t_R _23517_ (.A(_14704_),
    .B(net3523),
    .Y(_15123_));
 NAND2x1_ASAP7_75t_R _23518_ (.A(_14651_),
    .B(_14704_),
    .Y(_15124_));
 AND4x1_ASAP7_75t_R _23519_ (.A(_14706_),
    .B(_15123_),
    .C(_14950_),
    .D(_15124_),
    .Y(_15125_));
 OA211x2_ASAP7_75t_R _23520_ (.A1(_14620_),
    .A2(net3513),
    .B(_14704_),
    .C(net1989),
    .Y(_15126_));
 INVx1_ASAP7_75t_R _23521_ (.A(_15126_),
    .Y(_15127_));
 NAND2x1_ASAP7_75t_R _23522_ (.A(_14910_),
    .B(_14704_),
    .Y(_15128_));
 OA211x2_ASAP7_75t_R _23523_ (.A1(_14692_),
    .A2(_14712_),
    .B(_15127_),
    .C(_15128_),
    .Y(_15129_));
 NAND2x1_ASAP7_75t_R _23524_ (.A(net1985),
    .B(_14720_),
    .Y(_15130_));
 AO21x1_ASAP7_75t_R _23525_ (.A1(net1943),
    .A2(_14809_),
    .B(_14725_),
    .Y(_15131_));
 NAND2x1_ASAP7_75t_R _23526_ (.A(_14720_),
    .B(_14648_),
    .Y(_15132_));
 NAND2x1_ASAP7_75t_R _23527_ (.A(_14910_),
    .B(_14720_),
    .Y(_15133_));
 AND5x1_ASAP7_75t_R _23528_ (.A(_15130_),
    .B(_15131_),
    .C(_15132_),
    .D(_14932_),
    .E(_15133_),
    .Y(_15134_));
 AND5x2_ASAP7_75t_R _23529_ (.A(_15118_),
    .B(_15122_),
    .C(_15125_),
    .D(_15129_),
    .E(_15134_),
    .Y(_15135_));
 NAND2x2_ASAP7_75t_R _23530_ (.A(_15112_),
    .B(_15135_),
    .Y(_15136_));
 NOR2x2_ASAP7_75t_R _23531_ (.A(_15094_),
    .B(_15136_),
    .Y(_15137_));
 BUFx16f_ASAP7_75t_R load_slew396 (.A(_00528_),
    .Y(net396));
 XOR2x2_ASAP7_75t_R _23533_ (.A(_00473_),
    .B(_00517_),
    .Y(_15139_));
 BUFx16f_ASAP7_75t_R load_slew395 (.A(net396),
    .Y(net395));
 XOR2x1_ASAP7_75t_R _23535_ (.A(_00390_),
    .Y(_15141_),
    .B(_00441_));
 XNOR2x1_ASAP7_75t_R _23536_ (.B(_15141_),
    .Y(_15142_),
    .A(_15139_));
 XOR2x1_ASAP7_75t_R _23537_ (.A(_15137_),
    .Y(_15143_),
    .B(_15142_));
 AND2x2_ASAP7_75t_R _23538_ (.A(net404),
    .B(net4120),
    .Y(_15144_));
 AO21x1_ASAP7_75t_R _23539_ (.A1(_15143_),
    .A2(net399),
    .B(_15144_),
    .Y(_00355_));
 OR3x1_ASAP7_75t_R _23540_ (.A(_14906_),
    .B(_15096_),
    .C(_14690_),
    .Y(_15145_));
 NOR2x1_ASAP7_75t_R _23541_ (.A(_14735_),
    .B(_14657_),
    .Y(_15146_));
 AO21x1_ASAP7_75t_R _23542_ (.A1(_14651_),
    .A2(_14662_),
    .B(_15146_),
    .Y(_15147_));
 OA21x2_ASAP7_75t_R _23543_ (.A1(_14623_),
    .A2(_14870_),
    .B(_14662_),
    .Y(_15148_));
 OR3x1_ASAP7_75t_R _23544_ (.A(_15147_),
    .B(_15109_),
    .C(_15148_),
    .Y(_15149_));
 OA21x2_ASAP7_75t_R _23545_ (.A1(_14661_),
    .A2(_14819_),
    .B(_14684_),
    .Y(_15150_));
 NOR2x1_ASAP7_75t_R _23546_ (.A(_14667_),
    .B(_14686_),
    .Y(_15151_));
 AO21x1_ASAP7_75t_R _23547_ (.A1(_14626_),
    .A2(_14684_),
    .B(_15151_),
    .Y(_15152_));
 INVx1_ASAP7_75t_R _23548_ (.A(_14669_),
    .Y(_15153_));
 NAND2x1_ASAP7_75t_R _23549_ (.A(_14651_),
    .B(_14647_),
    .Y(_15154_));
 NAND2x1_ASAP7_75t_R _23550_ (.A(_15154_),
    .B(_14924_),
    .Y(_15155_));
 OR3x1_ASAP7_75t_R _23551_ (.A(_15153_),
    .B(_15022_),
    .C(_15155_),
    .Y(_15156_));
 OR5x1_ASAP7_75t_R _23552_ (.A(_15145_),
    .B(_15149_),
    .C(_15150_),
    .D(_15152_),
    .E(_15156_),
    .Y(_15157_));
 AO21x1_ASAP7_75t_R _23553_ (.A1(net3521),
    .A2(_14652_),
    .B(_14712_),
    .Y(_15158_));
 AO21x1_ASAP7_75t_R _23554_ (.A1(net3509),
    .A2(_14735_),
    .B(_14712_),
    .Y(_15159_));
 AND3x1_ASAP7_75t_R _23555_ (.A(_15158_),
    .B(_15159_),
    .C(_15123_),
    .Y(_15160_));
 AO21x1_ASAP7_75t_R _23556_ (.A1(_14606_),
    .A2(_15039_),
    .B(_14740_),
    .Y(_15161_));
 AND5x1_ASAP7_75t_R _23557_ (.A(_15114_),
    .B(_15160_),
    .C(_14718_),
    .D(_15128_),
    .E(_15161_),
    .Y(_15162_));
 AO21x1_ASAP7_75t_R _23558_ (.A1(_14744_),
    .A2(net2136),
    .B(_14725_),
    .Y(_15163_));
 OA211x2_ASAP7_75t_R _23559_ (.A1(_14809_),
    .A2(_14725_),
    .B(_15163_),
    .C(_15040_),
    .Y(_15164_));
 AO21x1_ASAP7_75t_R _23560_ (.A1(_14809_),
    .A2(_14652_),
    .B(_14730_),
    .Y(_15165_));
 OA211x2_ASAP7_75t_R _23561_ (.A1(_14620_),
    .A2(_14672_),
    .B(_14729_),
    .C(_14614_),
    .Y(_15166_));
 INVx1_ASAP7_75t_R _23562_ (.A(_15166_),
    .Y(_15167_));
 AND5x1_ASAP7_75t_R _23563_ (.A(_15034_),
    .B(_15164_),
    .C(_15029_),
    .D(_15165_),
    .E(_15167_),
    .Y(_15168_));
 NAND2x1_ASAP7_75t_R _23564_ (.A(_15162_),
    .B(_15168_),
    .Y(_15169_));
 NOR2x1_ASAP7_75t_R _23565_ (.A(_15157_),
    .B(_15169_),
    .Y(_15170_));
 INVx1_ASAP7_75t_R _23566_ (.A(_14674_),
    .Y(_15171_));
 NAND2x1_ASAP7_75t_R _23567_ (.A(net1986),
    .B(_14806_),
    .Y(_15172_));
 AO21x1_ASAP7_75t_R _23568_ (.A1(net3510),
    .A2(net3518),
    .B(_14807_),
    .Y(_15173_));
 AND4x1_ASAP7_75t_R _23569_ (.A(_14857_),
    .B(_15172_),
    .C(_14810_),
    .D(_15173_),
    .Y(_15174_));
 AO21x1_ASAP7_75t_R _23570_ (.A1(net1817),
    .A2(_14805_),
    .B(_14816_),
    .Y(_15175_));
 OA211x2_ASAP7_75t_R _23571_ (.A1(_14816_),
    .A2(_15171_),
    .B(_15174_),
    .C(_15175_),
    .Y(_15176_));
 AO21x1_ASAP7_75t_R _23572_ (.A1(_14804_),
    .A2(_14716_),
    .B(_14610_),
    .Y(_15177_));
 NAND2x1_ASAP7_75t_R _23573_ (.A(_14609_),
    .B(_14762_),
    .Y(_15178_));
 NAND2x1_ASAP7_75t_R _23574_ (.A(_14609_),
    .B(_14648_),
    .Y(_15179_));
 AND5x1_ASAP7_75t_R _23575_ (.A(_15177_),
    .B(_14639_),
    .C(_15178_),
    .D(_15179_),
    .E(_14619_),
    .Y(_15180_));
 AO21x1_ASAP7_75t_R _23576_ (.A1(_14733_),
    .A2(_14804_),
    .B(_14835_),
    .Y(_15181_));
 NOR2x1_ASAP7_75t_R _23577_ (.A(net1817),
    .B(_14835_),
    .Y(_15182_));
 INVx1_ASAP7_75t_R _23578_ (.A(_15182_),
    .Y(_15183_));
 NAND2x1_ASAP7_75t_R _23579_ (.A(_14834_),
    .B(_14661_),
    .Y(_15184_));
 NAND2x1_ASAP7_75t_R _23580_ (.A(_14834_),
    .B(_14674_),
    .Y(_15185_));
 AND4x1_ASAP7_75t_R _23581_ (.A(_15181_),
    .B(_15183_),
    .C(_15184_),
    .D(_15185_),
    .Y(_15186_));
 AND3x1_ASAP7_75t_R _23582_ (.A(_15176_),
    .B(_15180_),
    .C(_15186_),
    .Y(_15187_));
 AO21x1_ASAP7_75t_R _23583_ (.A1(_14870_),
    .A2(_14792_),
    .B(_14899_),
    .Y(_15188_));
 NOR2x1_ASAP7_75t_R _23584_ (.A(_14968_),
    .B(_15188_),
    .Y(_15189_));
 NAND2x1_ASAP7_75t_R _23585_ (.A(_14670_),
    .B(_14792_),
    .Y(_15190_));
 AO21x1_ASAP7_75t_R _23586_ (.A1(_14733_),
    .A2(_14860_),
    .B(_14783_),
    .Y(_15191_));
 AO21x1_ASAP7_75t_R _23587_ (.A1(_14654_),
    .A2(_14660_),
    .B(_14783_),
    .Y(_15192_));
 INVx1_ASAP7_75t_R _23588_ (.A(_14893_),
    .Y(_15193_));
 AND4x1_ASAP7_75t_R _23589_ (.A(_15191_),
    .B(_15069_),
    .C(_15192_),
    .D(_15193_),
    .Y(_15194_));
 AO21x1_ASAP7_75t_R _23590_ (.A1(_14654_),
    .A2(_14631_),
    .B(_14793_),
    .Y(_15195_));
 AND4x1_ASAP7_75t_R _23591_ (.A(_15189_),
    .B(_15190_),
    .C(_15194_),
    .D(_15195_),
    .Y(_15196_));
 AO21x1_ASAP7_75t_R _23592_ (.A1(_14636_),
    .A2(_14654_),
    .B(_14768_),
    .Y(_15197_));
 AO21x1_ASAP7_75t_R _23593_ (.A1(_14733_),
    .A2(net3507),
    .B(_14768_),
    .Y(_15198_));
 AND4x1_ASAP7_75t_R _23594_ (.A(_15197_),
    .B(_14769_),
    .C(_15002_),
    .D(_15198_),
    .Y(_15199_));
 AO21x1_ASAP7_75t_R _23595_ (.A1(_14744_),
    .A2(net2136),
    .B(_14776_),
    .Y(_15200_));
 AND5x1_ASAP7_75t_R _23596_ (.A(_14882_),
    .B(_15199_),
    .C(_14888_),
    .D(_14889_),
    .E(_15200_),
    .Y(_15201_));
 AND3x1_ASAP7_75t_R _23597_ (.A(_15187_),
    .B(_15196_),
    .C(_15201_),
    .Y(_15202_));
 NAND2x2_ASAP7_75t_R _23598_ (.A(_15170_),
    .B(_15202_),
    .Y(_15203_));
 BUFx16f_ASAP7_75t_R load_slew394 (.A(_00528_),
    .Y(net394));
 XOR2x1_ASAP7_75t_R _23600_ (.A(_00391_),
    .Y(_15205_),
    .B(_00440_));
 XNOR2x2_ASAP7_75t_R _23601_ (.A(_00472_),
    .B(_00516_),
    .Y(_15206_));
 XNOR2x1_ASAP7_75t_R _23602_ (.B(_15206_),
    .Y(_15207_),
    .A(_15205_));
 XOR2x1_ASAP7_75t_R _23603_ (.A(_15203_),
    .Y(_15208_),
    .B(_15207_));
 AND2x2_ASAP7_75t_R _23604_ (.A(net405),
    .B(net4052),
    .Y(_15209_));
 AO21x1_ASAP7_75t_R _23605_ (.A1(_15208_),
    .A2(net399),
    .B(_15209_),
    .Y(_00356_));
 AO21x1_ASAP7_75t_R _23606_ (.A1(_14804_),
    .A2(_14805_),
    .B(_14610_),
    .Y(_15210_));
 AND5x1_ASAP7_75t_R _23607_ (.A(_14639_),
    .B(_14855_),
    .C(_15210_),
    .D(_14619_),
    .E(_14627_),
    .Y(_15211_));
 AO21x1_ASAP7_75t_R _23608_ (.A1(_14744_),
    .A2(net3509),
    .B(_14835_),
    .Y(_15212_));
 AO21x1_ASAP7_75t_R _23609_ (.A1(net2178),
    .A2(_14625_),
    .B(_14835_),
    .Y(_15213_));
 AO21x1_ASAP7_75t_R _23610_ (.A1(_14733_),
    .A2(net2179),
    .B(_14835_),
    .Y(_15214_));
 AND4x1_ASAP7_75t_R _23611_ (.A(_15212_),
    .B(_15184_),
    .C(_15213_),
    .D(_15214_),
    .Y(_15215_));
 AO21x1_ASAP7_75t_R _23612_ (.A1(_14919_),
    .A2(_14625_),
    .B(_14807_),
    .Y(_15216_));
 AO21x1_ASAP7_75t_R _23613_ (.A1(_14809_),
    .A2(net1943),
    .B(_14807_),
    .Y(_15217_));
 AO21x1_ASAP7_75t_R _23614_ (.A1(_14733_),
    .A2(_14804_),
    .B(_14807_),
    .Y(_15218_));
 AND4x1_ASAP7_75t_R _23615_ (.A(_14857_),
    .B(_15216_),
    .C(_15217_),
    .D(_15218_),
    .Y(_15219_));
 AO21x1_ASAP7_75t_R _23616_ (.A1(_14805_),
    .A2(_14860_),
    .B(_14816_),
    .Y(_15220_));
 OA211x2_ASAP7_75t_R _23617_ (.A1(_14652_),
    .A2(_14816_),
    .B(_15220_),
    .C(_14862_),
    .Y(_15221_));
 AND4x2_ASAP7_75t_R _23618_ (.A(_15211_),
    .B(_15215_),
    .C(_15219_),
    .D(_15221_),
    .Y(_15222_));
 NOR2x1_ASAP7_75t_R _23619_ (.A(_14764_),
    .B(_14776_),
    .Y(_15223_));
 INVx1_ASAP7_75t_R _23620_ (.A(_15223_),
    .Y(_15224_));
 AND3x1_ASAP7_75t_R _23621_ (.A(_15224_),
    .B(_15004_),
    .C(_14998_),
    .Y(_15225_));
 OA211x2_ASAP7_75t_R _23622_ (.A1(net2201),
    .A2(net3517),
    .B(_14761_),
    .C(net2721),
    .Y(_15226_));
 INVx1_ASAP7_75t_R _23623_ (.A(_15226_),
    .Y(_15227_));
 AO21x1_ASAP7_75t_R _23624_ (.A1(net3506),
    .A2(net2178),
    .B(_14768_),
    .Y(_15228_));
 AND5x1_ASAP7_75t_R _23625_ (.A(_15001_),
    .B(_15225_),
    .C(_15227_),
    .D(_14778_),
    .E(_15228_),
    .Y(_15229_));
 AO21x1_ASAP7_75t_R _23626_ (.A1(_14774_),
    .A2(_15042_),
    .B(_14783_),
    .Y(_15230_));
 AND3x1_ASAP7_75t_R _23627_ (.A(_15068_),
    .B(_15193_),
    .C(_15230_),
    .Y(_15231_));
 AO21x1_ASAP7_75t_R _23628_ (.A1(net2136),
    .A2(net3509),
    .B(_14793_),
    .Y(_15232_));
 NAND2x1_ASAP7_75t_R _23629_ (.A(_14635_),
    .B(_14792_),
    .Y(_15233_));
 AND5x1_ASAP7_75t_R _23630_ (.A(_14799_),
    .B(_14800_),
    .C(_15232_),
    .D(_14969_),
    .E(_15233_),
    .Y(_15234_));
 AND3x1_ASAP7_75t_R _23631_ (.A(_15229_),
    .B(_15231_),
    .C(_15234_),
    .Y(_15235_));
 NAND2x2_ASAP7_75t_R _23632_ (.A(_15222_),
    .B(_15235_),
    .Y(_15236_));
 OA21x2_ASAP7_75t_R _23633_ (.A1(_14922_),
    .A2(_14819_),
    .B(_14720_),
    .Y(_15237_));
 AO21x1_ASAP7_75t_R _23634_ (.A1(_14637_),
    .A2(_14720_),
    .B(_15237_),
    .Y(_15238_));
 NOR2x1_ASAP7_75t_R _23635_ (.A(_14716_),
    .B(_14725_),
    .Y(_15239_));
 OA21x2_ASAP7_75t_R _23636_ (.A1(_14618_),
    .A2(_14870_),
    .B(_14720_),
    .Y(_15240_));
 AO21x1_ASAP7_75t_R _23637_ (.A1(_14637_),
    .A2(_14729_),
    .B(_15033_),
    .Y(_15241_));
 AO21x1_ASAP7_75t_R _23638_ (.A1(_14910_),
    .A2(_14729_),
    .B(_15119_),
    .Y(_15242_));
 OR5x2_ASAP7_75t_R _23639_ (.A(_15238_),
    .B(_15239_),
    .C(_15240_),
    .D(_15241_),
    .E(_15242_),
    .Y(_15243_));
 AND3x1_ASAP7_75t_R _23640_ (.A(_14739_),
    .B(_00452_),
    .C(net1989),
    .Y(_15244_));
 AO21x1_ASAP7_75t_R _23641_ (.A1(_14870_),
    .A2(_14739_),
    .B(_15244_),
    .Y(_15245_));
 OA21x2_ASAP7_75t_R _23642_ (.A1(_14797_),
    .A2(_14732_),
    .B(_14704_),
    .Y(_15246_));
 NOR2x1_ASAP7_75t_R _23643_ (.A(_14809_),
    .B(_14712_),
    .Y(_15247_));
 AO21x1_ASAP7_75t_R _23644_ (.A1(_14648_),
    .A2(_14704_),
    .B(_15247_),
    .Y(_15248_));
 NAND2x1_ASAP7_75t_R _23645_ (.A(_15117_),
    .B(_14952_),
    .Y(_15249_));
 OR5x2_ASAP7_75t_R _23646_ (.A(_14746_),
    .B(_15245_),
    .C(_15246_),
    .D(_15248_),
    .E(_15249_),
    .Y(_15250_));
 NOR2x2_ASAP7_75t_R _23647_ (.A(_15243_),
    .B(_15250_),
    .Y(_15251_));
 AO21x1_ASAP7_75t_R _23648_ (.A1(_14733_),
    .A2(net1874),
    .B(_14668_),
    .Y(_15252_));
 OA211x2_ASAP7_75t_R _23649_ (.A1(net3510),
    .A2(_14668_),
    .B(_15252_),
    .C(_15020_),
    .Y(_15253_));
 NAND2x1_ASAP7_75t_R _23650_ (.A(_14653_),
    .B(_14647_),
    .Y(_15254_));
 AND5x1_ASAP7_75t_R _23651_ (.A(_15253_),
    .B(_15154_),
    .C(_14924_),
    .D(_15024_),
    .E(_15254_),
    .Y(_15255_));
 OA211x2_ASAP7_75t_R _23652_ (.A1(_14654_),
    .A2(_14686_),
    .B(_14908_),
    .C(_15103_),
    .Y(_15256_));
 AO21x1_ASAP7_75t_R _23653_ (.A1(_14804_),
    .A2(net1874),
    .B(_14694_),
    .Y(_15257_));
 AND3x1_ASAP7_75t_R _23654_ (.A(_15257_),
    .B(_14928_),
    .C(_15097_),
    .Y(_15258_));
 OA211x2_ASAP7_75t_R _23655_ (.A1(_14694_),
    .A2(net1943),
    .B(_15256_),
    .C(_15258_),
    .Y(_15259_));
 OA211x2_ASAP7_75t_R _23656_ (.A1(_14620_),
    .A2(net3516),
    .B(_14662_),
    .C(net3525),
    .Y(_15260_));
 INVx1_ASAP7_75t_R _23657_ (.A(_15260_),
    .Y(_15261_));
 NAND2x1_ASAP7_75t_R _23658_ (.A(_15035_),
    .B(_14662_),
    .Y(_15262_));
 AO21x1_ASAP7_75t_R _23659_ (.A1(_14733_),
    .A2(_14860_),
    .B(_14657_),
    .Y(_15263_));
 AND4x1_ASAP7_75t_R _23660_ (.A(_15261_),
    .B(_14664_),
    .C(_15262_),
    .D(_15263_),
    .Y(_15264_));
 AND3x1_ASAP7_75t_R _23661_ (.A(_15255_),
    .B(_15259_),
    .C(_15264_),
    .Y(_15265_));
 NAND2x2_ASAP7_75t_R _23662_ (.A(_15251_),
    .B(_15265_),
    .Y(_15266_));
 NOR2x2_ASAP7_75t_R _23663_ (.A(_15236_),
    .B(_15266_),
    .Y(_15267_));
 NAND2x2_ASAP7_75t_R _23664_ (.A(_14905_),
    .B(_15267_),
    .Y(_15268_));
 BUFx16f_ASAP7_75t_R load_slew393 (.A(net397),
    .Y(net393));
 XNOR2x1_ASAP7_75t_R _23666_ (.B(_00471_),
    .Y(_15270_),
    .A(_00439_));
 BUFx16f_ASAP7_75t_R load_slew392 (.A(net393),
    .Y(net392));
 XNOR2x2_ASAP7_75t_R _23668_ (.A(_00494_),
    .B(_00515_),
    .Y(_15272_));
 XNOR2x1_ASAP7_75t_R _23669_ (.B(_15272_),
    .Y(_15273_),
    .A(_15270_));
 XOR2x1_ASAP7_75t_R _23670_ (.A(_15268_),
    .Y(_15274_),
    .B(_15273_));
 NAND2x2_ASAP7_75t_R _23671_ (.A(net402),
    .B(net4036),
    .Y(_15275_));
 OAI21x1_ASAP7_75t_R _23672_ (.A1(net405),
    .A2(_15274_),
    .B(_15275_),
    .Y(_00357_));
 BUFx16f_ASAP7_75t_R load_slew391 (.A(net397),
    .Y(net391));
 XNOR2x1_ASAP7_75t_R _23674_ (.B(_00470_),
    .Y(_15277_),
    .A(_00438_));
 XNOR2x2_ASAP7_75t_R _23675_ (.A(_00493_),
    .B(_00514_),
    .Y(_15278_));
 XNOR2x1_ASAP7_75t_R _23676_ (.B(_15278_),
    .Y(_15279_),
    .A(_15277_));
 NOR2x1_ASAP7_75t_R _23677_ (.A(_14814_),
    .B(_14816_),
    .Y(_15280_));
 INVx1_ASAP7_75t_R _23678_ (.A(_15280_),
    .Y(_15281_));
 AND4x1_ASAP7_75t_R _23679_ (.A(_15281_),
    .B(_14823_),
    .C(_15077_),
    .D(_14862_),
    .Y(_15282_));
 NOR2x1_ASAP7_75t_R _23680_ (.A(_14805_),
    .B(_14835_),
    .Y(_15283_));
 NOR2x1_ASAP7_75t_R _23681_ (.A(_14631_),
    .B(_14835_),
    .Y(_15284_));
 OR4x1_ASAP7_75t_R _23682_ (.A(_15079_),
    .B(_15283_),
    .C(_15182_),
    .D(_15284_),
    .Y(_15285_));
 INVx1_ASAP7_75t_R _23683_ (.A(_15285_),
    .Y(_15286_));
 AO21x1_ASAP7_75t_R _23684_ (.A1(_14764_),
    .A2(net3537),
    .B(_14807_),
    .Y(_15287_));
 AO21x1_ASAP7_75t_R _23685_ (.A1(_14625_),
    .A2(_14860_),
    .B(_14807_),
    .Y(_15288_));
 AND3x1_ASAP7_75t_R _23686_ (.A(_15287_),
    .B(_15288_),
    .C(_15089_),
    .Y(_15289_));
 AND5x2_ASAP7_75t_R _23687_ (.A(_14640_),
    .B(_15282_),
    .C(_15286_),
    .D(_14987_),
    .E(_15289_),
    .Y(_15290_));
 AO21x1_ASAP7_75t_R _23688_ (.A1(_14926_),
    .A2(net2178),
    .B(_14776_),
    .Y(_15291_));
 INVx1_ASAP7_75t_R _23689_ (.A(_14886_),
    .Y(_15292_));
 AND3x1_ASAP7_75t_R _23690_ (.A(_15291_),
    .B(_14880_),
    .C(_15292_),
    .Y(_15293_));
 AND5x2_ASAP7_75t_R _23691_ (.A(_15063_),
    .B(_15293_),
    .C(_15066_),
    .D(_14760_),
    .E(_15002_),
    .Y(_15294_));
 INVx1_ASAP7_75t_R _23692_ (.A(_15188_),
    .Y(_15295_));
 AO21x1_ASAP7_75t_R _23693_ (.A1(_14654_),
    .A2(_14652_),
    .B(_14793_),
    .Y(_15296_));
 OA211x2_ASAP7_75t_R _23694_ (.A1(net3509),
    .A2(_14793_),
    .B(_15295_),
    .C(_15296_),
    .Y(_15297_));
 AO21x1_ASAP7_75t_R _23695_ (.A1(_14744_),
    .A2(net1830),
    .B(_14783_),
    .Y(_15298_));
 AO21x1_ASAP7_75t_R _23696_ (.A1(_14636_),
    .A2(_14654_),
    .B(_14783_),
    .Y(_15299_));
 NAND2x1_ASAP7_75t_R _23697_ (.A(_14782_),
    .B(_14670_),
    .Y(_15300_));
 NAND2x1_ASAP7_75t_R _23698_ (.A(_14782_),
    .B(_14661_),
    .Y(_15301_));
 AND5x1_ASAP7_75t_R _23699_ (.A(_15298_),
    .B(_15299_),
    .C(_14789_),
    .D(_15300_),
    .E(_15301_),
    .Y(_15302_));
 AND2x2_ASAP7_75t_R _23700_ (.A(_15297_),
    .B(_15302_),
    .Y(_15303_));
 NAND3x2_ASAP7_75t_R _23701_ (.B(_15294_),
    .C(_15303_),
    .Y(_15304_),
    .A(_15290_));
 OA21x2_ASAP7_75t_R _23702_ (.A1(_14692_),
    .A2(_14712_),
    .B(_15050_),
    .Y(_15305_));
 INVx1_ASAP7_75t_R _23703_ (.A(_15247_),
    .Y(_15306_));
 OA211x2_ASAP7_75t_R _23704_ (.A1(_14620_),
    .A2(_14672_),
    .B(_14739_),
    .C(_14630_),
    .Y(_15307_));
 INVx1_ASAP7_75t_R _23705_ (.A(_15307_),
    .Y(_15308_));
 AO21x1_ASAP7_75t_R _23706_ (.A1(net2179),
    .A2(net2178),
    .B(_14740_),
    .Y(_15309_));
 AND5x2_ASAP7_75t_R _23707_ (.A(_14706_),
    .B(_15305_),
    .C(_15306_),
    .D(_15308_),
    .E(_15309_),
    .Y(_15310_));
 AO21x1_ASAP7_75t_R _23708_ (.A1(_14744_),
    .A2(net3538),
    .B(_14694_),
    .Y(_15311_));
 AO21x1_ASAP7_75t_R _23709_ (.A1(_14654_),
    .A2(_14660_),
    .B(_14694_),
    .Y(_15312_));
 AND2x2_ASAP7_75t_R _23710_ (.A(_15311_),
    .B(_15312_),
    .Y(_15313_));
 AO21x1_ASAP7_75t_R _23711_ (.A1(_14926_),
    .A2(net3520),
    .B(_14694_),
    .Y(_15314_));
 AO21x1_ASAP7_75t_R _23712_ (.A1(net1874),
    .A2(_14860_),
    .B(_14694_),
    .Y(_15315_));
 AO21x1_ASAP7_75t_R _23713_ (.A1(_14654_),
    .A2(_14638_),
    .B(_14686_),
    .Y(_15316_));
 AO21x1_ASAP7_75t_R _23714_ (.A1(_14919_),
    .A2(_14667_),
    .B(_14686_),
    .Y(_15317_));
 AND5x1_ASAP7_75t_R _23715_ (.A(_15313_),
    .B(_15314_),
    .C(_15315_),
    .D(_15316_),
    .E(_15317_),
    .Y(_15318_));
 AND5x1_ASAP7_75t_R _23716_ (.A(_15252_),
    .B(_14920_),
    .C(_15023_),
    .D(_14649_),
    .E(_15254_),
    .Y(_15319_));
 AO21x1_ASAP7_75t_R _23717_ (.A1(_14728_),
    .A2(_14860_),
    .B(_14657_),
    .Y(_15320_));
 AO21x1_ASAP7_75t_R _23718_ (.A1(_14636_),
    .A2(_14654_),
    .B(_14657_),
    .Y(_15321_));
 INVx1_ASAP7_75t_R _23719_ (.A(_15146_),
    .Y(_15322_));
 AND5x1_ASAP7_75t_R _23720_ (.A(_15320_),
    .B(_15321_),
    .C(_14663_),
    .D(_15322_),
    .E(_14916_),
    .Y(_15323_));
 AND3x2_ASAP7_75t_R _23721_ (.A(_15318_),
    .B(_15319_),
    .C(_15323_),
    .Y(_15324_));
 AO21x1_ASAP7_75t_R _23722_ (.A1(_14654_),
    .A2(net1943),
    .B(_14730_),
    .Y(_15325_));
 AND3x1_ASAP7_75t_R _23723_ (.A(_15325_),
    .B(_15034_),
    .C(_15121_),
    .Y(_15326_));
 AO21x1_ASAP7_75t_R _23724_ (.A1(_14636_),
    .A2(net3509),
    .B(_14725_),
    .Y(_15327_));
 AO21x1_ASAP7_75t_R _23725_ (.A1(_14926_),
    .A2(net2178),
    .B(_14730_),
    .Y(_15328_));
 OA21x2_ASAP7_75t_R _23726_ (.A1(net2179),
    .A2(_14730_),
    .B(_15328_),
    .Y(_15329_));
 AO21x1_ASAP7_75t_R _23727_ (.A1(_14926_),
    .A2(_14919_),
    .B(_14725_),
    .Y(_15330_));
 AND5x2_ASAP7_75t_R _23728_ (.A(_14937_),
    .B(_15326_),
    .C(_15327_),
    .D(_15329_),
    .E(_15330_),
    .Y(_15331_));
 NAND3x2_ASAP7_75t_R _23729_ (.B(_15324_),
    .C(_15331_),
    .Y(_15332_),
    .A(_15310_));
 NOR2x2_ASAP7_75t_R _23730_ (.A(_15304_),
    .B(_15332_),
    .Y(_15333_));
 NAND2x2_ASAP7_75t_R _23731_ (.A(_14905_),
    .B(_15333_),
    .Y(_15334_));
 XNOR2x1_ASAP7_75t_R _23732_ (.B(_15334_),
    .Y(_15335_),
    .A(_15279_));
 AND2x2_ASAP7_75t_R _23733_ (.A(net402),
    .B(net4170),
    .Y(_15336_));
 AO21x1_ASAP7_75t_R _23734_ (.A1(_15335_),
    .A2(net398),
    .B(_15336_),
    .Y(_00358_));
 XNOR2x2_ASAP7_75t_R _23735_ (.A(_00469_),
    .B(_00513_),
    .Y(_15337_));
 BUFx16f_ASAP7_75t_R load_slew390 (.A(_18753_),
    .Y(net390));
 XOR2x1_ASAP7_75t_R _23737_ (.A(_00392_),
    .Y(_15339_),
    .B(_00437_));
 XOR2x1_ASAP7_75t_R _23738_ (.A(_15337_),
    .Y(_15340_),
    .B(_15339_));
 AO21x1_ASAP7_75t_R _23739_ (.A1(_14744_),
    .A2(net3509),
    .B(_14610_),
    .Y(_15341_));
 OA211x2_ASAP7_75t_R _23740_ (.A1(_14733_),
    .A2(_14610_),
    .B(_15177_),
    .C(_15341_),
    .Y(_15342_));
 OA211x2_ASAP7_75t_R _23741_ (.A1(_14835_),
    .A2(_14652_),
    .B(_15212_),
    .C(_14853_),
    .Y(_15343_));
 NAND2x1_ASAP7_75t_R _23742_ (.A(_14834_),
    .B(_14762_),
    .Y(_15344_));
 OA211x2_ASAP7_75t_R _23743_ (.A1(_14728_),
    .A2(_14835_),
    .B(_14989_),
    .C(_15344_),
    .Y(_15345_));
 AND3x1_ASAP7_75t_R _23744_ (.A(_15342_),
    .B(_15343_),
    .C(_15345_),
    .Y(_15346_));
 AO21x1_ASAP7_75t_R _23745_ (.A1(net3524),
    .A2(_14805_),
    .B(_14783_),
    .Y(_15347_));
 OA211x2_ASAP7_75t_R _23746_ (.A1(_14633_),
    .A2(_14783_),
    .B(_15347_),
    .C(_14979_),
    .Y(_15348_));
 AND3x1_ASAP7_75t_R _23747_ (.A(_14792_),
    .B(_14650_),
    .C(net2722),
    .Y(_15349_));
 NOR2x1_ASAP7_75t_R _23748_ (.A(_14897_),
    .B(_15349_),
    .Y(_15350_));
 AND3x1_ASAP7_75t_R _23749_ (.A(_15189_),
    .B(_15348_),
    .C(_15350_),
    .Y(_15351_));
 AO21x1_ASAP7_75t_R _23750_ (.A1(net3510),
    .A2(_14926_),
    .B(_14816_),
    .Y(_15352_));
 AO21x1_ASAP7_75t_R _23751_ (.A1(_14733_),
    .A2(_14804_),
    .B(_14816_),
    .Y(_15353_));
 AND4x1_ASAP7_75t_R _23752_ (.A(_14865_),
    .B(_15352_),
    .C(_15353_),
    .D(_15281_),
    .Y(_15354_));
 AND4x1_ASAP7_75t_R _23753_ (.A(_14811_),
    .B(_14810_),
    .C(_15287_),
    .D(_15090_),
    .Y(_15355_));
 AND2x2_ASAP7_75t_R _23754_ (.A(_15354_),
    .B(_15355_),
    .Y(_15356_));
 AO21x1_ASAP7_75t_R _23755_ (.A1(_14926_),
    .A2(net3511),
    .B(_14776_),
    .Y(_15357_));
 AO21x1_ASAP7_75t_R _23756_ (.A1(net2179),
    .A2(net1874),
    .B(_14776_),
    .Y(_15358_));
 AND4x1_ASAP7_75t_R _23757_ (.A(_15357_),
    .B(_15358_),
    .C(_15224_),
    .D(_14884_),
    .Y(_15359_));
 AO21x1_ASAP7_75t_R _23758_ (.A1(_14636_),
    .A2(net1943),
    .B(_14768_),
    .Y(_15360_));
 AO21x1_ASAP7_75t_R _23759_ (.A1(net1830),
    .A2(net2136),
    .B(_14768_),
    .Y(_15361_));
 INVx1_ASAP7_75t_R _23760_ (.A(_14875_),
    .Y(_15362_));
 AND5x1_ASAP7_75t_R _23761_ (.A(_15000_),
    .B(_15360_),
    .C(_15361_),
    .D(_15362_),
    .E(_14763_),
    .Y(_15363_));
 AND5x2_ASAP7_75t_R _23762_ (.A(_15346_),
    .B(_15351_),
    .C(_15356_),
    .D(_15359_),
    .E(_15363_),
    .Y(_15364_));
 OA211x2_ASAP7_75t_R _23763_ (.A1(_14620_),
    .A2(_14672_),
    .B(_14704_),
    .C(_14630_),
    .Y(_15365_));
 INVx1_ASAP7_75t_R _23764_ (.A(_15365_),
    .Y(_15366_));
 AND5x1_ASAP7_75t_R _23765_ (.A(_15306_),
    .B(_15366_),
    .C(_14709_),
    .D(_14948_),
    .E(_15124_),
    .Y(_15367_));
 OA211x2_ASAP7_75t_R _23766_ (.A1(net2199),
    .A2(_00452_),
    .B(_14739_),
    .C(_14637_),
    .Y(_15368_));
 INVx1_ASAP7_75t_R _23767_ (.A(_15368_),
    .Y(_15369_));
 NOR2x1_ASAP7_75t_R _23768_ (.A(_14748_),
    .B(_15244_),
    .Y(_15370_));
 AND3x1_ASAP7_75t_R _23769_ (.A(_15369_),
    .B(_14952_),
    .C(_15370_),
    .Y(_15371_));
 AO21x1_ASAP7_75t_R _23770_ (.A1(_15035_),
    .A2(_14720_),
    .B(_15237_),
    .Y(_15372_));
 INVx1_ASAP7_75t_R _23771_ (.A(_15372_),
    .Y(_15373_));
 INVx1_ASAP7_75t_R _23772_ (.A(_15239_),
    .Y(_15374_));
 AND3x1_ASAP7_75t_R _23773_ (.A(_14936_),
    .B(_15133_),
    .C(_15374_),
    .Y(_15375_));
 OA211x2_ASAP7_75t_R _23774_ (.A1(_14654_),
    .A2(_14725_),
    .B(_15373_),
    .C(_15375_),
    .Y(_15376_));
 OA211x2_ASAP7_75t_R _23775_ (.A1(net2199),
    .A2(_14672_),
    .B(_14729_),
    .C(_14605_),
    .Y(_15377_));
 NOR2x1_ASAP7_75t_R _23776_ (.A(_15119_),
    .B(_15377_),
    .Y(_15378_));
 OA211x2_ASAP7_75t_R _23777_ (.A1(_14652_),
    .A2(_14730_),
    .B(_15378_),
    .C(_15034_),
    .Y(_15379_));
 AND4x1_ASAP7_75t_R _23778_ (.A(_15367_),
    .B(_15371_),
    .C(_15376_),
    .D(_15379_),
    .Y(_15380_));
 AO21x1_ASAP7_75t_R _23779_ (.A1(net3509),
    .A2(net2136),
    .B(_14686_),
    .Y(_15381_));
 AO21x1_ASAP7_75t_R _23780_ (.A1(net1819),
    .A2(net3520),
    .B(_14694_),
    .Y(_15382_));
 OA211x2_ASAP7_75t_R _23781_ (.A1(net1830),
    .A2(_14694_),
    .B(_15312_),
    .C(_15382_),
    .Y(_15383_));
 AO21x1_ASAP7_75t_R _23782_ (.A1(_14804_),
    .A2(net1874),
    .B(_14686_),
    .Y(_15384_));
 AO21x1_ASAP7_75t_R _23783_ (.A1(_14636_),
    .A2(net1943),
    .B(_14686_),
    .Y(_15385_));
 AND5x1_ASAP7_75t_R _23784_ (.A(_15381_),
    .B(_15383_),
    .C(_15103_),
    .D(_15384_),
    .E(_15385_),
    .Y(_15386_));
 AO221x1_ASAP7_75t_R _23785_ (.A1(_14620_),
    .A2(_14672_),
    .B1(_14728_),
    .B2(_14606_),
    .C(_14668_),
    .Y(_15387_));
 AO21x1_ASAP7_75t_R _23786_ (.A1(_14733_),
    .A2(net3506),
    .B(_14657_),
    .Y(_15388_));
 AND5x1_ASAP7_75t_R _23787_ (.A(_14675_),
    .B(_15387_),
    .C(_15388_),
    .D(_15254_),
    .E(_15321_),
    .Y(_15389_));
 AND3x1_ASAP7_75t_R _23788_ (.A(_15380_),
    .B(_15386_),
    .C(_15389_),
    .Y(_15390_));
 NAND2x2_ASAP7_75t_R _23789_ (.A(_15364_),
    .B(_15390_),
    .Y(_15391_));
 XNOR2x1_ASAP7_75t_R _23790_ (.B(_15391_),
    .Y(_15392_),
    .A(_15340_));
 BUFx16f_ASAP7_75t_R wire389 (.A(net390),
    .Y(net389));
 BUFx16f_ASAP7_75t_R load_slew388 (.A(_18753_),
    .Y(net388));
 AND2x2_ASAP7_75t_R _23793_ (.A(net402),
    .B(net4156),
    .Y(_15395_));
 AO21x1_ASAP7_75t_R _23794_ (.A1(_15392_),
    .A2(net398),
    .B(_15395_),
    .Y(_00359_));
 INVx3_ASAP7_75t_R _23795_ (.A(net3967),
    .Y(_15396_));
 NOR2x2_ASAP7_75t_R _23796_ (.A(_00443_),
    .B(net3548),
    .Y(_15397_));
 NOR2x2_ASAP7_75t_R _23797_ (.A(_00441_),
    .B(_00442_),
    .Y(_15398_));
 AND2x6_ASAP7_75t_R _23798_ (.A(_15397_),
    .B(_15398_),
    .Y(_15399_));
 INVx4_ASAP7_75t_R _23799_ (.A(_00440_),
    .Y(_15400_));
 NAND2x2_ASAP7_75t_R _23800_ (.A(_00439_),
    .B(_15400_),
    .Y(_15401_));
 INVx4_ASAP7_75t_R _23801_ (.A(_00438_),
    .Y(_15402_));
 NAND2x2_ASAP7_75t_R _23802_ (.A(_00437_),
    .B(_15402_),
    .Y(_15403_));
 NOR2x2_ASAP7_75t_R _23803_ (.A(_15401_),
    .B(_15403_),
    .Y(_15404_));
 BUFx2_ASAP7_75t_R output387 (.A(net387),
    .Y(text_out[9]));
 AND2x2_ASAP7_75t_R _23805_ (.A(_15399_),
    .B(_15404_),
    .Y(_15406_));
 BUFx2_ASAP7_75t_R output386 (.A(net386),
    .Y(text_out[99]));
 AND2x6_ASAP7_75t_R _23807_ (.A(net3546),
    .B(net3551),
    .Y(_15408_));
 NAND2x2_ASAP7_75t_R _23808_ (.A(_15398_),
    .B(_15408_),
    .Y(_15409_));
 NOR2x2_ASAP7_75t_R _23809_ (.A(_00439_),
    .B(_00440_),
    .Y(_15410_));
 CKINVDCx5p33_ASAP7_75t_R _23810_ (.A(_00437_),
    .Y(_15411_));
 AND3x4_ASAP7_75t_R _23811_ (.A(_15410_),
    .B(_15411_),
    .C(_00438_),
    .Y(_15412_));
 INVx5_ASAP7_75t_R _23812_ (.A(_15412_),
    .Y(_15413_));
 NOR2x1_ASAP7_75t_R _23813_ (.A(_15409_),
    .B(_15413_),
    .Y(_15414_));
 NAND2x2_ASAP7_75t_R _23814_ (.A(_00441_),
    .B(_00442_),
    .Y(_15415_));
 CKINVDCx8_ASAP7_75t_R _23815_ (.A(_15415_),
    .Y(_15416_));
 NAND2x2_ASAP7_75t_R _23816_ (.A(_15408_),
    .B(_15416_),
    .Y(_15417_));
 NAND2x2_ASAP7_75t_R _23817_ (.A(_00439_),
    .B(_00440_),
    .Y(_15418_));
 NAND2x2_ASAP7_75t_R _23818_ (.A(_00438_),
    .B(_15411_),
    .Y(_15419_));
 NOR2x2_ASAP7_75t_R _23819_ (.A(_15418_),
    .B(_15419_),
    .Y(_15420_));
 INVx5_ASAP7_75t_R _23820_ (.A(_15420_),
    .Y(_15421_));
 NOR2x1_ASAP7_75t_R _23821_ (.A(_15417_),
    .B(_15421_),
    .Y(_15422_));
 NAND2x2_ASAP7_75t_R _23822_ (.A(_00437_),
    .B(_00438_),
    .Y(_15423_));
 NOR2x2_ASAP7_75t_R _23823_ (.A(_15418_),
    .B(_15423_),
    .Y(_15424_));
 CKINVDCx20_ASAP7_75t_R _23824_ (.A(net3544),
    .Y(_15425_));
 BUFx2_ASAP7_75t_R output385 (.A(net385),
    .Y(text_out[98]));
 INVx3_ASAP7_75t_R _23826_ (.A(_00442_),
    .Y(_15427_));
 NAND2x2_ASAP7_75t_R _23827_ (.A(_00441_),
    .B(_15427_),
    .Y(_15428_));
 CKINVDCx9p33_ASAP7_75t_R _23828_ (.A(_15428_),
    .Y(_15429_));
 BUFx2_ASAP7_75t_R output384 (.A(net384),
    .Y(text_out[97]));
 AND3x1_ASAP7_75t_R _23830_ (.A(_15424_),
    .B(_15425_),
    .C(_15429_),
    .Y(_15431_));
 CKINVDCx9p33_ASAP7_75t_R _23831_ (.A(net3548),
    .Y(_15432_));
 INVx3_ASAP7_75t_R _23832_ (.A(_00441_),
    .Y(_15433_));
 NAND2x2_ASAP7_75t_R _23833_ (.A(_00442_),
    .B(_15433_),
    .Y(_15434_));
 INVx5_ASAP7_75t_R _23834_ (.A(net3553),
    .Y(_15435_));
 NAND2x2_ASAP7_75t_R _23835_ (.A(_15432_),
    .B(_15435_),
    .Y(_15436_));
 INVx4_ASAP7_75t_R _23836_ (.A(_15404_),
    .Y(_15437_));
 BUFx2_ASAP7_75t_R output383 (.A(net383),
    .Y(text_out[96]));
 NOR2x1_ASAP7_75t_R _23838_ (.A(_15436_),
    .B(_15437_),
    .Y(_15439_));
 OR4x1_ASAP7_75t_R _23839_ (.A(_15414_),
    .B(_15422_),
    .C(_15431_),
    .D(_15439_),
    .Y(_15440_));
 NAND2x2_ASAP7_75t_R _23840_ (.A(_00444_),
    .B(_15425_),
    .Y(_15441_));
 CKINVDCx8_ASAP7_75t_R _23841_ (.A(_15398_),
    .Y(_15442_));
 NOR2x2_ASAP7_75t_R _23842_ (.A(_15441_),
    .B(_15442_),
    .Y(_15443_));
 NOR2x1_ASAP7_75t_R _23843_ (.A(_00437_),
    .B(_00438_),
    .Y(_15444_));
 AND2x6_ASAP7_75t_R _23844_ (.A(_15444_),
    .B(_15410_),
    .Y(_15445_));
 BUFx2_ASAP7_75t_R output382 (.A(net382),
    .Y(text_out[95]));
 NAND2x2_ASAP7_75t_R _23846_ (.A(_15443_),
    .B(_15445_),
    .Y(_15447_));
 NAND2x2_ASAP7_75t_R _23847_ (.A(_15408_),
    .B(_15429_),
    .Y(_15448_));
 INVx4_ASAP7_75t_R _23848_ (.A(_15448_),
    .Y(_15449_));
 NAND2x1_ASAP7_75t_R _23849_ (.A(_15445_),
    .B(_15449_),
    .Y(_15450_));
 NAND2x1_ASAP7_75t_R _23850_ (.A(_15447_),
    .B(_15450_),
    .Y(_15451_));
 NOR2x2_ASAP7_75t_R _23851_ (.A(_00438_),
    .B(_15411_),
    .Y(_15452_));
 NAND2x2_ASAP7_75t_R _23852_ (.A(_15410_),
    .B(_15452_),
    .Y(_15453_));
 CKINVDCx5p33_ASAP7_75t_R _23853_ (.A(_15453_),
    .Y(_15454_));
 NAND2x1_ASAP7_75t_R _23854_ (.A(_15429_),
    .B(_15454_),
    .Y(_15455_));
 NOR2x1_ASAP7_75t_R _23855_ (.A(net3551),
    .B(_15455_),
    .Y(_15456_));
 INVx2_ASAP7_75t_R _23856_ (.A(_00439_),
    .Y(_15457_));
 NAND2x2_ASAP7_75t_R _23857_ (.A(_00440_),
    .B(_15457_),
    .Y(_15458_));
 NAND2x2_ASAP7_75t_R _23858_ (.A(_15411_),
    .B(_15402_),
    .Y(_15459_));
 NOR2x2_ASAP7_75t_R _23859_ (.A(_15458_),
    .B(_15459_),
    .Y(_15460_));
 BUFx2_ASAP7_75t_R output381 (.A(net381),
    .Y(text_out[94]));
 NOR2x2_ASAP7_75t_R _23861_ (.A(net3548),
    .B(_15425_),
    .Y(_15462_));
 NOR2x1_ASAP7_75t_R _23862_ (.A(_15415_),
    .B(_15462_),
    .Y(_15463_));
 AND3x1_ASAP7_75t_R _23863_ (.A(_15460_),
    .B(_15463_),
    .C(_15441_),
    .Y(_15464_));
 OR5x1_ASAP7_75t_R _23864_ (.A(_15406_),
    .B(_15440_),
    .C(_15451_),
    .D(_15456_),
    .E(_15464_),
    .Y(_15465_));
 INVx1_ASAP7_75t_R _23865_ (.A(_15465_),
    .Y(_15466_));
 NAND2x2_ASAP7_75t_R _23866_ (.A(net3546),
    .B(_15432_),
    .Y(_15467_));
 NOR2x2_ASAP7_75t_R _23867_ (.A(_15467_),
    .B(net3553),
    .Y(_15468_));
 CKINVDCx9p33_ASAP7_75t_R _23868_ (.A(_15468_),
    .Y(_15469_));
 BUFx2_ASAP7_75t_R output380 (.A(net380),
    .Y(text_out[93]));
 BUFx2_ASAP7_75t_R output379 (.A(net379),
    .Y(text_out[92]));
 NOR2x2_ASAP7_75t_R _23871_ (.A(net3544),
    .B(net3553),
    .Y(_15472_));
 INVx5_ASAP7_75t_R _23872_ (.A(_15472_),
    .Y(_15473_));
 BUFx2_ASAP7_75t_R output378 (.A(net378),
    .Y(text_out[91]));
 NOR2x2_ASAP7_75t_R _23874_ (.A(_15423_),
    .B(_15458_),
    .Y(_15475_));
 INVx6_ASAP7_75t_R _23875_ (.A(_15475_),
    .Y(_15476_));
 BUFx2_ASAP7_75t_R output377 (.A(net377),
    .Y(text_out[90]));
 AO21x1_ASAP7_75t_R _23877_ (.A1(_15469_),
    .A2(_15473_),
    .B(_15476_),
    .Y(_15478_));
 INVx5_ASAP7_75t_R _23878_ (.A(_15441_),
    .Y(_15479_));
 NOR2x2_ASAP7_75t_R _23879_ (.A(_15442_),
    .B(_15479_),
    .Y(_15480_));
 NOR2x2_ASAP7_75t_R _23880_ (.A(_15419_),
    .B(_15458_),
    .Y(_15481_));
 OA21x2_ASAP7_75t_R _23881_ (.A1(_15480_),
    .A2(_15468_),
    .B(_15481_),
    .Y(_15482_));
 CKINVDCx8_ASAP7_75t_R _23882_ (.A(_15399_),
    .Y(_15483_));
 AND3x4_ASAP7_75t_R _23883_ (.A(_15410_),
    .B(_00437_),
    .C(_00438_),
    .Y(_15484_));
 BUFx2_ASAP7_75t_R output376 (.A(net376),
    .Y(text_out[8]));
 INVx5_ASAP7_75t_R _23885_ (.A(_15484_),
    .Y(_15486_));
 BUFx2_ASAP7_75t_R output375 (.A(net375),
    .Y(text_out[89]));
 NOR2x1_ASAP7_75t_R _23887_ (.A(_15483_),
    .B(_15486_),
    .Y(_15488_));
 NOR2x1_ASAP7_75t_R _23888_ (.A(_15482_),
    .B(_15488_),
    .Y(_15489_));
 CKINVDCx5p33_ASAP7_75t_R _23889_ (.A(_15460_),
    .Y(_15490_));
 BUFx2_ASAP7_75t_R output374 (.A(net374),
    .Y(text_out[88]));
 OR3x1_ASAP7_75t_R _23891_ (.A(_15490_),
    .B(_15462_),
    .C(net3553),
    .Y(_15492_));
 NOR2x2_ASAP7_75t_R _23892_ (.A(net3556),
    .B(_15479_),
    .Y(_15493_));
 BUFx2_ASAP7_75t_R output373 (.A(net373),
    .Y(text_out[87]));
 NAND2x1_ASAP7_75t_R _23894_ (.A(_15493_),
    .B(_15412_),
    .Y(_15495_));
 NAND2x2_ASAP7_75t_R _23895_ (.A(_15462_),
    .B(_15416_),
    .Y(_15496_));
 BUFx2_ASAP7_75t_R output372 (.A(net372),
    .Y(text_out[86]));
 NOR2x2_ASAP7_75t_R _23897_ (.A(_15419_),
    .B(_15401_),
    .Y(_15498_));
 CKINVDCx5p33_ASAP7_75t_R _23898_ (.A(_15498_),
    .Y(_15499_));
 BUFx2_ASAP7_75t_R output371 (.A(net371),
    .Y(text_out[85]));
 NOR2x1_ASAP7_75t_R _23900_ (.A(_15496_),
    .B(_15499_),
    .Y(_15501_));
 NOR2x2_ASAP7_75t_R _23901_ (.A(_15423_),
    .B(_15401_),
    .Y(_15502_));
 CKINVDCx5p33_ASAP7_75t_R _23902_ (.A(_15502_),
    .Y(_15503_));
 NOR2x2_ASAP7_75t_R _23903_ (.A(_15428_),
    .B(_15441_),
    .Y(_15504_));
 INVx8_ASAP7_75t_R _23904_ (.A(_15504_),
    .Y(_15505_));
 NOR2x1_ASAP7_75t_R _23905_ (.A(_15503_),
    .B(_15505_),
    .Y(_15506_));
 NOR2x1_ASAP7_75t_R _23906_ (.A(_15501_),
    .B(_15506_),
    .Y(_15507_));
 AND5x1_ASAP7_75t_R _23907_ (.A(_15478_),
    .B(_15489_),
    .C(_15492_),
    .D(_15495_),
    .E(_15507_),
    .Y(_15508_));
 NOR2x2_ASAP7_75t_R _23908_ (.A(_15418_),
    .B(_15403_),
    .Y(_15509_));
 CKINVDCx6p67_ASAP7_75t_R _23909_ (.A(_15509_),
    .Y(_15510_));
 BUFx2_ASAP7_75t_R output370 (.A(net370),
    .Y(text_out[84]));
 NOR2x1_ASAP7_75t_R _23911_ (.A(net3553),
    .B(_15510_),
    .Y(_15512_));
 INVx1_ASAP7_75t_R _23912_ (.A(_15512_),
    .Y(_15513_));
 NOR2x2_ASAP7_75t_R _23913_ (.A(_15467_),
    .B(_15442_),
    .Y(_15514_));
 INVx8_ASAP7_75t_R _23914_ (.A(_15514_),
    .Y(_15515_));
 NAND2x2_ASAP7_75t_R _23915_ (.A(_15398_),
    .B(_15479_),
    .Y(_15516_));
 AO21x1_ASAP7_75t_R _23916_ (.A1(_15515_),
    .A2(_15516_),
    .B(_15510_),
    .Y(_15517_));
 NOR2x1_ASAP7_75t_R _23917_ (.A(_15409_),
    .B(_15510_),
    .Y(_15518_));
 INVx1_ASAP7_75t_R _23918_ (.A(_15518_),
    .Y(_15519_));
 OA211x2_ASAP7_75t_R _23919_ (.A1(net3547),
    .A2(_15513_),
    .B(_15517_),
    .C(_15519_),
    .Y(_15520_));
 BUFx2_ASAP7_75t_R output369 (.A(net369),
    .Y(text_out[83]));
 AND3x1_ASAP7_75t_R _23921_ (.A(_15484_),
    .B(_15432_),
    .C(_15416_),
    .Y(_15522_));
 NOR2x2_ASAP7_75t_R _23922_ (.A(_00439_),
    .B(_15400_),
    .Y(_15523_));
 NAND2x2_ASAP7_75t_R _23923_ (.A(_15452_),
    .B(_15523_),
    .Y(_15524_));
 NOR2x1_ASAP7_75t_R _23924_ (.A(_15524_),
    .B(_15516_),
    .Y(_15525_));
 AND3x1_ASAP7_75t_R _23925_ (.A(_15420_),
    .B(_15462_),
    .C(_15435_),
    .Y(_15526_));
 NOR2x2_ASAP7_75t_R _23926_ (.A(_15415_),
    .B(_15441_),
    .Y(_15527_));
 INVx5_ASAP7_75t_R _23927_ (.A(_15527_),
    .Y(_15528_));
 NOR2x1_ASAP7_75t_R _23928_ (.A(_15528_),
    .B(_15486_),
    .Y(_15529_));
 OR4x1_ASAP7_75t_R _23929_ (.A(_15522_),
    .B(_15525_),
    .C(_15526_),
    .D(_15529_),
    .Y(_15530_));
 INVx1_ASAP7_75t_R _23930_ (.A(_15530_),
    .Y(_15531_));
 AND3x1_ASAP7_75t_R _23931_ (.A(_15508_),
    .B(_15520_),
    .C(_15531_),
    .Y(_15532_));
 NAND2x2_ASAP7_75t_R _23932_ (.A(_15425_),
    .B(_15429_),
    .Y(_15533_));
 NOR2x1_ASAP7_75t_R _23933_ (.A(_15533_),
    .B(_15437_),
    .Y(_15534_));
 INVx1_ASAP7_75t_R _23934_ (.A(_15534_),
    .Y(_15535_));
 NOR2x2_ASAP7_75t_R _23935_ (.A(_15425_),
    .B(net3559),
    .Y(_15536_));
 INVx1_ASAP7_75t_R _23936_ (.A(_15536_),
    .Y(_15537_));
 AND3x1_ASAP7_75t_R _23937_ (.A(_15424_),
    .B(_15429_),
    .C(_15462_),
    .Y(_15538_));
 INVx1_ASAP7_75t_R _23938_ (.A(_15538_),
    .Y(_15539_));
 NAND2x2_ASAP7_75t_R _23939_ (.A(_15425_),
    .B(_15416_),
    .Y(_15540_));
 INVx4_ASAP7_75t_R _23940_ (.A(_15445_),
    .Y(_15541_));
 NOR2x1_ASAP7_75t_R _23941_ (.A(_15540_),
    .B(_15541_),
    .Y(_15542_));
 INVx1_ASAP7_75t_R _23942_ (.A(_15542_),
    .Y(_15543_));
 OA211x2_ASAP7_75t_R _23943_ (.A1(_15490_),
    .A2(_15537_),
    .B(_15539_),
    .C(_15543_),
    .Y(_15544_));
 BUFx2_ASAP7_75t_R output368 (.A(net368),
    .Y(text_out[82]));
 OR3x1_ASAP7_75t_R _23945_ (.A(_15413_),
    .B(_15462_),
    .C(net3561),
    .Y(_15546_));
 BUFx2_ASAP7_75t_R output367 (.A(net367),
    .Y(text_out[81]));
 INVx4_ASAP7_75t_R _23947_ (.A(_15397_),
    .Y(_15548_));
 NOR2x2_ASAP7_75t_R _23948_ (.A(net3553),
    .B(_15548_),
    .Y(_15549_));
 INVx5_ASAP7_75t_R _23949_ (.A(_15549_),
    .Y(_15550_));
 BUFx2_ASAP7_75t_R output366 (.A(net366),
    .Y(text_out[80]));
 NOR2x2_ASAP7_75t_R _23951_ (.A(_15401_),
    .B(_15459_),
    .Y(_15552_));
 BUFx2_ASAP7_75t_R output365 (.A(net365),
    .Y(text_out[7]));
 NAND2x1_ASAP7_75t_R _23953_ (.A(_15527_),
    .B(_15552_),
    .Y(_15554_));
 OA21x2_ASAP7_75t_R _23954_ (.A1(_15421_),
    .A2(_15550_),
    .B(_15554_),
    .Y(_15555_));
 BUFx2_ASAP7_75t_R output364 (.A(net364),
    .Y(text_out[79]));
 NOR2x1_ASAP7_75t_R _23956_ (.A(_15476_),
    .B(_15505_),
    .Y(_15557_));
 BUFx2_ASAP7_75t_R output363 (.A(net363),
    .Y(text_out[78]));
 AND2x2_ASAP7_75t_R _23958_ (.A(_15514_),
    .B(_15552_),
    .Y(_15559_));
 NOR2x1_ASAP7_75t_R _23959_ (.A(_15557_),
    .B(_15559_),
    .Y(_15560_));
 AND5x1_ASAP7_75t_R _23960_ (.A(_15535_),
    .B(_15544_),
    .C(_15546_),
    .D(_15555_),
    .E(_15560_),
    .Y(_15561_));
 AND3x1_ASAP7_75t_R _23961_ (.A(_15466_),
    .B(_15532_),
    .C(_15561_),
    .Y(_15562_));
 INVx8_ASAP7_75t_R _23962_ (.A(_15424_),
    .Y(_15563_));
 NOR2x1_ASAP7_75t_R _23963_ (.A(_15540_),
    .B(_15563_),
    .Y(_15564_));
 INVx1_ASAP7_75t_R _23964_ (.A(_15564_),
    .Y(_15565_));
 AO21x1_ASAP7_75t_R _23965_ (.A1(net3563),
    .A2(_15515_),
    .B(_15486_),
    .Y(_15566_));
 NOR2x2_ASAP7_75t_R _23966_ (.A(_15415_),
    .B(_15479_),
    .Y(_15567_));
 NAND2x1_ASAP7_75t_R _23967_ (.A(_15567_),
    .B(_15454_),
    .Y(_15568_));
 NAND2x1_ASAP7_75t_R _23968_ (.A(_15527_),
    .B(_15502_),
    .Y(_15569_));
 NOR2x2_ASAP7_75t_R _23969_ (.A(_15415_),
    .B(_15548_),
    .Y(_15570_));
 CKINVDCx8_ASAP7_75t_R _23970_ (.A(_15570_),
    .Y(_15571_));
 NOR2x1_ASAP7_75t_R _23971_ (.A(_15503_),
    .B(_15571_),
    .Y(_15572_));
 INVx1_ASAP7_75t_R _23972_ (.A(_15572_),
    .Y(_15573_));
 AND5x1_ASAP7_75t_R _23973_ (.A(_15565_),
    .B(_15566_),
    .C(_15568_),
    .D(_15569_),
    .E(_15573_),
    .Y(_15574_));
 NAND2x2_ASAP7_75t_R _23974_ (.A(_15408_),
    .B(_15435_),
    .Y(_15575_));
 INVx2_ASAP7_75t_R _23975_ (.A(_15575_),
    .Y(_15576_));
 NAND2x1_ASAP7_75t_R _23976_ (.A(_15576_),
    .B(_15484_),
    .Y(_15577_));
 NOR2x1_ASAP7_75t_R _23977_ (.A(_15496_),
    .B(_15510_),
    .Y(_15578_));
 INVx1_ASAP7_75t_R _23978_ (.A(_15578_),
    .Y(_15579_));
 NAND2x1_ASAP7_75t_R _23979_ (.A(_15424_),
    .B(_15443_),
    .Y(_15580_));
 NAND2x1_ASAP7_75t_R _23980_ (.A(_15527_),
    .B(_15498_),
    .Y(_15581_));
 AND4x1_ASAP7_75t_R _23981_ (.A(_15577_),
    .B(_15579_),
    .C(_15580_),
    .D(_15581_),
    .Y(_15582_));
 NOR2x2_ASAP7_75t_R _23982_ (.A(_15428_),
    .B(_15467_),
    .Y(_15583_));
 CKINVDCx9p33_ASAP7_75t_R _23983_ (.A(_15583_),
    .Y(_15584_));
 BUFx2_ASAP7_75t_R output362 (.A(net362),
    .Y(text_out[77]));
 BUFx2_ASAP7_75t_R output361 (.A(net361),
    .Y(text_out[76]));
 BUFx2_ASAP7_75t_R output360 (.A(net360),
    .Y(text_out[75]));
 AO21x1_ASAP7_75t_R _23987_ (.A1(_15483_),
    .A2(net3562),
    .B(_15476_),
    .Y(_15588_));
 NAND2x1_ASAP7_75t_R _23988_ (.A(_15502_),
    .B(_15583_),
    .Y(_15589_));
 OA211x2_ASAP7_75t_R _23989_ (.A1(_15584_),
    .A2(_15476_),
    .B(_15588_),
    .C(_15589_),
    .Y(_15590_));
 NAND2x1_ASAP7_75t_R _23990_ (.A(_15424_),
    .B(_15514_),
    .Y(_15591_));
 NAND2x1_ASAP7_75t_R _23991_ (.A(_15509_),
    .B(_15449_),
    .Y(_15592_));
 NOR2x1_ASAP7_75t_R _23992_ (.A(_15496_),
    .B(_15524_),
    .Y(_15593_));
 INVx1_ASAP7_75t_R _23993_ (.A(_15593_),
    .Y(_15594_));
 INVx3_ASAP7_75t_R _23994_ (.A(_15496_),
    .Y(_15595_));
 NAND2x1_ASAP7_75t_R _23995_ (.A(_15445_),
    .B(_15595_),
    .Y(_15596_));
 INVx3_ASAP7_75t_R _23996_ (.A(_15524_),
    .Y(_15597_));
 NAND2x1_ASAP7_75t_R _23997_ (.A(_15570_),
    .B(_15597_),
    .Y(_15598_));
 AND5x1_ASAP7_75t_R _23998_ (.A(_15591_),
    .B(_15592_),
    .C(_15594_),
    .D(_15596_),
    .E(_15598_),
    .Y(_15599_));
 AND4x1_ASAP7_75t_R _23999_ (.A(_15574_),
    .B(_15582_),
    .C(_15590_),
    .D(_15599_),
    .Y(_15600_));
 BUFx2_ASAP7_75t_R output359 (.A(net359),
    .Y(text_out[74]));
 NOR2x2_ASAP7_75t_R _24001_ (.A(_15418_),
    .B(_15459_),
    .Y(_15602_));
 INVx4_ASAP7_75t_R _24002_ (.A(_15602_),
    .Y(_15603_));
 AO21x1_ASAP7_75t_R _24003_ (.A1(_15515_),
    .A2(net3562),
    .B(_15603_),
    .Y(_15604_));
 BUFx2_ASAP7_75t_R output358 (.A(net358),
    .Y(text_out[73]));
 AO21x1_ASAP7_75t_R _24005_ (.A1(_15516_),
    .A2(_15436_),
    .B(_15603_),
    .Y(_15606_));
 NAND2x2_ASAP7_75t_R _24006_ (.A(_15432_),
    .B(_15398_),
    .Y(_15607_));
 NAND2x2_ASAP7_75t_R _24007_ (.A(_15425_),
    .B(_15398_),
    .Y(_15608_));
 AO21x1_ASAP7_75t_R _24008_ (.A1(_15607_),
    .A2(_15608_),
    .B(_15421_),
    .Y(_15609_));
 BUFx2_ASAP7_75t_R output357 (.A(net357),
    .Y(text_out[72]));
 NAND2x1_ASAP7_75t_R _24010_ (.A(net3540),
    .B(_15484_),
    .Y(_15611_));
 INVx3_ASAP7_75t_R _24011_ (.A(_15417_),
    .Y(_15612_));
 NAND2x1_ASAP7_75t_R _24012_ (.A(_15509_),
    .B(_15612_),
    .Y(_15613_));
 AND4x1_ASAP7_75t_R _24013_ (.A(_15606_),
    .B(_15609_),
    .C(_15611_),
    .D(_15613_),
    .Y(_15614_));
 NAND2x1_ASAP7_75t_R _24014_ (.A(_15429_),
    .B(_15597_),
    .Y(_15615_));
 BUFx2_ASAP7_75t_R output356 (.A(net356),
    .Y(text_out[71]));
 AO21x1_ASAP7_75t_R _24016_ (.A1(_15469_),
    .A2(_15473_),
    .B(_15563_),
    .Y(_15617_));
 INVx6_ASAP7_75t_R _24017_ (.A(_15552_),
    .Y(_15618_));
 BUFx2_ASAP7_75t_R output355 (.A(net355),
    .Y(text_out[70]));
 AO21x1_ASAP7_75t_R _24019_ (.A1(_15584_),
    .A2(net3553),
    .B(_15618_),
    .Y(_15620_));
 AND5x1_ASAP7_75t_R _24020_ (.A(_15604_),
    .B(_15614_),
    .C(_15615_),
    .D(_15617_),
    .E(_15620_),
    .Y(_15621_));
 BUFx2_ASAP7_75t_R output354 (.A(net354),
    .Y(text_out[6]));
 NOR2x1_ASAP7_75t_R _24022_ (.A(_15453_),
    .B(_15550_),
    .Y(_15623_));
 AO21x1_ASAP7_75t_R _24023_ (.A1(_15618_),
    .A2(_15476_),
    .B(_15516_),
    .Y(_15624_));
 INVx1_ASAP7_75t_R _24024_ (.A(_15624_),
    .Y(_15625_));
 NOR2x1_ASAP7_75t_R _24025_ (.A(_15607_),
    .B(_15490_),
    .Y(_15626_));
 OA21x2_ASAP7_75t_R _24026_ (.A1(_15493_),
    .A2(_15527_),
    .B(_15420_),
    .Y(_15627_));
 OA21x2_ASAP7_75t_R _24027_ (.A1(_15514_),
    .A2(_15443_),
    .B(_15454_),
    .Y(_15628_));
 OR5x1_ASAP7_75t_R _24028_ (.A(_15623_),
    .B(_15625_),
    .C(_15626_),
    .D(_15627_),
    .E(_15628_),
    .Y(_15629_));
 INVx1_ASAP7_75t_R _24029_ (.A(_15629_),
    .Y(_15630_));
 AO21x1_ASAP7_75t_R _24030_ (.A1(_15469_),
    .A2(_15473_),
    .B(_15541_),
    .Y(_15631_));
 NAND2x1_ASAP7_75t_R _24031_ (.A(_15445_),
    .B(_15576_),
    .Y(_15632_));
 AND2x2_ASAP7_75t_R _24032_ (.A(_15631_),
    .B(_15632_),
    .Y(_15633_));
 BUFx2_ASAP7_75t_R output353 (.A(net353),
    .Y(text_out[69]));
 NOR2x1_ASAP7_75t_R _24034_ (.A(net3561),
    .B(_15397_),
    .Y(_15635_));
 BUFx2_ASAP7_75t_R output352 (.A(net352),
    .Y(text_out[68]));
 NOR2x1_ASAP7_75t_R _24036_ (.A(_15608_),
    .B(_15499_),
    .Y(_15637_));
 AO21x1_ASAP7_75t_R _24037_ (.A1(_15602_),
    .A2(_15527_),
    .B(_15637_),
    .Y(_15638_));
 AO221x1_ASAP7_75t_R _24038_ (.A1(_15449_),
    .A2(_15481_),
    .B1(_15475_),
    .B2(_15635_),
    .C(_15638_),
    .Y(_15639_));
 INVx1_ASAP7_75t_R _24039_ (.A(_15639_),
    .Y(_15640_));
 OR3x2_ASAP7_75t_R _24040_ (.A(_15524_),
    .B(_15479_),
    .C(net3553),
    .Y(_15641_));
 BUFx2_ASAP7_75t_R output351 (.A(net351),
    .Y(text_out[67]));
 BUFx2_ASAP7_75t_R output350 (.A(net350),
    .Y(text_out[66]));
 AO21x1_ASAP7_75t_R _24043_ (.A1(_15550_),
    .A2(_15575_),
    .B(_15503_),
    .Y(_15644_));
 NAND2x1_ASAP7_75t_R _24044_ (.A(_15404_),
    .B(_15567_),
    .Y(_15645_));
 AND3x1_ASAP7_75t_R _24045_ (.A(_15641_),
    .B(_15644_),
    .C(_15645_),
    .Y(_15646_));
 AND4x1_ASAP7_75t_R _24046_ (.A(_15630_),
    .B(_15633_),
    .C(_15640_),
    .D(_15646_),
    .Y(_15647_));
 AND3x1_ASAP7_75t_R _24047_ (.A(_15600_),
    .B(_15621_),
    .C(_15647_),
    .Y(_15648_));
 NAND2x2_ASAP7_75t_R _24048_ (.A(_15562_),
    .B(_15648_),
    .Y(_15649_));
 AO21x1_ASAP7_75t_R _24049_ (.A1(_15496_),
    .A2(_15540_),
    .B(_15563_),
    .Y(_15650_));
 OA21x2_ASAP7_75t_R _24050_ (.A1(net3558),
    .A2(_15563_),
    .B(_15650_),
    .Y(_15651_));
 NAND2x1_ASAP7_75t_R _24051_ (.A(_15424_),
    .B(_15472_),
    .Y(_15652_));
 NOR2x1_ASAP7_75t_R _24052_ (.A(_15442_),
    .B(_15563_),
    .Y(_15653_));
 INVx1_ASAP7_75t_R _24053_ (.A(_15653_),
    .Y(_15654_));
 AO21x1_ASAP7_75t_R _24054_ (.A1(_15469_),
    .A2(_15575_),
    .B(_15563_),
    .Y(_15655_));
 AND4x1_ASAP7_75t_R _24055_ (.A(_15651_),
    .B(_15652_),
    .C(_15654_),
    .D(_15655_),
    .Y(_15656_));
 AND5x2_ASAP7_75t_R _24056_ (.A(_00437_),
    .B(_15656_),
    .C(_00438_),
    .D(_00439_),
    .E(_00440_),
    .Y(_15657_));
 BUFx2_ASAP7_75t_R output349 (.A(net349),
    .Y(text_out[65]));
 BUFx2_ASAP7_75t_R output348 (.A(net348),
    .Y(text_out[64]));
 XOR2x1_ASAP7_75t_R _24059_ (.A(_00413_),
    .Y(_15660_),
    .B(net2203));
 INVx4_ASAP7_75t_R _24060_ (.A(_00468_),
    .Y(_15661_));
 XOR2x1_ASAP7_75t_R _24061_ (.A(_15660_),
    .Y(_15662_),
    .B(_15661_));
 XOR2x1_ASAP7_75t_R _24062_ (.A(_15662_),
    .Y(_15663_),
    .B(_00492_));
 NOR3x1_ASAP7_75t_R _24063_ (.A(_15649_),
    .B(_15657_),
    .C(_15663_),
    .Y(_15664_));
 OA21x2_ASAP7_75t_R _24064_ (.A1(_15649_),
    .A2(_15657_),
    .B(_15663_),
    .Y(_15665_));
 OAI21x1_ASAP7_75t_R _24065_ (.A1(_15664_),
    .A2(_15665_),
    .B(_08823_),
    .Y(_15666_));
 OAI21x1_ASAP7_75t_R _24066_ (.A1(_08823_),
    .A2(net3968),
    .B(_15666_),
    .Y(_00360_));
 INVx2_ASAP7_75t_R _24067_ (.A(net3794),
    .Y(_15667_));
 AO21x1_ASAP7_75t_R _24068_ (.A1(_15473_),
    .A2(_15516_),
    .B(_15503_),
    .Y(_15668_));
 AO21x1_ASAP7_75t_R _24069_ (.A1(_15496_),
    .A2(_15417_),
    .B(_15503_),
    .Y(_15669_));
 NAND2x1_ASAP7_75t_R _24070_ (.A(_15502_),
    .B(_15449_),
    .Y(_15670_));
 INVx1_ASAP7_75t_R _24071_ (.A(_15506_),
    .Y(_15671_));
 AND4x1_ASAP7_75t_R _24072_ (.A(_15668_),
    .B(_15669_),
    .C(_15670_),
    .D(_15671_),
    .Y(_15672_));
 OA211x2_ASAP7_75t_R _24073_ (.A1(_00443_),
    .A2(_00444_),
    .B(_15424_),
    .C(_15429_),
    .Y(_15673_));
 INVx1_ASAP7_75t_R _24074_ (.A(_15673_),
    .Y(_15674_));
 AND5x1_ASAP7_75t_R _24075_ (.A(_15565_),
    .B(_15672_),
    .C(_15652_),
    .D(_15654_),
    .E(_15674_),
    .Y(_15675_));
 NAND2x1_ASAP7_75t_R _24076_ (.A(_15443_),
    .B(_15484_),
    .Y(_15676_));
 NAND2x1_ASAP7_75t_R _24077_ (.A(_15468_),
    .B(_15484_),
    .Y(_15677_));
 NAND2x1_ASAP7_75t_R _24078_ (.A(_15549_),
    .B(_15484_),
    .Y(_15678_));
 AND5x1_ASAP7_75t_R _24079_ (.A(_15566_),
    .B(_15577_),
    .C(_15676_),
    .D(_15677_),
    .E(_15678_),
    .Y(_15679_));
 AND3x1_ASAP7_75t_R _24080_ (.A(_15475_),
    .B(_15429_),
    .C(_15548_),
    .Y(_15680_));
 INVx1_ASAP7_75t_R _24081_ (.A(_15680_),
    .Y(_15681_));
 BUFx2_ASAP7_75t_R output347 (.A(net347),
    .Y(text_out[63]));
 OA211x2_ASAP7_75t_R _24083_ (.A1(_15425_),
    .A2(net3551),
    .B(_15475_),
    .C(_15416_),
    .Y(_15683_));
 INVx1_ASAP7_75t_R _24084_ (.A(_15683_),
    .Y(_15684_));
 INVx1_ASAP7_75t_R _24085_ (.A(_15522_),
    .Y(_15685_));
 INVx1_ASAP7_75t_R _24086_ (.A(_15529_),
    .Y(_15686_));
 NAND2x2_ASAP7_75t_R _24087_ (.A(_15397_),
    .B(_15429_),
    .Y(_15687_));
 BUFx2_ASAP7_75t_R output346 (.A(net346),
    .Y(text_out[62]));
 AO21x1_ASAP7_75t_R _24089_ (.A1(_15584_),
    .A2(_15687_),
    .B(_15486_),
    .Y(_15689_));
 AND3x1_ASAP7_75t_R _24090_ (.A(_15685_),
    .B(_15686_),
    .C(_15689_),
    .Y(_15690_));
 AND4x1_ASAP7_75t_R _24091_ (.A(_15679_),
    .B(_15681_),
    .C(_15684_),
    .D(_15690_),
    .Y(_15691_));
 NAND2x1_ASAP7_75t_R _24092_ (.A(_15675_),
    .B(_15691_),
    .Y(_15692_));
 AO21x1_ASAP7_75t_R _24093_ (.A1(_15483_),
    .A2(net3562),
    .B(_15437_),
    .Y(_15693_));
 NOR2x2_ASAP7_75t_R _24094_ (.A(_15441_),
    .B(net3553),
    .Y(_15694_));
 INVx8_ASAP7_75t_R _24095_ (.A(_15694_),
    .Y(_15695_));
 BUFx2_ASAP7_75t_R output345 (.A(net345),
    .Y(text_out[61]));
 NOR2x2_ASAP7_75t_R _24097_ (.A(_15425_),
    .B(net3554),
    .Y(_15697_));
 INVx3_ASAP7_75t_R _24098_ (.A(_15697_),
    .Y(_15698_));
 AO21x1_ASAP7_75t_R _24099_ (.A1(_15695_),
    .A2(_15698_),
    .B(_15437_),
    .Y(_15699_));
 BUFx2_ASAP7_75t_R output344 (.A(net344),
    .Y(text_out[60]));
 AO21x1_ASAP7_75t_R _24101_ (.A1(_15417_),
    .A2(_15687_),
    .B(_15437_),
    .Y(_15701_));
 AND3x1_ASAP7_75t_R _24102_ (.A(_15693_),
    .B(_15699_),
    .C(_15701_),
    .Y(_15702_));
 AND3x1_ASAP7_75t_R _24103_ (.A(_15509_),
    .B(_15429_),
    .C(_15548_),
    .Y(_15703_));
 INVx1_ASAP7_75t_R _24104_ (.A(_15703_),
    .Y(_15704_));
 BUFx2_ASAP7_75t_R output343 (.A(net343),
    .Y(text_out[5]));
 NOR2x1_ASAP7_75t_R _24106_ (.A(_15510_),
    .B(_15571_),
    .Y(_15706_));
 INVx1_ASAP7_75t_R _24107_ (.A(_15706_),
    .Y(_15707_));
 AND5x1_ASAP7_75t_R _24108_ (.A(_15513_),
    .B(_15704_),
    .C(_15517_),
    .D(_15579_),
    .E(_15707_),
    .Y(_15708_));
 NAND2x1_ASAP7_75t_R _24109_ (.A(_15702_),
    .B(_15708_),
    .Y(_15709_));
 NOR2x1_ASAP7_75t_R _24110_ (.A(net3561),
    .B(_15524_),
    .Y(_15710_));
 INVx1_ASAP7_75t_R _24111_ (.A(_15408_),
    .Y(_15711_));
 AND2x2_ASAP7_75t_R _24112_ (.A(_15710_),
    .B(_15711_),
    .Y(_15712_));
 INVx1_ASAP7_75t_R _24113_ (.A(_15712_),
    .Y(_15713_));
 BUFx2_ASAP7_75t_R output342 (.A(net342),
    .Y(text_out[59]));
 BUFx2_ASAP7_75t_R output341 (.A(net341),
    .Y(text_out[58]));
 AO21x1_ASAP7_75t_R _24116_ (.A1(_15505_),
    .A2(_15448_),
    .B(_15524_),
    .Y(_15716_));
 AO21x1_ASAP7_75t_R _24117_ (.A1(_15473_),
    .A2(_15516_),
    .B(_15524_),
    .Y(_15717_));
 AND3x1_ASAP7_75t_R _24118_ (.A(_15713_),
    .B(_15716_),
    .C(_15717_),
    .Y(_15718_));
 INVx1_ASAP7_75t_R _24119_ (.A(_15718_),
    .Y(_15719_));
 NAND2x1_ASAP7_75t_R _24120_ (.A(_15570_),
    .B(_15454_),
    .Y(_15720_));
 NOR2x1_ASAP7_75t_R _24121_ (.A(_15453_),
    .B(_15496_),
    .Y(_15721_));
 INVx1_ASAP7_75t_R _24122_ (.A(_15721_),
    .Y(_15722_));
 NAND2x1_ASAP7_75t_R _24123_ (.A(_15720_),
    .B(_15722_),
    .Y(_15723_));
 AO21x1_ASAP7_75t_R _24124_ (.A1(_15449_),
    .A2(_15454_),
    .B(_15723_),
    .Y(_15724_));
 AND3x2_ASAP7_75t_R _24125_ (.A(_15454_),
    .B(_15398_),
    .C(_15711_),
    .Y(_15725_));
 NAND2x1_ASAP7_75t_R _24126_ (.A(_15694_),
    .B(_15454_),
    .Y(_15726_));
 INVx1_ASAP7_75t_R _24127_ (.A(_15726_),
    .Y(_15727_));
 NOR2x1_ASAP7_75t_R _24128_ (.A(_15453_),
    .B(_15469_),
    .Y(_15728_));
 OR3x1_ASAP7_75t_R _24129_ (.A(_15725_),
    .B(_15727_),
    .C(_15728_),
    .Y(_15729_));
 OR4x2_ASAP7_75t_R _24130_ (.A(_15709_),
    .B(_15719_),
    .C(_15724_),
    .D(_15729_),
    .Y(_15730_));
 NOR2x1_ASAP7_75t_R _24131_ (.A(_15692_),
    .B(_15730_),
    .Y(_15731_));
 AO21x1_ASAP7_75t_R _24132_ (.A1(_15584_),
    .A2(_15687_),
    .B(_15603_),
    .Y(_15732_));
 NAND2x1_ASAP7_75t_R _24133_ (.A(_15602_),
    .B(_15612_),
    .Y(_15733_));
 NAND2x1_ASAP7_75t_R _24134_ (.A(_15602_),
    .B(_15570_),
    .Y(_15734_));
 AND3x1_ASAP7_75t_R _24135_ (.A(_15732_),
    .B(_15733_),
    .C(_15734_),
    .Y(_15735_));
 AO21x1_ASAP7_75t_R _24136_ (.A1(_15584_),
    .A2(_15533_),
    .B(_15618_),
    .Y(_15736_));
 AO21x1_ASAP7_75t_R _24137_ (.A1(_15483_),
    .A2(_15409_),
    .B(_15618_),
    .Y(_15737_));
 NAND2x1_ASAP7_75t_R _24138_ (.A(_15552_),
    .B(_15595_),
    .Y(_15738_));
 NAND2x1_ASAP7_75t_R _24139_ (.A(_15552_),
    .B(_15570_),
    .Y(_15739_));
 NAND2x1_ASAP7_75t_R _24140_ (.A(_15694_),
    .B(_15552_),
    .Y(_15740_));
 AND5x1_ASAP7_75t_R _24141_ (.A(_15736_),
    .B(_15737_),
    .C(_15738_),
    .D(_15739_),
    .E(_15740_),
    .Y(_15741_));
 NOR2x1_ASAP7_75t_R _24142_ (.A(_15608_),
    .B(_15603_),
    .Y(_15742_));
 INVx1_ASAP7_75t_R _24143_ (.A(_15742_),
    .Y(_15743_));
 INVx3_ASAP7_75t_R _24144_ (.A(_15409_),
    .Y(_15744_));
 NAND2x1_ASAP7_75t_R _24145_ (.A(_15602_),
    .B(_15744_),
    .Y(_15745_));
 NAND2x1_ASAP7_75t_R _24146_ (.A(_15602_),
    .B(_15549_),
    .Y(_15746_));
 AND3x1_ASAP7_75t_R _24147_ (.A(_15743_),
    .B(_15745_),
    .C(_15746_),
    .Y(_15747_));
 AO21x1_ASAP7_75t_R _24148_ (.A1(_15483_),
    .A2(_15409_),
    .B(_15490_),
    .Y(_15748_));
 NAND2x1_ASAP7_75t_R _24149_ (.A(_15504_),
    .B(_15460_),
    .Y(_15749_));
 NAND2x1_ASAP7_75t_R _24150_ (.A(net3542),
    .B(_15460_),
    .Y(_15750_));
 NAND2x1_ASAP7_75t_R _24151_ (.A(_15697_),
    .B(_15460_),
    .Y(_15751_));
 AND4x1_ASAP7_75t_R _24152_ (.A(_15748_),
    .B(_15749_),
    .C(_15750_),
    .D(_15751_),
    .Y(_15752_));
 AO21x1_ASAP7_75t_R _24153_ (.A1(_15505_),
    .A2(_15537_),
    .B(_15541_),
    .Y(_15753_));
 NAND2x1_ASAP7_75t_R _24154_ (.A(_15549_),
    .B(_15445_),
    .Y(_15754_));
 NAND2x1_ASAP7_75t_R _24155_ (.A(_15445_),
    .B(_15399_),
    .Y(_15755_));
 AND4x1_ASAP7_75t_R _24156_ (.A(_15753_),
    .B(_15754_),
    .C(_15447_),
    .D(_15755_),
    .Y(_15756_));
 AND5x1_ASAP7_75t_R _24157_ (.A(_15735_),
    .B(_15741_),
    .C(_15747_),
    .D(_15752_),
    .E(_15756_),
    .Y(_15757_));
 AO21x1_ASAP7_75t_R _24158_ (.A1(_15528_),
    .A2(_15417_),
    .B(_15413_),
    .Y(_15758_));
 AO21x1_ASAP7_75t_R _24159_ (.A1(_15469_),
    .A2(_15550_),
    .B(_15413_),
    .Y(_15759_));
 NAND2x1_ASAP7_75t_R _24160_ (.A(net2773),
    .B(_15412_),
    .Y(_15760_));
 NAND2x1_ASAP7_75t_R _24161_ (.A(_15514_),
    .B(_15412_),
    .Y(_15761_));
 NAND2x2_ASAP7_75t_R _24162_ (.A(_15443_),
    .B(_15412_),
    .Y(_15762_));
 AND5x1_ASAP7_75t_R _24163_ (.A(_15758_),
    .B(_15759_),
    .C(_15760_),
    .D(_15761_),
    .E(_15762_),
    .Y(_15763_));
 INVx1_ASAP7_75t_R _24164_ (.A(_15627_),
    .Y(_15764_));
 NAND2x1_ASAP7_75t_R _24165_ (.A(_15420_),
    .B(_15399_),
    .Y(_15765_));
 AO21x1_ASAP7_75t_R _24166_ (.A1(_15469_),
    .A2(_15695_),
    .B(_15421_),
    .Y(_15766_));
 AND3x1_ASAP7_75t_R _24167_ (.A(_15764_),
    .B(_15765_),
    .C(_15766_),
    .Y(_15767_));
 AO21x1_ASAP7_75t_R _24168_ (.A1(_15584_),
    .A2(_15448_),
    .B(_15499_),
    .Y(_15768_));
 NAND2x1_ASAP7_75t_R _24169_ (.A(_15398_),
    .B(_15498_),
    .Y(_15769_));
 NAND2x1_ASAP7_75t_R _24170_ (.A(_15697_),
    .B(_15498_),
    .Y(_15770_));
 AND4x1_ASAP7_75t_R _24171_ (.A(_15768_),
    .B(_15581_),
    .C(_15769_),
    .D(_15770_),
    .Y(_15771_));
 INVx4_ASAP7_75t_R _24172_ (.A(_15481_),
    .Y(_15772_));
 BUFx2_ASAP7_75t_R output340 (.A(net340),
    .Y(text_out[57]));
 AO21x1_ASAP7_75t_R _24174_ (.A1(_15550_),
    .A2(_15698_),
    .B(_15772_),
    .Y(_15774_));
 BUFx2_ASAP7_75t_R output339 (.A(net339),
    .Y(text_out[56]));
 AO21x1_ASAP7_75t_R _24176_ (.A1(_15540_),
    .A2(net3541),
    .B(_15772_),
    .Y(_15776_));
 OA211x2_ASAP7_75t_R _24177_ (.A1(_15584_),
    .A2(_15772_),
    .B(_15774_),
    .C(_15776_),
    .Y(_15777_));
 AND4x1_ASAP7_75t_R _24178_ (.A(_15763_),
    .B(_15767_),
    .C(_15771_),
    .D(_15777_),
    .Y(_15778_));
 AND2x2_ASAP7_75t_R _24179_ (.A(_15757_),
    .B(_15778_),
    .Y(_15779_));
 NAND2x2_ASAP7_75t_R _24180_ (.A(_15731_),
    .B(_15779_),
    .Y(_15780_));
 BUFx2_ASAP7_75t_R output338 (.A(net338),
    .Y(text_out[55]));
 BUFx2_ASAP7_75t_R output337 (.A(net337),
    .Y(text_out[54]));
 XOR2x1_ASAP7_75t_R _24183_ (.A(_00414_),
    .Y(_15783_),
    .B(net1854));
 INVx4_ASAP7_75t_R _24184_ (.A(_00467_),
    .Y(_15784_));
 XOR2x1_ASAP7_75t_R _24185_ (.A(_15783_),
    .Y(_15785_),
    .B(_15784_));
 BUFx2_ASAP7_75t_R output336 (.A(net336),
    .Y(text_out[53]));
 XOR2x1_ASAP7_75t_R _24187_ (.A(_15785_),
    .Y(_15787_),
    .B(_00491_));
 NOR3x1_ASAP7_75t_R _24188_ (.A(_15780_),
    .B(_15657_),
    .C(_15787_),
    .Y(_15788_));
 OA21x2_ASAP7_75t_R _24189_ (.A1(_15780_),
    .A2(_15657_),
    .B(_15787_),
    .Y(_15789_));
 OAI21x1_ASAP7_75t_R _24190_ (.A1(_15788_),
    .A2(_15789_),
    .B(_08823_),
    .Y(_15790_));
 OAI21x1_ASAP7_75t_R _24191_ (.A1(_08823_),
    .A2(net3795),
    .B(_15790_),
    .Y(_00361_));
 OA21x2_ASAP7_75t_R _24192_ (.A1(_15744_),
    .A2(_15514_),
    .B(_15420_),
    .Y(_15791_));
 INVx1_ASAP7_75t_R _24193_ (.A(_15791_),
    .Y(_15792_));
 AO21x1_ASAP7_75t_R _24194_ (.A1(_15515_),
    .A2(_15409_),
    .B(_15499_),
    .Y(_15793_));
 NAND2x1_ASAP7_75t_R _24195_ (.A(_15498_),
    .B(_15549_),
    .Y(_15794_));
 AND3x1_ASAP7_75t_R _24196_ (.A(_15793_),
    .B(_15770_),
    .C(_15794_),
    .Y(_15795_));
 NAND2x1_ASAP7_75t_R _24197_ (.A(_15435_),
    .B(_15420_),
    .Y(_15796_));
 NAND2x1_ASAP7_75t_R _24198_ (.A(_15420_),
    .B(_15567_),
    .Y(_15797_));
 OA21x2_ASAP7_75t_R _24199_ (.A1(_15421_),
    .A2(_15428_),
    .B(_15797_),
    .Y(_15798_));
 AO21x1_ASAP7_75t_R _24200_ (.A1(_15571_),
    .A2(_15528_),
    .B(_15499_),
    .Y(_15799_));
 AND5x2_ASAP7_75t_R _24201_ (.A(_15792_),
    .B(_15795_),
    .C(_15796_),
    .D(_15798_),
    .E(_15799_),
    .Y(_15800_));
 AND2x2_ASAP7_75t_R _24202_ (.A(net3542),
    .B(_15481_),
    .Y(_15801_));
 OA21x2_ASAP7_75t_R _24203_ (.A1(_15514_),
    .A2(_15443_),
    .B(_15481_),
    .Y(_15802_));
 AND2x2_ASAP7_75t_R _24204_ (.A(_15583_),
    .B(_15481_),
    .Y(_15803_));
 AND2x2_ASAP7_75t_R _24205_ (.A(net2773),
    .B(_15481_),
    .Y(_15804_));
 NOR2x1_ASAP7_75t_R _24206_ (.A(_15687_),
    .B(_15772_),
    .Y(_15805_));
 OR5x1_ASAP7_75t_R _24207_ (.A(_15801_),
    .B(_15802_),
    .C(_15803_),
    .D(_15804_),
    .E(_15805_),
    .Y(_15806_));
 OA211x2_ASAP7_75t_R _24208_ (.A1(_15425_),
    .A2(net3549),
    .B(_15412_),
    .C(_15416_),
    .Y(_15807_));
 INVx1_ASAP7_75t_R _24209_ (.A(_15762_),
    .Y(_15808_));
 OA21x2_ASAP7_75t_R _24210_ (.A1(net2773),
    .A2(_15536_),
    .B(_15412_),
    .Y(_15809_));
 OA21x2_ASAP7_75t_R _24211_ (.A1(net3542),
    .A2(_15697_),
    .B(_15412_),
    .Y(_15810_));
 OR5x1_ASAP7_75t_R _24212_ (.A(_15807_),
    .B(_15414_),
    .C(_15808_),
    .D(_15809_),
    .E(_15810_),
    .Y(_15811_));
 NOR2x1_ASAP7_75t_R _24213_ (.A(_15806_),
    .B(_15811_),
    .Y(_15812_));
 NAND2x2_ASAP7_75t_R _24214_ (.A(_15800_),
    .B(_15812_),
    .Y(_15813_));
 AND2x2_ASAP7_75t_R _24215_ (.A(_15602_),
    .B(_15504_),
    .Y(_15814_));
 INVx1_ASAP7_75t_R _24216_ (.A(_15814_),
    .Y(_15815_));
 AO21x1_ASAP7_75t_R _24217_ (.A1(_15571_),
    .A2(_15528_),
    .B(_15603_),
    .Y(_15816_));
 NOR2x1_ASAP7_75t_R _24218_ (.A(_00441_),
    .B(_15467_),
    .Y(_15817_));
 OA21x2_ASAP7_75t_R _24219_ (.A1(_15472_),
    .A2(_15817_),
    .B(_15602_),
    .Y(_15818_));
 INVx1_ASAP7_75t_R _24220_ (.A(_15818_),
    .Y(_15819_));
 NOR2x1_ASAP7_75t_R _24221_ (.A(_15448_),
    .B(_15603_),
    .Y(_15820_));
 INVx1_ASAP7_75t_R _24222_ (.A(_15820_),
    .Y(_15821_));
 AND5x1_ASAP7_75t_R _24223_ (.A(_15815_),
    .B(_15816_),
    .C(_15819_),
    .D(_15732_),
    .E(_15821_),
    .Y(_15822_));
 INVx1_ASAP7_75t_R _24224_ (.A(_15822_),
    .Y(_15823_));
 AND2x2_ASAP7_75t_R _24225_ (.A(_15445_),
    .B(_15694_),
    .Y(_15824_));
 INVx1_ASAP7_75t_R _24226_ (.A(_15824_),
    .Y(_15825_));
 AO21x1_ASAP7_75t_R _24227_ (.A1(_15483_),
    .A2(_15515_),
    .B(_15541_),
    .Y(_15826_));
 AO21x1_ASAP7_75t_R _24228_ (.A1(_15571_),
    .A2(_15417_),
    .B(_15541_),
    .Y(_15827_));
 NAND2x1_ASAP7_75t_R _24229_ (.A(_15536_),
    .B(_15445_),
    .Y(_15828_));
 AND5x1_ASAP7_75t_R _24230_ (.A(_15825_),
    .B(_15826_),
    .C(_15827_),
    .D(_15754_),
    .E(_15828_),
    .Y(_15829_));
 INVx1_ASAP7_75t_R _24231_ (.A(_15829_),
    .Y(_15830_));
 OA211x2_ASAP7_75t_R _24232_ (.A1(net3546),
    .A2(_15432_),
    .B(_15460_),
    .C(_15398_),
    .Y(_15831_));
 NOR2x1_ASAP7_75t_R _24233_ (.A(_15533_),
    .B(_15490_),
    .Y(_15832_));
 OA21x2_ASAP7_75t_R _24234_ (.A1(_15468_),
    .A2(net3542),
    .B(_15460_),
    .Y(_15833_));
 OR3x1_ASAP7_75t_R _24235_ (.A(_15831_),
    .B(_15832_),
    .C(_15833_),
    .Y(_15834_));
 AO21x1_ASAP7_75t_R _24236_ (.A1(_15571_),
    .A2(_15528_),
    .B(_15618_),
    .Y(_15835_));
 OA211x2_ASAP7_75t_R _24237_ (.A1(_15533_),
    .A2(_15618_),
    .B(_15835_),
    .C(_15738_),
    .Y(_15836_));
 AO21x1_ASAP7_75t_R _24238_ (.A1(_15469_),
    .A2(_15695_),
    .B(_15618_),
    .Y(_15837_));
 OA211x2_ASAP7_75t_R _24239_ (.A1(_15425_),
    .A2(net3549),
    .B(_15552_),
    .C(_15398_),
    .Y(_15838_));
 INVx1_ASAP7_75t_R _24240_ (.A(_15838_),
    .Y(_15839_));
 NAND3x1_ASAP7_75t_R _24241_ (.A(_15836_),
    .B(_15837_),
    .C(_15839_),
    .Y(_15840_));
 OR4x2_ASAP7_75t_R _24242_ (.A(_15823_),
    .B(_15830_),
    .C(_15834_),
    .D(_15840_),
    .Y(_15841_));
 NOR2x2_ASAP7_75t_R _24243_ (.A(_15813_),
    .B(_15841_),
    .Y(_15842_));
 OA211x2_ASAP7_75t_R _24244_ (.A1(_00443_),
    .A2(_15432_),
    .B(_15475_),
    .C(_15416_),
    .Y(_15843_));
 AO21x1_ASAP7_75t_R _24245_ (.A1(_15429_),
    .A2(_15475_),
    .B(_15843_),
    .Y(_15844_));
 NOR2x1_ASAP7_75t_R _24246_ (.A(_15476_),
    .B(_15483_),
    .Y(_15845_));
 NAND2x1_ASAP7_75t_R _24247_ (.A(_15697_),
    .B(_15475_),
    .Y(_15846_));
 INVx1_ASAP7_75t_R _24248_ (.A(_15846_),
    .Y(_15847_));
 AO21x1_ASAP7_75t_R _24249_ (.A1(net3542),
    .A2(_15475_),
    .B(_15847_),
    .Y(_15848_));
 OR3x1_ASAP7_75t_R _24250_ (.A(_15844_),
    .B(_15845_),
    .C(_15848_),
    .Y(_15849_));
 OA21x2_ASAP7_75t_R _24251_ (.A1(_15612_),
    .A2(_15595_),
    .B(_15484_),
    .Y(_15850_));
 INVx1_ASAP7_75t_R _24252_ (.A(_15850_),
    .Y(_15851_));
 AO21x1_ASAP7_75t_R _24253_ (.A1(_15505_),
    .A2(_15584_),
    .B(_15486_),
    .Y(_15852_));
 AO21x1_ASAP7_75t_R _24254_ (.A1(_15483_),
    .A2(_15515_),
    .B(_15486_),
    .Y(_15853_));
 AND4x1_ASAP7_75t_R _24255_ (.A(_15851_),
    .B(_15852_),
    .C(_15853_),
    .D(_15577_),
    .Y(_15854_));
 INVx1_ASAP7_75t_R _24256_ (.A(_15854_),
    .Y(_15855_));
 NOR2x1_ASAP7_75t_R _24257_ (.A(_15496_),
    .B(_15563_),
    .Y(_15856_));
 AO21x1_ASAP7_75t_R _24258_ (.A1(_15424_),
    .A2(_15527_),
    .B(_15856_),
    .Y(_15857_));
 INVx1_ASAP7_75t_R _24259_ (.A(_15480_),
    .Y(_15858_));
 AO21x1_ASAP7_75t_R _24260_ (.A1(_15858_),
    .A2(_15695_),
    .B(_15563_),
    .Y(_15859_));
 INVx1_ASAP7_75t_R _24261_ (.A(_15859_),
    .Y(_15860_));
 OR3x1_ASAP7_75t_R _24262_ (.A(_15857_),
    .B(_15860_),
    .C(_15431_),
    .Y(_15861_));
 AO21x1_ASAP7_75t_R _24263_ (.A1(_15515_),
    .A2(net3563),
    .B(_15503_),
    .Y(_15862_));
 AO21x1_ASAP7_75t_R _24264_ (.A1(_15550_),
    .A2(_15698_),
    .B(_15503_),
    .Y(_15863_));
 AND4x1_ASAP7_75t_R _24265_ (.A(_15862_),
    .B(_15863_),
    .C(_15671_),
    .D(_15573_),
    .Y(_15864_));
 INVx1_ASAP7_75t_R _24266_ (.A(_15864_),
    .Y(_15865_));
 OR4x2_ASAP7_75t_R _24267_ (.A(_15849_),
    .B(_15855_),
    .C(_15861_),
    .D(_15865_),
    .Y(_15866_));
 NOR2x1_ASAP7_75t_R _24268_ (.A(_15524_),
    .B(_15515_),
    .Y(_15867_));
 NOR2x1_ASAP7_75t_R _24269_ (.A(_15462_),
    .B(_15641_),
    .Y(_15868_));
 AO21x1_ASAP7_75t_R _24270_ (.A1(_15584_),
    .A2(_15687_),
    .B(_15524_),
    .Y(_15869_));
 INVx1_ASAP7_75t_R _24271_ (.A(_15869_),
    .Y(_15870_));
 OR5x1_ASAP7_75t_R _24272_ (.A(_15867_),
    .B(_15868_),
    .C(_15870_),
    .D(_15525_),
    .E(_15593_),
    .Y(_15871_));
 INVx1_ASAP7_75t_R _24273_ (.A(_15871_),
    .Y(_15872_));
 AND2x2_ASAP7_75t_R _24274_ (.A(_15694_),
    .B(_15404_),
    .Y(_15873_));
 AND2x2_ASAP7_75t_R _24275_ (.A(_15570_),
    .B(_15404_),
    .Y(_15874_));
 AND2x2_ASAP7_75t_R _24276_ (.A(_15514_),
    .B(_15404_),
    .Y(_15875_));
 AND2x2_ASAP7_75t_R _24277_ (.A(_15583_),
    .B(_15404_),
    .Y(_15876_));
 OR5x1_ASAP7_75t_R _24278_ (.A(_15873_),
    .B(_15874_),
    .C(_15406_),
    .D(_15875_),
    .E(_15876_),
    .Y(_15877_));
 NOR2x2_ASAP7_75t_R _24279_ (.A(_15510_),
    .B(_15695_),
    .Y(_15878_));
 INVx1_ASAP7_75t_R _24280_ (.A(_15878_),
    .Y(_15879_));
 NOR2x1_ASAP7_75t_R _24281_ (.A(_15516_),
    .B(_15510_),
    .Y(_15880_));
 INVx1_ASAP7_75t_R _24282_ (.A(_15880_),
    .Y(_15881_));
 NOR2x1_ASAP7_75t_R _24283_ (.A(_15510_),
    .B(_15483_),
    .Y(_15882_));
 INVx1_ASAP7_75t_R _24284_ (.A(_15882_),
    .Y(_15883_));
 NOR2x1_ASAP7_75t_R _24285_ (.A(_15510_),
    .B(_15584_),
    .Y(_15884_));
 INVx1_ASAP7_75t_R _24286_ (.A(_15884_),
    .Y(_15885_));
 AND2x2_ASAP7_75t_R _24287_ (.A(_15527_),
    .B(_15509_),
    .Y(_15886_));
 INVx1_ASAP7_75t_R _24288_ (.A(_15886_),
    .Y(_15887_));
 AND5x1_ASAP7_75t_R _24289_ (.A(_15879_),
    .B(_15881_),
    .C(_15883_),
    .D(_15885_),
    .E(_15887_),
    .Y(_15888_));
 INVx1_ASAP7_75t_R _24290_ (.A(_15888_),
    .Y(_15889_));
 NOR2x1_ASAP7_75t_R _24291_ (.A(_15877_),
    .B(_15889_),
    .Y(_15890_));
 AO21x1_ASAP7_75t_R _24292_ (.A1(_15469_),
    .A2(_15575_),
    .B(_15453_),
    .Y(_15891_));
 NOR2x1_ASAP7_75t_R _24293_ (.A(_15453_),
    .B(_15687_),
    .Y(_15892_));
 INVx1_ASAP7_75t_R _24294_ (.A(_15892_),
    .Y(_15893_));
 NAND2x1_ASAP7_75t_R _24295_ (.A(_15583_),
    .B(_15454_),
    .Y(_15894_));
 NAND2x1_ASAP7_75t_R _24296_ (.A(_15514_),
    .B(_15454_),
    .Y(_15895_));
 AND5x1_ASAP7_75t_R _24297_ (.A(_15891_),
    .B(_15720_),
    .C(_15893_),
    .D(_15894_),
    .E(_15895_),
    .Y(_15896_));
 AND3x1_ASAP7_75t_R _24298_ (.A(_15872_),
    .B(_15890_),
    .C(_15896_),
    .Y(_15897_));
 INVx1_ASAP7_75t_R _24299_ (.A(_15897_),
    .Y(_15898_));
 NOR2x1_ASAP7_75t_R _24300_ (.A(_15866_),
    .B(_15898_),
    .Y(_15899_));
 NAND2x2_ASAP7_75t_R _24301_ (.A(_15842_),
    .B(_15899_),
    .Y(_15900_));
 XOR2x2_ASAP7_75t_R _24302_ (.A(_00466_),
    .B(_00512_),
    .Y(_15901_));
 BUFx2_ASAP7_75t_R output335 (.A(net335),
    .Y(text_out[52]));
 XOR2x1_ASAP7_75t_R _24304_ (.A(_00393_),
    .Y(_15903_),
    .B(net3483));
 XOR2x1_ASAP7_75t_R _24305_ (.A(_15901_),
    .Y(_15904_),
    .B(_15903_));
 XOR2x1_ASAP7_75t_R _24306_ (.A(_15900_),
    .Y(_15905_),
    .B(_15904_));
 AND2x2_ASAP7_75t_R _24307_ (.A(net402),
    .B(net4144),
    .Y(_15906_));
 AO21x1_ASAP7_75t_R _24308_ (.A1(_15905_),
    .A2(net398),
    .B(_15906_),
    .Y(_00362_));
 AO21x1_ASAP7_75t_R _24309_ (.A1(_15515_),
    .A2(_15516_),
    .B(_15421_),
    .Y(_15907_));
 NAND2x1_ASAP7_75t_R _24310_ (.A(_15420_),
    .B(_15472_),
    .Y(_15908_));
 NAND2x1_ASAP7_75t_R _24311_ (.A(_15420_),
    .B(_15449_),
    .Y(_15909_));
 AND4x1_ASAP7_75t_R _24312_ (.A(_15907_),
    .B(_15908_),
    .C(_15797_),
    .D(_15909_),
    .Y(_15910_));
 AO21x1_ASAP7_75t_R _24313_ (.A1(_15571_),
    .A2(net3541),
    .B(_15413_),
    .Y(_15911_));
 INVx2_ASAP7_75t_R _24314_ (.A(_15687_),
    .Y(_15912_));
 NAND2x1_ASAP7_75t_R _24315_ (.A(_15912_),
    .B(_15412_),
    .Y(_15913_));
 NAND2x1_ASAP7_75t_R _24316_ (.A(_15449_),
    .B(_15412_),
    .Y(_15914_));
 AND4x1_ASAP7_75t_R _24317_ (.A(_15911_),
    .B(_15913_),
    .C(_15914_),
    .D(_15760_),
    .Y(_15915_));
 AO21x1_ASAP7_75t_R _24318_ (.A1(_15469_),
    .A2(_15695_),
    .B(_15499_),
    .Y(_15916_));
 BUFx2_ASAP7_75t_R output334 (.A(net334),
    .Y(text_out[51]));
 AO21x1_ASAP7_75t_R _24320_ (.A1(_15584_),
    .A2(_15687_),
    .B(_15499_),
    .Y(_15918_));
 AND4x1_ASAP7_75t_R _24321_ (.A(_15799_),
    .B(_15916_),
    .C(_15918_),
    .D(_15769_),
    .Y(_15919_));
 AO21x1_ASAP7_75t_R _24322_ (.A1(_15483_),
    .A2(_15695_),
    .B(_15772_),
    .Y(_15920_));
 AO21x1_ASAP7_75t_R _24323_ (.A1(_15687_),
    .A2(_15448_),
    .B(_15772_),
    .Y(_15921_));
 OA211x2_ASAP7_75t_R _24324_ (.A1(_15540_),
    .A2(_15772_),
    .B(_15920_),
    .C(_15921_),
    .Y(_15922_));
 AO21x1_ASAP7_75t_R _24325_ (.A1(_15607_),
    .A2(_15608_),
    .B(_15413_),
    .Y(_15923_));
 AO21x1_ASAP7_75t_R _24326_ (.A1(_15575_),
    .A2(_15550_),
    .B(_15413_),
    .Y(_15924_));
 AND2x2_ASAP7_75t_R _24327_ (.A(_15923_),
    .B(_15924_),
    .Y(_15925_));
 AND5x2_ASAP7_75t_R _24328_ (.A(_15910_),
    .B(_15915_),
    .C(_15919_),
    .D(_15922_),
    .E(_15925_),
    .Y(_15926_));
 AO21x1_ASAP7_75t_R _24329_ (.A1(_15528_),
    .A2(net3541),
    .B(_15490_),
    .Y(_15927_));
 OA211x2_ASAP7_75t_R _24330_ (.A1(_15490_),
    .A2(_15537_),
    .B(_15927_),
    .C(_15749_),
    .Y(_15928_));
 AO21x1_ASAP7_75t_R _24331_ (.A1(_15483_),
    .A2(net3562),
    .B(_15490_),
    .Y(_15929_));
 AO21x1_ASAP7_75t_R _24332_ (.A1(_15550_),
    .A2(_15516_),
    .B(_15490_),
    .Y(_15930_));
 AND3x1_ASAP7_75t_R _24333_ (.A(_15929_),
    .B(_15930_),
    .C(_15751_),
    .Y(_15931_));
 AO21x1_ASAP7_75t_R _24334_ (.A1(_15540_),
    .A2(_15417_),
    .B(_15541_),
    .Y(_15932_));
 NOR2x1_ASAP7_75t_R _24335_ (.A(_15687_),
    .B(_15541_),
    .Y(_15933_));
 INVx1_ASAP7_75t_R _24336_ (.A(_15933_),
    .Y(_15934_));
 AND3x1_ASAP7_75t_R _24337_ (.A(_15932_),
    .B(_15450_),
    .C(_15934_),
    .Y(_15935_));
 AND5x2_ASAP7_75t_R _24338_ (.A(_15631_),
    .B(_15928_),
    .C(_15447_),
    .D(_15931_),
    .E(_15935_),
    .Y(_15936_));
 AO21x1_ASAP7_75t_R _24339_ (.A1(_15483_),
    .A2(_15516_),
    .B(_15618_),
    .Y(_15937_));
 AO21x1_ASAP7_75t_R _24340_ (.A1(_15687_),
    .A2(_15448_),
    .B(_15618_),
    .Y(_15938_));
 NAND2x1_ASAP7_75t_R _24341_ (.A(_15552_),
    .B(_15549_),
    .Y(_15939_));
 AND4x1_ASAP7_75t_R _24342_ (.A(_15937_),
    .B(_15938_),
    .C(_15738_),
    .D(_15939_),
    .Y(_15940_));
 NAND2x1_ASAP7_75t_R _24343_ (.A(_15697_),
    .B(_15602_),
    .Y(_15941_));
 AND4x1_ASAP7_75t_R _24344_ (.A(_15604_),
    .B(_15743_),
    .C(_15941_),
    .D(_15746_),
    .Y(_15942_));
 NOR2x2_ASAP7_75t_R _24345_ (.A(_15425_),
    .B(net3560),
    .Y(_15943_));
 NAND2x1_ASAP7_75t_R _24346_ (.A(_15943_),
    .B(_15602_),
    .Y(_15944_));
 AND5x2_ASAP7_75t_R _24347_ (.A(_15821_),
    .B(_15940_),
    .C(_15942_),
    .D(_15734_),
    .E(_15944_),
    .Y(_15945_));
 NAND3x2_ASAP7_75t_R _24348_ (.B(_15936_),
    .C(_15945_),
    .Y(_15946_),
    .A(_15926_));
 NOR2x1_ASAP7_75t_R _24349_ (.A(_15409_),
    .B(_15486_),
    .Y(_15947_));
 INVx1_ASAP7_75t_R _24350_ (.A(_15947_),
    .Y(_15948_));
 NAND2x1_ASAP7_75t_R _24351_ (.A(_15502_),
    .B(_15744_),
    .Y(_15949_));
 AND2x2_ASAP7_75t_R _24352_ (.A(_15463_),
    .B(_15502_),
    .Y(_15950_));
 INVx1_ASAP7_75t_R _24353_ (.A(_15950_),
    .Y(_15951_));
 AND5x1_ASAP7_75t_R _24354_ (.A(_15949_),
    .B(_15644_),
    .C(_15589_),
    .D(_15951_),
    .E(_15670_),
    .Y(_15952_));
 AO21x1_ASAP7_75t_R _24355_ (.A1(_15571_),
    .A2(net3541),
    .B(_15563_),
    .Y(_15953_));
 AO21x1_ASAP7_75t_R _24356_ (.A1(_15584_),
    .A2(_15505_),
    .B(_15563_),
    .Y(_15954_));
 NAND2x1_ASAP7_75t_R _24357_ (.A(_15424_),
    .B(_15549_),
    .Y(_15955_));
 AO21x1_ASAP7_75t_R _24358_ (.A1(_15516_),
    .A2(net3562),
    .B(_15563_),
    .Y(_15956_));
 AND4x1_ASAP7_75t_R _24359_ (.A(_15953_),
    .B(_15954_),
    .C(_15955_),
    .D(_15956_),
    .Y(_15957_));
 AO21x1_ASAP7_75t_R _24360_ (.A1(_15584_),
    .A2(_15687_),
    .B(_15476_),
    .Y(_15958_));
 NOR2x1_ASAP7_75t_R _24361_ (.A(_15476_),
    .B(_15515_),
    .Y(_15959_));
 INVx1_ASAP7_75t_R _24362_ (.A(_15959_),
    .Y(_15960_));
 OA211x2_ASAP7_75t_R _24363_ (.A1(net3541),
    .A2(_15476_),
    .B(_15958_),
    .C(_15960_),
    .Y(_15961_));
 AO21x1_ASAP7_75t_R _24364_ (.A1(_15687_),
    .A2(_15448_),
    .B(_15486_),
    .Y(_15962_));
 AND5x2_ASAP7_75t_R _24365_ (.A(_15948_),
    .B(_15952_),
    .C(_15957_),
    .D(_15961_),
    .E(_15962_),
    .Y(_15963_));
 OA211x2_ASAP7_75t_R _24366_ (.A1(_15469_),
    .A2(_15510_),
    .B(_15881_),
    .C(_15519_),
    .Y(_15964_));
 AND5x1_ASAP7_75t_R _24367_ (.A(_15613_),
    .B(_15964_),
    .C(_15704_),
    .D(_15707_),
    .E(_15887_),
    .Y(_15965_));
 AO21x1_ASAP7_75t_R _24368_ (.A1(_15584_),
    .A2(_15687_),
    .B(_15437_),
    .Y(_15966_));
 INVx1_ASAP7_75t_R _24369_ (.A(_15874_),
    .Y(_15967_));
 AND2x2_ASAP7_75t_R _24370_ (.A(_15966_),
    .B(_15967_),
    .Y(_15968_));
 AO21x1_ASAP7_75t_R _24371_ (.A1(_15698_),
    .A2(_15442_),
    .B(_15437_),
    .Y(_15969_));
 OA211x2_ASAP7_75t_R _24372_ (.A1(_15473_),
    .A2(_15437_),
    .B(_15968_),
    .C(_15969_),
    .Y(_15970_));
 NAND2x1_ASAP7_75t_R _24373_ (.A(_15583_),
    .B(_15597_),
    .Y(_15971_));
 OA211x2_ASAP7_75t_R _24374_ (.A1(_15505_),
    .A2(_15453_),
    .B(_15894_),
    .C(_15720_),
    .Y(_15972_));
 OA211x2_ASAP7_75t_R _24375_ (.A1(_15575_),
    .A2(_15453_),
    .B(_15726_),
    .C(_15895_),
    .Y(_15973_));
 NOR2x2_ASAP7_75t_R _24376_ (.A(_15524_),
    .B(_15436_),
    .Y(_15974_));
 NOR2x1_ASAP7_75t_R _24377_ (.A(_15608_),
    .B(_15524_),
    .Y(_15975_));
 NOR3x1_ASAP7_75t_R _24378_ (.A(_15867_),
    .B(_15974_),
    .C(_15975_),
    .Y(_15976_));
 AND5x1_ASAP7_75t_R _24379_ (.A(_15971_),
    .B(_15972_),
    .C(_15973_),
    .D(_15713_),
    .E(_15976_),
    .Y(_15977_));
 AND3x1_ASAP7_75t_R _24380_ (.A(_15965_),
    .B(_15970_),
    .C(_15977_),
    .Y(_15978_));
 NAND2x2_ASAP7_75t_R _24381_ (.A(_15963_),
    .B(_15978_),
    .Y(_15979_));
 NOR2x2_ASAP7_75t_R _24382_ (.A(_15946_),
    .B(_15979_),
    .Y(_15980_));
 BUFx2_ASAP7_75t_R output333 (.A(net333),
    .Y(text_out[50]));
 XOR2x2_ASAP7_75t_R _24384_ (.A(_00465_),
    .B(_00511_),
    .Y(_15982_));
 BUFx2_ASAP7_75t_R output332 (.A(net332),
    .Y(text_out[4]));
 XOR2x1_ASAP7_75t_R _24386_ (.A(_00394_),
    .Y(_15984_),
    .B(net3492));
 XNOR2x1_ASAP7_75t_R _24387_ (.B(_15984_),
    .Y(_15985_),
    .A(_15982_));
 XOR2x1_ASAP7_75t_R _24388_ (.A(_15980_),
    .Y(_15986_),
    .B(_15985_));
 AND2x2_ASAP7_75t_R _24389_ (.A(net402),
    .B(net4154),
    .Y(_15987_));
 AO21x1_ASAP7_75t_R _24390_ (.A1(_15986_),
    .A2(net398),
    .B(_15987_),
    .Y(_00363_));
 AO21x1_ASAP7_75t_R _24391_ (.A1(_15571_),
    .A2(_15505_),
    .B(_15499_),
    .Y(_15988_));
 INVx1_ASAP7_75t_R _24392_ (.A(_15482_),
    .Y(_15989_));
 AO21x1_ASAP7_75t_R _24393_ (.A1(_15528_),
    .A2(_15496_),
    .B(_15772_),
    .Y(_15990_));
 OA211x2_ASAP7_75t_R _24394_ (.A1(_15687_),
    .A2(_15772_),
    .B(_15989_),
    .C(_15990_),
    .Y(_15991_));
 AND3x1_ASAP7_75t_R _24395_ (.A(_15764_),
    .B(_15908_),
    .C(_15609_),
    .Y(_15992_));
 NAND2x1_ASAP7_75t_R _24396_ (.A(_15498_),
    .B(_15480_),
    .Y(_15993_));
 OA211x2_ASAP7_75t_R _24397_ (.A1(_15695_),
    .A2(_15499_),
    .B(_15993_),
    .C(_15794_),
    .Y(_15994_));
 AO21x1_ASAP7_75t_R _24398_ (.A1(_15584_),
    .A2(_15528_),
    .B(_15413_),
    .Y(_15995_));
 AO21x1_ASAP7_75t_R _24399_ (.A1(_15469_),
    .A2(_15695_),
    .B(_15413_),
    .Y(_15996_));
 AND3x1_ASAP7_75t_R _24400_ (.A(_15995_),
    .B(_15996_),
    .C(_15761_),
    .Y(_15997_));
 AND5x1_ASAP7_75t_R _24401_ (.A(_15988_),
    .B(_15991_),
    .C(_15992_),
    .D(_15994_),
    .E(_15997_),
    .Y(_15998_));
 AO21x1_ASAP7_75t_R _24402_ (.A1(_15540_),
    .A2(net3541),
    .B(_15490_),
    .Y(_15999_));
 AND2x2_ASAP7_75t_R _24403_ (.A(_15460_),
    .B(_15583_),
    .Y(_16000_));
 INVx1_ASAP7_75t_R _24404_ (.A(_16000_),
    .Y(_16001_));
 OA211x2_ASAP7_75t_R _24405_ (.A1(_15687_),
    .A2(_15490_),
    .B(_15999_),
    .C(_16001_),
    .Y(_16002_));
 AO21x1_ASAP7_75t_R _24406_ (.A1(_15483_),
    .A2(_15515_),
    .B(_15490_),
    .Y(_16003_));
 AO21x1_ASAP7_75t_R _24407_ (.A1(_15469_),
    .A2(_15442_),
    .B(_15541_),
    .Y(_16004_));
 AND5x1_ASAP7_75t_R _24408_ (.A(_15450_),
    .B(_16002_),
    .C(_15751_),
    .D(_16003_),
    .E(_16004_),
    .Y(_16005_));
 AND2x2_ASAP7_75t_R _24409_ (.A(_15552_),
    .B(_15504_),
    .Y(_16006_));
 INVx1_ASAP7_75t_R _24410_ (.A(_16006_),
    .Y(_16007_));
 AND4x1_ASAP7_75t_R _24411_ (.A(_15819_),
    .B(_15821_),
    .C(_15815_),
    .D(_15944_),
    .Y(_16008_));
 INVx2_ASAP7_75t_R _24412_ (.A(_15943_),
    .Y(_16009_));
 AO21x1_ASAP7_75t_R _24413_ (.A1(_15528_),
    .A2(_16009_),
    .B(_15618_),
    .Y(_16010_));
 AO21x1_ASAP7_75t_R _24414_ (.A1(_15469_),
    .A2(_15473_),
    .B(_15618_),
    .Y(_16011_));
 AND5x1_ASAP7_75t_R _24415_ (.A(_16007_),
    .B(_16008_),
    .C(_15937_),
    .D(_16010_),
    .E(_16011_),
    .Y(_16012_));
 AND3x2_ASAP7_75t_R _24416_ (.A(_15998_),
    .B(_16005_),
    .C(_16012_),
    .Y(_16013_));
 NAND2x1_ASAP7_75t_R _24417_ (.A(_15509_),
    .B(net3540),
    .Y(_16014_));
 AND4x1_ASAP7_75t_R _24418_ (.A(_15707_),
    .B(_15513_),
    .C(_15592_),
    .D(_16014_),
    .Y(_16015_));
 AO21x1_ASAP7_75t_R _24419_ (.A1(_15515_),
    .A2(net3562),
    .B(_15524_),
    .Y(_16016_));
 AO21x1_ASAP7_75t_R _24420_ (.A1(_15571_),
    .A2(_15417_),
    .B(_15524_),
    .Y(_16017_));
 NOR2x1_ASAP7_75t_R _24421_ (.A(_15524_),
    .B(_15505_),
    .Y(_16018_));
 INVx1_ASAP7_75t_R _24422_ (.A(_16018_),
    .Y(_16019_));
 INVx1_ASAP7_75t_R _24423_ (.A(_15525_),
    .Y(_16020_));
 INVx1_ASAP7_75t_R _24424_ (.A(_15974_),
    .Y(_16021_));
 AND5x1_ASAP7_75t_R _24425_ (.A(_16016_),
    .B(_16017_),
    .C(_16019_),
    .D(_16020_),
    .E(_16021_),
    .Y(_16022_));
 AO21x1_ASAP7_75t_R _24426_ (.A1(_15417_),
    .A2(net3541),
    .B(_15437_),
    .Y(_16023_));
 OA211x2_ASAP7_75t_R _24427_ (.A1(_15584_),
    .A2(_15437_),
    .B(_16023_),
    .C(_15535_),
    .Y(_16024_));
 AO21x1_ASAP7_75t_R _24428_ (.A1(_15473_),
    .A2(_15516_),
    .B(_15437_),
    .Y(_16025_));
 AO21x1_ASAP7_75t_R _24429_ (.A1(_15695_),
    .A2(_15698_),
    .B(_15453_),
    .Y(_16026_));
 AO21x1_ASAP7_75t_R _24430_ (.A1(_15417_),
    .A2(net3557),
    .B(_15453_),
    .Y(_16027_));
 OA211x2_ASAP7_75t_R _24431_ (.A1(_15442_),
    .A2(_15453_),
    .B(_16026_),
    .C(_16027_),
    .Y(_16028_));
 AND5x1_ASAP7_75t_R _24432_ (.A(_16015_),
    .B(_16022_),
    .C(_16024_),
    .D(_16025_),
    .E(_16028_),
    .Y(_16029_));
 AO21x1_ASAP7_75t_R _24433_ (.A1(_15858_),
    .A2(_15575_),
    .B(_15563_),
    .Y(_16030_));
 OA211x2_ASAP7_75t_R _24434_ (.A1(_15448_),
    .A2(_15563_),
    .B(_16030_),
    .C(_15650_),
    .Y(_16031_));
 NOR2x1_ASAP7_75t_R _24435_ (.A(net3558),
    .B(_15503_),
    .Y(_16032_));
 NAND2x1_ASAP7_75t_R _24436_ (.A(_15441_),
    .B(_16032_),
    .Y(_16033_));
 NOR2x1_ASAP7_75t_R _24437_ (.A(_15503_),
    .B(_15469_),
    .Y(_16034_));
 INVx1_ASAP7_75t_R _24438_ (.A(_16034_),
    .Y(_16035_));
 NAND2x1_ASAP7_75t_R _24439_ (.A(_15502_),
    .B(_15443_),
    .Y(_16036_));
 AND3x1_ASAP7_75t_R _24440_ (.A(_16035_),
    .B(_15949_),
    .C(_16036_),
    .Y(_16037_));
 AND4x1_ASAP7_75t_R _24441_ (.A(_16031_),
    .B(_15573_),
    .C(_16033_),
    .D(_16037_),
    .Y(_16038_));
 NAND2x1_ASAP7_75t_R _24442_ (.A(_15398_),
    .B(_15475_),
    .Y(_16039_));
 INVx1_ASAP7_75t_R _24443_ (.A(_15493_),
    .Y(_16040_));
 NOR2x1_ASAP7_75t_R _24444_ (.A(_15608_),
    .B(_15486_),
    .Y(_16041_));
 INVx1_ASAP7_75t_R _24445_ (.A(_16041_),
    .Y(_16042_));
 OA211x2_ASAP7_75t_R _24446_ (.A1(_15486_),
    .A2(_16040_),
    .B(_16042_),
    .C(_15677_),
    .Y(_16043_));
 OA211x2_ASAP7_75t_R _24447_ (.A1(_00443_),
    .A2(net3547),
    .B(_15475_),
    .C(_15416_),
    .Y(_16044_));
 INVx1_ASAP7_75t_R _24448_ (.A(_16044_),
    .Y(_16045_));
 AO21x1_ASAP7_75t_R _24449_ (.A1(_15550_),
    .A2(_15575_),
    .B(_15476_),
    .Y(_16046_));
 AND5x1_ASAP7_75t_R _24450_ (.A(_16039_),
    .B(_16043_),
    .C(_15681_),
    .D(_16045_),
    .E(_16046_),
    .Y(_16047_));
 AND3x2_ASAP7_75t_R _24451_ (.A(_16029_),
    .B(_16038_),
    .C(_16047_),
    .Y(_16048_));
 NAND2x2_ASAP7_75t_R _24452_ (.A(_16013_),
    .B(_16048_),
    .Y(_16049_));
 XNOR2x2_ASAP7_75t_R _24453_ (.A(_00464_),
    .B(_00510_),
    .Y(_16050_));
 BUFx2_ASAP7_75t_R output331 (.A(net331),
    .Y(text_out[49]));
 XOR2x1_ASAP7_75t_R _24455_ (.A(_00395_),
    .Y(_16052_),
    .B(net3500));
 XOR2x1_ASAP7_75t_R _24456_ (.A(_16050_),
    .Y(_16053_),
    .B(_16052_));
 XOR2x1_ASAP7_75t_R _24457_ (.A(_16049_),
    .Y(_16054_),
    .B(_16053_));
 NAND2x2_ASAP7_75t_R _24458_ (.A(net405),
    .B(net3873),
    .Y(_16055_));
 OAI21x1_ASAP7_75t_R _24459_ (.A1(net405),
    .A2(_16054_),
    .B(net3874),
    .Y(_00365_));
 INVx1_ASAP7_75t_R _24460_ (.A(net3659),
    .Y(_16056_));
 BUFx2_ASAP7_75t_R output330 (.A(net330),
    .Y(text_out[48]));
 BUFx2_ASAP7_75t_R output329 (.A(net329),
    .Y(text_out[47]));
 XOR2x1_ASAP7_75t_R _24463_ (.A(_00415_),
    .Y(_16059_),
    .B(net3497));
 INVx3_ASAP7_75t_R _24464_ (.A(_00463_),
    .Y(_16060_));
 XOR2x1_ASAP7_75t_R _24465_ (.A(_16059_),
    .Y(_16061_),
    .B(_16060_));
 INVx2_ASAP7_75t_R _24466_ (.A(_00490_),
    .Y(_16062_));
 XOR2x1_ASAP7_75t_R _24467_ (.A(_16061_),
    .Y(_16063_),
    .B(_16062_));
 NAND2x1_ASAP7_75t_R _24468_ (.A(_15509_),
    .B(_15912_),
    .Y(_16064_));
 AND3x1_ASAP7_75t_R _24469_ (.A(_15885_),
    .B(_15887_),
    .C(_16064_),
    .Y(_16065_));
 OA21x2_ASAP7_75t_R _24470_ (.A1(_15576_),
    .A2(_15472_),
    .B(_15404_),
    .Y(_16066_));
 AND3x1_ASAP7_75t_R _24471_ (.A(_15404_),
    .B(_15429_),
    .C(_15548_),
    .Y(_16067_));
 NOR3x1_ASAP7_75t_R _24472_ (.A(_16066_),
    .B(_15874_),
    .C(_16067_),
    .Y(_16068_));
 AND3x1_ASAP7_75t_R _24473_ (.A(_15520_),
    .B(_16065_),
    .C(_16068_),
    .Y(_16069_));
 AOI21x1_ASAP7_75t_R _24474_ (.A1(_15607_),
    .A2(_15436_),
    .B(_15524_),
    .Y(_16070_));
 OR3x1_ASAP7_75t_R _24475_ (.A(_16070_),
    .B(_15712_),
    .C(_16018_),
    .Y(_16071_));
 INVx1_ASAP7_75t_R _24476_ (.A(_16071_),
    .Y(_16072_));
 INVx1_ASAP7_75t_R _24477_ (.A(_15628_),
    .Y(_16073_));
 INVx1_ASAP7_75t_R _24478_ (.A(_15623_),
    .Y(_16074_));
 AO21x1_ASAP7_75t_R _24479_ (.A1(_15533_),
    .A2(net3541),
    .B(_15453_),
    .Y(_16075_));
 AND4x1_ASAP7_75t_R _24480_ (.A(_16073_),
    .B(_15891_),
    .C(_16074_),
    .D(_16075_),
    .Y(_16076_));
 AND3x1_ASAP7_75t_R _24481_ (.A(_16069_),
    .B(_16072_),
    .C(_16076_),
    .Y(_16077_));
 AND3x1_ASAP7_75t_R _24482_ (.A(_15566_),
    .B(_16042_),
    .C(_15678_),
    .Y(_16078_));
 NAND2x1_ASAP7_75t_R _24483_ (.A(_15686_),
    .B(_16078_),
    .Y(_16079_));
 NOR2x1_ASAP7_75t_R _24484_ (.A(net3555),
    .B(_15476_),
    .Y(_16080_));
 AO21x1_ASAP7_75t_R _24485_ (.A1(_15516_),
    .A2(net3563),
    .B(_15476_),
    .Y(_16081_));
 INVx1_ASAP7_75t_R _24486_ (.A(_16081_),
    .Y(_16082_));
 OR4x1_ASAP7_75t_R _24487_ (.A(_15843_),
    .B(_16080_),
    .C(_15680_),
    .D(_16082_),
    .Y(_16083_));
 NOR2x1_ASAP7_75t_R _24488_ (.A(_16079_),
    .B(_16083_),
    .Y(_16084_));
 AO221x1_ASAP7_75t_R _24489_ (.A1(_00443_),
    .A2(_15432_),
    .B1(_15442_),
    .B2(net3555),
    .C(_15563_),
    .Y(_16085_));
 AND3x1_ASAP7_75t_R _24490_ (.A(_16085_),
    .B(_15650_),
    .C(_15674_),
    .Y(_16086_));
 AO21x1_ASAP7_75t_R _24491_ (.A1(_15515_),
    .A2(_15516_),
    .B(_15503_),
    .Y(_16087_));
 AO21x1_ASAP7_75t_R _24492_ (.A1(_15473_),
    .A2(_15575_),
    .B(_15503_),
    .Y(_16088_));
 AO21x1_ASAP7_75t_R _24493_ (.A1(_15687_),
    .A2(_15448_),
    .B(_15503_),
    .Y(_16089_));
 AND4x1_ASAP7_75t_R _24494_ (.A(_16087_),
    .B(_16088_),
    .C(_16089_),
    .D(_15573_),
    .Y(_16090_));
 AND3x1_ASAP7_75t_R _24495_ (.A(_16084_),
    .B(_16086_),
    .C(_16090_),
    .Y(_16091_));
 AND2x2_ASAP7_75t_R _24496_ (.A(_16077_),
    .B(_16091_),
    .Y(_16092_));
 OA211x2_ASAP7_75t_R _24497_ (.A1(_15417_),
    .A2(_15499_),
    .B(_15916_),
    .C(_15768_),
    .Y(_16093_));
 AO21x1_ASAP7_75t_R _24498_ (.A1(_15469_),
    .A2(_15473_),
    .B(_15421_),
    .Y(_16094_));
 OA211x2_ASAP7_75t_R _24499_ (.A1(net3562),
    .A2(_15421_),
    .B(_16094_),
    .C(_15765_),
    .Y(_16095_));
 OA211x2_ASAP7_75t_R _24500_ (.A1(_15421_),
    .A2(_15571_),
    .B(_16093_),
    .C(_16095_),
    .Y(_16096_));
 OA211x2_ASAP7_75t_R _24501_ (.A1(net3544),
    .A2(net3550),
    .B(_15481_),
    .C(_15416_),
    .Y(_16097_));
 AND3x1_ASAP7_75t_R _24502_ (.A(_15481_),
    .B(_15433_),
    .C(_15425_),
    .Y(_16098_));
 OR3x1_ASAP7_75t_R _24503_ (.A(_16097_),
    .B(_16098_),
    .C(_15804_),
    .Y(_16099_));
 OR3x1_ASAP7_75t_R _24504_ (.A(_15413_),
    .B(_15425_),
    .C(_15442_),
    .Y(_16100_));
 NAND2x1_ASAP7_75t_R _24505_ (.A(_15762_),
    .B(_16100_),
    .Y(_16101_));
 INVx1_ASAP7_75t_R _24506_ (.A(_15913_),
    .Y(_16102_));
 OA211x2_ASAP7_75t_R _24507_ (.A1(_15425_),
    .A2(net3549),
    .B(_15412_),
    .C(_15435_),
    .Y(_16103_));
 OR4x1_ASAP7_75t_R _24508_ (.A(_16101_),
    .B(_16102_),
    .C(_15807_),
    .D(_16103_),
    .Y(_16104_));
 NOR2x1_ASAP7_75t_R _24509_ (.A(_16099_),
    .B(_16104_),
    .Y(_16105_));
 NAND2x2_ASAP7_75t_R _24510_ (.A(_16096_),
    .B(_16105_),
    .Y(_16106_));
 AND3x1_ASAP7_75t_R _24511_ (.A(_15934_),
    .B(_15828_),
    .C(_15596_),
    .Y(_16107_));
 AND3x1_ASAP7_75t_R _24512_ (.A(_15445_),
    .B(net3549),
    .C(_15398_),
    .Y(_16108_));
 INVx1_ASAP7_75t_R _24513_ (.A(_16108_),
    .Y(_16109_));
 AO21x1_ASAP7_75t_R _24514_ (.A1(_15448_),
    .A2(_16009_),
    .B(_15490_),
    .Y(_16110_));
 AND5x1_ASAP7_75t_R _24515_ (.A(_15825_),
    .B(_16107_),
    .C(_15930_),
    .D(_16109_),
    .E(_16110_),
    .Y(_16111_));
 OA31x2_ASAP7_75t_R _24516_ (.A1(net3540),
    .A2(_15583_),
    .A3(_15416_),
    .B1(_15602_),
    .Y(_16112_));
 INVx1_ASAP7_75t_R _24517_ (.A(_16112_),
    .Y(_16113_));
 NAND2x1_ASAP7_75t_R _24518_ (.A(_15602_),
    .B(_15514_),
    .Y(_16114_));
 AO21x1_ASAP7_75t_R _24519_ (.A1(_15695_),
    .A2(_15575_),
    .B(_15603_),
    .Y(_16115_));
 AO21x1_ASAP7_75t_R _24520_ (.A1(_15505_),
    .A2(net3561),
    .B(_15618_),
    .Y(_16116_));
 AO21x1_ASAP7_75t_R _24521_ (.A1(_15550_),
    .A2(_15698_),
    .B(_15618_),
    .Y(_16117_));
 AND5x1_ASAP7_75t_R _24522_ (.A(_16113_),
    .B(_16114_),
    .C(_16115_),
    .D(_16116_),
    .E(_16117_),
    .Y(_16118_));
 AND2x2_ASAP7_75t_R _24523_ (.A(_16111_),
    .B(_16118_),
    .Y(_16119_));
 INVx1_ASAP7_75t_R _24524_ (.A(_16119_),
    .Y(_16120_));
 NOR2x2_ASAP7_75t_R _24525_ (.A(_16106_),
    .B(_16120_),
    .Y(_16121_));
 NAND2x1_ASAP7_75t_R _24526_ (.A(_16092_),
    .B(_16121_),
    .Y(_16122_));
 NOR2x2_ASAP7_75t_R _24527_ (.A(_15657_),
    .B(_16122_),
    .Y(_16123_));
 NOR2x1_ASAP7_75t_R _24528_ (.A(_16063_),
    .B(_16123_),
    .Y(_16124_));
 AND2x2_ASAP7_75t_R _24529_ (.A(_16123_),
    .B(_16063_),
    .Y(_16125_));
 OAI21x1_ASAP7_75t_R _24530_ (.A1(_16124_),
    .A2(_16125_),
    .B(net398),
    .Y(_16126_));
 OAI21x1_ASAP7_75t_R _24531_ (.A1(net398),
    .A2(net3660),
    .B(_16126_),
    .Y(_00366_));
 INVx2_ASAP7_75t_R _24532_ (.A(net3970),
    .Y(_16127_));
 BUFx2_ASAP7_75t_R output328 (.A(net328),
    .Y(text_out[46]));
 XOR2x1_ASAP7_75t_R _24534_ (.A(_00416_),
    .Y(_16129_),
    .B(_00430_));
 INVx4_ASAP7_75t_R _24535_ (.A(_00462_),
    .Y(_16130_));
 XOR2x1_ASAP7_75t_R _24536_ (.A(_16129_),
    .Y(_16131_),
    .B(_16130_));
 INVx3_ASAP7_75t_R _24537_ (.A(_00489_),
    .Y(_16132_));
 XOR2x1_ASAP7_75t_R _24538_ (.A(_16131_),
    .Y(_16133_),
    .B(_16132_));
 INVx1_ASAP7_75t_R _24539_ (.A(_16133_),
    .Y(_16134_));
 INVx1_ASAP7_75t_R _24540_ (.A(_15657_),
    .Y(_16135_));
 AND3x1_ASAP7_75t_R _24541_ (.A(_15966_),
    .B(_15969_),
    .C(_15645_),
    .Y(_16136_));
 NOR2x1_ASAP7_75t_R _24542_ (.A(_15510_),
    .B(_15515_),
    .Y(_16137_));
 AOI211x1_ASAP7_75t_R _24543_ (.A1(_15576_),
    .A2(_15509_),
    .B(_16137_),
    .C(_15878_),
    .Y(_16138_));
 AND4x1_ASAP7_75t_R _24544_ (.A(_16136_),
    .B(_15885_),
    .C(_16014_),
    .D(_16138_),
    .Y(_16139_));
 NAND2x1_ASAP7_75t_R _24545_ (.A(_15744_),
    .B(_15597_),
    .Y(_16140_));
 NAND2x1_ASAP7_75t_R _24546_ (.A(_15536_),
    .B(_15597_),
    .Y(_16141_));
 AO21x1_ASAP7_75t_R _24547_ (.A1(_15417_),
    .A2(_15496_),
    .B(_15524_),
    .Y(_16142_));
 AND5x1_ASAP7_75t_R _24548_ (.A(_16140_),
    .B(_15641_),
    .C(_16141_),
    .D(_16142_),
    .E(_15598_),
    .Y(_16143_));
 NOR2x1_ASAP7_75t_R _24549_ (.A(_15727_),
    .B(_15725_),
    .Y(_16144_));
 AO21x1_ASAP7_75t_R _24550_ (.A1(_15528_),
    .A2(_15417_),
    .B(_15453_),
    .Y(_16145_));
 AND3x1_ASAP7_75t_R _24551_ (.A(_16144_),
    .B(_15893_),
    .C(_16145_),
    .Y(_16146_));
 NAND3x1_ASAP7_75t_R _24552_ (.A(_16139_),
    .B(_16143_),
    .C(_16146_),
    .Y(_16147_));
 NOR2x1_ASAP7_75t_R _24553_ (.A(_16032_),
    .B(_15950_),
    .Y(_16148_));
 NAND2x1_ASAP7_75t_R _24554_ (.A(_15502_),
    .B(_15399_),
    .Y(_16149_));
 AND4x1_ASAP7_75t_R _24555_ (.A(_16148_),
    .B(_16036_),
    .C(_16149_),
    .D(_16035_),
    .Y(_16150_));
 AND3x1_ASAP7_75t_R _24556_ (.A(_16150_),
    .B(_15651_),
    .C(_15859_),
    .Y(_16151_));
 INVx1_ASAP7_75t_R _24557_ (.A(_16151_),
    .Y(_16152_));
 INVx1_ASAP7_75t_R _24558_ (.A(_15488_),
    .Y(_16153_));
 AND3x1_ASAP7_75t_R _24559_ (.A(_15948_),
    .B(_16153_),
    .C(_15678_),
    .Y(_16154_));
 NAND2x1_ASAP7_75t_R _24560_ (.A(_15685_),
    .B(_16154_),
    .Y(_16155_));
 OA31x2_ASAP7_75t_R _24561_ (.A1(_15514_),
    .A2(_15744_),
    .A3(_15472_),
    .B1(_15475_),
    .Y(_16156_));
 AO21x1_ASAP7_75t_R _24562_ (.A1(_15505_),
    .A2(_15687_),
    .B(_15476_),
    .Y(_16157_));
 INVx1_ASAP7_75t_R _24563_ (.A(_16157_),
    .Y(_16158_));
 AO21x1_ASAP7_75t_R _24564_ (.A1(_15595_),
    .A2(_15475_),
    .B(_16158_),
    .Y(_16159_));
 OR3x1_ASAP7_75t_R _24565_ (.A(_16155_),
    .B(_16156_),
    .C(_16159_),
    .Y(_16160_));
 OR3x2_ASAP7_75t_R _24566_ (.A(_16147_),
    .B(_16152_),
    .C(_16160_),
    .Y(_16161_));
 AO21x1_ASAP7_75t_R _24567_ (.A1(_15571_),
    .A2(_15417_),
    .B(_15421_),
    .Y(_16162_));
 OA211x2_ASAP7_75t_R _24568_ (.A1(_15505_),
    .A2(_15421_),
    .B(_16162_),
    .C(_15909_),
    .Y(_16163_));
 AO21x1_ASAP7_75t_R _24569_ (.A1(_15695_),
    .A2(_15575_),
    .B(_15421_),
    .Y(_16164_));
 AND3x1_ASAP7_75t_R _24570_ (.A(_15792_),
    .B(_15765_),
    .C(_16164_),
    .Y(_16165_));
 AO21x1_ASAP7_75t_R _24571_ (.A1(_15540_),
    .A2(_15417_),
    .B(_15499_),
    .Y(_16166_));
 AND3x1_ASAP7_75t_R _24572_ (.A(_16166_),
    .B(_15770_),
    .C(_15993_),
    .Y(_16167_));
 AND3x1_ASAP7_75t_R _24573_ (.A(_16163_),
    .B(_16165_),
    .C(_16167_),
    .Y(_16168_));
 AO21x1_ASAP7_75t_R _24574_ (.A1(_15483_),
    .A2(_15516_),
    .B(_15772_),
    .Y(_16169_));
 NAND2x1_ASAP7_75t_R _24575_ (.A(_15481_),
    .B(_15612_),
    .Y(_16170_));
 AND4x1_ASAP7_75t_R _24576_ (.A(_16169_),
    .B(_15774_),
    .C(_15921_),
    .D(_16170_),
    .Y(_16171_));
 NAND2x1_ASAP7_75t_R _24577_ (.A(_15435_),
    .B(_15412_),
    .Y(_16172_));
 AO21x1_ASAP7_75t_R _24578_ (.A1(_15571_),
    .A2(_16009_),
    .B(_15413_),
    .Y(_16173_));
 AO21x1_ASAP7_75t_R _24579_ (.A1(_15505_),
    .A2(_15584_),
    .B(_15413_),
    .Y(_16174_));
 AND4x1_ASAP7_75t_R _24580_ (.A(_16100_),
    .B(_16172_),
    .C(_16173_),
    .D(_16174_),
    .Y(_16175_));
 AND3x1_ASAP7_75t_R _24581_ (.A(_16168_),
    .B(_16171_),
    .C(_16175_),
    .Y(_16176_));
 INVx1_ASAP7_75t_R _24582_ (.A(_16176_),
    .Y(_16177_));
 AOI21x1_ASAP7_75t_R _24583_ (.A1(_15549_),
    .A2(_15460_),
    .B(_15831_),
    .Y(_16178_));
 AO21x1_ASAP7_75t_R _24584_ (.A1(_15537_),
    .A2(_16009_),
    .B(_15490_),
    .Y(_16179_));
 OA211x2_ASAP7_75t_R _24585_ (.A1(_15425_),
    .A2(_15432_),
    .B(_15445_),
    .C(_15429_),
    .Y(_16180_));
 INVx1_ASAP7_75t_R _24586_ (.A(_16180_),
    .Y(_16181_));
 AO21x1_ASAP7_75t_R _24587_ (.A1(_15515_),
    .A2(_15575_),
    .B(_15541_),
    .Y(_16182_));
 AND4x1_ASAP7_75t_R _24588_ (.A(_16178_),
    .B(_16179_),
    .C(_16181_),
    .D(_16182_),
    .Y(_16183_));
 INVx1_ASAP7_75t_R _24589_ (.A(_15559_),
    .Y(_16184_));
 AO21x1_ASAP7_75t_R _24590_ (.A1(_15505_),
    .A2(_15448_),
    .B(_15618_),
    .Y(_16185_));
 OA211x2_ASAP7_75t_R _24591_ (.A1(_15618_),
    .A2(_15417_),
    .B(_16185_),
    .C(_15739_),
    .Y(_16186_));
 AO21x1_ASAP7_75t_R _24592_ (.A1(_15687_),
    .A2(net3541),
    .B(_15603_),
    .Y(_16187_));
 OA211x2_ASAP7_75t_R _24593_ (.A1(_15603_),
    .A2(_15695_),
    .B(_15745_),
    .C(_15941_),
    .Y(_16188_));
 AO21x1_ASAP7_75t_R _24594_ (.A1(_15695_),
    .A2(_15575_),
    .B(_15618_),
    .Y(_16189_));
 AND5x2_ASAP7_75t_R _24595_ (.A(_16184_),
    .B(_16186_),
    .C(_16187_),
    .D(_16188_),
    .E(_16189_),
    .Y(_16190_));
 NAND2x2_ASAP7_75t_R _24596_ (.A(_16183_),
    .B(_16190_),
    .Y(_16191_));
 NOR3x2_ASAP7_75t_R _24597_ (.B(_16177_),
    .C(_16191_),
    .Y(_16192_),
    .A(_16161_));
 NAND2x2_ASAP7_75t_R _24598_ (.A(_16135_),
    .B(_16192_),
    .Y(_16193_));
 NOR2x1_ASAP7_75t_R _24599_ (.A(_16134_),
    .B(_16193_),
    .Y(_16194_));
 AND2x2_ASAP7_75t_R _24600_ (.A(_16193_),
    .B(_16134_),
    .Y(_16195_));
 OAI21x1_ASAP7_75t_R _24601_ (.A1(_16194_),
    .A2(_16195_),
    .B(net398),
    .Y(_16196_));
 OAI21x1_ASAP7_75t_R _24602_ (.A1(net398),
    .A2(net3971),
    .B(_16196_),
    .Y(_00367_));
 OA211x2_ASAP7_75t_R _24603_ (.A1(_15425_),
    .A2(net3549),
    .B(_15460_),
    .C(_15435_),
    .Y(_16197_));
 INVx1_ASAP7_75t_R _24604_ (.A(_15748_),
    .Y(_16198_));
 OA21x2_ASAP7_75t_R _24605_ (.A1(_15527_),
    .A2(_15943_),
    .B(_15460_),
    .Y(_16199_));
 OR5x1_ASAP7_75t_R _24606_ (.A(_16000_),
    .B(_16197_),
    .C(_15832_),
    .D(_16198_),
    .E(_16199_),
    .Y(_16200_));
 AO21x1_ASAP7_75t_R _24607_ (.A1(_15744_),
    .A2(_15552_),
    .B(_15559_),
    .Y(_16201_));
 AND2x2_ASAP7_75t_R _24608_ (.A(_15399_),
    .B(_15552_),
    .Y(_16202_));
 INVx1_ASAP7_75t_R _24609_ (.A(_15554_),
    .Y(_16203_));
 INVx1_ASAP7_75t_R _24610_ (.A(_15939_),
    .Y(_16204_));
 OR5x1_ASAP7_75t_R _24611_ (.A(_16201_),
    .B(_16006_),
    .C(_16202_),
    .D(_16203_),
    .E(_16204_),
    .Y(_16205_));
 NAND2x1_ASAP7_75t_R _24612_ (.A(_15815_),
    .B(_15732_),
    .Y(_16206_));
 INVx1_ASAP7_75t_R _24613_ (.A(_16114_),
    .Y(_16207_));
 INVx1_ASAP7_75t_R _24614_ (.A(_15941_),
    .Y(_16208_));
 INVx1_ASAP7_75t_R _24615_ (.A(_15733_),
    .Y(_16209_));
 OR5x1_ASAP7_75t_R _24616_ (.A(_16206_),
    .B(_16207_),
    .C(_15742_),
    .D(_16208_),
    .E(_16209_),
    .Y(_16210_));
 AO21x1_ASAP7_75t_R _24617_ (.A1(_15468_),
    .A2(_15445_),
    .B(_16108_),
    .Y(_16211_));
 INVx1_ASAP7_75t_R _24618_ (.A(_15828_),
    .Y(_16212_));
 OA21x2_ASAP7_75t_R _24619_ (.A1(_15527_),
    .A2(_15943_),
    .B(_15445_),
    .Y(_16213_));
 OR3x1_ASAP7_75t_R _24620_ (.A(_16211_),
    .B(_16212_),
    .C(_16213_),
    .Y(_16214_));
 OR4x2_ASAP7_75t_R _24621_ (.A(_16200_),
    .B(_16205_),
    .C(_16210_),
    .D(_16214_),
    .Y(_16215_));
 AO221x1_ASAP7_75t_R _24622_ (.A1(_15425_),
    .A2(_15432_),
    .B1(_15442_),
    .B2(net3553),
    .C(_15772_),
    .Y(_16216_));
 AO21x1_ASAP7_75t_R _24623_ (.A1(_15516_),
    .A2(_15473_),
    .B(_15413_),
    .Y(_16217_));
 AO21x1_ASAP7_75t_R _24624_ (.A1(_16009_),
    .A2(_16040_),
    .B(_15413_),
    .Y(_16218_));
 AND4x1_ASAP7_75t_R _24625_ (.A(_16216_),
    .B(_16170_),
    .C(_16217_),
    .D(_16218_),
    .Y(_16219_));
 AO21x1_ASAP7_75t_R _24626_ (.A1(_15469_),
    .A2(_15575_),
    .B(_15421_),
    .Y(_16220_));
 OA211x2_ASAP7_75t_R _24627_ (.A1(_15584_),
    .A2(_15421_),
    .B(_16220_),
    .C(_16162_),
    .Y(_16221_));
 AO21x1_ASAP7_75t_R _24628_ (.A1(_15483_),
    .A2(net3562),
    .B(_15499_),
    .Y(_16222_));
 AO21x1_ASAP7_75t_R _24629_ (.A1(_15505_),
    .A2(_15687_),
    .B(_15499_),
    .Y(_16223_));
 AO21x1_ASAP7_75t_R _24630_ (.A1(_15571_),
    .A2(net3541),
    .B(_15499_),
    .Y(_16224_));
 AND5x2_ASAP7_75t_R _24631_ (.A(_15916_),
    .B(_16221_),
    .C(_16222_),
    .D(_16223_),
    .E(_16224_),
    .Y(_16225_));
 NAND2x2_ASAP7_75t_R _24632_ (.A(_16219_),
    .B(_16225_),
    .Y(_16226_));
 NOR2x2_ASAP7_75t_R _24633_ (.A(_16215_),
    .B(_16226_),
    .Y(_16227_));
 OA211x2_ASAP7_75t_R _24634_ (.A1(net3555),
    .A2(_15503_),
    .B(_15862_),
    .C(_16149_),
    .Y(_16228_));
 AO21x1_ASAP7_75t_R _24635_ (.A1(_15515_),
    .A2(net3562),
    .B(_15563_),
    .Y(_16229_));
 AO21x1_ASAP7_75t_R _24636_ (.A1(_15448_),
    .A2(_15687_),
    .B(_15563_),
    .Y(_16230_));
 AND3x1_ASAP7_75t_R _24637_ (.A(_16229_),
    .B(_15580_),
    .C(_16230_),
    .Y(_16231_));
 AND5x1_ASAP7_75t_R _24638_ (.A(_15569_),
    .B(_16228_),
    .C(_15669_),
    .D(_16089_),
    .E(_16231_),
    .Y(_16232_));
 AND4x1_ASAP7_75t_R _24639_ (.A(_16045_),
    .B(_15960_),
    .C(_15478_),
    .D(_16157_),
    .Y(_16233_));
 AO21x1_ASAP7_75t_R _24640_ (.A1(_15550_),
    .A2(_15695_),
    .B(_15486_),
    .Y(_16234_));
 AND5x1_ASAP7_75t_R _24641_ (.A(_15685_),
    .B(_15948_),
    .C(_15689_),
    .D(_16234_),
    .E(_15676_),
    .Y(_16235_));
 NAND3x1_ASAP7_75t_R _24642_ (.A(_16232_),
    .B(_16233_),
    .C(_16235_),
    .Y(_16236_));
 AO21x1_ASAP7_75t_R _24643_ (.A1(_15549_),
    .A2(_15509_),
    .B(_15878_),
    .Y(_16237_));
 INVx1_ASAP7_75t_R _24644_ (.A(_16064_),
    .Y(_16238_));
 OR5x1_ASAP7_75t_R _24645_ (.A(_16237_),
    .B(_16137_),
    .C(_15882_),
    .D(_16238_),
    .E(_15578_),
    .Y(_16239_));
 AO21x1_ASAP7_75t_R _24646_ (.A1(_15404_),
    .A2(_15595_),
    .B(_15874_),
    .Y(_16240_));
 AO21x1_ASAP7_75t_R _24647_ (.A1(net3540),
    .A2(_15404_),
    .B(_15876_),
    .Y(_16241_));
 AO21x1_ASAP7_75t_R _24648_ (.A1(_15468_),
    .A2(_15404_),
    .B(_15873_),
    .Y(_16242_));
 OR4x1_ASAP7_75t_R _24649_ (.A(_16240_),
    .B(_16241_),
    .C(_16242_),
    .D(_15406_),
    .Y(_16243_));
 AO21x1_ASAP7_75t_R _24650_ (.A1(_15912_),
    .A2(_15597_),
    .B(_15710_),
    .Y(_16244_));
 AO21x1_ASAP7_75t_R _24651_ (.A1(_15468_),
    .A2(_15597_),
    .B(_15975_),
    .Y(_16245_));
 AO21x1_ASAP7_75t_R _24652_ (.A1(_15454_),
    .A2(_15536_),
    .B(_15892_),
    .Y(_16246_));
 INVx1_ASAP7_75t_R _24653_ (.A(_16026_),
    .Y(_16247_));
 OR4x1_ASAP7_75t_R _24654_ (.A(_16246_),
    .B(_16247_),
    .C(_15725_),
    .D(_15723_),
    .Y(_16248_));
 OR5x1_ASAP7_75t_R _24655_ (.A(_16239_),
    .B(_16243_),
    .C(_16244_),
    .D(_16245_),
    .E(_16248_),
    .Y(_16249_));
 NOR2x1_ASAP7_75t_R _24656_ (.A(_16236_),
    .B(_16249_),
    .Y(_16250_));
 NAND2x2_ASAP7_75t_R _24657_ (.A(_16227_),
    .B(_16250_),
    .Y(_16251_));
 BUFx2_ASAP7_75t_R output327 (.A(net327),
    .Y(text_out[45]));
 XOR2x1_ASAP7_75t_R _24659_ (.A(_00396_),
    .Y(_16253_),
    .B(_00429_));
 XNOR2x2_ASAP7_75t_R _24660_ (.A(_00461_),
    .B(_00509_),
    .Y(_16254_));
 XNOR2x1_ASAP7_75t_R _24661_ (.B(_16254_),
    .Y(_16255_),
    .A(_16253_));
 XOR2x1_ASAP7_75t_R _24662_ (.A(_16251_),
    .Y(_16256_),
    .B(_16255_));
 AND2x2_ASAP7_75t_R _24663_ (.A(net402),
    .B(net4122),
    .Y(_16257_));
 AO21x1_ASAP7_75t_R _24664_ (.A1(_16256_),
    .A2(net398),
    .B(_16257_),
    .Y(_00368_));
 XOR2x2_ASAP7_75t_R _24665_ (.A(_00460_),
    .B(_00508_),
    .Y(_16258_));
 XOR2x1_ASAP7_75t_R _24666_ (.A(_00398_),
    .Y(_16259_),
    .B(net2128));
 XOR2x1_ASAP7_75t_R _24667_ (.A(_16258_),
    .Y(_16260_),
    .B(_16259_));
 XNOR2x1_ASAP7_75t_R _24668_ (.B(_16260_),
    .Y(_16261_),
    .A(_00397_));
 CKINVDCx12_ASAP7_75t_R _24669_ (.A(net3479),
    .Y(_16262_));
 NAND2x2_ASAP7_75t_R _24670_ (.A(net2207),
    .B(_16262_),
    .Y(_16263_));
 BUFx2_ASAP7_75t_R output326 (.A(net326),
    .Y(text_out[44]));
 NOR2x2_ASAP7_75t_R _24672_ (.A(_00433_),
    .B(_00434_),
    .Y(_16265_));
 INVx8_ASAP7_75t_R _24673_ (.A(_16265_),
    .Y(_16266_));
 NOR2x2_ASAP7_75t_R _24674_ (.A(_16263_),
    .B(_16266_),
    .Y(_16267_));
 INVx2_ASAP7_75t_R _24675_ (.A(_00430_),
    .Y(_16268_));
 NAND2x2_ASAP7_75t_R _24676_ (.A(_16268_),
    .B(_00429_),
    .Y(_16269_));
 INVx3_ASAP7_75t_R _24677_ (.A(net3495),
    .Y(_16270_));
 NAND2x2_ASAP7_75t_R _24678_ (.A(net3501),
    .B(_16270_),
    .Y(_16271_));
 NOR2x2_ASAP7_75t_R _24679_ (.A(_16269_),
    .B(_16271_),
    .Y(_16272_));
 AND2x2_ASAP7_75t_R _24680_ (.A(_16267_),
    .B(_16272_),
    .Y(_16273_));
 INVx1_ASAP7_75t_R _24681_ (.A(_16273_),
    .Y(_16274_));
 NAND2x2_ASAP7_75t_R _24682_ (.A(net3479),
    .B(net2207),
    .Y(_16275_));
 INVx4_ASAP7_75t_R _24683_ (.A(net3489),
    .Y(_16276_));
 NAND2x2_ASAP7_75t_R _24684_ (.A(_00434_),
    .B(_16276_),
    .Y(_16277_));
 NOR2x2_ASAP7_75t_R _24685_ (.A(_16275_),
    .B(_16277_),
    .Y(_16278_));
 CKINVDCx6p67_ASAP7_75t_R _24686_ (.A(_16278_),
    .Y(_16279_));
 BUFx2_ASAP7_75t_R output325 (.A(net325),
    .Y(text_out[43]));
 NOR2x2_ASAP7_75t_R _24688_ (.A(net2207),
    .B(net2665),
    .Y(_16281_));
 INVx1_ASAP7_75t_R _24689_ (.A(_16281_),
    .Y(_16282_));
 INVx5_ASAP7_75t_R _24690_ (.A(_16272_),
    .Y(_16283_));
 AO21x1_ASAP7_75t_R _24691_ (.A1(_16279_),
    .A2(_16282_),
    .B(_16283_),
    .Y(_16284_));
 NAND2x1_ASAP7_75t_R _24692_ (.A(_16274_),
    .B(_16284_),
    .Y(_16285_));
 INVx3_ASAP7_75t_R _24693_ (.A(net3484),
    .Y(_16286_));
 CKINVDCx10_ASAP7_75t_R _24694_ (.A(net2207),
    .Y(_16287_));
 OA211x2_ASAP7_75t_R _24695_ (.A1(_16286_),
    .A2(_16287_),
    .B(_16272_),
    .C(_00433_),
    .Y(_16288_));
 OR2x2_ASAP7_75t_R _24696_ (.A(_16285_),
    .B(_16288_),
    .Y(_16289_));
 NOR2x2_ASAP7_75t_R _24697_ (.A(net3494),
    .B(_00432_),
    .Y(_16290_));
 CKINVDCx5p33_ASAP7_75t_R _24698_ (.A(_00429_),
    .Y(_16291_));
 NOR2x1_ASAP7_75t_R _24699_ (.A(_00430_),
    .B(_16291_),
    .Y(_16292_));
 NAND2x2_ASAP7_75t_R _24700_ (.A(_16290_),
    .B(_16292_),
    .Y(_16293_));
 INVx3_ASAP7_75t_R _24701_ (.A(_16293_),
    .Y(_16294_));
 NAND2x2_ASAP7_75t_R _24702_ (.A(_00433_),
    .B(_00434_),
    .Y(_16295_));
 CKINVDCx8_ASAP7_75t_R _24703_ (.A(_16295_),
    .Y(_16296_));
 BUFx2_ASAP7_75t_R output324 (.A(net324),
    .Y(text_out[42]));
 AND3x1_ASAP7_75t_R _24705_ (.A(_16294_),
    .B(net2158),
    .C(_16296_),
    .Y(_16298_));
 NOR2x2_ASAP7_75t_R _24706_ (.A(net3477),
    .B(net2204),
    .Y(_16299_));
 INVx6_ASAP7_75t_R _24707_ (.A(_16299_),
    .Y(_16300_));
 NAND2x2_ASAP7_75t_R _24708_ (.A(net2587),
    .B(_16300_),
    .Y(_16301_));
 NAND2x2_ASAP7_75t_R _24709_ (.A(_16265_),
    .B(_16294_),
    .Y(_16302_));
 NOR2x1_ASAP7_75t_R _24710_ (.A(_16301_),
    .B(_16302_),
    .Y(_16303_));
 NAND2x2_ASAP7_75t_R _24711_ (.A(net3489),
    .B(_16286_),
    .Y(_16304_));
 BUFx2_ASAP7_75t_R output323 (.A(net323),
    .Y(text_out[41]));
 INVx6_ASAP7_75t_R _24713_ (.A(net2765),
    .Y(_16306_));
 BUFx2_ASAP7_75t_R output322 (.A(net322),
    .Y(text_out[40]));
 NAND2x1_ASAP7_75t_R _24715_ (.A(_16306_),
    .B(_16294_),
    .Y(_16308_));
 NOR2x1_ASAP7_75t_R _24716_ (.A(net2206),
    .B(_16308_),
    .Y(_16309_));
 BUFx2_ASAP7_75t_R output321 (.A(net321),
    .Y(text_out[3]));
 NOR2x2_ASAP7_75t_R _24718_ (.A(_16277_),
    .B(_16300_),
    .Y(_16311_));
 INVx4_ASAP7_75t_R _24719_ (.A(_16311_),
    .Y(_16312_));
 NOR2x1_ASAP7_75t_R _24720_ (.A(_16293_),
    .B(_16312_),
    .Y(_16313_));
 OR4x1_ASAP7_75t_R _24721_ (.A(_16298_),
    .B(_16303_),
    .C(_16309_),
    .D(_16313_),
    .Y(_16314_));
 NOR2x1_ASAP7_75t_R _24722_ (.A(_16289_),
    .B(_16314_),
    .Y(_16315_));
 NAND2x2_ASAP7_75t_R _24723_ (.A(net3494),
    .B(_00432_),
    .Y(_16316_));
 NOR2x2_ASAP7_75t_R _24724_ (.A(_16316_),
    .B(_16269_),
    .Y(_16317_));
 NOR2x2_ASAP7_75t_R _24725_ (.A(_16275_),
    .B(_16304_),
    .Y(_16318_));
 AND2x2_ASAP7_75t_R _24726_ (.A(_16317_),
    .B(net2622),
    .Y(_16319_));
 BUFx2_ASAP7_75t_R output320 (.A(net320),
    .Y(text_out[39]));
 NAND2x2_ASAP7_75t_R _24728_ (.A(net3479),
    .B(_16287_),
    .Y(_16321_));
 NOR2x2_ASAP7_75t_R _24729_ (.A(_16295_),
    .B(_16321_),
    .Y(_16322_));
 AND2x2_ASAP7_75t_R _24730_ (.A(_16317_),
    .B(_16322_),
    .Y(_16323_));
 NOR2x2_ASAP7_75t_R _24731_ (.A(_16275_),
    .B(_16295_),
    .Y(_16324_));
 INVx11_ASAP7_75t_R _24732_ (.A(_16324_),
    .Y(_16325_));
 BUFx2_ASAP7_75t_R output319 (.A(net319),
    .Y(text_out[38]));
 CKINVDCx5p33_ASAP7_75t_R _24734_ (.A(_16317_),
    .Y(_16327_));
 BUFx2_ASAP7_75t_R output318 (.A(net318),
    .Y(text_out[37]));
 NOR2x1_ASAP7_75t_R _24736_ (.A(_16325_),
    .B(_16327_),
    .Y(_16329_));
 OR3x1_ASAP7_75t_R _24737_ (.A(_16319_),
    .B(_16323_),
    .C(_16329_),
    .Y(_16330_));
 BUFx2_ASAP7_75t_R output317 (.A(net317),
    .Y(text_out[36]));
 AND3x1_ASAP7_75t_R _24739_ (.A(_16317_),
    .B(net2205),
    .C(_16265_),
    .Y(_16332_));
 AND2x2_ASAP7_75t_R _24740_ (.A(_16317_),
    .B(_16281_),
    .Y(_16333_));
 NOR2x2_ASAP7_75t_R _24741_ (.A(net2277),
    .B(_16266_),
    .Y(_16334_));
 CKINVDCx8_ASAP7_75t_R _24742_ (.A(_16334_),
    .Y(_16335_));
 NOR2x1_ASAP7_75t_R _24743_ (.A(_16327_),
    .B(_16335_),
    .Y(_16336_));
 OR3x1_ASAP7_75t_R _24744_ (.A(_16332_),
    .B(_16333_),
    .C(_16336_),
    .Y(_16337_));
 NOR2x1_ASAP7_75t_R _24745_ (.A(_16330_),
    .B(_16337_),
    .Y(_16338_));
 INVx2_ASAP7_75t_R _24746_ (.A(_00432_),
    .Y(_16339_));
 NAND2x2_ASAP7_75t_R _24747_ (.A(net3494),
    .B(_16339_),
    .Y(_16340_));
 NOR2x2_ASAP7_75t_R _24748_ (.A(_16340_),
    .B(_16269_),
    .Y(_16341_));
 CKINVDCx5p33_ASAP7_75t_R _24749_ (.A(_16341_),
    .Y(_16342_));
 BUFx2_ASAP7_75t_R output316 (.A(net316),
    .Y(text_out[35]));
 NOR2x2_ASAP7_75t_R _24751_ (.A(net3480),
    .B(_16304_),
    .Y(_16344_));
 AND2x2_ASAP7_75t_R _24752_ (.A(_16341_),
    .B(_16344_),
    .Y(_16345_));
 AND3x1_ASAP7_75t_R _24753_ (.A(_16341_),
    .B(net2158),
    .C(_16296_),
    .Y(_16346_));
 NOR2x1_ASAP7_75t_R _24754_ (.A(_16345_),
    .B(_16346_),
    .Y(_16347_));
 AND2x6_ASAP7_75t_R _24755_ (.A(_16299_),
    .B(_16265_),
    .Y(_16348_));
 NAND2x1_ASAP7_75t_R _24756_ (.A(_16341_),
    .B(_16348_),
    .Y(_16349_));
 OA211x2_ASAP7_75t_R _24757_ (.A1(_16342_),
    .A2(_16282_),
    .B(_16347_),
    .C(_16349_),
    .Y(_16350_));
 AND3x1_ASAP7_75t_R _24758_ (.A(_16315_),
    .B(_16338_),
    .C(_16350_),
    .Y(_16351_));
 NAND2x2_ASAP7_75t_R _24759_ (.A(_00429_),
    .B(_00430_),
    .Y(_16352_));
 NOR2x2_ASAP7_75t_R _24760_ (.A(_16352_),
    .B(_16316_),
    .Y(_16353_));
 INVx6_ASAP7_75t_R _24761_ (.A(_16353_),
    .Y(_16354_));
 BUFx2_ASAP7_75t_R output315 (.A(net315),
    .Y(text_out[34]));
 NOR2x2_ASAP7_75t_R _24763_ (.A(net2278),
    .B(_16304_),
    .Y(_16356_));
 CKINVDCx11_ASAP7_75t_R _24764_ (.A(_16356_),
    .Y(_16357_));
 BUFx2_ASAP7_75t_R output314 (.A(net314),
    .Y(text_out[33]));
 BUFx2_ASAP7_75t_R output313 (.A(net313),
    .Y(text_out[32]));
 AND3x1_ASAP7_75t_R _24767_ (.A(_16353_),
    .B(_16262_),
    .C(_16306_),
    .Y(_16360_));
 INVx1_ASAP7_75t_R _24768_ (.A(_16360_),
    .Y(_16361_));
 NOR2x2_ASAP7_75t_R _24769_ (.A(net3479),
    .B(_16295_),
    .Y(_16362_));
 NAND2x1_ASAP7_75t_R _24770_ (.A(_16362_),
    .B(_16353_),
    .Y(_16363_));
 OA211x2_ASAP7_75t_R _24771_ (.A1(_16354_),
    .A2(_16357_),
    .B(_16361_),
    .C(_16363_),
    .Y(_16364_));
 BUFx2_ASAP7_75t_R output312 (.A(net312),
    .Y(text_out[31]));
 CKINVDCx9p33_ASAP7_75t_R _24773_ (.A(_16267_),
    .Y(_16366_));
 BUFx2_ASAP7_75t_R output311 (.A(net311),
    .Y(text_out[30]));
 AO21x1_ASAP7_75t_R _24775_ (.A1(_16335_),
    .A2(_16366_),
    .B(_16354_),
    .Y(_16368_));
 NOR2x2_ASAP7_75t_R _24776_ (.A(_00435_),
    .B(_16277_),
    .Y(_16369_));
 INVx4_ASAP7_75t_R _24777_ (.A(_16369_),
    .Y(_16370_));
 NOR2x1_ASAP7_75t_R _24778_ (.A(_16354_),
    .B(_16370_),
    .Y(_16371_));
 INVx1_ASAP7_75t_R _24779_ (.A(_16371_),
    .Y(_16372_));
 NOR2x2_ASAP7_75t_R _24780_ (.A(_16277_),
    .B(net2278),
    .Y(_16373_));
 NAND2x1_ASAP7_75t_R _24781_ (.A(_16353_),
    .B(_16373_),
    .Y(_16374_));
 AND3x1_ASAP7_75t_R _24782_ (.A(_16368_),
    .B(_16372_),
    .C(_16374_),
    .Y(_16375_));
 NOR2x2_ASAP7_75t_R _24783_ (.A(_16352_),
    .B(_16340_),
    .Y(_16376_));
 INVx1_ASAP7_75t_R _24784_ (.A(_16301_),
    .Y(_16377_));
 CKINVDCx8_ASAP7_75t_R _24785_ (.A(_16376_),
    .Y(_16378_));
 BUFx2_ASAP7_75t_R output310 (.A(net310),
    .Y(text_out[2]));
 NOR2x1_ASAP7_75t_R _24787_ (.A(net2766),
    .B(_16378_),
    .Y(_16380_));
 INVx5_ASAP7_75t_R _24788_ (.A(net2666),
    .Y(_16381_));
 NAND2x1_ASAP7_75t_R _24789_ (.A(_16381_),
    .B(_16376_),
    .Y(_16382_));
 NOR2x1_ASAP7_75t_R _24790_ (.A(_16377_),
    .B(_16382_),
    .Y(_16383_));
 AOI221x1_ASAP7_75t_R _24791_ (.A1(_16376_),
    .A2(_16362_),
    .B1(_16377_),
    .B2(_16380_),
    .C(_16383_),
    .Y(_16384_));
 AND3x1_ASAP7_75t_R _24792_ (.A(_16364_),
    .B(_16375_),
    .C(_16384_),
    .Y(_16385_));
 NOR2x2_ASAP7_75t_R _24793_ (.A(_16263_),
    .B(_16304_),
    .Y(_16386_));
 CKINVDCx8_ASAP7_75t_R _24794_ (.A(_16386_),
    .Y(_16387_));
 BUFx2_ASAP7_75t_R output309 (.A(net309),
    .Y(text_out[29]));
 BUFx2_ASAP7_75t_R output308 (.A(net308),
    .Y(text_out[28]));
 NOR2x2_ASAP7_75t_R _24797_ (.A(_16352_),
    .B(_16271_),
    .Y(_16390_));
 INVx5_ASAP7_75t_R _24798_ (.A(_16390_),
    .Y(_16391_));
 BUFx2_ASAP7_75t_R output307 (.A(net307),
    .Y(text_out[27]));
 AO21x1_ASAP7_75t_R _24800_ (.A1(_16387_),
    .A2(_16357_),
    .B(_16391_),
    .Y(_16393_));
 NOR2x2_ASAP7_75t_R _24801_ (.A(net2587),
    .B(_16266_),
    .Y(_16394_));
 CKINVDCx5p33_ASAP7_75t_R _24802_ (.A(_16394_),
    .Y(_16395_));
 BUFx2_ASAP7_75t_R output306 (.A(net306),
    .Y(text_out[26]));
 NOR2x2_ASAP7_75t_R _24804_ (.A(net3482),
    .B(_16266_),
    .Y(_16397_));
 CKINVDCx5p33_ASAP7_75t_R _24805_ (.A(_16397_),
    .Y(_16398_));
 BUFx2_ASAP7_75t_R output305 (.A(net305),
    .Y(text_out[25]));
 AO21x1_ASAP7_75t_R _24807_ (.A1(_16395_),
    .A2(_16398_),
    .B(_16391_),
    .Y(_16400_));
 BUFx2_ASAP7_75t_R output304 (.A(net304),
    .Y(text_out[24]));
 AND3x1_ASAP7_75t_R _24809_ (.A(_16390_),
    .B(_16300_),
    .C(_16296_),
    .Y(_16402_));
 INVx1_ASAP7_75t_R _24810_ (.A(_16402_),
    .Y(_16403_));
 INVx3_ASAP7_75t_R _24811_ (.A(net2587),
    .Y(_16404_));
 NAND2x1_ASAP7_75t_R _24812_ (.A(_16381_),
    .B(_16390_),
    .Y(_16405_));
 NOR2x1_ASAP7_75t_R _24813_ (.A(_16404_),
    .B(_16405_),
    .Y(_16406_));
 INVx1_ASAP7_75t_R _24814_ (.A(_16406_),
    .Y(_16407_));
 AND4x1_ASAP7_75t_R _24815_ (.A(_16393_),
    .B(_16400_),
    .C(_16403_),
    .D(_16407_),
    .Y(_16408_));
 AND3x4_ASAP7_75t_R _24816_ (.A(_16290_),
    .B(_00429_),
    .C(_00430_),
    .Y(_16409_));
 BUFx2_ASAP7_75t_R output303 (.A(net303),
    .Y(text_out[23]));
 INVx6_ASAP7_75t_R _24818_ (.A(_16409_),
    .Y(_16411_));
 BUFx2_ASAP7_75t_R output302 (.A(net302),
    .Y(text_out[22]));
 NOR2x1_ASAP7_75t_R _24820_ (.A(_16387_),
    .B(_16411_),
    .Y(_16413_));
 AND3x1_ASAP7_75t_R _24821_ (.A(_16409_),
    .B(_16287_),
    .C(_16296_),
    .Y(_16414_));
 INVx1_ASAP7_75t_R _24822_ (.A(_16414_),
    .Y(_16415_));
 NOR2x2_ASAP7_75t_R _24823_ (.A(net2840),
    .B(_16263_),
    .Y(_16416_));
 NAND2x1_ASAP7_75t_R _24824_ (.A(_16416_),
    .B(_16409_),
    .Y(_16417_));
 AND2x2_ASAP7_75t_R _24825_ (.A(_16415_),
    .B(_16417_),
    .Y(_16418_));
 INVx1_ASAP7_75t_R _24826_ (.A(_16418_),
    .Y(_16419_));
 NOR2x1_ASAP7_75t_R _24827_ (.A(_16413_),
    .B(_16419_),
    .Y(_16420_));
 CKINVDCx6p67_ASAP7_75t_R _24828_ (.A(_16348_),
    .Y(_16421_));
 BUFx2_ASAP7_75t_R output301 (.A(net301),
    .Y(text_out[21]));
 NOR2x1_ASAP7_75t_R _24830_ (.A(_16421_),
    .B(_16411_),
    .Y(_16423_));
 INVx1_ASAP7_75t_R _24831_ (.A(_16423_),
    .Y(_16424_));
 NOR2x2_ASAP7_75t_R _24832_ (.A(_16262_),
    .B(_16266_),
    .Y(_16425_));
 INVx2_ASAP7_75t_R _24833_ (.A(_16425_),
    .Y(_16426_));
 NOR2x1_ASAP7_75t_R _24834_ (.A(_16426_),
    .B(_16411_),
    .Y(_16427_));
 INVx1_ASAP7_75t_R _24835_ (.A(_16427_),
    .Y(_16428_));
 OA211x2_ASAP7_75t_R _24836_ (.A1(_16279_),
    .A2(_16411_),
    .B(_16424_),
    .C(_16428_),
    .Y(_16429_));
 AND3x1_ASAP7_75t_R _24837_ (.A(_16408_),
    .B(_16420_),
    .C(_16429_),
    .Y(_16430_));
 AND3x1_ASAP7_75t_R _24838_ (.A(_16351_),
    .B(_16385_),
    .C(_16430_),
    .Y(_16431_));
 INVx1_ASAP7_75t_R _24839_ (.A(_16431_),
    .Y(_16432_));
 NOR2x2_ASAP7_75t_R _24840_ (.A(_00429_),
    .B(_00430_),
    .Y(_16433_));
 AND2x6_ASAP7_75t_R _24841_ (.A(_16433_),
    .B(_16290_),
    .Y(_16434_));
 NAND2x1_ASAP7_75t_R _24842_ (.A(_16278_),
    .B(_16434_),
    .Y(_16435_));
 CKINVDCx5p33_ASAP7_75t_R _24843_ (.A(_16373_),
    .Y(_16436_));
 INVx5_ASAP7_75t_R _24844_ (.A(_16434_),
    .Y(_16437_));
 BUFx2_ASAP7_75t_R output300 (.A(net300),
    .Y(text_out[20]));
 AO21x1_ASAP7_75t_R _24846_ (.A1(_16436_),
    .A2(_16370_),
    .B(_16437_),
    .Y(_16439_));
 INVx11_ASAP7_75t_R _24847_ (.A(_16322_),
    .Y(_16440_));
 BUFx2_ASAP7_75t_R output299 (.A(net299),
    .Y(text_out[1]));
 BUFx2_ASAP7_75t_R output298 (.A(net298),
    .Y(text_out[19]));
 INVx5_ASAP7_75t_R _24850_ (.A(_16362_),
    .Y(_16443_));
 AO21x1_ASAP7_75t_R _24851_ (.A1(_16440_),
    .A2(_16443_),
    .B(_16437_),
    .Y(_16444_));
 CKINVDCx9p33_ASAP7_75t_R _24852_ (.A(_16318_),
    .Y(_16445_));
 NOR2x1_ASAP7_75t_R _24853_ (.A(_16445_),
    .B(_16437_),
    .Y(_16446_));
 INVx1_ASAP7_75t_R _24854_ (.A(_16446_),
    .Y(_16447_));
 AND2x2_ASAP7_75t_R _24855_ (.A(_16434_),
    .B(net3498),
    .Y(_16448_));
 INVx1_ASAP7_75t_R _24856_ (.A(_16448_),
    .Y(_16449_));
 AND5x1_ASAP7_75t_R _24857_ (.A(_16435_),
    .B(_16439_),
    .C(_16444_),
    .D(_16447_),
    .E(_16449_),
    .Y(_16450_));
 INVx3_ASAP7_75t_R _24858_ (.A(_16433_),
    .Y(_16451_));
 NOR2x2_ASAP7_75t_R _24859_ (.A(_16316_),
    .B(_16451_),
    .Y(_16452_));
 BUFx2_ASAP7_75t_R output297 (.A(net297),
    .Y(text_out[18]));
 OA211x2_ASAP7_75t_R _24861_ (.A1(net1854),
    .A2(net2209),
    .B(_16452_),
    .C(_16265_),
    .Y(_16454_));
 INVx1_ASAP7_75t_R _24862_ (.A(_16454_),
    .Y(_16455_));
 NAND2x1_ASAP7_75t_R _24863_ (.A(_16416_),
    .B(_16452_),
    .Y(_16456_));
 NAND2x1_ASAP7_75t_R _24864_ (.A(_16281_),
    .B(_16452_),
    .Y(_16457_));
 AND3x1_ASAP7_75t_R _24865_ (.A(_16455_),
    .B(_16456_),
    .C(_16457_),
    .Y(_16458_));
 NOR2x2_ASAP7_75t_R _24866_ (.A(_16340_),
    .B(_16451_),
    .Y(_16459_));
 CKINVDCx5p33_ASAP7_75t_R _24867_ (.A(_16459_),
    .Y(_16460_));
 BUFx2_ASAP7_75t_R output296 (.A(net296),
    .Y(text_out[17]));
 AO21x1_ASAP7_75t_R _24869_ (.A1(_16335_),
    .A2(_16366_),
    .B(_16460_),
    .Y(_16462_));
 INVx6_ASAP7_75t_R _24870_ (.A(_16416_),
    .Y(_16463_));
 BUFx2_ASAP7_75t_R output295 (.A(net295),
    .Y(text_out[16]));
 AO21x1_ASAP7_75t_R _24872_ (.A1(_16357_),
    .A2(_16463_),
    .B(_16460_),
    .Y(_16465_));
 OA211x2_ASAP7_75t_R _24873_ (.A1(net3493),
    .A2(_16460_),
    .B(_16462_),
    .C(_16465_),
    .Y(_16466_));
 NOR2x2_ASAP7_75t_R _24874_ (.A(_16271_),
    .B(_16451_),
    .Y(_16467_));
 BUFx2_ASAP7_75t_R output294 (.A(net294),
    .Y(text_out[15]));
 NAND2x2_ASAP7_75t_R _24876_ (.A(_16299_),
    .B(_16296_),
    .Y(_16469_));
 BUFx2_ASAP7_75t_R output293 (.A(net293),
    .Y(text_out[14]));
 INVx4_ASAP7_75t_R _24878_ (.A(_16467_),
    .Y(_16471_));
 NOR2x1_ASAP7_75t_R _24879_ (.A(_16469_),
    .B(_16471_),
    .Y(_16472_));
 AO21x1_ASAP7_75t_R _24880_ (.A1(_16324_),
    .A2(_16467_),
    .B(_16472_),
    .Y(_16473_));
 AND3x1_ASAP7_75t_R _24881_ (.A(_16467_),
    .B(_16381_),
    .C(net2278),
    .Y(_16474_));
 BUFx2_ASAP7_75t_R output292 (.A(net292),
    .Y(text_out[13]));
 AO21x1_ASAP7_75t_R _24883_ (.A1(_16357_),
    .A2(_16445_),
    .B(_16471_),
    .Y(_16476_));
 INVx1_ASAP7_75t_R _24884_ (.A(_16476_),
    .Y(_16477_));
 BUFx2_ASAP7_75t_R output291 (.A(net291),
    .Y(text_out[12]));
 AND3x1_ASAP7_75t_R _24886_ (.A(_16467_),
    .B(_16287_),
    .C(_16265_),
    .Y(_16479_));
 OR4x1_ASAP7_75t_R _24887_ (.A(_16473_),
    .B(_16474_),
    .C(_16477_),
    .D(_16479_),
    .Y(_16480_));
 INVx1_ASAP7_75t_R _24888_ (.A(_16480_),
    .Y(_16481_));
 AND4x1_ASAP7_75t_R _24889_ (.A(_16450_),
    .B(_16458_),
    .C(_16466_),
    .D(_16481_),
    .Y(_16482_));
 NAND2x2_ASAP7_75t_R _24890_ (.A(_00430_),
    .B(_16291_),
    .Y(_16483_));
 NOR2x2_ASAP7_75t_R _24891_ (.A(_16316_),
    .B(_16483_),
    .Y(_16484_));
 AND3x1_ASAP7_75t_R _24892_ (.A(_16484_),
    .B(net2588),
    .C(_16265_),
    .Y(_16485_));
 INVx1_ASAP7_75t_R _24893_ (.A(_16485_),
    .Y(_16486_));
 NOR2x2_ASAP7_75t_R _24894_ (.A(_16340_),
    .B(_16483_),
    .Y(_16487_));
 INVx5_ASAP7_75t_R _24895_ (.A(_16487_),
    .Y(_16488_));
 BUFx2_ASAP7_75t_R output290 (.A(net290),
    .Y(text_out[127]));
 AO21x1_ASAP7_75t_R _24897_ (.A1(_16440_),
    .A2(_16463_),
    .B(_16488_),
    .Y(_16490_));
 OA21x2_ASAP7_75t_R _24898_ (.A1(_16488_),
    .A2(_16398_),
    .B(_16490_),
    .Y(_16491_));
 BUFx2_ASAP7_75t_R output289 (.A(net289),
    .Y(text_out[126]));
 OA211x2_ASAP7_75t_R _24900_ (.A1(net1854),
    .A2(_16287_),
    .B(_16484_),
    .C(_16306_),
    .Y(_16493_));
 INVx1_ASAP7_75t_R _24901_ (.A(_16493_),
    .Y(_16494_));
 INVx4_ASAP7_75t_R _24902_ (.A(_16484_),
    .Y(_16495_));
 BUFx2_ASAP7_75t_R output288 (.A(net288),
    .Y(text_out[125]));
 AO21x1_ASAP7_75t_R _24904_ (.A1(_16312_),
    .A2(_16436_),
    .B(_16495_),
    .Y(_16497_));
 BUFx2_ASAP7_75t_R output287 (.A(net287),
    .Y(text_out[124]));
 AO21x1_ASAP7_75t_R _24906_ (.A1(_16463_),
    .A2(_16325_),
    .B(_16495_),
    .Y(_16499_));
 AND5x1_ASAP7_75t_R _24907_ (.A(_16486_),
    .B(_16491_),
    .C(_16494_),
    .D(_16497_),
    .E(_16499_),
    .Y(_16500_));
 AND3x4_ASAP7_75t_R _24908_ (.A(_16290_),
    .B(_16291_),
    .C(_00430_),
    .Y(_16501_));
 BUFx2_ASAP7_75t_R output286 (.A(net286),
    .Y(text_out[123]));
 NAND2x1_ASAP7_75t_R _24910_ (.A(_16394_),
    .B(_16501_),
    .Y(_16503_));
 INVx5_ASAP7_75t_R _24911_ (.A(_16501_),
    .Y(_16504_));
 AO21x1_ASAP7_75t_R _24912_ (.A1(_16325_),
    .A2(_16443_),
    .B(_16504_),
    .Y(_16505_));
 AND2x2_ASAP7_75t_R _24913_ (.A(_16306_),
    .B(net2157),
    .Y(_16506_));
 AND2x2_ASAP7_75t_R _24914_ (.A(_16501_),
    .B(_16506_),
    .Y(_16507_));
 INVx1_ASAP7_75t_R _24915_ (.A(_16507_),
    .Y(_16508_));
 NOR2x2_ASAP7_75t_R _24916_ (.A(_16483_),
    .B(_16271_),
    .Y(_16509_));
 NAND2x1_ASAP7_75t_R _24917_ (.A(_16318_),
    .B(_16509_),
    .Y(_16510_));
 NAND2x2_ASAP7_75t_R _24918_ (.A(_16265_),
    .B(net2158),
    .Y(_16511_));
 CKINVDCx6p67_ASAP7_75t_R _24919_ (.A(_16509_),
    .Y(_16512_));
 AO21x1_ASAP7_75t_R _24920_ (.A1(_16436_),
    .A2(_16511_),
    .B(_16512_),
    .Y(_16513_));
 AND5x1_ASAP7_75t_R _24921_ (.A(_16503_),
    .B(_16505_),
    .C(_16508_),
    .D(_16510_),
    .E(_16513_),
    .Y(_16514_));
 NAND3x1_ASAP7_75t_R _24922_ (.A(_16482_),
    .B(_16500_),
    .C(_16514_),
    .Y(_16515_));
 NOR2x1_ASAP7_75t_R _24923_ (.A(_16432_),
    .B(_16515_),
    .Y(_16516_));
 AO21x1_ASAP7_75t_R _24924_ (.A1(_16440_),
    .A2(_16443_),
    .B(_16354_),
    .Y(_16517_));
 OA21x2_ASAP7_75t_R _24925_ (.A1(_16354_),
    .A2(net2766),
    .B(_16517_),
    .Y(_16518_));
 NAND2x1_ASAP7_75t_R _24926_ (.A(_16353_),
    .B(_16278_),
    .Y(_16519_));
 NOR2x1_ASAP7_75t_R _24927_ (.A(_16266_),
    .B(_16354_),
    .Y(_16520_));
 INVx1_ASAP7_75t_R _24928_ (.A(_16520_),
    .Y(_16521_));
 AND5x1_ASAP7_75t_R _24929_ (.A(_16372_),
    .B(_16518_),
    .C(_16519_),
    .D(_16521_),
    .E(_16374_),
    .Y(_16522_));
 AND5x2_ASAP7_75t_R _24930_ (.A(_16269_),
    .B(_16522_),
    .C(_16411_),
    .D(_16378_),
    .E(_16391_),
    .Y(_16523_));
 NAND2x2_ASAP7_75t_R _24931_ (.A(_00429_),
    .B(_16523_),
    .Y(_16524_));
 NAND2x2_ASAP7_75t_R _24932_ (.A(_16516_),
    .B(_16524_),
    .Y(_16525_));
 XNOR2x1_ASAP7_75t_R _24933_ (.B(_16525_),
    .Y(_16526_),
    .A(_16261_));
 NAND2x2_ASAP7_75t_R _24934_ (.A(net403),
    .B(net4142),
    .Y(_16527_));
 OAI21x1_ASAP7_75t_R _24935_ (.A1(net405),
    .A2(_16526_),
    .B(_16527_),
    .Y(_00369_));
 BUFx2_ASAP7_75t_R output285 (.A(net285),
    .Y(text_out[122]));
 NAND2x1_ASAP7_75t_R _24937_ (.A(net3498),
    .B(_16501_),
    .Y(_16529_));
 NOR2x1_ASAP7_75t_R _24938_ (.A(_16463_),
    .B(_16504_),
    .Y(_16530_));
 NOR2x1_ASAP7_75t_R _24939_ (.A(_16387_),
    .B(_16504_),
    .Y(_16531_));
 AOI211x1_ASAP7_75t_R _24940_ (.A1(_16324_),
    .A2(_16501_),
    .B(_16530_),
    .C(_16531_),
    .Y(_16532_));
 NAND2x1_ASAP7_75t_R _24941_ (.A(_16373_),
    .B(_16501_),
    .Y(_16533_));
 NOR2x1_ASAP7_75t_R _24942_ (.A(_16312_),
    .B(_16504_),
    .Y(_16534_));
 INVx1_ASAP7_75t_R _24943_ (.A(_16534_),
    .Y(_16535_));
 NAND2x1_ASAP7_75t_R _24944_ (.A(_16334_),
    .B(_16501_),
    .Y(_16536_));
 AND5x1_ASAP7_75t_R _24945_ (.A(_16529_),
    .B(_16532_),
    .C(_16533_),
    .D(_16535_),
    .E(_16536_),
    .Y(_16537_));
 NOR2x2_ASAP7_75t_R _24946_ (.A(_16262_),
    .B(net2664),
    .Y(_16538_));
 INVx3_ASAP7_75t_R _24947_ (.A(_16538_),
    .Y(_16539_));
 AO21x1_ASAP7_75t_R _24948_ (.A1(_16539_),
    .A2(_16266_),
    .B(_16488_),
    .Y(_16540_));
 NOR2x2_ASAP7_75t_R _24949_ (.A(_16277_),
    .B(_16263_),
    .Y(_16541_));
 CKINVDCx10_ASAP7_75t_R _24950_ (.A(_16541_),
    .Y(_16542_));
 BUFx2_ASAP7_75t_R output284 (.A(net284),
    .Y(text_out[121]));
 NAND2x1_ASAP7_75t_R _24952_ (.A(_16484_),
    .B(_16348_),
    .Y(_16544_));
 NAND2x1_ASAP7_75t_R _24953_ (.A(_16484_),
    .B(_16373_),
    .Y(_16545_));
 OA211x2_ASAP7_75t_R _24954_ (.A1(net3499),
    .A2(_16495_),
    .B(_16544_),
    .C(_16545_),
    .Y(_16546_));
 NAND2x1_ASAP7_75t_R _24955_ (.A(_16416_),
    .B(_16487_),
    .Y(_16547_));
 AND3x1_ASAP7_75t_R _24956_ (.A(_16487_),
    .B(net1854),
    .C(_16306_),
    .Y(_16548_));
 INVx1_ASAP7_75t_R _24957_ (.A(_16548_),
    .Y(_16549_));
 OAI21x1_ASAP7_75t_R _24958_ (.A1(_16416_),
    .A2(_16506_),
    .B(_16484_),
    .Y(_16550_));
 AND5x1_ASAP7_75t_R _24959_ (.A(_16540_),
    .B(_16546_),
    .C(_16547_),
    .D(_16549_),
    .E(_16550_),
    .Y(_16551_));
 BUFx2_ASAP7_75t_R output283 (.A(net283),
    .Y(text_out[120]));
 AND3x1_ASAP7_75t_R _24961_ (.A(_16509_),
    .B(_16381_),
    .C(net2157),
    .Y(_16553_));
 INVx1_ASAP7_75t_R _24962_ (.A(_16553_),
    .Y(_16554_));
 AO21x1_ASAP7_75t_R _24963_ (.A1(_16440_),
    .A2(_16443_),
    .B(_16512_),
    .Y(_16555_));
 OA211x2_ASAP7_75t_R _24964_ (.A1(_16357_),
    .A2(_16512_),
    .B(_16554_),
    .C(_16555_),
    .Y(_16556_));
 AND3x2_ASAP7_75t_R _24965_ (.A(_16537_),
    .B(_16551_),
    .C(_16556_),
    .Y(_16557_));
 AND2x2_ASAP7_75t_R _24966_ (.A(_16311_),
    .B(_16452_),
    .Y(_16558_));
 INVx1_ASAP7_75t_R _24967_ (.A(_16558_),
    .Y(_16559_));
 NOR2x2_ASAP7_75t_R _24968_ (.A(_16304_),
    .B(_16300_),
    .Y(_16560_));
 CKINVDCx8_ASAP7_75t_R _24969_ (.A(_16560_),
    .Y(_16561_));
 BUFx2_ASAP7_75t_R output282 (.A(net282),
    .Y(text_out[11]));
 INVx5_ASAP7_75t_R _24971_ (.A(_16452_),
    .Y(_16563_));
 BUFx2_ASAP7_75t_R output281 (.A(net281),
    .Y(text_out[119]));
 AO21x1_ASAP7_75t_R _24973_ (.A1(_16561_),
    .A2(_16357_),
    .B(_16563_),
    .Y(_16565_));
 AO21x1_ASAP7_75t_R _24974_ (.A1(_16325_),
    .A2(_16469_),
    .B(_16563_),
    .Y(_16566_));
 AND2x2_ASAP7_75t_R _24975_ (.A(_16394_),
    .B(_16452_),
    .Y(_16567_));
 INVx1_ASAP7_75t_R _24976_ (.A(_16567_),
    .Y(_16568_));
 AND2x2_ASAP7_75t_R _24977_ (.A(_16452_),
    .B(_16397_),
    .Y(_16569_));
 INVx1_ASAP7_75t_R _24978_ (.A(_16569_),
    .Y(_16570_));
 AND5x1_ASAP7_75t_R _24979_ (.A(_16559_),
    .B(_16565_),
    .C(_16566_),
    .D(_16568_),
    .E(_16570_),
    .Y(_16571_));
 BUFx2_ASAP7_75t_R output280 (.A(net280),
    .Y(text_out[118]));
 AND2x2_ASAP7_75t_R _24981_ (.A(_16459_),
    .B(_16541_),
    .Y(_16573_));
 INVx1_ASAP7_75t_R _24982_ (.A(_16573_),
    .Y(_16574_));
 AO21x1_ASAP7_75t_R _24983_ (.A1(_16421_),
    .A2(_16395_),
    .B(_16460_),
    .Y(_16575_));
 OR3x1_ASAP7_75t_R _24984_ (.A(_16460_),
    .B(_16404_),
    .C(net2769),
    .Y(_16576_));
 NOR2x1_ASAP7_75t_R _24985_ (.A(_16440_),
    .B(_16460_),
    .Y(_16577_));
 INVx1_ASAP7_75t_R _24986_ (.A(_16577_),
    .Y(_16578_));
 OA211x2_ASAP7_75t_R _24987_ (.A1(_16460_),
    .A2(_16469_),
    .B(_16576_),
    .C(_16578_),
    .Y(_16579_));
 AND4x2_ASAP7_75t_R _24988_ (.A(_16571_),
    .B(_16574_),
    .C(_16575_),
    .D(_16579_),
    .Y(_16580_));
 AO21x1_ASAP7_75t_R _24989_ (.A1(_16436_),
    .A2(_16279_),
    .B(_16471_),
    .Y(_16581_));
 AO21x1_ASAP7_75t_R _24990_ (.A1(_16421_),
    .A2(_16366_),
    .B(_16437_),
    .Y(_16582_));
 AO21x1_ASAP7_75t_R _24991_ (.A1(_16357_),
    .A2(_16445_),
    .B(_16437_),
    .Y(_16583_));
 NAND2x1_ASAP7_75t_R _24992_ (.A(_16311_),
    .B(_16434_),
    .Y(_16584_));
 NAND2x1_ASAP7_75t_R _24993_ (.A(net1744),
    .B(_16434_),
    .Y(_16585_));
 AND4x1_ASAP7_75t_R _24994_ (.A(_16582_),
    .B(_16583_),
    .C(_16584_),
    .D(_16585_),
    .Y(_16586_));
 NAND2x1_ASAP7_75t_R _24995_ (.A(_16541_),
    .B(_16467_),
    .Y(_16587_));
 AND3x1_ASAP7_75t_R _24996_ (.A(_16467_),
    .B(_16301_),
    .C(_16265_),
    .Y(_16588_));
 INVx1_ASAP7_75t_R _24997_ (.A(_16588_),
    .Y(_16589_));
 NAND2x1_ASAP7_75t_R _24998_ (.A(net1745),
    .B(_16467_),
    .Y(_16590_));
 AND5x2_ASAP7_75t_R _24999_ (.A(_16581_),
    .B(_16586_),
    .C(_16587_),
    .D(_16589_),
    .E(_16590_),
    .Y(_16591_));
 NAND3x2_ASAP7_75t_R _25000_ (.B(_16580_),
    .C(_16591_),
    .Y(_16592_),
    .A(_16557_));
 NOR2x1_ASAP7_75t_R _25001_ (.A(_16327_),
    .B(_16366_),
    .Y(_16593_));
 BUFx2_ASAP7_75t_R output279 (.A(net279),
    .Y(text_out[117]));
 NOR2x1_ASAP7_75t_R _25003_ (.A(_16469_),
    .B(_16327_),
    .Y(_16595_));
 AO21x1_ASAP7_75t_R _25004_ (.A1(_16317_),
    .A2(_16322_),
    .B(_16595_),
    .Y(_16596_));
 AND3x1_ASAP7_75t_R _25005_ (.A(_16317_),
    .B(_16300_),
    .C(_16306_),
    .Y(_16597_));
 NAND2x1_ASAP7_75t_R _25006_ (.A(_16381_),
    .B(_16317_),
    .Y(_16598_));
 INVx1_ASAP7_75t_R _25007_ (.A(_16598_),
    .Y(_16599_));
 OR5x1_ASAP7_75t_R _25008_ (.A(_16593_),
    .B(_16596_),
    .C(_16336_),
    .D(_16597_),
    .E(_16599_),
    .Y(_16600_));
 INVx1_ASAP7_75t_R _25009_ (.A(_16600_),
    .Y(_16601_));
 AO21x1_ASAP7_75t_R _25010_ (.A1(_16421_),
    .A2(_16395_),
    .B(_16342_),
    .Y(_16602_));
 AO21x1_ASAP7_75t_R _25011_ (.A1(_16561_),
    .A2(_16325_),
    .B(_16342_),
    .Y(_16603_));
 AO21x1_ASAP7_75t_R _25012_ (.A1(net3499),
    .A2(_16539_),
    .B(_16342_),
    .Y(_16604_));
 AND3x1_ASAP7_75t_R _25013_ (.A(_16602_),
    .B(_16603_),
    .C(_16604_),
    .Y(_16605_));
 AND3x1_ASAP7_75t_R _25014_ (.A(_16272_),
    .B(_16275_),
    .C(_16296_),
    .Y(_16606_));
 INVx1_ASAP7_75t_R _25015_ (.A(_16606_),
    .Y(_16607_));
 BUFx2_ASAP7_75t_R output278 (.A(net278),
    .Y(text_out[116]));
 AO21x1_ASAP7_75t_R _25017_ (.A1(_16387_),
    .A2(_16445_),
    .B(_16283_),
    .Y(_16609_));
 AO21x1_ASAP7_75t_R _25018_ (.A1(_16366_),
    .A2(_16370_),
    .B(_16283_),
    .Y(_16610_));
 AND3x1_ASAP7_75t_R _25019_ (.A(_16607_),
    .B(_16609_),
    .C(_16610_),
    .Y(_16611_));
 NOR2x2_ASAP7_75t_R _25020_ (.A(_16404_),
    .B(_16302_),
    .Y(_16612_));
 NOR2x1_ASAP7_75t_R _25021_ (.A(_16293_),
    .B(_16542_),
    .Y(_16613_));
 NOR2x1_ASAP7_75t_R _25022_ (.A(_16293_),
    .B(_16436_),
    .Y(_16614_));
 OR3x1_ASAP7_75t_R _25023_ (.A(_16612_),
    .B(_16613_),
    .C(_16614_),
    .Y(_16615_));
 AO21x1_ASAP7_75t_R _25024_ (.A1(_16440_),
    .A2(_16469_),
    .B(_16293_),
    .Y(_16616_));
 INVx1_ASAP7_75t_R _25025_ (.A(_16616_),
    .Y(_16617_));
 AOI211x1_ASAP7_75t_R _25026_ (.A1(net2622),
    .A2(_16294_),
    .B(_16615_),
    .C(_16617_),
    .Y(_16618_));
 AND4x1_ASAP7_75t_R _25027_ (.A(_16601_),
    .B(_16605_),
    .C(_16611_),
    .D(_16618_),
    .Y(_16619_));
 INVx1_ASAP7_75t_R _25028_ (.A(_16619_),
    .Y(_16620_));
 NAND2x2_ASAP7_75t_R _25029_ (.A(net3479),
    .B(_16296_),
    .Y(_16621_));
 AO21x1_ASAP7_75t_R _25030_ (.A1(_16366_),
    .A2(_16370_),
    .B(_16378_),
    .Y(_16622_));
 AO21x1_ASAP7_75t_R _25031_ (.A1(_16387_),
    .A2(_16445_),
    .B(_16378_),
    .Y(_16623_));
 OA211x2_ASAP7_75t_R _25032_ (.A1(_16378_),
    .A2(_16621_),
    .B(_16622_),
    .C(_16623_),
    .Y(_16624_));
 OR3x1_ASAP7_75t_R _25033_ (.A(_16354_),
    .B(_16299_),
    .C(net2768),
    .Y(_16625_));
 AND5x1_ASAP7_75t_R _25034_ (.A(_16372_),
    .B(_16624_),
    .C(_16521_),
    .D(_16363_),
    .E(_16625_),
    .Y(_16626_));
 AO21x1_ASAP7_75t_R _25035_ (.A1(_16312_),
    .A2(_16539_),
    .B(_16411_),
    .Y(_16627_));
 OA211x2_ASAP7_75t_R _25036_ (.A1(_16411_),
    .A2(_16366_),
    .B(_16627_),
    .C(_16428_),
    .Y(_16628_));
 NOR2x1_ASAP7_75t_R _25037_ (.A(_16357_),
    .B(_16411_),
    .Y(_16629_));
 AO21x1_ASAP7_75t_R _25038_ (.A1(_16409_),
    .A2(net2492),
    .B(_16629_),
    .Y(_16630_));
 INVx1_ASAP7_75t_R _25039_ (.A(_16630_),
    .Y(_16631_));
 OR3x2_ASAP7_75t_R _25040_ (.A(_16391_),
    .B(_16299_),
    .C(net2768),
    .Y(_16632_));
 AO21x1_ASAP7_75t_R _25041_ (.A1(_16325_),
    .A2(_16443_),
    .B(_16391_),
    .Y(_16633_));
 AND5x1_ASAP7_75t_R _25042_ (.A(_16418_),
    .B(_16628_),
    .C(_16631_),
    .D(_16632_),
    .E(_16633_),
    .Y(_16634_));
 NAND2x1_ASAP7_75t_R _25043_ (.A(_16626_),
    .B(_16634_),
    .Y(_16635_));
 NOR2x1_ASAP7_75t_R _25044_ (.A(_16620_),
    .B(_16635_),
    .Y(_16636_));
 INVx1_ASAP7_75t_R _25045_ (.A(_16636_),
    .Y(_16637_));
 NOR2x2_ASAP7_75t_R _25046_ (.A(_16592_),
    .B(_16637_),
    .Y(_16638_));
 BUFx2_ASAP7_75t_R output277 (.A(net277),
    .Y(text_out[115]));
 XOR2x2_ASAP7_75t_R _25048_ (.A(_00459_),
    .B(_00507_),
    .Y(_16640_));
 XOR2x1_ASAP7_75t_R _25049_ (.A(_00400_),
    .Y(_16641_),
    .B(net1146));
 XOR2x1_ASAP7_75t_R _25050_ (.A(_16640_),
    .Y(_16642_),
    .B(_16641_));
 XNOR2x1_ASAP7_75t_R _25051_ (.B(_16642_),
    .Y(_16643_),
    .A(_00399_));
 INVx1_ASAP7_75t_R _25052_ (.A(_16643_),
    .Y(_16644_));
 NAND3x1_ASAP7_75t_R _25053_ (.A(_16638_),
    .B(_16524_),
    .C(_16644_),
    .Y(_16645_));
 AO21x1_ASAP7_75t_R _25054_ (.A1(_16638_),
    .A2(_16524_),
    .B(_16644_),
    .Y(_16646_));
 NAND2x1_ASAP7_75t_R _25055_ (.A(_16645_),
    .B(_16646_),
    .Y(_16647_));
 BUFx2_ASAP7_75t_R output276 (.A(net276),
    .Y(text_out[114]));
 NOR2x1_ASAP7_75t_R _25057_ (.A(net4160),
    .B(net399),
    .Y(_16649_));
 AOI21x1_ASAP7_75t_R _25058_ (.A1(net399),
    .A2(_16647_),
    .B(_16649_),
    .Y(_00370_));
 BUFx2_ASAP7_75t_R output275 (.A(net275),
    .Y(text_out[113]));
 BUFx2_ASAP7_75t_R output274 (.A(net274),
    .Y(text_out[112]));
 AO21x1_ASAP7_75t_R _25061_ (.A1(_16348_),
    .A2(_16317_),
    .B(_16593_),
    .Y(_16652_));
 NOR2x1_ASAP7_75t_R _25062_ (.A(_16327_),
    .B(_16357_),
    .Y(_16653_));
 NOR2x1_ASAP7_75t_R _25063_ (.A(_16327_),
    .B(_16542_),
    .Y(_16654_));
 AND2x2_ASAP7_75t_R _25064_ (.A(_16317_),
    .B(_16416_),
    .Y(_16655_));
 OR4x1_ASAP7_75t_R _25065_ (.A(_16652_),
    .B(_16653_),
    .C(_16654_),
    .D(_16655_),
    .Y(_16656_));
 INVx1_ASAP7_75t_R _25066_ (.A(_16349_),
    .Y(_16657_));
 AO21x1_ASAP7_75t_R _25067_ (.A1(_16341_),
    .A2(_16334_),
    .B(_16657_),
    .Y(_16658_));
 NAND2x1_ASAP7_75t_R _25068_ (.A(_16541_),
    .B(_16341_),
    .Y(_16659_));
 INVx1_ASAP7_75t_R _25069_ (.A(_16659_),
    .Y(_16660_));
 NOR2x1_ASAP7_75t_R _25070_ (.A(_16469_),
    .B(_16342_),
    .Y(_16661_));
 AND2x2_ASAP7_75t_R _25071_ (.A(_16341_),
    .B(_16356_),
    .Y(_16662_));
 OR4x1_ASAP7_75t_R _25072_ (.A(_16658_),
    .B(_16660_),
    .C(_16661_),
    .D(_16662_),
    .Y(_16663_));
 NOR2x1_ASAP7_75t_R _25073_ (.A(_16656_),
    .B(_16663_),
    .Y(_16664_));
 NOR2x1_ASAP7_75t_R _25074_ (.A(_16440_),
    .B(_16283_),
    .Y(_16665_));
 INVx1_ASAP7_75t_R _25075_ (.A(_16665_),
    .Y(_16666_));
 OA21x2_ASAP7_75t_R _25076_ (.A1(_16311_),
    .A2(_16278_),
    .B(_16272_),
    .Y(_16667_));
 INVx1_ASAP7_75t_R _25077_ (.A(_16667_),
    .Y(_16668_));
 AO21x1_ASAP7_75t_R _25078_ (.A1(_16561_),
    .A2(_16357_),
    .B(_16283_),
    .Y(_16669_));
 AND2x2_ASAP7_75t_R _25079_ (.A(_16334_),
    .B(_16272_),
    .Y(_16670_));
 INVx1_ASAP7_75t_R _25080_ (.A(_16670_),
    .Y(_16671_));
 AND5x1_ASAP7_75t_R _25081_ (.A(_16666_),
    .B(_16668_),
    .C(_16669_),
    .D(_16671_),
    .E(_16274_),
    .Y(_16672_));
 NOR2x1_ASAP7_75t_R _25082_ (.A(net3503),
    .B(_16469_),
    .Y(_16673_));
 NOR2x1_ASAP7_75t_R _25083_ (.A(_16293_),
    .B(_16539_),
    .Y(_16674_));
 NOR2x1_ASAP7_75t_R _25084_ (.A(net3503),
    .B(_16335_),
    .Y(_16675_));
 OR4x1_ASAP7_75t_R _25085_ (.A(_16309_),
    .B(_16673_),
    .C(_16674_),
    .D(_16675_),
    .Y(_16676_));
 INVx1_ASAP7_75t_R _25086_ (.A(_16676_),
    .Y(_16677_));
 AND3x1_ASAP7_75t_R _25087_ (.A(_16664_),
    .B(_16672_),
    .C(_16677_),
    .Y(_16678_));
 AO21x1_ASAP7_75t_R _25088_ (.A1(_16542_),
    .A2(_16511_),
    .B(_16354_),
    .Y(_16679_));
 AO21x1_ASAP7_75t_R _25089_ (.A1(_16440_),
    .A2(_16463_),
    .B(_16354_),
    .Y(_16680_));
 AND3x1_ASAP7_75t_R _25090_ (.A(_16361_),
    .B(_16679_),
    .C(_16680_),
    .Y(_16681_));
 INVx1_ASAP7_75t_R _25091_ (.A(_16681_),
    .Y(_16682_));
 NOR2x1_ASAP7_75t_R _25092_ (.A(_16378_),
    .B(_16426_),
    .Y(_16683_));
 NOR2x1_ASAP7_75t_R _25093_ (.A(_16469_),
    .B(_16378_),
    .Y(_16684_));
 AO21x1_ASAP7_75t_R _25094_ (.A1(_16386_),
    .A2(_16376_),
    .B(_16684_),
    .Y(_16685_));
 OA211x2_ASAP7_75t_R _25095_ (.A1(net1854),
    .A2(_16287_),
    .B(_16376_),
    .C(_16381_),
    .Y(_16686_));
 OR4x2_ASAP7_75t_R _25096_ (.A(_16682_),
    .B(_16683_),
    .C(_16685_),
    .D(_16686_),
    .Y(_16687_));
 NAND2x1_ASAP7_75t_R _25097_ (.A(_16538_),
    .B(_16390_),
    .Y(_16688_));
 INVx1_ASAP7_75t_R _25098_ (.A(_16688_),
    .Y(_16689_));
 AO21x1_ASAP7_75t_R _25099_ (.A1(_16541_),
    .A2(_16390_),
    .B(_16689_),
    .Y(_16690_));
 NOR2x1_ASAP7_75t_R _25100_ (.A(_16391_),
    .B(_16421_),
    .Y(_16691_));
 NAND2x1_ASAP7_75t_R _25101_ (.A(_16306_),
    .B(_16390_),
    .Y(_16692_));
 INVx1_ASAP7_75t_R _25102_ (.A(_16692_),
    .Y(_16693_));
 AND3x1_ASAP7_75t_R _25103_ (.A(_16390_),
    .B(net2159),
    .C(_16296_),
    .Y(_16694_));
 OR4x2_ASAP7_75t_R _25104_ (.A(_16690_),
    .B(_16691_),
    .C(_16693_),
    .D(_16694_),
    .Y(_16695_));
 OA21x2_ASAP7_75t_R _25105_ (.A1(_16324_),
    .A2(_16322_),
    .B(_16409_),
    .Y(_16696_));
 OA21x2_ASAP7_75t_R _25106_ (.A1(_16334_),
    .A2(_16348_),
    .B(_16409_),
    .Y(_16697_));
 NOR2x1_ASAP7_75t_R _25107_ (.A(_16279_),
    .B(_16411_),
    .Y(_16698_));
 OR5x2_ASAP7_75t_R _25108_ (.A(_16413_),
    .B(_16696_),
    .C(_16697_),
    .D(_16698_),
    .E(_16629_),
    .Y(_16699_));
 NOR3x2_ASAP7_75t_R _25109_ (.B(_16695_),
    .C(_16699_),
    .Y(_16700_),
    .A(_16687_));
 NAND2x2_ASAP7_75t_R _25110_ (.A(_16678_),
    .B(_16700_),
    .Y(_16701_));
 INVx1_ASAP7_75t_R _25111_ (.A(_16701_),
    .Y(_16702_));
 NOR2x1_ASAP7_75t_R _25112_ (.A(_16279_),
    .B(_16504_),
    .Y(_16703_));
 INVx1_ASAP7_75t_R _25113_ (.A(_16703_),
    .Y(_16704_));
 NAND2x1_ASAP7_75t_R _25114_ (.A(_16541_),
    .B(_16501_),
    .Y(_16705_));
 AND5x1_ASAP7_75t_R _25115_ (.A(_16704_),
    .B(_16529_),
    .C(_16533_),
    .D(_16705_),
    .E(_16503_),
    .Y(_16706_));
 OR3x1_ASAP7_75t_R _25116_ (.A(_16512_),
    .B(_16404_),
    .C(net2769),
    .Y(_16707_));
 AO21x1_ASAP7_75t_R _25117_ (.A1(_16335_),
    .A2(_16366_),
    .B(_16512_),
    .Y(_16708_));
 OA211x2_ASAP7_75t_R _25118_ (.A1(net3499),
    .A2(_16512_),
    .B(_16707_),
    .C(_16708_),
    .Y(_16709_));
 INVx1_ASAP7_75t_R _25119_ (.A(_16531_),
    .Y(_16710_));
 NOR2x1_ASAP7_75t_R _25120_ (.A(_16445_),
    .B(_16504_),
    .Y(_16711_));
 INVx1_ASAP7_75t_R _25121_ (.A(_16711_),
    .Y(_16712_));
 NAND2x1_ASAP7_75t_R _25122_ (.A(_16356_),
    .B(_16501_),
    .Y(_16713_));
 AND4x1_ASAP7_75t_R _25123_ (.A(_16505_),
    .B(_16710_),
    .C(_16712_),
    .D(_16713_),
    .Y(_16714_));
 AND3x2_ASAP7_75t_R _25124_ (.A(_16706_),
    .B(_16709_),
    .C(_16714_),
    .Y(_16715_));
 AO21x1_ASAP7_75t_R _25125_ (.A1(_16312_),
    .A2(_16542_),
    .B(_16437_),
    .Y(_16716_));
 AO21x1_ASAP7_75t_R _25126_ (.A1(_16421_),
    .A2(_16335_),
    .B(_16437_),
    .Y(_16717_));
 AO21x1_ASAP7_75t_R _25127_ (.A1(_16325_),
    .A2(_16469_),
    .B(_16437_),
    .Y(_16718_));
 AND4x1_ASAP7_75t_R _25128_ (.A(_16716_),
    .B(_16717_),
    .C(_16583_),
    .D(_16718_),
    .Y(_16719_));
 AO21x1_ASAP7_75t_R _25129_ (.A1(_16436_),
    .A2(_16542_),
    .B(_16471_),
    .Y(_16720_));
 NOR2x1_ASAP7_75t_R _25130_ (.A(_16511_),
    .B(_16471_),
    .Y(_16721_));
 INVx1_ASAP7_75t_R _25131_ (.A(_16721_),
    .Y(_16722_));
 NAND2x1_ASAP7_75t_R _25132_ (.A(_16344_),
    .B(_16467_),
    .Y(_16723_));
 AND3x1_ASAP7_75t_R _25133_ (.A(_16720_),
    .B(_16722_),
    .C(_16723_),
    .Y(_16724_));
 AND2x2_ASAP7_75t_R _25134_ (.A(_16719_),
    .B(_16724_),
    .Y(_16725_));
 OR3x1_ASAP7_75t_R _25135_ (.A(_16262_),
    .B(net3487),
    .C(net2210),
    .Y(_16726_));
 AO21x1_ASAP7_75t_R _25136_ (.A1(_16726_),
    .A2(_16370_),
    .B(_16563_),
    .Y(_16727_));
 AO21x1_ASAP7_75t_R _25137_ (.A1(_16463_),
    .A2(_16469_),
    .B(_16563_),
    .Y(_16728_));
 OA211x2_ASAP7_75t_R _25138_ (.A1(net2769),
    .A2(_16563_),
    .B(_16727_),
    .C(_16728_),
    .Y(_16729_));
 AO21x1_ASAP7_75t_R _25139_ (.A1(_16463_),
    .A2(_16469_),
    .B(_16460_),
    .Y(_16730_));
 NAND2x2_ASAP7_75t_R _25140_ (.A(net1744),
    .B(_16459_),
    .Y(_16731_));
 AND2x2_ASAP7_75t_R _25141_ (.A(_16459_),
    .B(_16560_),
    .Y(_16732_));
 INVx1_ASAP7_75t_R _25142_ (.A(_16732_),
    .Y(_16733_));
 AND4x1_ASAP7_75t_R _25143_ (.A(_16730_),
    .B(_16731_),
    .C(_16733_),
    .D(_16578_),
    .Y(_16734_));
 AO21x1_ASAP7_75t_R _25144_ (.A1(_16395_),
    .A2(_16398_),
    .B(_16460_),
    .Y(_16735_));
 NAND2x1_ASAP7_75t_R _25145_ (.A(_16373_),
    .B(_16459_),
    .Y(_16736_));
 AND3x1_ASAP7_75t_R _25146_ (.A(_16735_),
    .B(_16736_),
    .C(_16574_),
    .Y(_16737_));
 AND2x2_ASAP7_75t_R _25147_ (.A(_16734_),
    .B(_16737_),
    .Y(_16738_));
 AND3x2_ASAP7_75t_R _25148_ (.A(_16725_),
    .B(_16729_),
    .C(_16738_),
    .Y(_16739_));
 OR3x1_ASAP7_75t_R _25149_ (.A(_16495_),
    .B(_16416_),
    .C(_16397_),
    .Y(_16740_));
 NAND2x1_ASAP7_75t_R _25150_ (.A(_16362_),
    .B(_16487_),
    .Y(_16741_));
 NAND2x1_ASAP7_75t_R _25151_ (.A(_16487_),
    .B(_16425_),
    .Y(_16742_));
 AO21x1_ASAP7_75t_R _25152_ (.A1(_16312_),
    .A2(_16539_),
    .B(_16488_),
    .Y(_16743_));
 AND4x2_ASAP7_75t_R _25153_ (.A(_16740_),
    .B(_16741_),
    .C(_16742_),
    .D(_16743_),
    .Y(_16744_));
 NAND3x2_ASAP7_75t_R _25154_ (.B(_16739_),
    .C(_16744_),
    .Y(_16745_),
    .A(_16715_));
 INVx1_ASAP7_75t_R _25155_ (.A(_16745_),
    .Y(_16746_));
 NAND2x2_ASAP7_75t_R _25156_ (.A(_16702_),
    .B(_16746_),
    .Y(_16747_));
 XNOR2x1_ASAP7_75t_R _25157_ (.B(_00506_),
    .Y(_16748_),
    .A(_00488_));
 XNOR2x1_ASAP7_75t_R _25158_ (.B(_00458_),
    .Y(_16749_),
    .A(net3397));
 XOR2x1_ASAP7_75t_R _25159_ (.A(_16748_),
    .Y(_16750_),
    .B(_16749_));
 XOR2x1_ASAP7_75t_R _25160_ (.A(_16750_),
    .Y(_16751_),
    .B(_00401_));
 XOR2x1_ASAP7_75t_R _25161_ (.A(_16747_),
    .Y(_16752_),
    .B(_16751_));
 NOR2x1_ASAP7_75t_R _25162_ (.A(net401),
    .B(_16752_),
    .Y(_16753_));
 AO21x1_ASAP7_75t_R _25163_ (.A1(net401),
    .A2(net3864),
    .B(_16753_),
    .Y(_00371_));
 XNOR2x2_ASAP7_75t_R _25164_ (.A(_00487_),
    .B(_00505_),
    .Y(_16754_));
 XOR2x1_ASAP7_75t_R _25165_ (.A(net3399),
    .Y(_16755_),
    .B(_00457_));
 XOR2x1_ASAP7_75t_R _25166_ (.A(_16754_),
    .Y(_16756_),
    .B(_16755_));
 INVx3_ASAP7_75t_R _25167_ (.A(_00402_),
    .Y(_16757_));
 XOR2x1_ASAP7_75t_R _25168_ (.A(_16756_),
    .Y(_16758_),
    .B(_16757_));
 AO21x1_ASAP7_75t_R _25169_ (.A1(_16440_),
    .A2(_16469_),
    .B(_16504_),
    .Y(_16759_));
 NAND2x1_ASAP7_75t_R _25170_ (.A(_16560_),
    .B(_16501_),
    .Y(_16760_));
 AND4x2_ASAP7_75t_R _25171_ (.A(_16759_),
    .B(_16710_),
    .C(_16760_),
    .D(_16712_),
    .Y(_16761_));
 AO21x1_ASAP7_75t_R _25172_ (.A1(_16335_),
    .A2(_16398_),
    .B(_16504_),
    .Y(_16762_));
 AND3x2_ASAP7_75t_R _25173_ (.A(_16762_),
    .B(_16704_),
    .C(_16535_),
    .Y(_16763_));
 AO21x1_ASAP7_75t_R _25174_ (.A1(_16421_),
    .A2(_16542_),
    .B(_16512_),
    .Y(_16764_));
 INVx1_ASAP7_75t_R _25175_ (.A(_16764_),
    .Y(_16765_));
 AO21x1_ASAP7_75t_R _25176_ (.A1(_16561_),
    .A2(_16445_),
    .B(_16512_),
    .Y(_16766_));
 INVx1_ASAP7_75t_R _25177_ (.A(_16766_),
    .Y(_16767_));
 NOR2x1_ASAP7_75t_R _25178_ (.A(_16443_),
    .B(_16512_),
    .Y(_16768_));
 OR3x1_ASAP7_75t_R _25179_ (.A(_16765_),
    .B(_16767_),
    .C(_16768_),
    .Y(_16769_));
 INVx1_ASAP7_75t_R _25180_ (.A(_16769_),
    .Y(_16770_));
 NAND3x2_ASAP7_75t_R _25181_ (.B(_16763_),
    .C(_16770_),
    .Y(_16771_),
    .A(_16761_));
 NOR2x1_ASAP7_75t_R _25182_ (.A(_16495_),
    .B(_16366_),
    .Y(_16772_));
 AO21x1_ASAP7_75t_R _25183_ (.A1(_16334_),
    .A2(_16484_),
    .B(_16772_),
    .Y(_16773_));
 AND2x2_ASAP7_75t_R _25184_ (.A(_16369_),
    .B(_16484_),
    .Y(_16774_));
 AND2x2_ASAP7_75t_R _25185_ (.A(_16318_),
    .B(_16484_),
    .Y(_16775_));
 AND3x1_ASAP7_75t_R _25186_ (.A(_16484_),
    .B(net2157),
    .C(_16296_),
    .Y(_16776_));
 OR4x2_ASAP7_75t_R _25187_ (.A(_16773_),
    .B(_16774_),
    .C(_16775_),
    .D(_16776_),
    .Y(_16777_));
 AND3x1_ASAP7_75t_R _25188_ (.A(_16377_),
    .B(_16381_),
    .C(_16487_),
    .Y(_16778_));
 AO21x1_ASAP7_75t_R _25189_ (.A1(_16487_),
    .A2(_16265_),
    .B(_16778_),
    .Y(_16779_));
 INVx1_ASAP7_75t_R _25190_ (.A(_16741_),
    .Y(_16780_));
 AND2x2_ASAP7_75t_R _25191_ (.A(_16487_),
    .B(_16356_),
    .Y(_16781_));
 AO21x1_ASAP7_75t_R _25192_ (.A1(_16487_),
    .A2(net2492),
    .B(_16781_),
    .Y(_16782_));
 OR3x2_ASAP7_75t_R _25193_ (.A(_16779_),
    .B(_16780_),
    .C(_16782_),
    .Y(_16783_));
 NOR3x2_ASAP7_75t_R _25194_ (.B(_16777_),
    .C(_16783_),
    .Y(_16784_),
    .A(_16771_));
 OA211x2_ASAP7_75t_R _25195_ (.A1(_16460_),
    .A2(_16445_),
    .B(_16733_),
    .C(_16578_),
    .Y(_16785_));
 NAND2x1_ASAP7_75t_R _25196_ (.A(_16538_),
    .B(_16452_),
    .Y(_16786_));
 OA211x2_ASAP7_75t_R _25197_ (.A1(_16266_),
    .A2(_16563_),
    .B(_16559_),
    .C(_16786_),
    .Y(_16787_));
 AO21x1_ASAP7_75t_R _25198_ (.A1(_16469_),
    .A2(_16621_),
    .B(_16563_),
    .Y(_16788_));
 OA21x2_ASAP7_75t_R _25199_ (.A1(_16445_),
    .A2(_16563_),
    .B(_16788_),
    .Y(_16789_));
 AO21x1_ASAP7_75t_R _25200_ (.A1(_16312_),
    .A2(_16398_),
    .B(_16460_),
    .Y(_16790_));
 AND4x1_ASAP7_75t_R _25201_ (.A(_16785_),
    .B(_16787_),
    .C(_16789_),
    .D(_16790_),
    .Y(_16791_));
 INVx1_ASAP7_75t_R _25202_ (.A(_16791_),
    .Y(_16792_));
 AO21x1_ASAP7_75t_R _25203_ (.A1(_16325_),
    .A2(_16443_),
    .B(_16437_),
    .Y(_16793_));
 NAND2x1_ASAP7_75t_R _25204_ (.A(_16560_),
    .B(_16434_),
    .Y(_16794_));
 AND5x1_ASAP7_75t_R _25205_ (.A(_16439_),
    .B(_16793_),
    .C(_16449_),
    .D(_16447_),
    .E(_16794_),
    .Y(_16795_));
 AO21x1_ASAP7_75t_R _25206_ (.A1(_16440_),
    .A2(_16463_),
    .B(_16471_),
    .Y(_16796_));
 AND3x1_ASAP7_75t_R _25207_ (.A(_16476_),
    .B(_16796_),
    .C(_16590_),
    .Y(_16797_));
 OA211x2_ASAP7_75t_R _25208_ (.A1(_16262_),
    .A2(net2209),
    .B(_16467_),
    .C(_16265_),
    .Y(_16798_));
 INVx1_ASAP7_75t_R _25209_ (.A(_16798_),
    .Y(_16799_));
 AND2x2_ASAP7_75t_R _25210_ (.A(_16311_),
    .B(_16467_),
    .Y(_16800_));
 INVx1_ASAP7_75t_R _25211_ (.A(_16800_),
    .Y(_16801_));
 AND3x1_ASAP7_75t_R _25212_ (.A(_16799_),
    .B(_16581_),
    .C(_16801_),
    .Y(_16802_));
 NAND3x1_ASAP7_75t_R _25213_ (.A(_16795_),
    .B(_16797_),
    .C(_16802_),
    .Y(_16803_));
 NOR2x1_ASAP7_75t_R _25214_ (.A(_16792_),
    .B(_16803_),
    .Y(_16804_));
 NAND2x2_ASAP7_75t_R _25215_ (.A(_16784_),
    .B(_16804_),
    .Y(_16805_));
 NAND2x1_ASAP7_75t_R _25216_ (.A(_16322_),
    .B(_16390_),
    .Y(_16806_));
 AO21x1_ASAP7_75t_R _25217_ (.A1(_16561_),
    .A2(_16445_),
    .B(_16411_),
    .Y(_16807_));
 NAND2x1_ASAP7_75t_R _25218_ (.A(_16394_),
    .B(_16409_),
    .Y(_16808_));
 NOR2x1_ASAP7_75t_R _25219_ (.A(_16391_),
    .B(_16335_),
    .Y(_16809_));
 INVx1_ASAP7_75t_R _25220_ (.A(_16809_),
    .Y(_16810_));
 AO21x1_ASAP7_75t_R _25221_ (.A1(_16561_),
    .A2(_16357_),
    .B(_16391_),
    .Y(_16811_));
 AND5x1_ASAP7_75t_R _25222_ (.A(_16806_),
    .B(_16807_),
    .C(_16808_),
    .D(_16810_),
    .E(_16811_),
    .Y(_16812_));
 AO21x1_ASAP7_75t_R _25223_ (.A1(_16366_),
    .A2(_16395_),
    .B(_16354_),
    .Y(_16813_));
 AO21x1_ASAP7_75t_R _25224_ (.A1(_16387_),
    .A2(_16357_),
    .B(_16354_),
    .Y(_16814_));
 AO21x1_ASAP7_75t_R _25225_ (.A1(_16440_),
    .A2(_16469_),
    .B(_16354_),
    .Y(_16815_));
 NAND2x1_ASAP7_75t_R _25226_ (.A(_16353_),
    .B(_16311_),
    .Y(_16816_));
 AND4x1_ASAP7_75t_R _25227_ (.A(_16813_),
    .B(_16814_),
    .C(_16815_),
    .D(_16816_),
    .Y(_16817_));
 INVx1_ASAP7_75t_R _25228_ (.A(_16383_),
    .Y(_16818_));
 OA21x2_ASAP7_75t_R _25229_ (.A1(_16356_),
    .A2(net2622),
    .B(_16376_),
    .Y(_16819_));
 INVx1_ASAP7_75t_R _25230_ (.A(_16819_),
    .Y(_16820_));
 NOR2x1_ASAP7_75t_R _25231_ (.A(_16378_),
    .B(_16395_),
    .Y(_16821_));
 INVx1_ASAP7_75t_R _25232_ (.A(_16821_),
    .Y(_16822_));
 AO21x1_ASAP7_75t_R _25233_ (.A1(_16325_),
    .A2(_16443_),
    .B(_16378_),
    .Y(_16823_));
 AND4x1_ASAP7_75t_R _25234_ (.A(_16818_),
    .B(_16820_),
    .C(_16822_),
    .D(_16823_),
    .Y(_16824_));
 AND3x2_ASAP7_75t_R _25235_ (.A(_16812_),
    .B(_16817_),
    .C(_16824_),
    .Y(_16825_));
 AO21x1_ASAP7_75t_R _25236_ (.A1(_16387_),
    .A2(_16357_),
    .B(net3504),
    .Y(_16826_));
 AO21x1_ASAP7_75t_R _25237_ (.A1(net3499),
    .A2(_16279_),
    .B(net3503),
    .Y(_16827_));
 INVx1_ASAP7_75t_R _25238_ (.A(_16673_),
    .Y(_16828_));
 INVx1_ASAP7_75t_R _25239_ (.A(_16675_),
    .Y(_16829_));
 AND4x1_ASAP7_75t_R _25240_ (.A(_16826_),
    .B(_16827_),
    .C(_16828_),
    .D(_16829_),
    .Y(_16830_));
 NOR2x1_ASAP7_75t_R _25241_ (.A(_16282_),
    .B(_16283_),
    .Y(_16831_));
 INVx1_ASAP7_75t_R _25242_ (.A(_16831_),
    .Y(_16832_));
 OA211x2_ASAP7_75t_R _25243_ (.A1(_16283_),
    .A2(_16398_),
    .B(_16671_),
    .C(_16832_),
    .Y(_16833_));
 OA211x2_ASAP7_75t_R _25244_ (.A1(_16283_),
    .A2(_16357_),
    .B(_16833_),
    .C(_16607_),
    .Y(_16834_));
 NAND2x1_ASAP7_75t_R _25245_ (.A(_16830_),
    .B(_16834_),
    .Y(_16835_));
 NOR2x1_ASAP7_75t_R _25246_ (.A(_16370_),
    .B(_16342_),
    .Y(_16836_));
 OR4x1_ASAP7_75t_R _25247_ (.A(_16597_),
    .B(_16329_),
    .C(_16595_),
    .D(_16655_),
    .Y(_16837_));
 AO21x1_ASAP7_75t_R _25248_ (.A1(_16262_),
    .A2(_00434_),
    .B(_00433_),
    .Y(_16838_));
 NOR2x1_ASAP7_75t_R _25249_ (.A(_16838_),
    .B(_16342_),
    .Y(_16839_));
 AO21x1_ASAP7_75t_R _25250_ (.A1(_16373_),
    .A2(_16317_),
    .B(_16332_),
    .Y(_16840_));
 INVx1_ASAP7_75t_R _25251_ (.A(_16661_),
    .Y(_16841_));
 AO21x1_ASAP7_75t_R _25252_ (.A1(_16561_),
    .A2(_16357_),
    .B(_16342_),
    .Y(_16842_));
 NAND2x1_ASAP7_75t_R _25253_ (.A(_16841_),
    .B(_16842_),
    .Y(_16843_));
 OR5x2_ASAP7_75t_R _25254_ (.A(_16836_),
    .B(_16837_),
    .C(_16839_),
    .D(_16840_),
    .E(_16843_),
    .Y(_16844_));
 NOR2x2_ASAP7_75t_R _25255_ (.A(_16835_),
    .B(_16844_),
    .Y(_16845_));
 NAND2x2_ASAP7_75t_R _25256_ (.A(_16825_),
    .B(_16845_),
    .Y(_16846_));
 OR2x2_ASAP7_75t_R _25257_ (.A(_16805_),
    .B(_16846_),
    .Y(_16847_));
 XNOR2x1_ASAP7_75t_R _25258_ (.B(_16847_),
    .Y(_16848_),
    .A(_16758_));
 AND2x2_ASAP7_75t_R _25259_ (.A(net402),
    .B(net48),
    .Y(_16849_));
 AO21x1_ASAP7_75t_R _25260_ (.A1(_16848_),
    .A2(net398),
    .B(_16849_),
    .Y(_00372_));
 BUFx2_ASAP7_75t_R output273 (.A(net273),
    .Y(text_out[111]));
 XNOR2x2_ASAP7_75t_R _25262_ (.A(_00486_),
    .B(_00504_),
    .Y(_16851_));
 XNOR2x1_ASAP7_75t_R _25263_ (.B(_00456_),
    .Y(_16852_),
    .A(_00424_));
 XOR2x1_ASAP7_75t_R _25264_ (.A(_16851_),
    .Y(_16853_),
    .B(_16852_));
 BUFx2_ASAP7_75t_R output272 (.A(net272),
    .Y(text_out[110]));
 XOR2x1_ASAP7_75t_R _25266_ (.A(_16853_),
    .Y(_16855_),
    .B(_00403_));
 AND2x2_ASAP7_75t_R _25267_ (.A(_16311_),
    .B(_16459_),
    .Y(_16856_));
 INVx1_ASAP7_75t_R _25268_ (.A(_16856_),
    .Y(_16857_));
 NAND2x1_ASAP7_75t_R _25269_ (.A(_16459_),
    .B(_16397_),
    .Y(_16858_));
 AND4x1_ASAP7_75t_R _25270_ (.A(_16857_),
    .B(_16574_),
    .C(_16736_),
    .D(_16858_),
    .Y(_16859_));
 AO21x1_ASAP7_75t_R _25271_ (.A1(_16440_),
    .A2(_16325_),
    .B(_16460_),
    .Y(_16860_));
 AO21x1_ASAP7_75t_R _25272_ (.A1(_16387_),
    .A2(_16445_),
    .B(_16563_),
    .Y(_16861_));
 AO21x1_ASAP7_75t_R _25273_ (.A1(_16440_),
    .A2(_16325_),
    .B(_16563_),
    .Y(_16862_));
 AND3x1_ASAP7_75t_R _25274_ (.A(_16727_),
    .B(_16861_),
    .C(_16862_),
    .Y(_16863_));
 NAND2x1_ASAP7_75t_R _25275_ (.A(_16416_),
    .B(_16459_),
    .Y(_16864_));
 AND5x2_ASAP7_75t_R _25276_ (.A(_16731_),
    .B(_16859_),
    .C(_16860_),
    .D(_16863_),
    .E(_16864_),
    .Y(_16865_));
 OA211x2_ASAP7_75t_R _25277_ (.A1(_16262_),
    .A2(_16287_),
    .B(_16467_),
    .C(_16296_),
    .Y(_16866_));
 INVx1_ASAP7_75t_R _25278_ (.A(_16866_),
    .Y(_16867_));
 INVx1_ASAP7_75t_R _25279_ (.A(_16479_),
    .Y(_16868_));
 AO21x1_ASAP7_75t_R _25280_ (.A1(net2279),
    .A2(_00434_),
    .B(net3491),
    .Y(_16869_));
 AO21x1_ASAP7_75t_R _25281_ (.A1(_16869_),
    .A2(_16445_),
    .B(_16437_),
    .Y(_16870_));
 AO21x1_ASAP7_75t_R _25282_ (.A1(_16561_),
    .A2(_16357_),
    .B(_16471_),
    .Y(_16871_));
 AND5x2_ASAP7_75t_R _25283_ (.A(_16581_),
    .B(_16867_),
    .C(_16868_),
    .D(_16870_),
    .E(_16871_),
    .Y(_16872_));
 INVx1_ASAP7_75t_R _25284_ (.A(_16774_),
    .Y(_16873_));
 NOR2x1_ASAP7_75t_R _25285_ (.A(_16511_),
    .B(_16488_),
    .Y(_16874_));
 OA21x2_ASAP7_75t_R _25286_ (.A1(_16311_),
    .A2(_16541_),
    .B(_16487_),
    .Y(_16875_));
 NOR2x1_ASAP7_75t_R _25287_ (.A(_16874_),
    .B(_16875_),
    .Y(_16876_));
 AO21x1_ASAP7_75t_R _25288_ (.A1(_16387_),
    .A2(_16469_),
    .B(_16488_),
    .Y(_16877_));
 AND5x1_ASAP7_75t_R _25289_ (.A(_16873_),
    .B(_16876_),
    .C(_16877_),
    .D(_16486_),
    .E(_16550_),
    .Y(_16878_));
 AND3x1_ASAP7_75t_R _25290_ (.A(_16533_),
    .B(_16705_),
    .C(_16536_),
    .Y(_16879_));
 AO21x1_ASAP7_75t_R _25291_ (.A1(_16440_),
    .A2(_16463_),
    .B(_16512_),
    .Y(_16880_));
 OA21x2_ASAP7_75t_R _25292_ (.A1(_16561_),
    .A2(_16512_),
    .B(_16880_),
    .Y(_16881_));
 AO21x1_ASAP7_75t_R _25293_ (.A1(_16357_),
    .A2(_16463_),
    .B(_16504_),
    .Y(_16882_));
 AND4x1_ASAP7_75t_R _25294_ (.A(_16879_),
    .B(_16513_),
    .C(_16881_),
    .D(_16882_),
    .Y(_16883_));
 AND2x2_ASAP7_75t_R _25295_ (.A(_16878_),
    .B(_16883_),
    .Y(_16884_));
 NAND3x2_ASAP7_75t_R _25296_ (.B(_16872_),
    .C(_16884_),
    .Y(_16885_),
    .A(_16865_));
 INVx1_ASAP7_75t_R _25297_ (.A(_16885_),
    .Y(_16886_));
 AO21x1_ASAP7_75t_R _25298_ (.A1(_16317_),
    .A2(_16386_),
    .B(_16319_),
    .Y(_16887_));
 OR3x1_ASAP7_75t_R _25299_ (.A(_16887_),
    .B(_16599_),
    .C(_16595_),
    .Y(_16888_));
 AO21x1_ASAP7_75t_R _25300_ (.A1(_16341_),
    .A2(_16267_),
    .B(_16836_),
    .Y(_16889_));
 NOR2x1_ASAP7_75t_R _25301_ (.A(_16621_),
    .B(_16342_),
    .Y(_16890_));
 OR4x1_ASAP7_75t_R _25302_ (.A(_16889_),
    .B(_16890_),
    .C(_16345_),
    .D(_16662_),
    .Y(_16891_));
 NOR2x1_ASAP7_75t_R _25303_ (.A(_16888_),
    .B(_16891_),
    .Y(_16892_));
 AO21x1_ASAP7_75t_R _25304_ (.A1(_16335_),
    .A2(_16395_),
    .B(_16283_),
    .Y(_16893_));
 AND2x2_ASAP7_75t_R _25305_ (.A(_16272_),
    .B(_16386_),
    .Y(_16894_));
 INVx1_ASAP7_75t_R _25306_ (.A(_16894_),
    .Y(_16895_));
 AO21x1_ASAP7_75t_R _25307_ (.A1(_16325_),
    .A2(_16469_),
    .B(_16283_),
    .Y(_16896_));
 AND5x1_ASAP7_75t_R _25308_ (.A(_16893_),
    .B(_16895_),
    .C(_16896_),
    .D(_16274_),
    .E(_16832_),
    .Y(_16897_));
 AO21x1_ASAP7_75t_R _25309_ (.A1(net3499),
    .A2(_16539_),
    .B(_16293_),
    .Y(_16898_));
 AO21x1_ASAP7_75t_R _25310_ (.A1(_16325_),
    .A2(net2767),
    .B(_16293_),
    .Y(_16899_));
 AND3x1_ASAP7_75t_R _25311_ (.A(_16898_),
    .B(_16302_),
    .C(_16899_),
    .Y(_16900_));
 AND3x1_ASAP7_75t_R _25312_ (.A(_16892_),
    .B(_16897_),
    .C(_16900_),
    .Y(_16901_));
 AO21x1_ASAP7_75t_R _25313_ (.A1(_16279_),
    .A2(_16511_),
    .B(_16354_),
    .Y(_16902_));
 OA211x2_ASAP7_75t_R _25314_ (.A1(_16354_),
    .A2(_16445_),
    .B(_16517_),
    .C(_16902_),
    .Y(_16903_));
 INVx1_ASAP7_75t_R _25315_ (.A(_16684_),
    .Y(_16904_));
 AO21x1_ASAP7_75t_R _25316_ (.A1(net2492),
    .A2(_16376_),
    .B(_16819_),
    .Y(_16905_));
 INVx1_ASAP7_75t_R _25317_ (.A(_16905_),
    .Y(_16906_));
 NOR2x1_ASAP7_75t_R _25318_ (.A(_16378_),
    .B(_16436_),
    .Y(_16907_));
 INVx1_ASAP7_75t_R _25319_ (.A(_16907_),
    .Y(_16908_));
 OA211x2_ASAP7_75t_R _25320_ (.A1(_16366_),
    .A2(_16378_),
    .B(_16822_),
    .C(_16908_),
    .Y(_16909_));
 AND4x1_ASAP7_75t_R _25321_ (.A(_16903_),
    .B(_16904_),
    .C(_16906_),
    .D(_16909_),
    .Y(_16910_));
 NOR2x1_ASAP7_75t_R _25322_ (.A(_16391_),
    .B(_16398_),
    .Y(_16911_));
 INVx1_ASAP7_75t_R _25323_ (.A(_16911_),
    .Y(_16912_));
 AND3x1_ASAP7_75t_R _25324_ (.A(_16301_),
    .B(_16390_),
    .C(_16381_),
    .Y(_16913_));
 INVx1_ASAP7_75t_R _25325_ (.A(_16913_),
    .Y(_16914_));
 AO21x1_ASAP7_75t_R _25326_ (.A1(_16395_),
    .A2(_16335_),
    .B(_16391_),
    .Y(_16915_));
 AND5x1_ASAP7_75t_R _25327_ (.A(_16912_),
    .B(_16632_),
    .C(_16403_),
    .D(_16914_),
    .E(_16915_),
    .Y(_16916_));
 AO21x1_ASAP7_75t_R _25328_ (.A1(_16436_),
    .A2(_16398_),
    .B(_16411_),
    .Y(_16917_));
 AND2x2_ASAP7_75t_R _25329_ (.A(_16409_),
    .B(_16506_),
    .Y(_16918_));
 INVx1_ASAP7_75t_R _25330_ (.A(_16918_),
    .Y(_16919_));
 AND2x2_ASAP7_75t_R _25331_ (.A(_16917_),
    .B(_16919_),
    .Y(_16920_));
 AND3x1_ASAP7_75t_R _25332_ (.A(_16910_),
    .B(_16916_),
    .C(_16920_),
    .Y(_16921_));
 NAND2x1_ASAP7_75t_R _25333_ (.A(_16901_),
    .B(_16921_),
    .Y(_16922_));
 INVx1_ASAP7_75t_R _25334_ (.A(_16922_),
    .Y(_16923_));
 NAND2x2_ASAP7_75t_R _25335_ (.A(_16886_),
    .B(_16923_),
    .Y(_16924_));
 XNOR2x1_ASAP7_75t_R _25336_ (.B(_16924_),
    .Y(_16925_),
    .A(_16855_));
 AND2x2_ASAP7_75t_R _25337_ (.A(net402),
    .B(net49),
    .Y(_16926_));
 AO21x1_ASAP7_75t_R _25338_ (.A1(_16925_),
    .A2(net398),
    .B(_16926_),
    .Y(_00373_));
 NOR2x1_ASAP7_75t_R _25339_ (.A(_16469_),
    .B(_16495_),
    .Y(_16927_));
 OA21x2_ASAP7_75t_R _25340_ (.A1(_16348_),
    .A2(_16394_),
    .B(_16484_),
    .Y(_16928_));
 INVx1_ASAP7_75t_R _25341_ (.A(_16545_),
    .Y(_16929_));
 OR3x1_ASAP7_75t_R _25342_ (.A(_16928_),
    .B(_16929_),
    .C(_16774_),
    .Y(_16930_));
 NOR2x1_ASAP7_75t_R _25343_ (.A(_16325_),
    .B(_16488_),
    .Y(_16931_));
 OR5x1_ASAP7_75t_R _25344_ (.A(_16927_),
    .B(_16930_),
    .C(_16931_),
    .D(_16548_),
    .E(_16778_),
    .Y(_16932_));
 OR3x1_ASAP7_75t_R _25345_ (.A(_16512_),
    .B(net3488),
    .C(net1854),
    .Y(_16933_));
 AO21x1_ASAP7_75t_R _25346_ (.A1(_16463_),
    .A2(_16621_),
    .B(_16512_),
    .Y(_16934_));
 OA211x2_ASAP7_75t_R _25347_ (.A1(_16387_),
    .A2(_16512_),
    .B(_16933_),
    .C(_16934_),
    .Y(_16935_));
 OA211x2_ASAP7_75t_R _25348_ (.A1(net1854),
    .A2(net2210),
    .B(_16501_),
    .C(_16265_),
    .Y(_16936_));
 INVx1_ASAP7_75t_R _25349_ (.A(_16936_),
    .Y(_16937_));
 OA21x2_ASAP7_75t_R _25350_ (.A1(_16541_),
    .A2(_16311_),
    .B(_16501_),
    .Y(_16938_));
 INVx1_ASAP7_75t_R _25351_ (.A(_16938_),
    .Y(_16939_));
 AND5x1_ASAP7_75t_R _25352_ (.A(_16704_),
    .B(_16937_),
    .C(_16939_),
    .D(_16760_),
    .E(_16505_),
    .Y(_16940_));
 NAND2x1_ASAP7_75t_R _25353_ (.A(_16935_),
    .B(_16940_),
    .Y(_16941_));
 NOR2x1_ASAP7_75t_R _25354_ (.A(_16932_),
    .B(_16941_),
    .Y(_16942_));
 AO21x1_ASAP7_75t_R _25355_ (.A1(_16395_),
    .A2(_16398_),
    .B(_16354_),
    .Y(_16943_));
 AND5x1_ASAP7_75t_R _25356_ (.A(_16372_),
    .B(_16625_),
    .C(_16943_),
    .D(_16517_),
    .E(_16519_),
    .Y(_16944_));
 AO21x1_ASAP7_75t_R _25357_ (.A1(_16335_),
    .A2(_16366_),
    .B(_16378_),
    .Y(_16945_));
 AO21x1_ASAP7_75t_R _25358_ (.A1(_16561_),
    .A2(_16445_),
    .B(_16378_),
    .Y(_16946_));
 AO21x1_ASAP7_75t_R _25359_ (.A1(_16279_),
    .A2(_16370_),
    .B(_16378_),
    .Y(_16947_));
 AND4x1_ASAP7_75t_R _25360_ (.A(_16945_),
    .B(_16946_),
    .C(_16947_),
    .D(_16904_),
    .Y(_16948_));
 INVx1_ASAP7_75t_R _25361_ (.A(_16694_),
    .Y(_16949_));
 AO21x1_ASAP7_75t_R _25362_ (.A1(_16366_),
    .A2(_16395_),
    .B(_16391_),
    .Y(_16950_));
 AND4x1_ASAP7_75t_R _25363_ (.A(_16632_),
    .B(_16405_),
    .C(_16949_),
    .D(_16950_),
    .Y(_16951_));
 AO21x1_ASAP7_75t_R _25364_ (.A1(_16398_),
    .A2(_16426_),
    .B(_16411_),
    .Y(_16952_));
 NAND2x1_ASAP7_75t_R _25365_ (.A(_16311_),
    .B(_16409_),
    .Y(_16953_));
 AND3x1_ASAP7_75t_R _25366_ (.A(_16952_),
    .B(_16953_),
    .C(_16417_),
    .Y(_16954_));
 AND4x1_ASAP7_75t_R _25367_ (.A(_16944_),
    .B(_16948_),
    .C(_16951_),
    .D(_16954_),
    .Y(_16955_));
 AO21x1_ASAP7_75t_R _25368_ (.A1(_16278_),
    .A2(_16341_),
    .B(_16836_),
    .Y(_16956_));
 AND3x1_ASAP7_75t_R _25369_ (.A(_16341_),
    .B(_16300_),
    .C(_16306_),
    .Y(_16957_));
 OR3x1_ASAP7_75t_R _25370_ (.A(_16956_),
    .B(_16661_),
    .C(_16957_),
    .Y(_16958_));
 AO21x1_ASAP7_75t_R _25371_ (.A1(_16317_),
    .A2(_16560_),
    .B(_16653_),
    .Y(_16959_));
 OR4x2_ASAP7_75t_R _25372_ (.A(_16958_),
    .B(_16337_),
    .C(_16655_),
    .D(_16959_),
    .Y(_16960_));
 AND3x1_ASAP7_75t_R _25373_ (.A(_16272_),
    .B(_16287_),
    .C(_16265_),
    .Y(_16961_));
 OR4x2_ASAP7_75t_R _25374_ (.A(_16606_),
    .B(_16961_),
    .C(_16894_),
    .D(_16831_),
    .Y(_16962_));
 NOR2x1_ASAP7_75t_R _25375_ (.A(net3503),
    .B(_16440_),
    .Y(_16963_));
 NOR2x1_ASAP7_75t_R _25376_ (.A(_16293_),
    .B(_16561_),
    .Y(_16964_));
 AO21x1_ASAP7_75t_R _25377_ (.A1(_16386_),
    .A2(_16294_),
    .B(_16964_),
    .Y(_16965_));
 OR5x2_ASAP7_75t_R _25378_ (.A(_16963_),
    .B(_16965_),
    .C(_16313_),
    .D(_16303_),
    .E(_16674_),
    .Y(_16966_));
 NOR3x2_ASAP7_75t_R _25379_ (.B(_16962_),
    .C(_16966_),
    .Y(_16967_),
    .A(_16960_));
 AND3x1_ASAP7_75t_R _25380_ (.A(_16452_),
    .B(_16275_),
    .C(_16306_),
    .Y(_16968_));
 AOI22x1_ASAP7_75t_R _25381_ (.A1(_16968_),
    .A2(_16300_),
    .B1(_16452_),
    .B2(_16296_),
    .Y(_16969_));
 AND2x2_ASAP7_75t_R _25382_ (.A(_16334_),
    .B(_16452_),
    .Y(_16970_));
 INVx1_ASAP7_75t_R _25383_ (.A(_16970_),
    .Y(_16971_));
 AO21x1_ASAP7_75t_R _25384_ (.A1(_16542_),
    .A2(_16279_),
    .B(_16563_),
    .Y(_16972_));
 AND3x1_ASAP7_75t_R _25385_ (.A(_16969_),
    .B(_16971_),
    .C(_16972_),
    .Y(_16973_));
 AO21x1_ASAP7_75t_R _25386_ (.A1(_16445_),
    .A2(_16621_),
    .B(_16471_),
    .Y(_16974_));
 OA211x2_ASAP7_75t_R _25387_ (.A1(_16366_),
    .A2(_16471_),
    .B(_16974_),
    .C(_16801_),
    .Y(_16975_));
 AO21x1_ASAP7_75t_R _25388_ (.A1(_16387_),
    .A2(_16295_),
    .B(_16460_),
    .Y(_16976_));
 NOR2x1_ASAP7_75t_R _25389_ (.A(_16279_),
    .B(_16460_),
    .Y(_16977_));
 INVx1_ASAP7_75t_R _25390_ (.A(_16977_),
    .Y(_16978_));
 AND4x1_ASAP7_75t_R _25391_ (.A(_16976_),
    .B(_16978_),
    .C(_16736_),
    .D(_16857_),
    .Y(_16979_));
 OA211x2_ASAP7_75t_R _25392_ (.A1(_16437_),
    .A2(_16440_),
    .B(_16583_),
    .C(_16794_),
    .Y(_16980_));
 AND3x1_ASAP7_75t_R _25393_ (.A(_16434_),
    .B(net2209),
    .C(_16265_),
    .Y(_16981_));
 INVx1_ASAP7_75t_R _25394_ (.A(_16981_),
    .Y(_16982_));
 OA21x2_ASAP7_75t_R _25395_ (.A1(_16437_),
    .A2(net3499),
    .B(_16982_),
    .Y(_16983_));
 AND5x1_ASAP7_75t_R _25396_ (.A(_16973_),
    .B(_16975_),
    .C(_16979_),
    .D(_16980_),
    .E(_16983_),
    .Y(_16984_));
 AND4x1_ASAP7_75t_R _25397_ (.A(_16942_),
    .B(_16955_),
    .C(_16967_),
    .D(_16984_),
    .Y(_16985_));
 NAND2x2_ASAP7_75t_R _25398_ (.A(_16985_),
    .B(_16524_),
    .Y(_16986_));
 XOR2x2_ASAP7_75t_R _25399_ (.A(_00455_),
    .B(_00503_),
    .Y(_16987_));
 XOR2x1_ASAP7_75t_R _25400_ (.A(_00405_),
    .Y(_16988_),
    .B(_00423_));
 XOR2x1_ASAP7_75t_R _25401_ (.A(_16987_),
    .Y(_16989_),
    .B(_16988_));
 XOR2x1_ASAP7_75t_R _25402_ (.A(_16989_),
    .Y(_16990_),
    .B(_00404_));
 XOR2x2_ASAP7_75t_R _25403_ (.A(_16986_),
    .B(_16990_),
    .Y(_16991_));
 NAND2x1_ASAP7_75t_R _25404_ (.A(net404),
    .B(net3881),
    .Y(_16992_));
 OAI21x1_ASAP7_75t_R _25405_ (.A1(net404),
    .A2(_16991_),
    .B(net3882),
    .Y(_00374_));
 NAND2x1_ASAP7_75t_R _25406_ (.A(_16369_),
    .B(_16390_),
    .Y(_16993_));
 NAND2x1_ASAP7_75t_R _25407_ (.A(_16344_),
    .B(_16390_),
    .Y(_16994_));
 AND4x1_ASAP7_75t_R _25408_ (.A(_16915_),
    .B(_16806_),
    .C(_16993_),
    .D(_16994_),
    .Y(_16995_));
 AND5x1_ASAP7_75t_R _25409_ (.A(_16953_),
    .B(_16995_),
    .C(_16424_),
    .D(_16808_),
    .E(_16415_),
    .Y(_16996_));
 AO21x1_ASAP7_75t_R _25410_ (.A1(_16421_),
    .A2(_16366_),
    .B(_16378_),
    .Y(_16997_));
 NAND2x1_ASAP7_75t_R _25411_ (.A(_16306_),
    .B(_16376_),
    .Y(_16998_));
 AND4x1_ASAP7_75t_R _25412_ (.A(_16997_),
    .B(_16998_),
    .C(_16823_),
    .D(_16908_),
    .Y(_16999_));
 AND3x1_ASAP7_75t_R _25413_ (.A(_16999_),
    .B(_16518_),
    .C(_16679_),
    .Y(_17000_));
 AND2x2_ASAP7_75t_R _25414_ (.A(_16996_),
    .B(_17000_),
    .Y(_17001_));
 AO21x1_ASAP7_75t_R _25415_ (.A1(_16440_),
    .A2(_16325_),
    .B(_16283_),
    .Y(_17002_));
 AO21x1_ASAP7_75t_R _25416_ (.A1(_16357_),
    .A2(_16445_),
    .B(_16283_),
    .Y(_17003_));
 INVx1_ASAP7_75t_R _25417_ (.A(_16469_),
    .Y(_17004_));
 NAND2x1_ASAP7_75t_R _25418_ (.A(_16272_),
    .B(_17004_),
    .Y(_17005_));
 NAND2x1_ASAP7_75t_R _25419_ (.A(_16272_),
    .B(_16394_),
    .Y(_17006_));
 AND5x1_ASAP7_75t_R _25420_ (.A(_17002_),
    .B(_17003_),
    .C(_16284_),
    .D(_17005_),
    .E(_17006_),
    .Y(_17007_));
 AO21x1_ASAP7_75t_R _25421_ (.A1(_16387_),
    .A2(_16357_),
    .B(_16327_),
    .Y(_17008_));
 AO21x1_ASAP7_75t_R _25422_ (.A1(net3499),
    .A2(_16279_),
    .B(_16327_),
    .Y(_17009_));
 OA211x2_ASAP7_75t_R _25423_ (.A1(_16335_),
    .A2(_16327_),
    .B(_17008_),
    .C(_17009_),
    .Y(_17010_));
 INVx1_ASAP7_75t_R _25424_ (.A(_16346_),
    .Y(_17011_));
 OA211x2_ASAP7_75t_R _25425_ (.A1(_16342_),
    .A2(_16838_),
    .B(_17011_),
    .C(_16842_),
    .Y(_17012_));
 NOR2x1_ASAP7_75t_R _25426_ (.A(_16613_),
    .B(_16612_),
    .Y(_17013_));
 AO21x1_ASAP7_75t_R _25427_ (.A1(_16463_),
    .A2(_16325_),
    .B(_16293_),
    .Y(_17014_));
 OA211x2_ASAP7_75t_R _25428_ (.A1(_16561_),
    .A2(_16293_),
    .B(_17013_),
    .C(_17014_),
    .Y(_17015_));
 AND4x1_ASAP7_75t_R _25429_ (.A(_17007_),
    .B(_17010_),
    .C(_17012_),
    .D(_17015_),
    .Y(_17016_));
 OA211x2_ASAP7_75t_R _25430_ (.A1(_16542_),
    .A2(_16563_),
    .B(_16568_),
    .C(_16786_),
    .Y(_17017_));
 OA211x2_ASAP7_75t_R _25431_ (.A1(_16335_),
    .A2(_16460_),
    .B(_16574_),
    .C(_16978_),
    .Y(_17018_));
 AND2x2_ASAP7_75t_R _25432_ (.A(_16459_),
    .B(_16301_),
    .Y(_17019_));
 OA21x2_ASAP7_75t_R _25433_ (.A1(net1744),
    .A2(_16318_),
    .B(_16459_),
    .Y(_17020_));
 AOI21x1_ASAP7_75t_R _25434_ (.A1(_16296_),
    .A2(_17019_),
    .B(_17020_),
    .Y(_17021_));
 AO21x1_ASAP7_75t_R _25435_ (.A1(_16561_),
    .A2(_16440_),
    .B(_16563_),
    .Y(_17022_));
 AND4x1_ASAP7_75t_R _25436_ (.A(_17017_),
    .B(_17018_),
    .C(_17021_),
    .D(_17022_),
    .Y(_17023_));
 NOR2x1_ASAP7_75t_R _25437_ (.A(_16621_),
    .B(_16471_),
    .Y(_17024_));
 INVx1_ASAP7_75t_R _25438_ (.A(_17024_),
    .Y(_17025_));
 AND4x1_ASAP7_75t_R _25439_ (.A(_16476_),
    .B(_16801_),
    .C(_17025_),
    .D(_16722_),
    .Y(_17026_));
 OA211x2_ASAP7_75t_R _25440_ (.A1(_16262_),
    .A2(_16287_),
    .B(_16434_),
    .C(_16306_),
    .Y(_17027_));
 INVx1_ASAP7_75t_R _25441_ (.A(_17027_),
    .Y(_17028_));
 OA211x2_ASAP7_75t_R _25442_ (.A1(_16437_),
    .A2(_16335_),
    .B(_17028_),
    .C(_16435_),
    .Y(_17029_));
 AND3x1_ASAP7_75t_R _25443_ (.A(_17023_),
    .B(_17026_),
    .C(_17029_),
    .Y(_17030_));
 AO21x1_ASAP7_75t_R _25444_ (.A1(_16387_),
    .A2(_16445_),
    .B(_16495_),
    .Y(_17031_));
 AO21x1_ASAP7_75t_R _25445_ (.A1(_16325_),
    .A2(_16469_),
    .B(_16495_),
    .Y(_17032_));
 AND2x2_ASAP7_75t_R _25446_ (.A(_17031_),
    .B(_17032_),
    .Y(_17033_));
 AO21x1_ASAP7_75t_R _25447_ (.A1(net3499),
    .A2(_16279_),
    .B(_16495_),
    .Y(_17034_));
 AO21x1_ASAP7_75t_R _25448_ (.A1(_16421_),
    .A2(_16426_),
    .B(_16495_),
    .Y(_17035_));
 AO21x1_ASAP7_75t_R _25449_ (.A1(_16325_),
    .A2(_16443_),
    .B(_16488_),
    .Y(_17036_));
 AO21x1_ASAP7_75t_R _25450_ (.A1(_16539_),
    .A2(_16511_),
    .B(_16488_),
    .Y(_17037_));
 AND5x1_ASAP7_75t_R _25451_ (.A(_17033_),
    .B(_17034_),
    .C(_17035_),
    .D(_17036_),
    .E(_17037_),
    .Y(_17038_));
 NOR2x1_ASAP7_75t_R _25452_ (.A(_16325_),
    .B(_16512_),
    .Y(_17039_));
 INVx1_ASAP7_75t_R _25453_ (.A(_17039_),
    .Y(_17040_));
 AO21x1_ASAP7_75t_R _25454_ (.A1(_16421_),
    .A2(_16366_),
    .B(_16512_),
    .Y(_17041_));
 AND4x1_ASAP7_75t_R _25455_ (.A(_16554_),
    .B(_17040_),
    .C(_17041_),
    .D(_16766_),
    .Y(_17042_));
 NOR2x1_ASAP7_75t_R _25456_ (.A(_16621_),
    .B(_16504_),
    .Y(_17043_));
 AO21x1_ASAP7_75t_R _25457_ (.A1(_17004_),
    .A2(_16501_),
    .B(_17043_),
    .Y(_17044_));
 OA21x2_ASAP7_75t_R _25458_ (.A1(_16381_),
    .A2(_16425_),
    .B(_16501_),
    .Y(_17045_));
 NAND2x1_ASAP7_75t_R _25459_ (.A(_16713_),
    .B(_16710_),
    .Y(_17046_));
 OR3x1_ASAP7_75t_R _25460_ (.A(_17044_),
    .B(_17045_),
    .C(_17046_),
    .Y(_17047_));
 INVx1_ASAP7_75t_R _25461_ (.A(_17047_),
    .Y(_17048_));
 AND3x1_ASAP7_75t_R _25462_ (.A(_17038_),
    .B(_17042_),
    .C(_17048_),
    .Y(_17049_));
 AND2x2_ASAP7_75t_R _25463_ (.A(_17030_),
    .B(_17049_),
    .Y(_17050_));
 AND3x4_ASAP7_75t_R _25464_ (.A(_17001_),
    .B(_17016_),
    .C(_17050_),
    .Y(_17051_));
 NAND2x2_ASAP7_75t_R _25465_ (.A(_17051_),
    .B(_16524_),
    .Y(_17052_));
 XOR2x2_ASAP7_75t_R _25466_ (.A(_00407_),
    .B(_00406_),
    .Y(_17053_));
 XOR2x1_ASAP7_75t_R _25467_ (.A(_17053_),
    .Y(_17054_),
    .B(_06342_));
 BUFx2_ASAP7_75t_R output271 (.A(net271),
    .Y(text_out[10]));
 XOR2x2_ASAP7_75t_R _25469_ (.A(_00454_),
    .B(_00502_),
    .Y(_17056_));
 INVx1_ASAP7_75t_R _25470_ (.A(_17056_),
    .Y(_17057_));
 XOR2x1_ASAP7_75t_R _25471_ (.A(_17054_),
    .Y(_17058_),
    .B(_17057_));
 XOR2x1_ASAP7_75t_R _25472_ (.A(_17052_),
    .Y(_17059_),
    .B(_17058_));
 NOR2x1_ASAP7_75t_R _25473_ (.A(net4152),
    .B(net400),
    .Y(_17060_));
 AOI21x1_ASAP7_75t_R _25474_ (.A1(net400),
    .A2(_17059_),
    .B(_17060_),
    .Y(_00376_));
 BUFx2_ASAP7_75t_R output270 (.A(net270),
    .Y(text_out[109]));
 XNOR2x1_ASAP7_75t_R _25476_ (.B(_00501_),
    .Y(_17062_),
    .A(_00485_));
 XNOR2x1_ASAP7_75t_R _25477_ (.B(_00453_),
    .Y(_17063_),
    .A(net3385));
 XOR2x1_ASAP7_75t_R _25478_ (.A(_17062_),
    .Y(_17064_),
    .B(_17063_));
 XOR2x1_ASAP7_75t_R _25479_ (.A(_17064_),
    .Y(_17065_),
    .B(_00408_));
 OA211x2_ASAP7_75t_R _25480_ (.A1(net1854),
    .A2(_16287_),
    .B(_16459_),
    .C(_16265_),
    .Y(_17066_));
 NAND2x1_ASAP7_75t_R _25481_ (.A(_16864_),
    .B(_16731_),
    .Y(_17067_));
 OR3x1_ASAP7_75t_R _25482_ (.A(_17066_),
    .B(_16856_),
    .C(_17067_),
    .Y(_17068_));
 INVx1_ASAP7_75t_R _25483_ (.A(_16786_),
    .Y(_17069_));
 NOR2x1_ASAP7_75t_R _25484_ (.A(_16325_),
    .B(_16563_),
    .Y(_17070_));
 OR5x1_ASAP7_75t_R _25485_ (.A(_17069_),
    .B(_16968_),
    .C(_17070_),
    .D(_16970_),
    .E(_16569_),
    .Y(_17071_));
 NOR2x1_ASAP7_75t_R _25486_ (.A(_17068_),
    .B(_17071_),
    .Y(_17072_));
 AO21x1_ASAP7_75t_R _25487_ (.A1(_16416_),
    .A2(_16467_),
    .B(_17024_),
    .Y(_17073_));
 OA21x2_ASAP7_75t_R _25488_ (.A1(_16356_),
    .A2(_16344_),
    .B(_16467_),
    .Y(_17074_));
 OR4x1_ASAP7_75t_R _25489_ (.A(_17073_),
    .B(_16474_),
    .C(_16588_),
    .D(_17074_),
    .Y(_17075_));
 OA211x2_ASAP7_75t_R _25490_ (.A1(net3481),
    .A2(net2209),
    .B(_16434_),
    .C(_16296_),
    .Y(_17076_));
 INVx1_ASAP7_75t_R _25491_ (.A(_17076_),
    .Y(_17077_));
 AND2x2_ASAP7_75t_R _25492_ (.A(_16434_),
    .B(_16373_),
    .Y(_17078_));
 INVx1_ASAP7_75t_R _25493_ (.A(_17078_),
    .Y(_17079_));
 AND4x1_ASAP7_75t_R _25494_ (.A(_17077_),
    .B(_17079_),
    .C(_16583_),
    .D(_16982_),
    .Y(_17080_));
 INVx1_ASAP7_75t_R _25495_ (.A(_17080_),
    .Y(_17081_));
 NOR2x2_ASAP7_75t_R _25496_ (.A(_17075_),
    .B(_17081_),
    .Y(_17082_));
 NAND2x2_ASAP7_75t_R _25497_ (.A(_17072_),
    .B(_17082_),
    .Y(_17083_));
 INVx1_ASAP7_75t_R _25498_ (.A(_16778_),
    .Y(_17084_));
 AO21x1_ASAP7_75t_R _25499_ (.A1(_16440_),
    .A2(_16469_),
    .B(_16488_),
    .Y(_17085_));
 AO21x1_ASAP7_75t_R _25500_ (.A1(_16421_),
    .A2(_16395_),
    .B(_16488_),
    .Y(_17086_));
 AO21x1_ASAP7_75t_R _25501_ (.A1(_16561_),
    .A2(_16387_),
    .B(_16488_),
    .Y(_17087_));
 AND4x1_ASAP7_75t_R _25502_ (.A(_17084_),
    .B(_17085_),
    .C(_17086_),
    .D(_17087_),
    .Y(_17088_));
 NAND2x1_ASAP7_75t_R _25503_ (.A(_16538_),
    .B(_16484_),
    .Y(_17089_));
 OA211x2_ASAP7_75t_R _25504_ (.A1(_16357_),
    .A2(_16495_),
    .B(_17032_),
    .C(_17089_),
    .Y(_17090_));
 AND2x2_ASAP7_75t_R _25505_ (.A(_17088_),
    .B(_17090_),
    .Y(_17091_));
 INVx1_ASAP7_75t_R _25506_ (.A(_17091_),
    .Y(_17092_));
 NAND2x1_ASAP7_75t_R _25507_ (.A(_16529_),
    .B(_16939_),
    .Y(_17093_));
 AOI221x1_ASAP7_75t_R _25508_ (.A1(_16262_),
    .A2(_16287_),
    .B1(net3493),
    .B2(_16266_),
    .C(_16512_),
    .Y(_17094_));
 OR5x2_ASAP7_75t_R _25509_ (.A(_17039_),
    .B(_17093_),
    .C(_17043_),
    .D(_16507_),
    .E(_17094_),
    .Y(_17095_));
 NOR3x2_ASAP7_75t_R _25510_ (.B(_17092_),
    .C(_17095_),
    .Y(_17096_),
    .A(_17083_));
 OA21x2_ASAP7_75t_R _25511_ (.A1(net2492),
    .A2(_16318_),
    .B(_16353_),
    .Y(_17097_));
 AOI221x1_ASAP7_75t_R _25512_ (.A1(net1854),
    .A2(_16520_),
    .B1(_16353_),
    .B2(_16267_),
    .C(_17097_),
    .Y(_17098_));
 AND4x1_ASAP7_75t_R _25513_ (.A(_16403_),
    .B(_16407_),
    .C(_16994_),
    .D(_16810_),
    .Y(_17099_));
 AO21x1_ASAP7_75t_R _25514_ (.A1(_16421_),
    .A2(_16426_),
    .B(_16378_),
    .Y(_17100_));
 AO21x1_ASAP7_75t_R _25515_ (.A1(_16463_),
    .A2(_16621_),
    .B(_16378_),
    .Y(_17101_));
 AND4x1_ASAP7_75t_R _25516_ (.A(_17100_),
    .B(_16946_),
    .C(_17101_),
    .D(_16382_),
    .Y(_17102_));
 NOR2x1_ASAP7_75t_R _25517_ (.A(_16414_),
    .B(_16630_),
    .Y(_17103_));
 AO21x1_ASAP7_75t_R _25518_ (.A1(_16366_),
    .A2(_16395_),
    .B(_16411_),
    .Y(_17104_));
 NAND2x1_ASAP7_75t_R _25519_ (.A(_16369_),
    .B(_16409_),
    .Y(_17105_));
 AND2x2_ASAP7_75t_R _25520_ (.A(_17104_),
    .B(_17105_),
    .Y(_17106_));
 AND5x1_ASAP7_75t_R _25521_ (.A(_17098_),
    .B(_17099_),
    .C(_17102_),
    .D(_17103_),
    .E(_17106_),
    .Y(_17107_));
 AO21x1_ASAP7_75t_R _25522_ (.A1(_16421_),
    .A2(_16335_),
    .B(_16327_),
    .Y(_17108_));
 AO21x1_ASAP7_75t_R _25523_ (.A1(_16561_),
    .A2(_16440_),
    .B(_16327_),
    .Y(_17109_));
 OA211x2_ASAP7_75t_R _25524_ (.A1(_16370_),
    .A2(_16327_),
    .B(_17108_),
    .C(_17109_),
    .Y(_17110_));
 OR3x1_ASAP7_75t_R _25525_ (.A(_16612_),
    .B(_16613_),
    .C(_16674_),
    .Y(_17111_));
 AND3x1_ASAP7_75t_R _25526_ (.A(_16294_),
    .B(net3478),
    .C(_16306_),
    .Y(_17112_));
 OR3x1_ASAP7_75t_R _25527_ (.A(_17112_),
    .B(_16617_),
    .C(_16964_),
    .Y(_17113_));
 NOR2x1_ASAP7_75t_R _25528_ (.A(_17111_),
    .B(_17113_),
    .Y(_17114_));
 AO21x1_ASAP7_75t_R _25529_ (.A1(_16387_),
    .A2(_16357_),
    .B(_16342_),
    .Y(_17115_));
 AO21x1_ASAP7_75t_R _25530_ (.A1(_16436_),
    .A2(_16542_),
    .B(_16342_),
    .Y(_17116_));
 AO21x1_ASAP7_75t_R _25531_ (.A1(_16440_),
    .A2(_16469_),
    .B(_16342_),
    .Y(_17117_));
 AND4x1_ASAP7_75t_R _25532_ (.A(_17115_),
    .B(_17116_),
    .C(_17117_),
    .D(_16349_),
    .Y(_17118_));
 AO21x1_ASAP7_75t_R _25533_ (.A1(_16561_),
    .A2(_16295_),
    .B(_16283_),
    .Y(_17119_));
 AO21x1_ASAP7_75t_R _25534_ (.A1(_16398_),
    .A2(_16436_),
    .B(_16283_),
    .Y(_17120_));
 AND5x2_ASAP7_75t_R _25535_ (.A(_17110_),
    .B(_17114_),
    .C(_17118_),
    .D(_17119_),
    .E(_17120_),
    .Y(_17121_));
 NAND2x2_ASAP7_75t_R _25536_ (.A(_17107_),
    .B(_17121_),
    .Y(_17122_));
 INVx1_ASAP7_75t_R _25537_ (.A(_17122_),
    .Y(_17123_));
 NAND2x2_ASAP7_75t_R _25538_ (.A(_17096_),
    .B(_17123_),
    .Y(_17124_));
 XNOR2x1_ASAP7_75t_R _25539_ (.B(_17124_),
    .Y(_17125_),
    .A(_17065_));
 AND2x2_ASAP7_75t_R _25540_ (.A(net401),
    .B(net53),
    .Y(_17126_));
 AO21x1_ASAP7_75t_R _25541_ (.A1(_17125_),
    .A2(net399),
    .B(_17126_),
    .Y(_00377_));
 NAND2x2_ASAP7_75t_R _25542_ (.A(_06375_),
    .B(_08724_),
    .Y(_17127_));
 XOR2x2_ASAP7_75t_R _25543_ (.A(_00409_),
    .B(_00500_),
    .Y(_17128_));
 XOR2x1_ASAP7_75t_R _25544_ (.A(_17128_),
    .Y(_17129_),
    .B(_00484_));
 XOR2x1_ASAP7_75t_R _25545_ (.A(_17127_),
    .Y(_17130_),
    .B(_17129_));
 NOR2x1_ASAP7_75t_R _25546_ (.A(net4104),
    .B(net400),
    .Y(_17131_));
 AOI21x1_ASAP7_75t_R _25547_ (.A1(net400),
    .A2(_17130_),
    .B(_17131_),
    .Y(_00321_));
 BUFx2_ASAP7_75t_R output269 (.A(net269),
    .Y(text_out[108]));
 NOR2x2_ASAP7_75t_R _25549_ (.A(_10127_),
    .B(_10116_),
    .Y(_17133_));
 XOR2x2_ASAP7_75t_R _25550_ (.A(_00410_),
    .B(_00499_),
    .Y(_17134_));
 XOR2x1_ASAP7_75t_R _25551_ (.A(_17134_),
    .Y(_17135_),
    .B(_10171_));
 XOR2x1_ASAP7_75t_R _25552_ (.A(_17133_),
    .Y(_17136_),
    .B(_17135_));
 NOR2x1_ASAP7_75t_R _25553_ (.A(net4102),
    .B(net400),
    .Y(_17137_));
 AOI21x1_ASAP7_75t_R _25554_ (.A1(net400),
    .A2(_17136_),
    .B(_17137_),
    .Y(_00332_));
 NAND2x1_ASAP7_75t_R _25555_ (.A(net403),
    .B(net4066),
    .Y(_17138_));
 INVx5_ASAP7_75t_R _25556_ (.A(_00385_),
    .Y(_17139_));
 XOR2x1_ASAP7_75t_R _25557_ (.A(_11247_),
    .Y(_17140_),
    .B(_17139_));
 NOR2x1_ASAP7_75t_R _25558_ (.A(_17140_),
    .B(_11214_),
    .Y(_17141_));
 AND2x2_ASAP7_75t_R _25559_ (.A(_11214_),
    .B(_17140_),
    .Y(_17142_));
 OAI21x1_ASAP7_75t_R _25560_ (.A1(_17141_),
    .A2(_17142_),
    .B(net400),
    .Y(_17143_));
 NAND2x1_ASAP7_75t_R _25561_ (.A(_17138_),
    .B(_17143_),
    .Y(_00343_));
 INVx2_ASAP7_75t_R _25562_ (.A(net4084),
    .Y(_17144_));
 INVx4_ASAP7_75t_R _25563_ (.A(_00386_),
    .Y(_17145_));
 XOR2x1_ASAP7_75t_R _25564_ (.A(_12234_),
    .Y(_17146_),
    .B(_17145_));
 INVx1_ASAP7_75t_R _25565_ (.A(_17146_),
    .Y(_17147_));
 NOR2x1_ASAP7_75t_R _25566_ (.A(_17147_),
    .B(_12212_),
    .Y(_17148_));
 AND2x2_ASAP7_75t_R _25567_ (.A(_12212_),
    .B(_17147_),
    .Y(_17149_));
 BUFx2_ASAP7_75t_R output268 (.A(net268),
    .Y(text_out[107]));
 OAI21x1_ASAP7_75t_R _25569_ (.A1(_17148_),
    .A2(_17149_),
    .B(net399),
    .Y(_17151_));
 OAI21x1_ASAP7_75t_R _25570_ (.A1(net399),
    .A2(_17144_),
    .B(_17151_),
    .Y(_00346_));
 INVx1_ASAP7_75t_R _25571_ (.A(net4092),
    .Y(_17152_));
 XOR2x1_ASAP7_75t_R _25572_ (.A(_13023_),
    .Y(_17153_),
    .B(_00387_));
 INVx1_ASAP7_75t_R _25573_ (.A(_17153_),
    .Y(_17154_));
 NOR2x1_ASAP7_75t_R _25574_ (.A(_17154_),
    .B(_13001_),
    .Y(_17155_));
 AND2x2_ASAP7_75t_R _25575_ (.A(_13001_),
    .B(_17154_),
    .Y(_17156_));
 OAI21x1_ASAP7_75t_R _25576_ (.A1(_17155_),
    .A2(_17156_),
    .B(net399),
    .Y(_17157_));
 OAI21x1_ASAP7_75t_R _25577_ (.A1(net399),
    .A2(_17152_),
    .B(_17157_),
    .Y(_00347_));
 NAND2x2_ASAP7_75t_R _25578_ (.A(net403),
    .B(net4110),
    .Y(_17158_));
 XOR2x1_ASAP7_75t_R _25579_ (.A(_00479_),
    .Y(_17159_),
    .B(_00521_));
 INVx1_ASAP7_75t_R _25580_ (.A(_00498_),
    .Y(_17160_));
 XOR2x1_ASAP7_75t_R _25581_ (.A(_17159_),
    .Y(_17161_),
    .B(_17160_));
 NOR2x1_ASAP7_75t_R _25582_ (.A(_17161_),
    .B(_13790_),
    .Y(_17162_));
 AND2x2_ASAP7_75t_R _25583_ (.A(_13790_),
    .B(_17161_),
    .Y(_17163_));
 OAI21x1_ASAP7_75t_R _25584_ (.A1(_17162_),
    .A2(_17163_),
    .B(net400),
    .Y(_17164_));
 NAND2x1_ASAP7_75t_R _25585_ (.A(_17158_),
    .B(_17164_),
    .Y(_00348_));
 NAND2x2_ASAP7_75t_R _25586_ (.A(_14355_),
    .B(_06375_),
    .Y(_17165_));
 XOR2x2_ASAP7_75t_R _25587_ (.A(_00411_),
    .B(_00497_),
    .Y(_17166_));
 XOR2x1_ASAP7_75t_R _25588_ (.A(_17166_),
    .Y(_17167_),
    .B(_14358_));
 XOR2x2_ASAP7_75t_R _25589_ (.A(_17165_),
    .B(_17167_),
    .Y(_17168_));
 AND2x2_ASAP7_75t_R _25590_ (.A(net403),
    .B(net60),
    .Y(_17169_));
 AO21x1_ASAP7_75t_R _25591_ (.A1(_17168_),
    .A2(net400),
    .B(_17169_),
    .Y(_00349_));
 NAND2x1_ASAP7_75t_R _25592_ (.A(net405),
    .B(net4116),
    .Y(_17170_));
 INVx4_ASAP7_75t_R _25593_ (.A(_00388_),
    .Y(_17171_));
 XOR2x1_ASAP7_75t_R _25594_ (.A(_14590_),
    .Y(_17172_),
    .B(_17171_));
 OR3x1_ASAP7_75t_R _25595_ (.A(_14588_),
    .B(_14536_),
    .C(_17172_),
    .Y(_17173_));
 OAI21x1_ASAP7_75t_R _25596_ (.A1(_14536_),
    .A2(_14588_),
    .B(_17172_),
    .Y(_17174_));
 BUFx2_ASAP7_75t_R output267 (.A(net267),
    .Y(text_out[106]));
 AO21x1_ASAP7_75t_R _25598_ (.A1(_17173_),
    .A2(_17174_),
    .B(net405),
    .Y(_17176_));
 NAND2x1_ASAP7_75t_R _25599_ (.A(_17170_),
    .B(_17176_),
    .Y(_00350_));
 BUFx2_ASAP7_75t_R output266 (.A(net266),
    .Y(text_out[105]));
 XOR2x2_ASAP7_75t_R _25601_ (.A(_00412_),
    .B(_00496_),
    .Y(_17178_));
 XOR2x1_ASAP7_75t_R _25602_ (.A(_17178_),
    .Y(_17179_),
    .B(_14601_));
 XOR2x1_ASAP7_75t_R _25603_ (.A(_14844_),
    .Y(_17180_),
    .B(_17179_));
 NAND2x1_ASAP7_75t_R _25604_ (.A(net400),
    .B(_17180_),
    .Y(_17181_));
 OA21x2_ASAP7_75t_R _25605_ (.A1(net400),
    .A2(net4042),
    .B(_17181_),
    .Y(_00351_));
 INVx2_ASAP7_75t_R _25606_ (.A(net4058),
    .Y(_17182_));
 XOR2x1_ASAP7_75t_R _25607_ (.A(_00475_),
    .Y(_17183_),
    .B(_00519_));
 INVx3_ASAP7_75t_R _25608_ (.A(_00495_),
    .Y(_17184_));
 XOR2x1_ASAP7_75t_R _25609_ (.A(_17183_),
    .Y(_17185_),
    .B(_17184_));
 AND4x1_ASAP7_75t_R _25610_ (.A(_14904_),
    .B(_14905_),
    .C(_14958_),
    .D(_17185_),
    .Y(_17186_));
 NOR2x1_ASAP7_75t_R _25611_ (.A(_17185_),
    .B(_14959_),
    .Y(_17187_));
 OAI21x1_ASAP7_75t_R _25612_ (.A1(_17186_),
    .A2(_17187_),
    .B(net399),
    .Y(_17188_));
 OAI21x1_ASAP7_75t_R _25613_ (.A1(net399),
    .A2(_17182_),
    .B(_17188_),
    .Y(_00352_));
 XOR2x1_ASAP7_75t_R _25614_ (.A(_15054_),
    .Y(_17189_),
    .B(_00389_));
 OAI21x1_ASAP7_75t_R _25615_ (.A1(_15009_),
    .A2(_15052_),
    .B(_17189_),
    .Y(_17190_));
 OR3x1_ASAP7_75t_R _25616_ (.A(_15052_),
    .B(_15009_),
    .C(_17189_),
    .Y(_17191_));
 AOI21x1_ASAP7_75t_R _25617_ (.A1(_17190_),
    .A2(_17191_),
    .B(net405),
    .Y(_17192_));
 AO21x1_ASAP7_75t_R _25618_ (.A1(net405),
    .A2(net4100),
    .B(_17192_),
    .Y(_00322_));
 NAND2x2_ASAP7_75t_R _25619_ (.A(net404),
    .B(net3999),
    .Y(_17193_));
 XOR2x1_ASAP7_75t_R _25620_ (.A(_15139_),
    .Y(_17194_),
    .B(_00390_));
 OR3x1_ASAP7_75t_R _25621_ (.A(_15136_),
    .B(_15094_),
    .C(_17194_),
    .Y(_17195_));
 OAI21x1_ASAP7_75t_R _25622_ (.A1(_15094_),
    .A2(_15136_),
    .B(_17194_),
    .Y(_17196_));
 AO21x1_ASAP7_75t_R _25623_ (.A1(_17195_),
    .A2(_17196_),
    .B(net405),
    .Y(_17197_));
 NAND2x1_ASAP7_75t_R _25624_ (.A(net4000),
    .B(_17197_),
    .Y(_00323_));
 INVx1_ASAP7_75t_R _25625_ (.A(net3890),
    .Y(_17198_));
 INVx2_ASAP7_75t_R _25626_ (.A(_00391_),
    .Y(_17199_));
 XOR2x1_ASAP7_75t_R _25627_ (.A(_15206_),
    .Y(_17200_),
    .B(_17199_));
 NOR2x1_ASAP7_75t_R _25628_ (.A(_17200_),
    .B(_15203_),
    .Y(_17201_));
 AND2x2_ASAP7_75t_R _25629_ (.A(_15203_),
    .B(_17200_),
    .Y(_17202_));
 OAI21x1_ASAP7_75t_R _25630_ (.A1(_17201_),
    .A2(_17202_),
    .B(net399),
    .Y(_17203_));
 OAI21x1_ASAP7_75t_R _25631_ (.A1(net399),
    .A2(net3891),
    .B(_17203_),
    .Y(_00324_));
 NAND2x2_ASAP7_75t_R _25632_ (.A(net402),
    .B(net4064),
    .Y(_17204_));
 XOR2x1_ASAP7_75t_R _25633_ (.A(_00471_),
    .Y(_17205_),
    .B(_00515_));
 INVx2_ASAP7_75t_R _25634_ (.A(_00494_),
    .Y(_17206_));
 XOR2x1_ASAP7_75t_R _25635_ (.A(_17205_),
    .Y(_17207_),
    .B(_17206_));
 AOI21x1_ASAP7_75t_R _25636_ (.A1(_14905_),
    .A2(_15267_),
    .B(_17207_),
    .Y(_17208_));
 INVx1_ASAP7_75t_R _25637_ (.A(_17207_),
    .Y(_17209_));
 NOR2x1_ASAP7_75t_R _25638_ (.A(_17209_),
    .B(_15268_),
    .Y(_17210_));
 OAI21x1_ASAP7_75t_R _25639_ (.A1(_17208_),
    .A2(_17210_),
    .B(net398),
    .Y(_17211_));
 NAND2x1_ASAP7_75t_R _25640_ (.A(_17204_),
    .B(_17211_),
    .Y(_00325_));
 INVx1_ASAP7_75t_R _25641_ (.A(net4050),
    .Y(_17212_));
 XOR2x1_ASAP7_75t_R _25642_ (.A(_00470_),
    .Y(_17213_),
    .B(_00514_));
 INVx2_ASAP7_75t_R _25643_ (.A(_00493_),
    .Y(_17214_));
 XOR2x1_ASAP7_75t_R _25644_ (.A(_17213_),
    .Y(_17215_),
    .B(_17214_));
 AOI21x1_ASAP7_75t_R _25645_ (.A1(_14905_),
    .A2(_15333_),
    .B(_17215_),
    .Y(_17216_));
 AND3x1_ASAP7_75t_R _25646_ (.A(_15333_),
    .B(_14905_),
    .C(_17215_),
    .Y(_17217_));
 OAI21x1_ASAP7_75t_R _25647_ (.A1(_17216_),
    .A2(_17217_),
    .B(net398),
    .Y(_17218_));
 OAI21x1_ASAP7_75t_R _25648_ (.A1(net398),
    .A2(_17212_),
    .B(_17218_),
    .Y(_00326_));
 INVx1_ASAP7_75t_R _25649_ (.A(net3982),
    .Y(_17219_));
 INVx2_ASAP7_75t_R _25650_ (.A(_00392_),
    .Y(_17220_));
 XOR2x1_ASAP7_75t_R _25651_ (.A(_15337_),
    .Y(_17221_),
    .B(_17220_));
 NOR2x1_ASAP7_75t_R _25652_ (.A(_17221_),
    .B(_15391_),
    .Y(_17222_));
 AND2x2_ASAP7_75t_R _25653_ (.A(_15391_),
    .B(_17221_),
    .Y(_17223_));
 OAI21x1_ASAP7_75t_R _25654_ (.A1(_17222_),
    .A2(_17223_),
    .B(net398),
    .Y(_17224_));
 OAI21x1_ASAP7_75t_R _25655_ (.A1(net398),
    .A2(net3983),
    .B(_17224_),
    .Y(_00327_));
 NOR2x2_ASAP7_75t_R _25656_ (.A(_15657_),
    .B(_15649_),
    .Y(_17225_));
 XOR2x2_ASAP7_75t_R _25657_ (.A(_00413_),
    .B(_00492_),
    .Y(_17226_));
 XOR2x1_ASAP7_75t_R _25658_ (.A(_17226_),
    .Y(_17227_),
    .B(_15661_));
 XOR2x1_ASAP7_75t_R _25659_ (.A(_17225_),
    .Y(_17228_),
    .B(_17227_));
 NOR2x1_ASAP7_75t_R _25660_ (.A(net4019),
    .B(_08823_),
    .Y(_17229_));
 AOI21x1_ASAP7_75t_R _25661_ (.A1(_08823_),
    .A2(_17228_),
    .B(net4020),
    .Y(_00328_));
 NOR2x2_ASAP7_75t_R _25662_ (.A(_15657_),
    .B(_15780_),
    .Y(_17230_));
 XOR2x2_ASAP7_75t_R _25663_ (.A(_00414_),
    .B(_00491_),
    .Y(_17231_));
 XOR2x1_ASAP7_75t_R _25664_ (.A(_17231_),
    .Y(_17232_),
    .B(_15784_));
 XOR2x1_ASAP7_75t_R _25665_ (.A(_17230_),
    .Y(_17233_),
    .B(_17232_));
 NOR2x1_ASAP7_75t_R _25666_ (.A(net4038),
    .B(net400),
    .Y(_17234_));
 AOI21x1_ASAP7_75t_R _25667_ (.A1(net400),
    .A2(_17233_),
    .B(_17234_),
    .Y(_00329_));
 XOR2x1_ASAP7_75t_R _25668_ (.A(_15901_),
    .Y(_17235_),
    .B(_00393_));
 AND2x2_ASAP7_75t_R _25669_ (.A(_15900_),
    .B(_17235_),
    .Y(_17236_));
 NOR2x1_ASAP7_75t_R _25670_ (.A(_17235_),
    .B(_15900_),
    .Y(_17237_));
 OA21x2_ASAP7_75t_R _25671_ (.A1(_17236_),
    .A2(_17237_),
    .B(net398),
    .Y(_17238_));
 AO21x1_ASAP7_75t_R _25672_ (.A1(net402),
    .A2(net3651),
    .B(_17238_),
    .Y(_00330_));
 XOR2x1_ASAP7_75t_R _25673_ (.A(_15982_),
    .Y(_17239_),
    .B(_00394_));
 OAI21x1_ASAP7_75t_R _25674_ (.A1(_15946_),
    .A2(_15979_),
    .B(_17239_),
    .Y(_17240_));
 OR3x1_ASAP7_75t_R _25675_ (.A(_15979_),
    .B(_15946_),
    .C(_17239_),
    .Y(_17241_));
 AOI21x1_ASAP7_75t_R _25676_ (.A1(_17240_),
    .A2(_17241_),
    .B(net405),
    .Y(_17242_));
 AO21x1_ASAP7_75t_R _25677_ (.A1(net405),
    .A2(net3940),
    .B(_17242_),
    .Y(_00331_));
 INVx2_ASAP7_75t_R _25678_ (.A(net4060),
    .Y(_17243_));
 INVx2_ASAP7_75t_R _25679_ (.A(_00395_),
    .Y(_17244_));
 XOR2x1_ASAP7_75t_R _25680_ (.A(_16050_),
    .Y(_17245_),
    .B(_17244_));
 INVx1_ASAP7_75t_R _25681_ (.A(_17245_),
    .Y(_17246_));
 AOI21x1_ASAP7_75t_R _25682_ (.A1(_16013_),
    .A2(_16048_),
    .B(_17246_),
    .Y(_17247_));
 NOR2x1_ASAP7_75t_R _25683_ (.A(_17245_),
    .B(_16049_),
    .Y(_17248_));
 OAI21x1_ASAP7_75t_R _25684_ (.A1(_17247_),
    .A2(_17248_),
    .B(net398),
    .Y(_17249_));
 OAI21x1_ASAP7_75t_R _25685_ (.A1(net398),
    .A2(_17243_),
    .B(_17249_),
    .Y(_00333_));
 XOR2x2_ASAP7_75t_R _25686_ (.A(_00415_),
    .B(_00490_),
    .Y(_17250_));
 XOR2x1_ASAP7_75t_R _25687_ (.A(_17250_),
    .Y(_17251_),
    .B(_16060_));
 XNOR2x1_ASAP7_75t_R _25688_ (.B(_16123_),
    .Y(_17252_),
    .A(_17251_));
 AND2x2_ASAP7_75t_R _25689_ (.A(net402),
    .B(net4082),
    .Y(_17253_));
 AO21x1_ASAP7_75t_R _25690_ (.A1(_17252_),
    .A2(net398),
    .B(_17253_),
    .Y(_00334_));
 XOR2x2_ASAP7_75t_R _25691_ (.A(_00416_),
    .B(_00489_),
    .Y(_17254_));
 XOR2x1_ASAP7_75t_R _25692_ (.A(_17254_),
    .Y(_17255_),
    .B(_16130_));
 XOR2x1_ASAP7_75t_R _25693_ (.A(_16193_),
    .Y(_17256_),
    .B(_17255_));
 AND2x2_ASAP7_75t_R _25694_ (.A(net402),
    .B(net78),
    .Y(_17257_));
 AO21x1_ASAP7_75t_R _25695_ (.A1(_17256_),
    .A2(net398),
    .B(_17257_),
    .Y(_00335_));
 XOR2x1_ASAP7_75t_R _25696_ (.A(_16254_),
    .Y(_17258_),
    .B(_00396_));
 XOR2x1_ASAP7_75t_R _25697_ (.A(_16251_),
    .Y(_17259_),
    .B(_17258_));
 BUFx2_ASAP7_75t_R output265 (.A(net265),
    .Y(text_out[104]));
 BUFx2_ASAP7_75t_R output264 (.A(net264),
    .Y(text_out[103]));
 AND2x2_ASAP7_75t_R _25700_ (.A(net402),
    .B(net4112),
    .Y(_17262_));
 AO21x1_ASAP7_75t_R _25701_ (.A1(_17259_),
    .A2(net398),
    .B(_17262_),
    .Y(_00336_));
 XOR2x1_ASAP7_75t_R _25702_ (.A(_00398_),
    .Y(_17263_),
    .B(_00397_));
 XNOR2x1_ASAP7_75t_R _25703_ (.B(_16258_),
    .Y(_17264_),
    .A(_17263_));
 XOR2x2_ASAP7_75t_R _25704_ (.A(_16525_),
    .B(_17264_),
    .Y(_17265_));
 NOR2x1_ASAP7_75t_R _25705_ (.A(net4046),
    .B(net400),
    .Y(_17266_));
 AOI21x1_ASAP7_75t_R _25706_ (.A1(net400),
    .A2(_17265_),
    .B(_17266_),
    .Y(_00337_));
 XOR2x1_ASAP7_75t_R _25707_ (.A(_00400_),
    .Y(_17267_),
    .B(_00399_));
 XNOR2x1_ASAP7_75t_R _25708_ (.B(_16640_),
    .Y(_17268_),
    .A(_17267_));
 NAND3x1_ASAP7_75t_R _25709_ (.A(_16638_),
    .B(_16524_),
    .C(_17268_),
    .Y(_17269_));
 AO21x1_ASAP7_75t_R _25710_ (.A1(_16638_),
    .A2(_16524_),
    .B(_17268_),
    .Y(_17270_));
 NAND2x1_ASAP7_75t_R _25711_ (.A(_17269_),
    .B(_17270_),
    .Y(_17271_));
 NOR2x1_ASAP7_75t_R _25712_ (.A(net4072),
    .B(net399),
    .Y(_17272_));
 AOI21x1_ASAP7_75t_R _25713_ (.A1(net399),
    .A2(_17271_),
    .B(_17272_),
    .Y(_00338_));
 INVx2_ASAP7_75t_R _25714_ (.A(net3861),
    .Y(_17273_));
 XOR2x1_ASAP7_75t_R _25715_ (.A(_00458_),
    .Y(_17274_),
    .B(_00506_));
 INVx4_ASAP7_75t_R _25716_ (.A(_00488_),
    .Y(_17275_));
 XOR2x1_ASAP7_75t_R _25717_ (.A(_17274_),
    .Y(_17276_),
    .B(_17275_));
 NAND2x1_ASAP7_75t_R _25718_ (.A(_17276_),
    .B(_16747_),
    .Y(_17277_));
 OR3x1_ASAP7_75t_R _25719_ (.A(_16745_),
    .B(_16701_),
    .C(_17276_),
    .Y(_17278_));
 AOI21x1_ASAP7_75t_R _25720_ (.A1(_17277_),
    .A2(_17278_),
    .B(_00401_),
    .Y(_17279_));
 AND3x1_ASAP7_75t_R _25721_ (.A(_17278_),
    .B(_17277_),
    .C(_00401_),
    .Y(_17280_));
 OAI21x1_ASAP7_75t_R _25722_ (.A1(_17279_),
    .A2(_17280_),
    .B(net400),
    .Y(_17281_));
 OAI21x1_ASAP7_75t_R _25723_ (.A1(net400),
    .A2(net3862),
    .B(_17281_),
    .Y(_00339_));
 NAND2x2_ASAP7_75t_R _25724_ (.A(net402),
    .B(net4090),
    .Y(_17282_));
 XOR2x1_ASAP7_75t_R _25725_ (.A(_00457_),
    .Y(_17283_),
    .B(_00505_));
 INVx3_ASAP7_75t_R _25726_ (.A(_00487_),
    .Y(_17284_));
 XOR2x2_ASAP7_75t_R _25727_ (.A(_17283_),
    .B(_17284_),
    .Y(_17285_));
 OA21x2_ASAP7_75t_R _25728_ (.A1(_16846_),
    .A2(_16805_),
    .B(_17285_),
    .Y(_17286_));
 NOR3x2_ASAP7_75t_R _25729_ (.B(_16805_),
    .C(_17285_),
    .Y(_17287_),
    .A(_16846_));
 OA21x2_ASAP7_75t_R _25730_ (.A1(_17286_),
    .A2(_17287_),
    .B(_16757_),
    .Y(_17288_));
 NOR3x1_ASAP7_75t_R _25731_ (.A(_17286_),
    .B(_17287_),
    .C(_16757_),
    .Y(_17289_));
 OAI21x1_ASAP7_75t_R _25732_ (.A1(_17288_),
    .A2(_17289_),
    .B(net398),
    .Y(_17290_));
 NAND2x1_ASAP7_75t_R _25733_ (.A(_17282_),
    .B(_17290_),
    .Y(_00340_));
 NAND2x2_ASAP7_75t_R _25734_ (.A(net402),
    .B(net4088),
    .Y(_17291_));
 XOR2x1_ASAP7_75t_R _25735_ (.A(_00456_),
    .Y(_17292_),
    .B(_00504_));
 INVx2_ASAP7_75t_R _25736_ (.A(_00486_),
    .Y(_17293_));
 XOR2x1_ASAP7_75t_R _25737_ (.A(_17292_),
    .Y(_17294_),
    .B(_17293_));
 NAND2x1_ASAP7_75t_R _25738_ (.A(_17294_),
    .B(_16924_),
    .Y(_17295_));
 OR3x1_ASAP7_75t_R _25739_ (.A(_16922_),
    .B(_16885_),
    .C(_17294_),
    .Y(_17296_));
 AOI21x1_ASAP7_75t_R _25740_ (.A1(_17295_),
    .A2(_17296_),
    .B(_00403_),
    .Y(_17297_));
 INVx1_ASAP7_75t_R _25741_ (.A(_00403_),
    .Y(_17298_));
 NAND2x1_ASAP7_75t_R _25742_ (.A(_17295_),
    .B(_17296_),
    .Y(_17299_));
 NOR2x1_ASAP7_75t_R _25743_ (.A(_17298_),
    .B(_17299_),
    .Y(_17300_));
 OAI21x1_ASAP7_75t_R _25744_ (.A1(_17297_),
    .A2(_17300_),
    .B(net398),
    .Y(_17301_));
 NAND2x1_ASAP7_75t_R _25745_ (.A(_17291_),
    .B(_17301_),
    .Y(_00341_));
 XOR2x2_ASAP7_75t_R _25746_ (.A(_00405_),
    .B(_00404_),
    .Y(_17302_));
 XNOR2x1_ASAP7_75t_R _25747_ (.B(_16987_),
    .Y(_17303_),
    .A(_17302_));
 XOR2x1_ASAP7_75t_R _25748_ (.A(_16986_),
    .Y(_17304_),
    .B(_17303_));
 BUFx2_ASAP7_75t_R output263 (.A(net263),
    .Y(text_out[102]));
 NOR2x1_ASAP7_75t_R _25750_ (.A(net4150),
    .B(net399),
    .Y(_17306_));
 AOI21x1_ASAP7_75t_R _25751_ (.A1(net399),
    .A2(_17304_),
    .B(_17306_),
    .Y(_00342_));
 XOR2x1_ASAP7_75t_R _25752_ (.A(_17056_),
    .Y(_17307_),
    .B(_17053_));
 XNOR2x1_ASAP7_75t_R _25753_ (.B(_17052_),
    .Y(_17308_),
    .A(_17307_));
 NOR2x1_ASAP7_75t_R _25754_ (.A(net87),
    .B(net400),
    .Y(_17309_));
 AOI21x1_ASAP7_75t_R _25755_ (.A1(net400),
    .A2(_17308_),
    .B(_17309_),
    .Y(_00344_));
 NAND2x2_ASAP7_75t_R _25756_ (.A(net405),
    .B(net4124),
    .Y(_17310_));
 XOR2x1_ASAP7_75t_R _25757_ (.A(_00453_),
    .Y(_17311_),
    .B(_00501_));
 INVx3_ASAP7_75t_R _25758_ (.A(_00485_),
    .Y(_17312_));
 XOR2x1_ASAP7_75t_R _25759_ (.A(_17311_),
    .Y(_17313_),
    .B(_17312_));
 NOR2x1_ASAP7_75t_R _25760_ (.A(_17313_),
    .B(_17124_),
    .Y(_17314_));
 INVx2_ASAP7_75t_R _25761_ (.A(_00408_),
    .Y(_17315_));
 INVx1_ASAP7_75t_R _25762_ (.A(_17096_),
    .Y(_17316_));
 OA21x2_ASAP7_75t_R _25763_ (.A1(_17122_),
    .A2(_17316_),
    .B(_17313_),
    .Y(_17317_));
 NOR3x1_ASAP7_75t_R _25764_ (.A(_17314_),
    .B(_17315_),
    .C(_17317_),
    .Y(_17318_));
 OA21x2_ASAP7_75t_R _25765_ (.A1(_17314_),
    .A2(_17317_),
    .B(_17315_),
    .Y(_17319_));
 OAI21x1_ASAP7_75t_R _25766_ (.A1(_17318_),
    .A2(_17319_),
    .B(net399),
    .Y(_17320_));
 NAND2x1_ASAP7_75t_R _25767_ (.A(_17310_),
    .B(_17320_),
    .Y(_00345_));
 XNOR2x1_ASAP7_75t_R _25768_ (.B(_17127_),
    .Y(_17321_),
    .A(_17128_));
 NOR2x1_ASAP7_75t_R _25769_ (.A(net4096),
    .B(net400),
    .Y(_17322_));
 AOI21x1_ASAP7_75t_R _25770_ (.A1(net400),
    .A2(_17321_),
    .B(_17322_),
    .Y(_00289_));
 XOR2x1_ASAP7_75t_R _25771_ (.A(_17133_),
    .Y(_17323_),
    .B(_17134_));
 NOR2x1_ASAP7_75t_R _25772_ (.A(net4078),
    .B(net400),
    .Y(_17324_));
 AOI21x1_ASAP7_75t_R _25773_ (.A1(net400),
    .A2(_17323_),
    .B(_17324_),
    .Y(_00300_));
 XNOR2x1_ASAP7_75t_R _25774_ (.B(_00524_),
    .Y(_17325_),
    .A(_00385_));
 XNOR2x1_ASAP7_75t_R _25775_ (.B(_11214_),
    .Y(_17326_),
    .A(_17325_));
 AND2x2_ASAP7_75t_R _25776_ (.A(net403),
    .B(net4132),
    .Y(_17327_));
 AO21x1_ASAP7_75t_R _25777_ (.A1(_17326_),
    .A2(net400),
    .B(_17327_),
    .Y(_00311_));
 XNOR2x1_ASAP7_75t_R _25778_ (.B(_00523_),
    .Y(_17328_),
    .A(_00386_));
 XOR2x1_ASAP7_75t_R _25779_ (.A(_12212_),
    .Y(_17329_),
    .B(_17328_));
 AND2x2_ASAP7_75t_R _25780_ (.A(net404),
    .B(net4138),
    .Y(_17330_));
 AO21x1_ASAP7_75t_R _25781_ (.A1(_17329_),
    .A2(net399),
    .B(_17330_),
    .Y(_00314_));
 XOR2x1_ASAP7_75t_R _25782_ (.A(_00387_),
    .Y(_17331_),
    .B(_00522_));
 XNOR2x1_ASAP7_75t_R _25783_ (.B(_13001_),
    .Y(_17332_),
    .A(_17331_));
 AND2x2_ASAP7_75t_R _25784_ (.A(net403),
    .B(net93),
    .Y(_17333_));
 AO21x1_ASAP7_75t_R _25785_ (.A1(_17332_),
    .A2(net400),
    .B(_17333_),
    .Y(_00315_));
 XOR2x1_ASAP7_75t_R _25786_ (.A(_13790_),
    .Y(_17334_),
    .B(_13143_));
 AND2x2_ASAP7_75t_R _25787_ (.A(net403),
    .B(net94),
    .Y(_17335_));
 AO21x1_ASAP7_75t_R _25788_ (.A1(_17334_),
    .A2(net400),
    .B(_17335_),
    .Y(_00316_));
 XOR2x1_ASAP7_75t_R _25789_ (.A(_17165_),
    .Y(_17336_),
    .B(_17166_));
 AND2x2_ASAP7_75t_R _25790_ (.A(net404),
    .B(net96),
    .Y(_17337_));
 AO21x1_ASAP7_75t_R _25791_ (.A1(_17336_),
    .A2(net399),
    .B(_17337_),
    .Y(_00317_));
 XNOR2x1_ASAP7_75t_R _25792_ (.B(_00520_),
    .Y(_17338_),
    .A(_00388_));
 XOR2x1_ASAP7_75t_R _25793_ (.A(_14589_),
    .Y(_17339_),
    .B(_17338_));
 AND2x2_ASAP7_75t_R _25794_ (.A(net404),
    .B(net97),
    .Y(_17340_));
 AO21x1_ASAP7_75t_R _25795_ (.A1(_17339_),
    .A2(net399),
    .B(_17340_),
    .Y(_00318_));
 XOR2x1_ASAP7_75t_R _25796_ (.A(_14844_),
    .Y(_17341_),
    .B(_17178_));
 NAND2x1_ASAP7_75t_R _25797_ (.A(net399),
    .B(_17341_),
    .Y(_17342_));
 OA21x2_ASAP7_75t_R _25798_ (.A1(net399),
    .A2(net4098),
    .B(_17342_),
    .Y(_00319_));
 XOR2x1_ASAP7_75t_R _25799_ (.A(_14959_),
    .Y(_17343_),
    .B(_14963_));
 AND2x2_ASAP7_75t_R _25800_ (.A(net404),
    .B(net99),
    .Y(_17344_));
 AO21x1_ASAP7_75t_R _25801_ (.A1(_17343_),
    .A2(net399),
    .B(_17344_),
    .Y(_00320_));
 XOR2x1_ASAP7_75t_R _25802_ (.A(_15053_),
    .Y(_17345_),
    .B(_00518_));
 XOR2x1_ASAP7_75t_R _25803_ (.A(_17345_),
    .Y(_17346_),
    .B(_00389_));
 NOR2x1_ASAP7_75t_R _25804_ (.A(net4008),
    .B(net399),
    .Y(_17347_));
 AOI21x1_ASAP7_75t_R _25805_ (.A1(net399),
    .A2(_17346_),
    .B(net4009),
    .Y(_00290_));
 XOR2x1_ASAP7_75t_R _25806_ (.A(_00390_),
    .Y(_17348_),
    .B(_00517_));
 XNOR2x1_ASAP7_75t_R _25807_ (.B(_15137_),
    .Y(_17349_),
    .A(_17348_));
 AND2x2_ASAP7_75t_R _25808_ (.A(net404),
    .B(net4106),
    .Y(_17350_));
 AO21x1_ASAP7_75t_R _25809_ (.A1(_17349_),
    .A2(net399),
    .B(_17350_),
    .Y(_00291_));
 XNOR2x1_ASAP7_75t_R _25810_ (.B(_00516_),
    .Y(_17351_),
    .A(_00391_));
 XNOR2x1_ASAP7_75t_R _25811_ (.B(_15203_),
    .Y(_17352_),
    .A(_17351_));
 AND2x2_ASAP7_75t_R _25812_ (.A(net405),
    .B(net4126),
    .Y(_17353_));
 AO21x1_ASAP7_75t_R _25813_ (.A1(_17352_),
    .A2(net399),
    .B(_17353_),
    .Y(_00292_));
 BUFx2_ASAP7_75t_R output262 (.A(net262),
    .Y(text_out[101]));
 XOR2x1_ASAP7_75t_R _25815_ (.A(_15268_),
    .Y(_17355_),
    .B(_15272_));
 NOR2x1_ASAP7_75t_R _25816_ (.A(net4068),
    .B(net398),
    .Y(_17356_));
 AOI21x1_ASAP7_75t_R _25817_ (.A1(net398),
    .A2(_17355_),
    .B(_17356_),
    .Y(_00293_));
 XNOR2x1_ASAP7_75t_R _25818_ (.B(_15334_),
    .Y(_17357_),
    .A(_15278_));
 BUFx2_ASAP7_75t_R output261 (.A(net261),
    .Y(text_out[100]));
 BUFx2_ASAP7_75t_R output260 (.A(net260),
    .Y(text_out[0]));
 AND2x2_ASAP7_75t_R _25821_ (.A(net402),
    .B(net4168),
    .Y(_17360_));
 AO21x1_ASAP7_75t_R _25822_ (.A1(_17357_),
    .A2(net398),
    .B(_17360_),
    .Y(_00294_));
 XNOR2x1_ASAP7_75t_R _25823_ (.B(_00513_),
    .Y(_17361_),
    .A(_00392_));
 XNOR2x1_ASAP7_75t_R _25824_ (.B(_15391_),
    .Y(_17362_),
    .A(_17361_));
 AND2x2_ASAP7_75t_R _25825_ (.A(net402),
    .B(net4128),
    .Y(_17363_));
 AO21x1_ASAP7_75t_R _25826_ (.A1(_17362_),
    .A2(net398),
    .B(_17363_),
    .Y(_00295_));
 XOR2x1_ASAP7_75t_R _25827_ (.A(_17225_),
    .Y(_17364_),
    .B(_17226_));
 NOR2x1_ASAP7_75t_R _25828_ (.A(net4024),
    .B(_08823_),
    .Y(_17365_));
 AOI21x1_ASAP7_75t_R _25829_ (.A1(_08823_),
    .A2(_17364_),
    .B(net4025),
    .Y(_00296_));
 XOR2x1_ASAP7_75t_R _25830_ (.A(_17230_),
    .Y(_17366_),
    .B(_17231_));
 NOR2x1_ASAP7_75t_R _25831_ (.A(net4031),
    .B(_08823_),
    .Y(_17367_));
 AOI21x1_ASAP7_75t_R _25832_ (.A1(_08823_),
    .A2(_17366_),
    .B(net4032),
    .Y(_00297_));
 XOR2x2_ASAP7_75t_R _25833_ (.A(_15900_),
    .B(_00512_),
    .Y(_17368_));
 INVx2_ASAP7_75t_R _25834_ (.A(_00393_),
    .Y(_17369_));
 XOR2x1_ASAP7_75t_R _25835_ (.A(_17368_),
    .Y(_17370_),
    .B(_17369_));
 NOR2x1_ASAP7_75t_R _25836_ (.A(net3770),
    .B(net398),
    .Y(_17371_));
 AOI21x1_ASAP7_75t_R _25837_ (.A1(net398),
    .A2(_17370_),
    .B(net3771),
    .Y(_00298_));
 XOR2x1_ASAP7_75t_R _25838_ (.A(_00394_),
    .Y(_17372_),
    .B(_00511_));
 XNOR2x1_ASAP7_75t_R _25839_ (.B(_15980_),
    .Y(_17373_),
    .A(_17372_));
 AND2x2_ASAP7_75t_R _25840_ (.A(net402),
    .B(net4070),
    .Y(_17374_));
 AO21x1_ASAP7_75t_R _25841_ (.A1(_17373_),
    .A2(net398),
    .B(_17374_),
    .Y(_00299_));
 XNOR2x1_ASAP7_75t_R _25842_ (.B(_00510_),
    .Y(_17375_),
    .A(_00395_));
 XOR2x1_ASAP7_75t_R _25843_ (.A(_16049_),
    .Y(_17376_),
    .B(_17375_));
 NOR2x2_ASAP7_75t_R _25844_ (.A(net4040),
    .B(net398),
    .Y(_17377_));
 AOI21x1_ASAP7_75t_R _25845_ (.A1(net398),
    .A2(_17376_),
    .B(_17377_),
    .Y(_00301_));
 XNOR2x1_ASAP7_75t_R _25846_ (.B(_16123_),
    .Y(_17378_),
    .A(_17250_));
 AND2x2_ASAP7_75t_R _25847_ (.A(net402),
    .B(net4148),
    .Y(_17379_));
 AO21x1_ASAP7_75t_R _25848_ (.A1(_17378_),
    .A2(net398),
    .B(_17379_),
    .Y(_00302_));
 XOR2x1_ASAP7_75t_R _25849_ (.A(_16193_),
    .Y(_17380_),
    .B(_17254_));
 AND2x2_ASAP7_75t_R _25850_ (.A(net402),
    .B(net4178),
    .Y(_17381_));
 AO21x1_ASAP7_75t_R _25851_ (.A1(_17380_),
    .A2(net398),
    .B(_17381_),
    .Y(_00303_));
 XNOR2x1_ASAP7_75t_R _25852_ (.B(_00509_),
    .Y(_17382_),
    .A(_00396_));
 XNOR2x1_ASAP7_75t_R _25853_ (.B(_16251_),
    .Y(_17383_),
    .A(_17382_));
 AND2x2_ASAP7_75t_R _25854_ (.A(net402),
    .B(net4114),
    .Y(_17384_));
 AO21x1_ASAP7_75t_R _25855_ (.A1(_17383_),
    .A2(net398),
    .B(_17384_),
    .Y(_00304_));
 XOR2x2_ASAP7_75t_R _25856_ (.A(_00397_),
    .B(_00508_),
    .Y(_17385_));
 INVx3_ASAP7_75t_R _25857_ (.A(_00398_),
    .Y(_17386_));
 XOR2x1_ASAP7_75t_R _25858_ (.A(_17385_),
    .Y(_17387_),
    .B(_17386_));
 XNOR2x1_ASAP7_75t_R _25859_ (.B(_16525_),
    .Y(_17388_),
    .A(_17387_));
 BUFx2_ASAP7_75t_R output259 (.A(net259),
    .Y(done));
 NOR2x1_ASAP7_75t_R _25861_ (.A(net4134),
    .B(net399),
    .Y(_17390_));
 AOI21x1_ASAP7_75t_R _25862_ (.A1(net399),
    .A2(_17388_),
    .B(_17390_),
    .Y(_00305_));
 XOR2x1_ASAP7_75t_R _25863_ (.A(_00399_),
    .Y(_17391_),
    .B(_00507_));
 XOR2x1_ASAP7_75t_R _25864_ (.A(_17391_),
    .Y(_17392_),
    .B(_00400_));
 NAND3x1_ASAP7_75t_R _25865_ (.A(_16638_),
    .B(_16524_),
    .C(_17392_),
    .Y(_17393_));
 AO21x1_ASAP7_75t_R _25866_ (.A1(_16638_),
    .A2(_16524_),
    .B(_17392_),
    .Y(_17394_));
 NAND2x1_ASAP7_75t_R _25867_ (.A(_17393_),
    .B(_17394_),
    .Y(_17395_));
 NOR2x1_ASAP7_75t_R _25868_ (.A(net4054),
    .B(net399),
    .Y(_17396_));
 AOI21x1_ASAP7_75t_R _25869_ (.A1(net399),
    .A2(_17395_),
    .B(_17396_),
    .Y(_00306_));
 INVx2_ASAP7_75t_R _25870_ (.A(net3855),
    .Y(_17397_));
 XNOR2x2_ASAP7_75t_R _25871_ (.A(_00401_),
    .B(_00506_),
    .Y(_17398_));
 AND2x2_ASAP7_75t_R _25872_ (.A(_16747_),
    .B(_17398_),
    .Y(_17399_));
 NOR2x2_ASAP7_75t_R _25873_ (.A(_17398_),
    .B(_16747_),
    .Y(_17400_));
 NOR3x1_ASAP7_75t_R _25874_ (.A(_17399_),
    .B(_00488_),
    .C(_17400_),
    .Y(_17401_));
 OA21x2_ASAP7_75t_R _25875_ (.A1(_17399_),
    .A2(_17400_),
    .B(_00488_),
    .Y(_17402_));
 OAI21x1_ASAP7_75t_R _25876_ (.A1(_17401_),
    .A2(_17402_),
    .B(net400),
    .Y(_17403_));
 OAI21x1_ASAP7_75t_R _25877_ (.A1(net400),
    .A2(net3856),
    .B(_17403_),
    .Y(_00307_));
 NAND2x2_ASAP7_75t_R _25878_ (.A(net402),
    .B(net4080),
    .Y(_17404_));
 INVx1_ASAP7_75t_R _25879_ (.A(_16805_),
    .Y(_17405_));
 AND4x1_ASAP7_75t_R _25880_ (.A(_16845_),
    .B(_17405_),
    .C(_16825_),
    .D(_16754_),
    .Y(_17406_));
 INVx1_ASAP7_75t_R _25881_ (.A(_16754_),
    .Y(_17407_));
 OA21x2_ASAP7_75t_R _25882_ (.A1(_16846_),
    .A2(_16805_),
    .B(_17407_),
    .Y(_17408_));
 NOR3x1_ASAP7_75t_R _25883_ (.A(_17406_),
    .B(_17408_),
    .C(_16757_),
    .Y(_17409_));
 OA21x2_ASAP7_75t_R _25884_ (.A1(_17406_),
    .A2(_17408_),
    .B(_16757_),
    .Y(_17410_));
 OAI21x1_ASAP7_75t_R _25885_ (.A1(_17409_),
    .A2(_17410_),
    .B(net398),
    .Y(_17411_));
 NAND2x1_ASAP7_75t_R _25886_ (.A(_17404_),
    .B(_17411_),
    .Y(_00308_));
 NAND2x2_ASAP7_75t_R _25887_ (.A(net402),
    .B(net4086),
    .Y(_17412_));
 AO21x1_ASAP7_75t_R _25888_ (.A1(_16923_),
    .A2(_16886_),
    .B(_16851_),
    .Y(_17413_));
 INVx1_ASAP7_75t_R _25889_ (.A(_16851_),
    .Y(_17414_));
 OR3x1_ASAP7_75t_R _25890_ (.A(_16922_),
    .B(_16885_),
    .C(_17414_),
    .Y(_17415_));
 AOI21x1_ASAP7_75t_R _25891_ (.A1(_17413_),
    .A2(_17415_),
    .B(_00403_),
    .Y(_17416_));
 NAND2x1_ASAP7_75t_R _25892_ (.A(_17413_),
    .B(_17415_),
    .Y(_17417_));
 NOR2x1_ASAP7_75t_R _25893_ (.A(_17298_),
    .B(_17417_),
    .Y(_17418_));
 OAI21x1_ASAP7_75t_R _25894_ (.A1(_17416_),
    .A2(_17418_),
    .B(net398),
    .Y(_17419_));
 NAND2x1_ASAP7_75t_R _25895_ (.A(_17412_),
    .B(_17419_),
    .Y(_00309_));
 XOR2x1_ASAP7_75t_R _25896_ (.A(_17302_),
    .Y(_17420_),
    .B(_00503_));
 XOR2x1_ASAP7_75t_R _25897_ (.A(_16986_),
    .Y(_17421_),
    .B(_17420_));
 NOR2x1_ASAP7_75t_R _25898_ (.A(net4162),
    .B(net399),
    .Y(_17422_));
 AOI21x1_ASAP7_75t_R _25899_ (.A1(net399),
    .A2(_17421_),
    .B(_17422_),
    .Y(_00310_));
 XOR2x1_ASAP7_75t_R _25900_ (.A(_17053_),
    .Y(_17423_),
    .B(_00502_));
 XOR2x1_ASAP7_75t_R _25901_ (.A(_17052_),
    .Y(_17424_),
    .B(_17423_));
 NOR2x1_ASAP7_75t_R _25902_ (.A(net122),
    .B(net400),
    .Y(_17425_));
 AOI21x1_ASAP7_75t_R _25903_ (.A1(net400),
    .A2(_17424_),
    .B(_17425_),
    .Y(_00312_));
 NAND2x2_ASAP7_75t_R _25904_ (.A(net402),
    .B(net4034),
    .Y(_17426_));
 INVx1_ASAP7_75t_R _25905_ (.A(_17062_),
    .Y(_17427_));
 NOR2x1_ASAP7_75t_R _25906_ (.A(_17427_),
    .B(_17124_),
    .Y(_17428_));
 OA21x2_ASAP7_75t_R _25907_ (.A1(_17122_),
    .A2(_17316_),
    .B(_17427_),
    .Y(_17429_));
 NOR3x1_ASAP7_75t_R _25908_ (.A(_17428_),
    .B(_17315_),
    .C(_17429_),
    .Y(_17430_));
 OA21x2_ASAP7_75t_R _25909_ (.A1(_17428_),
    .A2(_17429_),
    .B(_17315_),
    .Y(_17431_));
 OAI21x1_ASAP7_75t_R _25910_ (.A1(_17430_),
    .A2(_17431_),
    .B(net399),
    .Y(_17432_));
 NAND2x1_ASAP7_75t_R _25911_ (.A(_17426_),
    .B(_17432_),
    .Y(_00313_));
 XOR2x1_ASAP7_75t_R _25912_ (.A(_17127_),
    .Y(_17433_),
    .B(_00409_));
 NAND2x2_ASAP7_75t_R _25913_ (.A(net403),
    .B(net4014),
    .Y(_17434_));
 OAI21x1_ASAP7_75t_R _25914_ (.A1(net404),
    .A2(_17433_),
    .B(net4015),
    .Y(_00257_));
 INVx1_ASAP7_75t_R _25915_ (.A(_00410_),
    .Y(_17435_));
 XOR2x1_ASAP7_75t_R _25916_ (.A(_17133_),
    .Y(_17436_),
    .B(_17435_));
 NAND2x2_ASAP7_75t_R _25917_ (.A(net403),
    .B(net4011),
    .Y(_17437_));
 OAI21x1_ASAP7_75t_R _25918_ (.A1(net404),
    .A2(_17436_),
    .B(net4012),
    .Y(_00268_));
 INVx1_ASAP7_75t_R _25919_ (.A(_00524_),
    .Y(_17438_));
 XOR2x1_ASAP7_75t_R _25920_ (.A(_11214_),
    .Y(_17439_),
    .B(_17438_));
 AND2x2_ASAP7_75t_R _25921_ (.A(net403),
    .B(net4136),
    .Y(_17440_));
 AO21x1_ASAP7_75t_R _25922_ (.A1(_17439_),
    .A2(net400),
    .B(_17440_),
    .Y(_00279_));
 XOR2x1_ASAP7_75t_R _25923_ (.A(_12212_),
    .Y(_17441_),
    .B(_00523_));
 AND2x2_ASAP7_75t_R _25924_ (.A(net403),
    .B(net127),
    .Y(_17442_));
 AO21x1_ASAP7_75t_R _25925_ (.A1(_17441_),
    .A2(net400),
    .B(_17442_),
    .Y(_00282_));
 XOR2x1_ASAP7_75t_R _25926_ (.A(_13001_),
    .Y(_17443_),
    .B(_00522_));
 AND2x2_ASAP7_75t_R _25927_ (.A(net403),
    .B(net2),
    .Y(_17444_));
 AO21x1_ASAP7_75t_R _25928_ (.A1(_17443_),
    .A2(net400),
    .B(_17444_),
    .Y(_00283_));
 INVx1_ASAP7_75t_R _25929_ (.A(net4076),
    .Y(_17445_));
 INVx2_ASAP7_75t_R _25930_ (.A(_00521_),
    .Y(_17446_));
 NOR2x1_ASAP7_75t_R _25931_ (.A(_17446_),
    .B(_13790_),
    .Y(_17447_));
 AND4x1_ASAP7_75t_R _25932_ (.A(_06375_),
    .B(_13768_),
    .C(_17446_),
    .D(_13461_),
    .Y(_17448_));
 OAI21x1_ASAP7_75t_R _25933_ (.A1(_17447_),
    .A2(_17448_),
    .B(net400),
    .Y(_17449_));
 OAI21x1_ASAP7_75t_R _25934_ (.A1(net400),
    .A2(_17445_),
    .B(_17449_),
    .Y(_00284_));
 INVx1_ASAP7_75t_R _25935_ (.A(_00411_),
    .Y(_17450_));
 XOR2x1_ASAP7_75t_R _25936_ (.A(_17165_),
    .Y(_17451_),
    .B(_17450_));
 AND2x2_ASAP7_75t_R _25937_ (.A(net403),
    .B(net4),
    .Y(_17452_));
 AO21x1_ASAP7_75t_R _25938_ (.A1(_17451_),
    .A2(net400),
    .B(_17452_),
    .Y(_00285_));
 XOR2x1_ASAP7_75t_R _25939_ (.A(_14589_),
    .Y(_17453_),
    .B(_00520_));
 BUFx2_ASAP7_75t_R input258 (.A(net3573),
    .Y(net258));
 BUFx2_ASAP7_75t_R input257 (.A(net3918),
    .Y(net257));
 AND2x2_ASAP7_75t_R _25942_ (.A(net404),
    .B(net5),
    .Y(_17456_));
 AO21x1_ASAP7_75t_R _25943_ (.A1(_17453_),
    .A2(net399),
    .B(_17456_),
    .Y(_00286_));
 XOR2x2_ASAP7_75t_R _25944_ (.A(_14844_),
    .B(_00412_),
    .Y(_17457_));
 AND2x2_ASAP7_75t_R _25945_ (.A(net403),
    .B(net6),
    .Y(_17458_));
 AO21x1_ASAP7_75t_R _25946_ (.A1(_17457_),
    .A2(net400),
    .B(_17458_),
    .Y(_00287_));
 XOR2x2_ASAP7_75t_R _25947_ (.A(_14959_),
    .B(_00519_),
    .Y(_17459_));
 AND2x2_ASAP7_75t_R _25948_ (.A(net403),
    .B(net4172),
    .Y(_17460_));
 AO21x1_ASAP7_75t_R _25949_ (.A1(_17459_),
    .A2(net400),
    .B(_17460_),
    .Y(_00288_));
 AND2x2_ASAP7_75t_R _25950_ (.A(net402),
    .B(net8),
    .Y(_17461_));
 AO21x1_ASAP7_75t_R _25951_ (.A1(_17345_),
    .A2(net399),
    .B(_17461_),
    .Y(_00258_));
 XOR2x1_ASAP7_75t_R _25952_ (.A(_15137_),
    .Y(_17462_),
    .B(_00517_));
 AND2x2_ASAP7_75t_R _25953_ (.A(net404),
    .B(net4108),
    .Y(_17463_));
 AO21x1_ASAP7_75t_R _25954_ (.A1(_17462_),
    .A2(net399),
    .B(_17463_),
    .Y(_00259_));
 INVx2_ASAP7_75t_R _25955_ (.A(_00516_),
    .Y(_17464_));
 XOR2x1_ASAP7_75t_R _25956_ (.A(_15203_),
    .Y(_17465_),
    .B(_17464_));
 AND2x2_ASAP7_75t_R _25957_ (.A(net403),
    .B(net4176),
    .Y(_17466_));
 AO21x1_ASAP7_75t_R _25958_ (.A1(_17465_),
    .A2(net400),
    .B(_17466_),
    .Y(_00260_));
 XOR2x1_ASAP7_75t_R _25959_ (.A(_15268_),
    .Y(_17467_),
    .B(_00515_));
 NAND2x1_ASAP7_75t_R _25960_ (.A(net405),
    .B(net4005),
    .Y(_17468_));
 OAI21x1_ASAP7_75t_R _25961_ (.A1(net405),
    .A2(_17467_),
    .B(net4006),
    .Y(_00261_));
 INVx5_ASAP7_75t_R _25962_ (.A(_00514_),
    .Y(_17469_));
 XOR2x1_ASAP7_75t_R _25963_ (.A(_15334_),
    .Y(_17470_),
    .B(_17469_));
 AND2x2_ASAP7_75t_R _25964_ (.A(net402),
    .B(net4158),
    .Y(_17471_));
 AO21x1_ASAP7_75t_R _25965_ (.A1(_17470_),
    .A2(net398),
    .B(_17471_),
    .Y(_00262_));
 INVx2_ASAP7_75t_R _25966_ (.A(_00513_),
    .Y(_17472_));
 XOR2x1_ASAP7_75t_R _25967_ (.A(_15391_),
    .Y(_17473_),
    .B(_17472_));
 AND2x2_ASAP7_75t_R _25968_ (.A(net403),
    .B(net4182),
    .Y(_17474_));
 AO21x1_ASAP7_75t_R _25969_ (.A1(_17473_),
    .A2(net400),
    .B(_17474_),
    .Y(_00263_));
 CKINVDCx5p33_ASAP7_75t_R _25970_ (.A(_00413_),
    .Y(_17475_));
 XOR2x1_ASAP7_75t_R _25971_ (.A(_17225_),
    .Y(_17476_),
    .B(_17475_));
 NAND2x2_ASAP7_75t_R _25972_ (.A(net401),
    .B(net3893),
    .Y(_17477_));
 OAI21x1_ASAP7_75t_R _25973_ (.A1(net401),
    .A2(_17476_),
    .B(net3894),
    .Y(_00264_));
 INVx5_ASAP7_75t_R _25974_ (.A(_00414_),
    .Y(_17478_));
 XOR2x1_ASAP7_75t_R _25975_ (.A(_17230_),
    .Y(_17479_),
    .B(_17478_));
 NAND2x2_ASAP7_75t_R _25976_ (.A(net401),
    .B(net3916),
    .Y(_17480_));
 OAI21x1_ASAP7_75t_R _25977_ (.A1(net401),
    .A2(_17479_),
    .B(net3917),
    .Y(_00265_));
 NOR2x1_ASAP7_75t_R _25978_ (.A(net402),
    .B(_17368_),
    .Y(_17481_));
 AO21x1_ASAP7_75t_R _25979_ (.A1(net402),
    .A2(net3592),
    .B(_17481_),
    .Y(_00266_));
 XOR2x1_ASAP7_75t_R _25980_ (.A(_15980_),
    .Y(_17482_),
    .B(_00511_));
 AND2x2_ASAP7_75t_R _25981_ (.A(net405),
    .B(net4062),
    .Y(_17483_));
 AO21x1_ASAP7_75t_R _25982_ (.A1(_17482_),
    .A2(net398),
    .B(_17483_),
    .Y(_00267_));
 CKINVDCx5p33_ASAP7_75t_R _25983_ (.A(_00510_),
    .Y(_17484_));
 XOR2x1_ASAP7_75t_R _25984_ (.A(_16049_),
    .Y(_17485_),
    .B(_17484_));
 AND2x2_ASAP7_75t_R _25985_ (.A(net402),
    .B(net4174),
    .Y(_17486_));
 AO21x1_ASAP7_75t_R _25986_ (.A1(_17485_),
    .A2(net398),
    .B(_17486_),
    .Y(_00269_));
 XOR2x1_ASAP7_75t_R _25987_ (.A(_16123_),
    .Y(_17487_),
    .B(_00415_));
 BUFx2_ASAP7_75t_R input256 (.A(net3948),
    .Y(net256));
 AND2x2_ASAP7_75t_R _25989_ (.A(net402),
    .B(net4140),
    .Y(_17489_));
 AO21x1_ASAP7_75t_R _25990_ (.A1(_17487_),
    .A2(net398),
    .B(_17489_),
    .Y(_00270_));
 INVx4_ASAP7_75t_R _25991_ (.A(_00416_),
    .Y(_17490_));
 XOR2x1_ASAP7_75t_R _25992_ (.A(_16193_),
    .Y(_17491_),
    .B(_17490_));
 AND2x2_ASAP7_75t_R _25993_ (.A(net402),
    .B(net21),
    .Y(_17492_));
 AO21x1_ASAP7_75t_R _25994_ (.A1(_17491_),
    .A2(net398),
    .B(_17492_),
    .Y(_00271_));
 INVx5_ASAP7_75t_R _25995_ (.A(_00509_),
    .Y(_17493_));
 XOR2x1_ASAP7_75t_R _25996_ (.A(_16251_),
    .Y(_17494_),
    .B(_17493_));
 AND2x2_ASAP7_75t_R _25997_ (.A(net402),
    .B(net4118),
    .Y(_17495_));
 AO21x1_ASAP7_75t_R _25998_ (.A1(_17494_),
    .A2(net398),
    .B(_17495_),
    .Y(_00272_));
 XNOR2x1_ASAP7_75t_R _25999_ (.B(_16525_),
    .Y(_17496_),
    .A(_17385_));
 NOR2x2_ASAP7_75t_R _26000_ (.A(net4180),
    .B(net400),
    .Y(_17497_));
 AOI21x1_ASAP7_75t_R _26001_ (.A1(net399),
    .A2(_17496_),
    .B(_17497_),
    .Y(_00273_));
 INVx1_ASAP7_75t_R _26002_ (.A(_17391_),
    .Y(_17498_));
 NAND3x1_ASAP7_75t_R _26003_ (.A(_16638_),
    .B(_16524_),
    .C(_17498_),
    .Y(_17499_));
 AO21x1_ASAP7_75t_R _26004_ (.A1(_16638_),
    .A2(_16524_),
    .B(_17498_),
    .Y(_17500_));
 NAND2x1_ASAP7_75t_R _26005_ (.A(_17499_),
    .B(_17500_),
    .Y(_17501_));
 NOR2x1_ASAP7_75t_R _26006_ (.A(net4048),
    .B(net399),
    .Y(_17502_));
 AOI21x1_ASAP7_75t_R _26007_ (.A1(net399),
    .A2(_17501_),
    .B(_17502_),
    .Y(_00274_));
 OA21x2_ASAP7_75t_R _26008_ (.A1(_17399_),
    .A2(_17400_),
    .B(net400),
    .Y(_17503_));
 AO21x1_ASAP7_75t_R _26009_ (.A1(net401),
    .A2(net3876),
    .B(_17503_),
    .Y(_00275_));
 BUFx2_ASAP7_75t_R input255 (.A(net3790),
    .Y(net255));
 XNOR2x1_ASAP7_75t_R _26011_ (.B(_00505_),
    .Y(_17505_),
    .A(_00402_));
 OR3x1_ASAP7_75t_R _26012_ (.A(_16846_),
    .B(_16805_),
    .C(_17505_),
    .Y(_17506_));
 NAND2x1_ASAP7_75t_R _26013_ (.A(_17505_),
    .B(_16847_),
    .Y(_17507_));
 AOI21x1_ASAP7_75t_R _26014_ (.A1(_17506_),
    .A2(_17507_),
    .B(net405),
    .Y(_17508_));
 AO21x1_ASAP7_75t_R _26015_ (.A1(net405),
    .A2(net3991),
    .B(_17508_),
    .Y(_00276_));
 XNOR2x1_ASAP7_75t_R _26016_ (.B(_00504_),
    .Y(_17509_),
    .A(_00403_));
 AND2x2_ASAP7_75t_R _26017_ (.A(_16924_),
    .B(_17509_),
    .Y(_17510_));
 NOR2x1_ASAP7_75t_R _26018_ (.A(_17509_),
    .B(_16924_),
    .Y(_17511_));
 OA21x2_ASAP7_75t_R _26019_ (.A1(_17510_),
    .A2(_17511_),
    .B(net398),
    .Y(_17512_));
 AO21x1_ASAP7_75t_R _26020_ (.A1(net405),
    .A2(net3908),
    .B(_17512_),
    .Y(_00277_));
 XNOR2x1_ASAP7_75t_R _26021_ (.B(_00503_),
    .Y(_17513_),
    .A(_00404_));
 XOR2x1_ASAP7_75t_R _26022_ (.A(_16986_),
    .Y(_17514_),
    .B(_17513_));
 NOR2x1_ASAP7_75t_R _26023_ (.A(net4166),
    .B(net399),
    .Y(_17515_));
 AOI21x1_ASAP7_75t_R _26024_ (.A1(net399),
    .A2(_17514_),
    .B(_17515_),
    .Y(_00278_));
 XOR2x1_ASAP7_75t_R _26025_ (.A(_00406_),
    .Y(_17516_),
    .B(_00502_));
 XNOR2x1_ASAP7_75t_R _26026_ (.B(_17052_),
    .Y(_17517_),
    .A(_17516_));
 NOR2x1_ASAP7_75t_R _26027_ (.A(net4146),
    .B(net400),
    .Y(_17518_));
 AOI21x1_ASAP7_75t_R _26028_ (.A1(net400),
    .A2(_17517_),
    .B(_17518_),
    .Y(_00280_));
 XNOR2x1_ASAP7_75t_R _26029_ (.B(_00501_),
    .Y(_17519_),
    .A(_00408_));
 AND2x2_ASAP7_75t_R _26030_ (.A(_17124_),
    .B(_17519_),
    .Y(_17520_));
 NOR2x1_ASAP7_75t_R _26031_ (.A(_17519_),
    .B(_17124_),
    .Y(_17521_));
 OA21x2_ASAP7_75t_R _26032_ (.A1(_17520_),
    .A2(_17521_),
    .B(net399),
    .Y(_17522_));
 AO21x1_ASAP7_75t_R _26033_ (.A1(net401),
    .A2(net4022),
    .B(_17522_),
    .Y(_00281_));
 AND2x2_ASAP7_75t_R _26034_ (.A(_22106_),
    .B(_00785_),
    .Y(_17523_));
 INVx1_ASAP7_75t_R _26035_ (.A(_00787_),
    .Y(_17524_));
 AND4x1_ASAP7_75t_R _26036_ (.A(_17523_),
    .B(net398),
    .C(_00786_),
    .D(_17524_),
    .Y(_00000_));
 BUFx2_ASAP7_75t_R input254 (.A(net3817),
    .Y(net254));
 BUFx2_ASAP7_75t_R input253 (.A(net3602),
    .Y(net253));
 NOR2x1_ASAP7_75t_R _26039_ (.A(net397),
    .B(_00915_),
    .Y(_17527_));
 INVx1_ASAP7_75t_R _26040_ (.A(_17527_),
    .Y(_17528_));
 INVx3_ASAP7_75t_R _26041_ (.A(_00557_),
    .Y(_17529_));
 NAND2x2_ASAP7_75t_R _26042_ (.A(net2910),
    .B(net3311),
    .Y(_17530_));
 BUFx2_ASAP7_75t_R input252 (.A(net3857),
    .Y(net252));
 BUFx2_ASAP7_75t_R input251 (.A(net3599),
    .Y(net251));
 CKINVDCx20_ASAP7_75t_R _26045_ (.A(net1188),
    .Y(_17533_));
 NAND2x2_ASAP7_75t_R _26046_ (.A(net1535),
    .B(_17533_),
    .Y(_17534_));
 NOR2x2_ASAP7_75t_R _26047_ (.A(net2902),
    .B(net1088),
    .Y(_17535_));
 NOR2x2_ASAP7_75t_R _26048_ (.A(_00557_),
    .B(_00558_),
    .Y(_17536_));
 BUFx2_ASAP7_75t_R input250 (.A(net3676),
    .Y(net250));
 NAND2x2_ASAP7_75t_R _26050_ (.A(net1535),
    .B(net1007),
    .Y(_17538_));
 INVx1_ASAP7_75t_R _26051_ (.A(_17538_),
    .Y(_17539_));
 BUFx2_ASAP7_75t_R input249 (.A(net3904),
    .Y(net249));
 BUFx2_ASAP7_75t_R input248 (.A(net3673),
    .Y(net248));
 INVx2_ASAP7_75t_R _26054_ (.A(_00556_),
    .Y(_17542_));
 NOR2x2_ASAP7_75t_R _26055_ (.A(_00555_),
    .B(_17542_),
    .Y(_17543_));
 BUFx2_ASAP7_75t_R input247 (.A(net3564),
    .Y(net247));
 INVx4_ASAP7_75t_R _26057_ (.A(_00554_),
    .Y(_17545_));
 NOR2x2_ASAP7_75t_R _26058_ (.A(_00553_),
    .B(_17545_),
    .Y(_17546_));
 NAND2x2_ASAP7_75t_R _26059_ (.A(_17543_),
    .B(_17546_),
    .Y(_17547_));
 INVx4_ASAP7_75t_R _26060_ (.A(_17547_),
    .Y(_17548_));
 OAI21x1_ASAP7_75t_R _26061_ (.A1(net2906),
    .A2(_17539_),
    .B(_17548_),
    .Y(_17549_));
 NOR2x2_ASAP7_75t_R _26062_ (.A(net1536),
    .B(net1191),
    .Y(_17550_));
 NAND2x2_ASAP7_75t_R _26063_ (.A(_17550_),
    .B(net1006),
    .Y(_17551_));
 BUFx2_ASAP7_75t_R input246 (.A(net3588),
    .Y(net246));
 INVx2_ASAP7_75t_R _26065_ (.A(_17551_),
    .Y(_17553_));
 NAND2x1_ASAP7_75t_R _26066_ (.A(_17553_),
    .B(_17548_),
    .Y(_17554_));
 NAND2x2_ASAP7_75t_R _26067_ (.A(net1534),
    .B(net1184),
    .Y(_17555_));
 INVx2_ASAP7_75t_R _26068_ (.A(_00558_),
    .Y(_17556_));
 NAND2x2_ASAP7_75t_R _26069_ (.A(_00557_),
    .B(_17556_),
    .Y(_17557_));
 NOR2x2_ASAP7_75t_R _26070_ (.A(_17555_),
    .B(_17557_),
    .Y(_17558_));
 NAND2x1_ASAP7_75t_R _26071_ (.A(_17558_),
    .B(_17548_),
    .Y(_17559_));
 NAND3x1_ASAP7_75t_R _26072_ (.A(_17549_),
    .B(_17554_),
    .C(_17559_),
    .Y(_17560_));
 NOR2x2_ASAP7_75t_R _26073_ (.A(_00558_),
    .B(_17529_),
    .Y(_17561_));
 NAND2x2_ASAP7_75t_R _26074_ (.A(net1538),
    .B(_17561_),
    .Y(_17562_));
 NAND2x2_ASAP7_75t_R _26075_ (.A(_17550_),
    .B(_17561_),
    .Y(_17563_));
 BUFx2_ASAP7_75t_R input245 (.A(net3626),
    .Y(net245));
 NOR2x2_ASAP7_75t_R _26077_ (.A(_00555_),
    .B(_00556_),
    .Y(_17565_));
 NAND2x2_ASAP7_75t_R _26078_ (.A(_17565_),
    .B(_17546_),
    .Y(_17566_));
 BUFx2_ASAP7_75t_R input244 (.A(net3841),
    .Y(net244));
 AO21x1_ASAP7_75t_R _26080_ (.A1(_17562_),
    .A2(net1380),
    .B(_17566_),
    .Y(_17568_));
 INVx3_ASAP7_75t_R _26081_ (.A(_17566_),
    .Y(_17569_));
 NAND2x2_ASAP7_75t_R _26082_ (.A(_00557_),
    .B(_00558_),
    .Y(_17570_));
 INVx6_ASAP7_75t_R _26083_ (.A(net1609),
    .Y(_17571_));
 NAND2x2_ASAP7_75t_R _26084_ (.A(net1089),
    .B(_17571_),
    .Y(_17572_));
 INVx2_ASAP7_75t_R _26085_ (.A(_17572_),
    .Y(_17573_));
 NAND2x2_ASAP7_75t_R _26086_ (.A(_17569_),
    .B(_17573_),
    .Y(_17574_));
 CKINVDCx14_ASAP7_75t_R _26087_ (.A(net1005),
    .Y(_17575_));
 NOR2x2_ASAP7_75t_R _26088_ (.A(_17555_),
    .B(_17575_),
    .Y(_17576_));
 NAND2x1_ASAP7_75t_R _26089_ (.A(_17576_),
    .B(_17569_),
    .Y(_17577_));
 NAND3x1_ASAP7_75t_R _26090_ (.A(_17568_),
    .B(_17574_),
    .C(_17577_),
    .Y(_17578_));
 NOR2x1_ASAP7_75t_R _26091_ (.A(_17560_),
    .B(_17578_),
    .Y(_17579_));
 CKINVDCx20_ASAP7_75t_R _26092_ (.A(net1537),
    .Y(_17580_));
 NOR2x2_ASAP7_75t_R _26093_ (.A(net1190),
    .B(_17580_),
    .Y(_17581_));
 NAND2x2_ASAP7_75t_R _26094_ (.A(net1003),
    .B(_17581_),
    .Y(_17582_));
 BUFx2_ASAP7_75t_R input243 (.A(net3877),
    .Y(net243));
 BUFx2_ASAP7_75t_R input242 (.A(net3796),
    .Y(net242));
 BUFx2_ASAP7_75t_R input241 (.A(net3596),
    .Y(net241));
 NAND2x2_ASAP7_75t_R _26098_ (.A(_17580_),
    .B(net1003),
    .Y(_17586_));
 BUFx2_ASAP7_75t_R input240 (.A(net3611),
    .Y(net240));
 AND2x4_ASAP7_75t_R _26100_ (.A(_00555_),
    .B(_00556_),
    .Y(_17588_));
 NAND2x2_ASAP7_75t_R _26101_ (.A(_17546_),
    .B(_17588_),
    .Y(_17589_));
 BUFx2_ASAP7_75t_R input239 (.A(net3826),
    .Y(net239));
 AO21x2_ASAP7_75t_R _26103_ (.A1(net2013),
    .A2(_17586_),
    .B(_17589_),
    .Y(_17591_));
 NOR2x2_ASAP7_75t_R _26104_ (.A(_00557_),
    .B(_17556_),
    .Y(_17592_));
 NAND2x2_ASAP7_75t_R _26105_ (.A(net2086),
    .B(_17581_),
    .Y(_17593_));
 BUFx2_ASAP7_75t_R input238 (.A(net3652),
    .Y(net238));
 BUFx2_ASAP7_75t_R input237 (.A(net3629),
    .Y(net237));
 NAND2x2_ASAP7_75t_R _26108_ (.A(_17550_),
    .B(net2086),
    .Y(_17596_));
 BUFx2_ASAP7_75t_R input236 (.A(net3620),
    .Y(net236));
 AO21x1_ASAP7_75t_R _26110_ (.A1(net1098),
    .A2(net2892),
    .B(_17589_),
    .Y(_17598_));
 NAND2x2_ASAP7_75t_R _26111_ (.A(_17591_),
    .B(_17598_),
    .Y(_17599_));
 NOR2x2_ASAP7_75t_R _26112_ (.A(net1534),
    .B(_17533_),
    .Y(_17600_));
 NAND2x2_ASAP7_75t_R _26113_ (.A(_00555_),
    .B(_00556_),
    .Y(_17601_));
 INVx4_ASAP7_75t_R _26114_ (.A(_00553_),
    .Y(_17602_));
 NAND2x2_ASAP7_75t_R _26115_ (.A(_00554_),
    .B(_17602_),
    .Y(_17603_));
 NOR2x2_ASAP7_75t_R _26116_ (.A(_17601_),
    .B(_17603_),
    .Y(_17604_));
 NAND2x2_ASAP7_75t_R _26117_ (.A(net2826),
    .B(_17604_),
    .Y(_17605_));
 BUFx2_ASAP7_75t_R input235 (.A(net3775),
    .Y(net235));
 NOR2x2_ASAP7_75t_R _26119_ (.A(_17555_),
    .B(net1607),
    .Y(_17607_));
 NAND2x2_ASAP7_75t_R _26120_ (.A(net1184),
    .B(_17580_),
    .Y(_17608_));
 NOR2x2_ASAP7_75t_R _26121_ (.A(net1607),
    .B(_17608_),
    .Y(_17609_));
 OAI21x1_ASAP7_75t_R _26122_ (.A1(_17607_),
    .A2(_17609_),
    .B(_17604_),
    .Y(_17610_));
 OAI21x1_ASAP7_75t_R _26123_ (.A1(net1832),
    .A2(_17605_),
    .B(_17610_),
    .Y(_17611_));
 INVx2_ASAP7_75t_R _26124_ (.A(_00555_),
    .Y(_17612_));
 NOR2x2_ASAP7_75t_R _26125_ (.A(_00556_),
    .B(_17612_),
    .Y(_17613_));
 NAND2x2_ASAP7_75t_R _26126_ (.A(_17613_),
    .B(_17546_),
    .Y(_17614_));
 BUFx2_ASAP7_75t_R input234 (.A(net3811),
    .Y(net234));
 NOR2x2_ASAP7_75t_R _26128_ (.A(net1607),
    .B(_17534_),
    .Y(_17616_));
 NAND2x2_ASAP7_75t_R _26129_ (.A(_00555_),
    .B(_17542_),
    .Y(_17617_));
 NOR2x2_ASAP7_75t_R _26130_ (.A(_17617_),
    .B(_17603_),
    .Y(_17618_));
 OAI21x1_ASAP7_75t_R _26131_ (.A1(net2640),
    .A2(_17609_),
    .B(_17618_),
    .Y(_17619_));
 OAI21x1_ASAP7_75t_R _26132_ (.A1(_17614_),
    .A2(_17586_),
    .B(_17619_),
    .Y(_17620_));
 NOR3x2_ASAP7_75t_R _26133_ (.B(_17611_),
    .C(_17620_),
    .Y(_17621_),
    .A(_17599_));
 NAND2x2_ASAP7_75t_R _26134_ (.A(_17579_),
    .B(_17621_),
    .Y(_17622_));
 INVx1_ASAP7_75t_R _26135_ (.A(_17622_),
    .Y(_17623_));
 NAND2x2_ASAP7_75t_R _26136_ (.A(_17550_),
    .B(_17571_),
    .Y(_17624_));
 BUFx2_ASAP7_75t_R input233 (.A(net3605),
    .Y(net233));
 CKINVDCx9p33_ASAP7_75t_R _26138_ (.A(_17607_),
    .Y(_17626_));
 BUFx2_ASAP7_75t_R input232 (.A(net3727),
    .Y(net232));
 NOR2x2_ASAP7_75t_R _26140_ (.A(_00553_),
    .B(_00554_),
    .Y(_17628_));
 NAND2x2_ASAP7_75t_R _26141_ (.A(_17628_),
    .B(_17543_),
    .Y(_17629_));
 BUFx2_ASAP7_75t_R input231 (.A(net3742),
    .Y(net231));
 AOI21x1_ASAP7_75t_R _26143_ (.A1(net2899),
    .A2(_17626_),
    .B(_17629_),
    .Y(_17631_));
 NAND2x2_ASAP7_75t_R _26144_ (.A(net2891),
    .B(net1004),
    .Y(_17632_));
 NAND2x1_ASAP7_75t_R _26145_ (.A(_17534_),
    .B(net2086),
    .Y(_17633_));
 AOI21x1_ASAP7_75t_R _26146_ (.A1(_17632_),
    .A2(_17633_),
    .B(_17629_),
    .Y(_17634_));
 BUFx2_ASAP7_75t_R input230 (.A(net3912),
    .Y(net230));
 NOR2x2_ASAP7_75t_R _26148_ (.A(_17629_),
    .B(_17562_),
    .Y(_17636_));
 NOR3x2_ASAP7_75t_R _26149_ (.B(_17634_),
    .C(_17636_),
    .Y(_17637_),
    .A(_17631_));
 AND2x4_ASAP7_75t_R _26150_ (.A(net1534),
    .B(net1184),
    .Y(_17638_));
 NAND2x2_ASAP7_75t_R _26151_ (.A(net2088),
    .B(_17638_),
    .Y(_17639_));
 BUFx2_ASAP7_75t_R input229 (.A(net3844),
    .Y(net229));
 NAND2x2_ASAP7_75t_R _26153_ (.A(_17628_),
    .B(_17565_),
    .Y(_17641_));
 BUFx2_ASAP7_75t_R input228 (.A(net3661),
    .Y(net228));
 BUFx2_ASAP7_75t_R input227 (.A(net3898),
    .Y(net227));
 AOI21x1_ASAP7_75t_R _26156_ (.A1(net2488),
    .A2(_17639_),
    .B(net2484),
    .Y(_17644_));
 NAND2x2_ASAP7_75t_R _26157_ (.A(net1001),
    .B(_17600_),
    .Y(_17645_));
 NOR2x2_ASAP7_75t_R _26158_ (.A(_17641_),
    .B(_17645_),
    .Y(_17646_));
 NAND2x2_ASAP7_75t_R _26159_ (.A(_17580_),
    .B(net2086),
    .Y(_17647_));
 NOR2x2_ASAP7_75t_R _26160_ (.A(_17641_),
    .B(_17647_),
    .Y(_17648_));
 NOR3x2_ASAP7_75t_R _26161_ (.B(_17646_),
    .C(_17648_),
    .Y(_17649_),
    .A(_17644_));
 INVx3_ASAP7_75t_R _26162_ (.A(_17641_),
    .Y(_17650_));
 BUFx2_ASAP7_75t_R input226 (.A(net3805),
    .Y(net226));
 BUFx2_ASAP7_75t_R input225 (.A(net3570),
    .Y(net225));
 BUFx2_ASAP7_75t_R input224 (.A(net3787),
    .Y(net224));
 AOI211x1_ASAP7_75t_R _26166_ (.A1(net1123),
    .A2(net1188),
    .B(net2484),
    .C(net1103),
    .Y(_17654_));
 AOI21x1_ASAP7_75t_R _26167_ (.A1(_17558_),
    .A2(_17650_),
    .B(_17654_),
    .Y(_17655_));
 NAND3x2_ASAP7_75t_R _26168_ (.B(_17649_),
    .C(_17655_),
    .Y(_17656_),
    .A(_17637_));
 NAND2x2_ASAP7_75t_R _26169_ (.A(_17628_),
    .B(_17588_),
    .Y(_17657_));
 BUFx2_ASAP7_75t_R input223 (.A(net3835),
    .Y(net223));
 NOR2x2_ASAP7_75t_R _26171_ (.A(_17575_),
    .B(_17657_),
    .Y(_17659_));
 NAND2x2_ASAP7_75t_R _26172_ (.A(_17580_),
    .B(_17533_),
    .Y(_17660_));
 NOR2x2_ASAP7_75t_R _26173_ (.A(net2902),
    .B(_17660_),
    .Y(_17661_));
 INVx2_ASAP7_75t_R _26174_ (.A(_17657_),
    .Y(_17662_));
 OA21x2_ASAP7_75t_R _26175_ (.A1(net2906),
    .A2(_17661_),
    .B(_17662_),
    .Y(_17663_));
 BUFx2_ASAP7_75t_R input222 (.A(net3848),
    .Y(net222));
 NAND2x2_ASAP7_75t_R _26177_ (.A(net1831),
    .B(_17571_),
    .Y(_17665_));
 NOR2x1_ASAP7_75t_R _26178_ (.A(net2847),
    .B(_17665_),
    .Y(_17666_));
 AOI211x1_ASAP7_75t_R _26179_ (.A1(_17659_),
    .A2(_17660_),
    .B(_17663_),
    .C(_17666_),
    .Y(_17667_));
 BUFx2_ASAP7_75t_R input221 (.A(net3670),
    .Y(net221));
 NOR2x2_ASAP7_75t_R _26181_ (.A(_17555_),
    .B(net2905),
    .Y(_17669_));
 NAND2x2_ASAP7_75t_R _26182_ (.A(_17628_),
    .B(_17613_),
    .Y(_17670_));
 INVx5_ASAP7_75t_R _26183_ (.A(_17670_),
    .Y(_17671_));
 OAI21x1_ASAP7_75t_R _26184_ (.A1(_17669_),
    .A2(net2906),
    .B(_17671_),
    .Y(_17672_));
 NOR2x2_ASAP7_75t_R _26185_ (.A(net2902),
    .B(_17608_),
    .Y(_17673_));
 OAI21x1_ASAP7_75t_R _26186_ (.A1(_17673_),
    .A2(_17661_),
    .B(_17671_),
    .Y(_17674_));
 NAND2x2_ASAP7_75t_R _26187_ (.A(_17672_),
    .B(_17674_),
    .Y(_17675_));
 NOR2x2_ASAP7_75t_R _26188_ (.A(net3323),
    .B(net1973),
    .Y(_17676_));
 OA21x2_ASAP7_75t_R _26189_ (.A1(net1901),
    .A2(_17609_),
    .B(_17671_),
    .Y(_17677_));
 INVx4_ASAP7_75t_R _26190_ (.A(_17582_),
    .Y(_17678_));
 NOR2x2_ASAP7_75t_R _26191_ (.A(_17608_),
    .B(_17575_),
    .Y(_17679_));
 OA21x2_ASAP7_75t_R _26192_ (.A1(_17678_),
    .A2(_17679_),
    .B(_17671_),
    .Y(_17680_));
 NOR3x2_ASAP7_75t_R _26193_ (.B(_17677_),
    .C(_17680_),
    .Y(_17681_),
    .A(_17675_));
 NAND2x2_ASAP7_75t_R _26194_ (.A(_17667_),
    .B(_17681_),
    .Y(_17682_));
 NOR2x1_ASAP7_75t_R _26195_ (.A(_17656_),
    .B(_17682_),
    .Y(_17683_));
 NAND2x1_ASAP7_75t_R _26196_ (.A(_17623_),
    .B(_17683_),
    .Y(_17684_));
 NAND2x2_ASAP7_75t_R _26197_ (.A(_17600_),
    .B(_17561_),
    .Y(_17685_));
 BUFx2_ASAP7_75t_R input220 (.A(net3614),
    .Y(net220));
 NAND2x2_ASAP7_75t_R _26199_ (.A(_17581_),
    .B(_17561_),
    .Y(_17687_));
 BUFx2_ASAP7_75t_R input219 (.A(net3582),
    .Y(net219));
 NAND2x2_ASAP7_75t_R _26201_ (.A(_00553_),
    .B(_00554_),
    .Y(_17689_));
 INVx3_ASAP7_75t_R _26202_ (.A(_17689_),
    .Y(_17690_));
 NAND2x2_ASAP7_75t_R _26203_ (.A(_17613_),
    .B(_17690_),
    .Y(_17691_));
 AOI21x1_ASAP7_75t_R _26204_ (.A1(net998),
    .A2(net2598),
    .B(_17691_),
    .Y(_17692_));
 AOI21x1_ASAP7_75t_R _26205_ (.A1(_17596_),
    .A2(_17639_),
    .B(_17691_),
    .Y(_17693_));
 NOR2x2_ASAP7_75t_R _26206_ (.A(net1535),
    .B(net1607),
    .Y(_17694_));
 CKINVDCx6p67_ASAP7_75t_R _26207_ (.A(_17694_),
    .Y(_17695_));
 BUFx2_ASAP7_75t_R input218 (.A(net3655),
    .Y(net218));
 NOR2x2_ASAP7_75t_R _26209_ (.A(_17695_),
    .B(net3088),
    .Y(_17697_));
 NOR3x2_ASAP7_75t_R _26210_ (.B(_17693_),
    .C(_17697_),
    .Y(_17698_),
    .A(_17692_));
 BUFx2_ASAP7_75t_R input217 (.A(net3688),
    .Y(net217));
 NOR2x2_ASAP7_75t_R _26212_ (.A(_17601_),
    .B(_17689_),
    .Y(_17700_));
 CKINVDCx6p67_ASAP7_75t_R _26213_ (.A(_17700_),
    .Y(_17701_));
 BUFx2_ASAP7_75t_R input216 (.A(net3954),
    .Y(net216));
 AO21x1_ASAP7_75t_R _26215_ (.A1(net1098),
    .A2(_17647_),
    .B(_17701_),
    .Y(_17703_));
 BUFx2_ASAP7_75t_R input215 (.A(net3617),
    .Y(net215));
 AO21x1_ASAP7_75t_R _26217_ (.A1(_17582_),
    .A2(net2385),
    .B(_17701_),
    .Y(_17705_));
 AND2x2_ASAP7_75t_R _26218_ (.A(_17703_),
    .B(_17705_),
    .Y(_17706_));
 NOR2x1_ASAP7_75t_R _26219_ (.A(_17695_),
    .B(_17701_),
    .Y(_17707_));
 BUFx2_ASAP7_75t_R input214 (.A(net4026),
    .Y(net214));
 AOI211x1_ASAP7_75t_R _26221_ (.A1(net1123),
    .A2(net2770),
    .B(_17701_),
    .C(net1976),
    .Y(_17709_));
 NOR2x2_ASAP7_75t_R _26222_ (.A(_17707_),
    .B(_17709_),
    .Y(_17710_));
 NAND3x1_ASAP7_75t_R _26223_ (.A(_17698_),
    .B(_17706_),
    .C(_17710_),
    .Y(_17711_));
 NAND2x2_ASAP7_75t_R _26224_ (.A(_17565_),
    .B(_17690_),
    .Y(_17712_));
 NOR2x2_ASAP7_75t_R _26225_ (.A(net2884),
    .B(net999),
    .Y(_17713_));
 INVx4_ASAP7_75t_R _26226_ (.A(_17712_),
    .Y(_17714_));
 OAI21x1_ASAP7_75t_R _26227_ (.A1(_17616_),
    .A2(_17694_),
    .B(_17714_),
    .Y(_17715_));
 INVx1_ASAP7_75t_R _26228_ (.A(_17715_),
    .Y(_17716_));
 NOR2x1_ASAP7_75t_R _26229_ (.A(_17716_),
    .B(_17713_),
    .Y(_17717_));
 NOR2x1_ASAP7_75t_R _26230_ (.A(net2884),
    .B(_17639_),
    .Y(_17718_));
 BUFx2_ASAP7_75t_R input213 (.A(net3703),
    .Y(net213));
 AOI211x1_ASAP7_75t_R _26232_ (.A1(net2862),
    .A2(net1194),
    .B(net2884),
    .C(_17575_),
    .Y(_17720_));
 NOR2x1_ASAP7_75t_R _26233_ (.A(_17718_),
    .B(_17720_),
    .Y(_17721_));
 NAND2x1_ASAP7_75t_R _26234_ (.A(_17717_),
    .B(_17721_),
    .Y(_17722_));
 INVx1_ASAP7_75t_R _26235_ (.A(_17722_),
    .Y(_17723_));
 BUFx2_ASAP7_75t_R input212 (.A(net3647),
    .Y(net212));
 NAND2x2_ASAP7_75t_R _26237_ (.A(_17543_),
    .B(_17690_),
    .Y(_17725_));
 BUFx2_ASAP7_75t_R input211 (.A(net3706),
    .Y(net211));
 AO21x1_ASAP7_75t_R _26239_ (.A1(net998),
    .A2(net2598),
    .B(_17725_),
    .Y(_17727_));
 NOR2x1_ASAP7_75t_R _26240_ (.A(net1610),
    .B(_17725_),
    .Y(_17728_));
 NAND2x1_ASAP7_75t_R _26241_ (.A(_17660_),
    .B(_17728_),
    .Y(_17729_));
 NAND2x1_ASAP7_75t_R _26242_ (.A(_17727_),
    .B(_17729_),
    .Y(_17730_));
 NOR2x2_ASAP7_75t_R _26243_ (.A(net1539),
    .B(net2902),
    .Y(_17731_));
 NAND2x2_ASAP7_75t_R _26244_ (.A(_00556_),
    .B(_17612_),
    .Y(_17732_));
 NOR2x2_ASAP7_75t_R _26245_ (.A(_17689_),
    .B(_17732_),
    .Y(_17733_));
 OAI21x1_ASAP7_75t_R _26246_ (.A1(_17731_),
    .A2(_17535_),
    .B(_17733_),
    .Y(_17734_));
 INVx1_ASAP7_75t_R _26247_ (.A(_17734_),
    .Y(_17735_));
 BUFx2_ASAP7_75t_R input210 (.A(net3745),
    .Y(net210));
 AOI211x1_ASAP7_75t_R _26249_ (.A1(net1123),
    .A2(net2879),
    .B(_17725_),
    .C(_17575_),
    .Y(_17737_));
 NOR2x1_ASAP7_75t_R _26250_ (.A(_17735_),
    .B(_17737_),
    .Y(_17738_));
 INVx1_ASAP7_75t_R _26251_ (.A(_17738_),
    .Y(_17739_));
 NOR2x1_ASAP7_75t_R _26252_ (.A(_17730_),
    .B(_17739_),
    .Y(_17740_));
 NAND2x1_ASAP7_75t_R _26253_ (.A(_17723_),
    .B(_17740_),
    .Y(_17741_));
 NOR2x1_ASAP7_75t_R _26254_ (.A(_17711_),
    .B(_17741_),
    .Y(_17742_));
 NOR2x2_ASAP7_75t_R _26255_ (.A(_00554_),
    .B(_17602_),
    .Y(_17743_));
 NAND2x2_ASAP7_75t_R _26256_ (.A(_17613_),
    .B(_17743_),
    .Y(_17744_));
 NOR2x2_ASAP7_75t_R _26257_ (.A(net1607),
    .B(net1831),
    .Y(_17745_));
 INVx2_ASAP7_75t_R _26258_ (.A(_17745_),
    .Y(_17746_));
 NOR2x1_ASAP7_75t_R _26259_ (.A(_17744_),
    .B(_17746_),
    .Y(_17747_));
 BUFx2_ASAP7_75t_R input209 (.A(net3579),
    .Y(net209));
 AOI21x1_ASAP7_75t_R _26261_ (.A1(net1383),
    .A2(_17685_),
    .B(_17744_),
    .Y(_17749_));
 NOR2x1_ASAP7_75t_R _26262_ (.A(_17747_),
    .B(_17749_),
    .Y(_17750_));
 BUFx2_ASAP7_75t_R input208 (.A(net3632),
    .Y(net208));
 BUFx2_ASAP7_75t_R input207 (.A(net3593),
    .Y(net207));
 BUFx2_ASAP7_75t_R input206 (.A(net3942),
    .Y(net206));
 AO31x2_ASAP7_75t_R _26266_ (.A1(net2630),
    .A2(net2893),
    .A3(net1082),
    .B(_17744_),
    .Y(_17754_));
 NAND2x1_ASAP7_75t_R _26267_ (.A(_17750_),
    .B(_17754_),
    .Y(_17755_));
 NAND2x2_ASAP7_75t_R _26268_ (.A(_17561_),
    .B(_17638_),
    .Y(_17756_));
 NOR2x2_ASAP7_75t_R _26269_ (.A(_17580_),
    .B(net1607),
    .Y(_17757_));
 INVx4_ASAP7_75t_R _26270_ (.A(_17757_),
    .Y(_17758_));
 NAND2x2_ASAP7_75t_R _26271_ (.A(_17743_),
    .B(_17588_),
    .Y(_17759_));
 BUFx2_ASAP7_75t_R input205 (.A(net3694),
    .Y(net205));
 AO21x1_ASAP7_75t_R _26273_ (.A1(_17756_),
    .A2(_17758_),
    .B(_17759_),
    .Y(_17761_));
 AO21x2_ASAP7_75t_R _26274_ (.A1(net2532),
    .A2(net2892),
    .B(_17759_),
    .Y(_17762_));
 BUFx2_ASAP7_75t_R input204 (.A(net3608),
    .Y(net204));
 AO21x2_ASAP7_75t_R _26276_ (.A1(net2385),
    .A2(_17538_),
    .B(_17759_),
    .Y(_17764_));
 NAND3x1_ASAP7_75t_R _26277_ (.A(_17761_),
    .B(_17762_),
    .C(_17764_),
    .Y(_17765_));
 NOR2x1_ASAP7_75t_R _26278_ (.A(_17765_),
    .B(_17755_),
    .Y(_17766_));
 INVx1_ASAP7_75t_R _26279_ (.A(_17766_),
    .Y(_17767_));
 AO21x1_ASAP7_75t_R _26280_ (.A1(net1089),
    .A2(_17608_),
    .B(_17575_),
    .Y(_17768_));
 NAND2x1_ASAP7_75t_R _26281_ (.A(net1082),
    .B(_17768_),
    .Y(_17769_));
 NAND2x2_ASAP7_75t_R _26282_ (.A(_17565_),
    .B(_17743_),
    .Y(_17770_));
 INVx4_ASAP7_75t_R _26283_ (.A(_17770_),
    .Y(_17771_));
 BUFx2_ASAP7_75t_R input203 (.A(net3641),
    .Y(net203));
 AOI211x1_ASAP7_75t_R _26285_ (.A1(net2862),
    .A2(net1192),
    .B(net2909),
    .C(net1103),
    .Y(_17773_));
 NOR2x2_ASAP7_75t_R _26286_ (.A(net1973),
    .B(_17660_),
    .Y(_17774_));
 OA21x2_ASAP7_75t_R _26287_ (.A1(net1901),
    .A2(_17774_),
    .B(_17771_),
    .Y(_17775_));
 AOI211x1_ASAP7_75t_R _26288_ (.A1(_17769_),
    .A2(_17771_),
    .B(_17773_),
    .C(_17775_),
    .Y(_17776_));
 NAND2x2_ASAP7_75t_R _26289_ (.A(_17743_),
    .B(_17543_),
    .Y(_17777_));
 BUFx2_ASAP7_75t_R input202 (.A(net3667),
    .Y(net202));
 NOR2x1_ASAP7_75t_R _26291_ (.A(net2385),
    .B(_17777_),
    .Y(_17779_));
 NOR2x2_ASAP7_75t_R _26292_ (.A(net2907),
    .B(net2902),
    .Y(_17780_));
 NAND2x2_ASAP7_75t_R _26293_ (.A(_00553_),
    .B(_17545_),
    .Y(_17781_));
 NOR2x2_ASAP7_75t_R _26294_ (.A(_17781_),
    .B(_17732_),
    .Y(_17782_));
 OA21x2_ASAP7_75t_R _26295_ (.A1(_17661_),
    .A2(_17780_),
    .B(_17782_),
    .Y(_17783_));
 OR2x2_ASAP7_75t_R _26296_ (.A(_17779_),
    .B(_17783_),
    .Y(_17784_));
 AO21x1_ASAP7_75t_R _26297_ (.A1(net936),
    .A2(net941),
    .B(_17777_),
    .Y(_17785_));
 INVx2_ASAP7_75t_R _26298_ (.A(_17562_),
    .Y(_17786_));
 NAND2x2_ASAP7_75t_R _26299_ (.A(_17782_),
    .B(_17786_),
    .Y(_17787_));
 NOR2x2_ASAP7_75t_R _26300_ (.A(net1608),
    .B(_17660_),
    .Y(_17788_));
 BUFx2_ASAP7_75t_R input201 (.A(net3682),
    .Y(net201));
 OAI21x1_ASAP7_75t_R _26302_ (.A1(net2641),
    .A2(_17788_),
    .B(_17782_),
    .Y(_17790_));
 NAND3x2_ASAP7_75t_R _26303_ (.B(_17787_),
    .C(_17790_),
    .Y(_17791_),
    .A(_17785_));
 NOR2x2_ASAP7_75t_R _26304_ (.A(_17784_),
    .B(_17791_),
    .Y(_17792_));
 NAND2x1_ASAP7_75t_R _26305_ (.A(_17776_),
    .B(_17792_),
    .Y(_17793_));
 NOR2x1_ASAP7_75t_R _26306_ (.A(_17767_),
    .B(_17793_),
    .Y(_17794_));
 NAND2x1_ASAP7_75t_R _26307_ (.A(_17742_),
    .B(_17794_),
    .Y(_17795_));
 NOR2x2_ASAP7_75t_R _26308_ (.A(_17684_),
    .B(_17795_),
    .Y(_17796_));
 OA21x2_ASAP7_75t_R _26309_ (.A1(_17774_),
    .A2(_17558_),
    .B(net3086),
    .Y(_17797_));
 BUFx2_ASAP7_75t_R input200 (.A(net4001),
    .Y(net200));
 AOI211x1_ASAP7_75t_R _26311_ (.A1(net2862),
    .A2(net2891),
    .B(_17701_),
    .C(_17575_),
    .Y(_17799_));
 NOR2x2_ASAP7_75t_R _26312_ (.A(_17797_),
    .B(_17799_),
    .Y(_17800_));
 NOR2x2_ASAP7_75t_R _26313_ (.A(_17689_),
    .B(_17617_),
    .Y(_17801_));
 OA21x2_ASAP7_75t_R _26314_ (.A1(_17780_),
    .A2(_17731_),
    .B(_17801_),
    .Y(_17802_));
 AOI211x1_ASAP7_75t_R _26315_ (.A1(net2907),
    .A2(net1194),
    .B(_17691_),
    .C(_17575_),
    .Y(_17803_));
 NOR2x2_ASAP7_75t_R _26316_ (.A(_17802_),
    .B(_17803_),
    .Y(_17804_));
 OA21x2_ASAP7_75t_R _26317_ (.A1(_17609_),
    .A2(_17757_),
    .B(_17801_),
    .Y(_17805_));
 OA21x2_ASAP7_75t_R _26318_ (.A1(_17774_),
    .A2(_17558_),
    .B(_17801_),
    .Y(_17806_));
 NOR2x2_ASAP7_75t_R _26319_ (.A(_17805_),
    .B(_17806_),
    .Y(_17807_));
 NAND3x2_ASAP7_75t_R _26320_ (.B(_17804_),
    .C(_17807_),
    .Y(_17808_),
    .A(_17800_));
 NOR2x2_ASAP7_75t_R _26321_ (.A(net1193),
    .B(net1611),
    .Y(_17809_));
 NAND2x2_ASAP7_75t_R _26322_ (.A(_17809_),
    .B(_17714_),
    .Y(_17810_));
 AO21x1_ASAP7_75t_R _26323_ (.A1(net2598),
    .A2(_17563_),
    .B(net2884),
    .Y(_17811_));
 NAND2x1_ASAP7_75t_R _26324_ (.A(_17810_),
    .B(_17811_),
    .Y(_17812_));
 NAND2x2_ASAP7_75t_R _26325_ (.A(net2871),
    .B(_17638_),
    .Y(_17813_));
 AO21x1_ASAP7_75t_R _26326_ (.A1(_17813_),
    .A2(net2385),
    .B(net2882),
    .Y(_17814_));
 NAND2x2_ASAP7_75t_R _26327_ (.A(net2086),
    .B(_17600_),
    .Y(_17815_));
 BUFx2_ASAP7_75t_R input199 (.A(net3901),
    .Y(net199));
 AO21x1_ASAP7_75t_R _26329_ (.A1(net2236),
    .A2(_17596_),
    .B(_17712_),
    .Y(_17817_));
 NAND2x1_ASAP7_75t_R _26330_ (.A(_17817_),
    .B(_17814_),
    .Y(_17818_));
 NOR2x1_ASAP7_75t_R _26331_ (.A(_17812_),
    .B(_17818_),
    .Y(_17819_));
 NAND2x2_ASAP7_75t_R _26332_ (.A(_17733_),
    .B(_17678_),
    .Y(_17820_));
 NAND2x2_ASAP7_75t_R _26333_ (.A(_17820_),
    .B(_17734_),
    .Y(_17821_));
 AND3x2_ASAP7_75t_R _26334_ (.A(_17733_),
    .B(_17660_),
    .C(_17571_),
    .Y(_17822_));
 AND3x1_ASAP7_75t_R _26335_ (.A(_17733_),
    .B(net2907),
    .C(_17561_),
    .Y(_17823_));
 NOR3x1_ASAP7_75t_R _26336_ (.A(_17821_),
    .B(_17822_),
    .C(_17823_),
    .Y(_17824_));
 NAND2x1_ASAP7_75t_R _26337_ (.A(_17819_),
    .B(_17824_),
    .Y(_17825_));
 NOR2x2_ASAP7_75t_R _26338_ (.A(_17808_),
    .B(_17825_),
    .Y(_17826_));
 AO21x1_ASAP7_75t_R _26339_ (.A1(net941),
    .A2(net1103),
    .B(_17777_),
    .Y(_17827_));
 AO21x1_ASAP7_75t_R _26340_ (.A1(net2532),
    .A2(_17586_),
    .B(_17777_),
    .Y(_17828_));
 NAND2x1_ASAP7_75t_R _26341_ (.A(_17827_),
    .B(_17828_),
    .Y(_17829_));
 INVx1_ASAP7_75t_R _26342_ (.A(_17829_),
    .Y(_17830_));
 INVx2_ASAP7_75t_R _26343_ (.A(_17809_),
    .Y(_17831_));
 AO21x1_ASAP7_75t_R _26344_ (.A1(_17562_),
    .A2(net1382),
    .B(_17770_),
    .Y(_17832_));
 OAI21x1_ASAP7_75t_R _26345_ (.A1(_17831_),
    .A2(_17770_),
    .B(_17832_),
    .Y(_17833_));
 NAND2x2_ASAP7_75t_R _26346_ (.A(net1537),
    .B(net2086),
    .Y(_17834_));
 AO21x1_ASAP7_75t_R _26347_ (.A1(net2236),
    .A2(_17834_),
    .B(_17770_),
    .Y(_17835_));
 NAND3x2_ASAP7_75t_R _26348_ (.B(net1003),
    .C(_17555_),
    .Y(_17836_),
    .A(_17771_));
 NAND2x2_ASAP7_75t_R _26349_ (.A(_17835_),
    .B(_17836_),
    .Y(_17837_));
 NOR2x1_ASAP7_75t_R _26350_ (.A(_17833_),
    .B(_17837_),
    .Y(_17838_));
 NAND2x1_ASAP7_75t_R _26351_ (.A(_17830_),
    .B(_17838_),
    .Y(_17839_));
 BUFx2_ASAP7_75t_R input198 (.A(net3623),
    .Y(net198));
 AO31x2_ASAP7_75t_R _26353_ (.A1(_17831_),
    .A2(net997),
    .A3(net2599),
    .B(_17744_),
    .Y(_17841_));
 AO31x2_ASAP7_75t_R _26354_ (.A1(net3195),
    .A2(net2532),
    .A3(net2238),
    .B(_17744_),
    .Y(_17842_));
 NAND2x1_ASAP7_75t_R _26355_ (.A(_17841_),
    .B(_17842_),
    .Y(_17843_));
 AO21x1_ASAP7_75t_R _26356_ (.A1(net2236),
    .A2(net2892),
    .B(_17759_),
    .Y(_17844_));
 NAND2x2_ASAP7_75t_R _26357_ (.A(_17581_),
    .B(_17571_),
    .Y(_17845_));
 BUFx2_ASAP7_75t_R input197 (.A(net3635),
    .Y(net197));
 AO21x1_ASAP7_75t_R _26359_ (.A1(_17845_),
    .A2(net1382),
    .B(_17759_),
    .Y(_17847_));
 AO21x1_ASAP7_75t_R _26360_ (.A1(net2013),
    .A2(net3195),
    .B(_17759_),
    .Y(_17848_));
 NAND3x1_ASAP7_75t_R _26361_ (.A(_17844_),
    .B(_17847_),
    .C(_17848_),
    .Y(_17849_));
 NOR2x1_ASAP7_75t_R _26362_ (.A(_17843_),
    .B(_17849_),
    .Y(_17850_));
 INVx1_ASAP7_75t_R _26363_ (.A(_17850_),
    .Y(_17851_));
 NOR2x1_ASAP7_75t_R _26364_ (.A(_17839_),
    .B(_17851_),
    .Y(_17852_));
 NAND2x2_ASAP7_75t_R _26365_ (.A(_17826_),
    .B(_17852_),
    .Y(_17853_));
 AO21x1_ASAP7_75t_R _26366_ (.A1(_17813_),
    .A2(net3194),
    .B(_17614_),
    .Y(_17854_));
 AO21x1_ASAP7_75t_R _26367_ (.A1(net2895),
    .A2(_17815_),
    .B(_17614_),
    .Y(_17855_));
 NAND2x1_ASAP7_75t_R _26368_ (.A(_17854_),
    .B(_17855_),
    .Y(_17856_));
 AO21x1_ASAP7_75t_R _26369_ (.A1(net997),
    .A2(net1380),
    .B(_17614_),
    .Y(_17857_));
 AO21x1_ASAP7_75t_R _26370_ (.A1(_17845_),
    .A2(net2901),
    .B(_17614_),
    .Y(_17858_));
 NAND2x1_ASAP7_75t_R _26371_ (.A(_17857_),
    .B(_17858_),
    .Y(_17859_));
 NOR2x1_ASAP7_75t_R _26372_ (.A(_17856_),
    .B(_17859_),
    .Y(_17860_));
 AO21x2_ASAP7_75t_R _26373_ (.A1(_17626_),
    .A2(net2901),
    .B(_17589_),
    .Y(_17861_));
 AO21x1_ASAP7_75t_R _26374_ (.A1(net2895),
    .A2(_17639_),
    .B(_17589_),
    .Y(_17862_));
 NAND2x2_ASAP7_75t_R _26375_ (.A(_17604_),
    .B(net1901),
    .Y(_17863_));
 NAND3x2_ASAP7_75t_R _26376_ (.B(_17862_),
    .C(_17863_),
    .Y(_17864_),
    .A(_17861_));
 INVx1_ASAP7_75t_R _26377_ (.A(_17864_),
    .Y(_17865_));
 NAND2x1_ASAP7_75t_R _26378_ (.A(_17860_),
    .B(_17865_),
    .Y(_17866_));
 BUFx2_ASAP7_75t_R input196 (.A(net3644),
    .Y(net196));
 AO21x1_ASAP7_75t_R _26380_ (.A1(net1788),
    .A2(_17834_),
    .B(_17547_),
    .Y(_17868_));
 AO21x1_ASAP7_75t_R _26381_ (.A1(_17645_),
    .A2(_17538_),
    .B(_17547_),
    .Y(_17869_));
 NAND2x1_ASAP7_75t_R _26382_ (.A(_17607_),
    .B(_17548_),
    .Y(_17870_));
 NAND3x1_ASAP7_75t_R _26383_ (.A(_17868_),
    .B(_17869_),
    .C(_17870_),
    .Y(_17871_));
 AO21x1_ASAP7_75t_R _26384_ (.A1(_17626_),
    .A2(_17845_),
    .B(_17566_),
    .Y(_17872_));
 AO21x1_ASAP7_75t_R _26385_ (.A1(_17647_),
    .A2(_17645_),
    .B(_17566_),
    .Y(_17873_));
 NAND3x1_ASAP7_75t_R _26386_ (.A(_17872_),
    .B(_17873_),
    .C(_17568_),
    .Y(_17874_));
 NOR2x1_ASAP7_75t_R _26387_ (.A(_17871_),
    .B(_17874_),
    .Y(_17875_));
 INVx1_ASAP7_75t_R _26388_ (.A(_17875_),
    .Y(_17876_));
 NOR2x1_ASAP7_75t_R _26389_ (.A(_17866_),
    .B(_17876_),
    .Y(_17877_));
 BUFx2_ASAP7_75t_R input195 (.A(net3697),
    .Y(net195));
 AOI21x1_ASAP7_75t_R _26391_ (.A1(net997),
    .A2(_17665_),
    .B(net2889),
    .Y(_17879_));
 AOI21x1_ASAP7_75t_R _26392_ (.A1(net3194),
    .A2(_17538_),
    .B(net2889),
    .Y(_17880_));
 NOR2x2_ASAP7_75t_R _26393_ (.A(net1816),
    .B(net2890),
    .Y(_17881_));
 NOR3x2_ASAP7_75t_R _26394_ (.B(_17880_),
    .C(_17881_),
    .Y(_17882_),
    .A(_17879_));
 NOR2x1_ASAP7_75t_R _26395_ (.A(_17657_),
    .B(_17626_),
    .Y(_17883_));
 AOI211x1_ASAP7_75t_R _26396_ (.A1(net1123),
    .A2(net1185),
    .B(_17657_),
    .C(_17557_),
    .Y(_17884_));
 NOR2x2_ASAP7_75t_R _26397_ (.A(_17883_),
    .B(_17884_),
    .Y(_17885_));
 INVx1_ASAP7_75t_R _26398_ (.A(_17586_),
    .Y(_17886_));
 NOR2x2_ASAP7_75t_R _26399_ (.A(_17834_),
    .B(_17657_),
    .Y(_17887_));
 NOR2x1_ASAP7_75t_R _26400_ (.A(_17582_),
    .B(_17657_),
    .Y(_17888_));
 AOI211x1_ASAP7_75t_R _26401_ (.A1(_17886_),
    .A2(_17662_),
    .B(_17887_),
    .C(_17888_),
    .Y(_17889_));
 NAND3x2_ASAP7_75t_R _26402_ (.B(_17885_),
    .C(_17889_),
    .Y(_17890_),
    .A(_17882_));
 AOI211x1_ASAP7_75t_R _26403_ (.A1(net2907),
    .A2(net2891),
    .B(_17641_),
    .C(net1103),
    .Y(_17891_));
 NAND2x2_ASAP7_75t_R _26404_ (.A(net2770),
    .B(net1003),
    .Y(_17892_));
 AOI21x1_ASAP7_75t_R _26405_ (.A1(_17892_),
    .A2(net2532),
    .B(net2484),
    .Y(_17893_));
 NOR2x2_ASAP7_75t_R _26406_ (.A(_17641_),
    .B(_17562_),
    .Y(_17894_));
 NOR3x2_ASAP7_75t_R _26407_ (.B(_17893_),
    .C(_17894_),
    .Y(_17895_),
    .A(_17891_));
 AOI211x1_ASAP7_75t_R _26408_ (.A1(net2862),
    .A2(_17533_),
    .B(net1103),
    .C(_17629_),
    .Y(_17896_));
 AOI211x1_ASAP7_75t_R _26409_ (.A1(net1123),
    .A2(net1187),
    .B(net1974),
    .C(_17629_),
    .Y(_17897_));
 NOR2x2_ASAP7_75t_R _26410_ (.A(_17896_),
    .B(_17897_),
    .Y(_17898_));
 AO21x1_ASAP7_75t_R _26411_ (.A1(_17639_),
    .A2(_17647_),
    .B(_17629_),
    .Y(_17899_));
 AO21x1_ASAP7_75t_R _26412_ (.A1(_17813_),
    .A2(_17551_),
    .B(_17629_),
    .Y(_17900_));
 AND2x2_ASAP7_75t_R _26413_ (.A(_17899_),
    .B(_17900_),
    .Y(_17901_));
 NAND3x2_ASAP7_75t_R _26414_ (.B(_17898_),
    .C(_17901_),
    .Y(_17902_),
    .A(_17895_));
 NOR2x2_ASAP7_75t_R _26415_ (.A(_17890_),
    .B(_17902_),
    .Y(_17903_));
 NAND2x2_ASAP7_75t_R _26416_ (.A(_17877_),
    .B(_17903_),
    .Y(_17904_));
 NOR2x2_ASAP7_75t_R _26417_ (.A(_17853_),
    .B(_17904_),
    .Y(_17905_));
 OAI21x1_ASAP7_75t_R _26418_ (.A1(_17669_),
    .A2(_17535_),
    .B(_17700_),
    .Y(_17906_));
 NAND2x2_ASAP7_75t_R _26419_ (.A(net1008),
    .B(net3086),
    .Y(_17907_));
 NAND2x2_ASAP7_75t_R _26420_ (.A(net3085),
    .B(_17731_),
    .Y(_17908_));
 NAND3x2_ASAP7_75t_R _26421_ (.B(_17907_),
    .C(_17908_),
    .Y(_17909_),
    .A(_17906_));
 AO21x2_ASAP7_75t_R _26422_ (.A1(_17685_),
    .A2(_17563_),
    .B(_17701_),
    .Y(_17910_));
 OAI21x1_ASAP7_75t_R _26423_ (.A1(_17558_),
    .A2(_17676_),
    .B(_17700_),
    .Y(_17911_));
 OAI21x1_ASAP7_75t_R _26424_ (.A1(_17694_),
    .A2(_17616_),
    .B(_17700_),
    .Y(_17912_));
 NAND3x2_ASAP7_75t_R _26425_ (.B(_17911_),
    .C(_17912_),
    .Y(_17913_),
    .A(_17910_));
 NOR2x2_ASAP7_75t_R _26426_ (.A(_17909_),
    .B(_17913_),
    .Y(_17914_));
 OR3x2_ASAP7_75t_R _26427_ (.A(_17602_),
    .B(_17545_),
    .C(_00555_),
    .Y(_17915_));
 NAND3x2_ASAP7_75t_R _26428_ (.B(net3089),
    .C(_17915_),
    .Y(_17916_),
    .A(_17914_));
 NOR2x1_ASAP7_75t_R _26429_ (.A(_17743_),
    .B(_17916_),
    .Y(_17917_));
 NAND2x2_ASAP7_75t_R _26430_ (.A(_00553_),
    .B(_17917_),
    .Y(_17918_));
 NAND3x2_ASAP7_75t_R _26431_ (.B(_17905_),
    .C(_17918_),
    .Y(_17919_),
    .A(_17796_));
 NOR2x2_ASAP7_75t_R _26432_ (.A(_17905_),
    .B(_17796_),
    .Y(_17920_));
 INVx2_ASAP7_75t_R _26433_ (.A(_17920_),
    .Y(_17921_));
 BUFx2_ASAP7_75t_R input194 (.A(net3679),
    .Y(net194));
 INVx6_ASAP7_75t_R _26435_ (.A(net1956),
    .Y(_17923_));
 NAND2x2_ASAP7_75t_R _26436_ (.A(net2155),
    .B(_17923_),
    .Y(_17924_));
 NOR2x2_ASAP7_75t_R _26437_ (.A(net1060),
    .B(net1365),
    .Y(_17925_));
 BUFx2_ASAP7_75t_R input193 (.A(net3691),
    .Y(net193));
 BUFx2_ASAP7_75t_R input192 (.A(net3992),
    .Y(net192));
 AND2x6_ASAP7_75t_R _26440_ (.A(_00641_),
    .B(_00642_),
    .Y(_17928_));
 BUFx2_ASAP7_75t_R input191 (.A(net3718),
    .Y(net191));
 AND2x4_ASAP7_75t_R _26442_ (.A(net2797),
    .B(net3179),
    .Y(_17930_));
 NAND2x2_ASAP7_75t_R _26443_ (.A(_17928_),
    .B(_17930_),
    .Y(_17931_));
 INVx3_ASAP7_75t_R _26444_ (.A(_17931_),
    .Y(_17932_));
 INVx2_ASAP7_75t_R _26445_ (.A(net2154),
    .Y(_17933_));
 NOR2x2_ASAP7_75t_R _26446_ (.A(net1957),
    .B(_17933_),
    .Y(_17934_));
 BUFx2_ASAP7_75t_R input190 (.A(net3739),
    .Y(net190));
 NAND2x2_ASAP7_75t_R _26448_ (.A(net1058),
    .B(net1643),
    .Y(_17936_));
 CKINVDCx9p33_ASAP7_75t_R _26449_ (.A(_17936_),
    .Y(_17937_));
 NAND2x2_ASAP7_75t_R _26450_ (.A(net1790),
    .B(_17937_),
    .Y(_17938_));
 BUFx2_ASAP7_75t_R input189 (.A(net4028),
    .Y(net189));
 BUFx2_ASAP7_75t_R input188 (.A(net3975),
    .Y(net188));
 CKINVDCx20_ASAP7_75t_R _26453_ (.A(net1064),
    .Y(_17941_));
 NOR2x2_ASAP7_75t_R _26454_ (.A(net1643),
    .B(_17941_),
    .Y(_17942_));
 NAND2x2_ASAP7_75t_R _26455_ (.A(net1790),
    .B(_17942_),
    .Y(_17943_));
 BUFx2_ASAP7_75t_R input187 (.A(net3638),
    .Y(net187));
 AOI21x1_ASAP7_75t_R _26457_ (.A1(_17938_),
    .A2(net3307),
    .B(_17931_),
    .Y(_17945_));
 NOR2x2_ASAP7_75t_R _26458_ (.A(net1956),
    .B(net2154),
    .Y(_17946_));
 CKINVDCx20_ASAP7_75t_R _26459_ (.A(net1235),
    .Y(_17947_));
 NOR2x2_ASAP7_75t_R _26460_ (.A(_17947_),
    .B(_17931_),
    .Y(_17948_));
 AOI211x1_ASAP7_75t_R _26461_ (.A1(_17925_),
    .A2(_17932_),
    .B(_17945_),
    .C(_17948_),
    .Y(_17949_));
 BUFx2_ASAP7_75t_R input186 (.A(net3733),
    .Y(net186));
 NAND2x2_ASAP7_75t_R _26463_ (.A(net1956),
    .B(_17933_),
    .Y(_17951_));
 NOR2x2_ASAP7_75t_R _26464_ (.A(_17941_),
    .B(_17951_),
    .Y(_17952_));
 INVx13_ASAP7_75t_R _26465_ (.A(net1647),
    .Y(_17953_));
 NOR2x2_ASAP7_75t_R _26466_ (.A(net1058),
    .B(_17953_),
    .Y(_17954_));
 NOR2x2_ASAP7_75t_R _26467_ (.A(net2154),
    .B(_17923_),
    .Y(_17955_));
 NAND2x2_ASAP7_75t_R _26468_ (.A(_17954_),
    .B(_17955_),
    .Y(_17956_));
 NOR2x2_ASAP7_75t_R _26469_ (.A(net1058),
    .B(net1643),
    .Y(_17957_));
 NAND2x2_ASAP7_75t_R _26470_ (.A(_17957_),
    .B(_17955_),
    .Y(_17958_));
 AOI21x1_ASAP7_75t_R _26471_ (.A1(net2944),
    .A2(_17958_),
    .B(_17931_),
    .Y(_17959_));
 NAND2x2_ASAP7_75t_R _26472_ (.A(net1956),
    .B(net2154),
    .Y(_17960_));
 CKINVDCx11_ASAP7_75t_R _26473_ (.A(net1070),
    .Y(_17961_));
 NAND2x2_ASAP7_75t_R _26474_ (.A(_17941_),
    .B(_17961_),
    .Y(_17962_));
 NAND2x2_ASAP7_75t_R _26475_ (.A(_17942_),
    .B(_17961_),
    .Y(_17963_));
 AOI21x1_ASAP7_75t_R _26476_ (.A1(_17962_),
    .A2(_17963_),
    .B(_17931_),
    .Y(_17964_));
 AOI211x1_ASAP7_75t_R _26477_ (.A1(_17932_),
    .A2(_17952_),
    .B(_17959_),
    .C(_17964_),
    .Y(_17965_));
 INVx3_ASAP7_75t_R _26478_ (.A(net2797),
    .Y(_17966_));
 NOR2x2_ASAP7_75t_R _26479_ (.A(net3179),
    .B(_17966_),
    .Y(_17967_));
 NAND2x2_ASAP7_75t_R _26480_ (.A(_17967_),
    .B(_17928_),
    .Y(_17968_));
 BUFx2_ASAP7_75t_R input185 (.A(net3715),
    .Y(net185));
 INVx5_ASAP7_75t_R _26482_ (.A(net2019),
    .Y(_17970_));
 INVx2_ASAP7_75t_R _26483_ (.A(_00642_),
    .Y(_17971_));
 OR3x1_ASAP7_75t_R _26484_ (.A(_17970_),
    .B(_17971_),
    .C(net2797),
    .Y(_17972_));
 AND4x2_ASAP7_75t_R _26485_ (.A(_17949_),
    .B(_17965_),
    .C(_17968_),
    .D(_17972_),
    .Y(_17973_));
 NAND3x2_ASAP7_75t_R _26486_ (.B(net2018),
    .C(net2749),
    .Y(_17974_),
    .A(_17973_));
 NOR2x2_ASAP7_75t_R _26487_ (.A(net2797),
    .B(net3179),
    .Y(_17975_));
 NOR2x2_ASAP7_75t_R _26488_ (.A(net2019),
    .B(_17971_),
    .Y(_17976_));
 NAND2x2_ASAP7_75t_R _26489_ (.A(_17975_),
    .B(_17976_),
    .Y(_17977_));
 BUFx2_ASAP7_75t_R input184 (.A(net3748),
    .Y(net184));
 BUFx2_ASAP7_75t_R input183 (.A(net3772),
    .Y(net183));
 NAND2x2_ASAP7_75t_R _26492_ (.A(net1235),
    .B(_17937_),
    .Y(_17980_));
 BUFx2_ASAP7_75t_R input182 (.A(net3778),
    .Y(net182));
 NOR2x1_ASAP7_75t_R _26494_ (.A(net1955),
    .B(net3224),
    .Y(_17982_));
 NAND2x2_ASAP7_75t_R _26495_ (.A(net1058),
    .B(_17953_),
    .Y(_17983_));
 NAND2x2_ASAP7_75t_R _26496_ (.A(_17983_),
    .B(_17961_),
    .Y(_17984_));
 NOR2x1_ASAP7_75t_R _26497_ (.A(_17977_),
    .B(_17984_),
    .Y(_17985_));
 INVx1_ASAP7_75t_R _26498_ (.A(_17985_),
    .Y(_17986_));
 NAND2x2_ASAP7_75t_R _26499_ (.A(net1063),
    .B(net2725),
    .Y(_17987_));
 BUFx2_ASAP7_75t_R input181 (.A(net3757),
    .Y(net181));
 BUFx2_ASAP7_75t_R input180 (.A(net3933),
    .Y(net180));
 AO21x1_ASAP7_75t_R _26502_ (.A1(_17987_),
    .A2(net1622),
    .B(_17977_),
    .Y(_17990_));
 NAND2x1_ASAP7_75t_R _26503_ (.A(_17986_),
    .B(_17990_),
    .Y(_17991_));
 NOR2x1_ASAP7_75t_R _26504_ (.A(_17982_),
    .B(_17991_),
    .Y(_17992_));
 NAND2x2_ASAP7_75t_R _26505_ (.A(net3197),
    .B(_17937_),
    .Y(_17993_));
 BUFx2_ASAP7_75t_R input179 (.A(net3799),
    .Y(net179));
 INVx2_ASAP7_75t_R _26507_ (.A(net3179),
    .Y(_17995_));
 NOR2x2_ASAP7_75t_R _26508_ (.A(net2797),
    .B(_17995_),
    .Y(_17996_));
 NAND2x2_ASAP7_75t_R _26509_ (.A(_17976_),
    .B(_17996_),
    .Y(_17997_));
 BUFx2_ASAP7_75t_R input178 (.A(net3927),
    .Y(net178));
 NAND2x2_ASAP7_75t_R _26511_ (.A(net1232),
    .B(_17957_),
    .Y(_17999_));
 INVx6_ASAP7_75t_R _26512_ (.A(_17999_),
    .Y(_18000_));
 BUFx2_ASAP7_75t_R input177 (.A(net3766),
    .Y(net177));
 NAND2x2_ASAP7_75t_R _26514_ (.A(net3204),
    .B(net1236),
    .Y(_18002_));
 NAND2x1_ASAP7_75t_R _26515_ (.A(_18002_),
    .B(net1690),
    .Y(_18003_));
 NAND2x2_ASAP7_75t_R _26516_ (.A(net2750),
    .B(_17970_),
    .Y(_18004_));
 NAND2x2_ASAP7_75t_R _26517_ (.A(net3179),
    .B(_17966_),
    .Y(_18005_));
 NOR2x2_ASAP7_75t_R _26518_ (.A(_18004_),
    .B(_18005_),
    .Y(_18006_));
 OAI21x1_ASAP7_75t_R _26519_ (.A1(_18000_),
    .A2(_18003_),
    .B(_18006_),
    .Y(_18007_));
 OA21x2_ASAP7_75t_R _26520_ (.A1(net2908),
    .A2(_17997_),
    .B(_18007_),
    .Y(_18008_));
 NAND2x1_ASAP7_75t_R _26521_ (.A(_17992_),
    .B(_18008_),
    .Y(_18009_));
 NAND2x2_ASAP7_75t_R _26522_ (.A(_17954_),
    .B(_17961_),
    .Y(_18010_));
 BUFx2_ASAP7_75t_R input176 (.A(net3951),
    .Y(net176));
 NAND2x2_ASAP7_75t_R _26524_ (.A(_17976_),
    .B(_17967_),
    .Y(_18012_));
 AO21x1_ASAP7_75t_R _26525_ (.A1(_18010_),
    .A2(net1531),
    .B(net3216),
    .Y(_18013_));
 NAND2x2_ASAP7_75t_R _26526_ (.A(net1234),
    .B(_17954_),
    .Y(_18014_));
 BUFx2_ASAP7_75t_R input175 (.A(net3869),
    .Y(net175));
 BUFx2_ASAP7_75t_R input174 (.A(net3685),
    .Y(net174));
 AO21x1_ASAP7_75t_R _26529_ (.A1(net1121),
    .A2(net1068),
    .B(net3216),
    .Y(_18017_));
 AND2x2_ASAP7_75t_R _26530_ (.A(_18013_),
    .B(_18017_),
    .Y(_18018_));
 NAND2x2_ASAP7_75t_R _26531_ (.A(net2797),
    .B(net3179),
    .Y(_18019_));
 NOR2x2_ASAP7_75t_R _26532_ (.A(_18019_),
    .B(_18004_),
    .Y(_18020_));
 NAND2x1_ASAP7_75t_R _26533_ (.A(net1235),
    .B(net3196),
    .Y(_18021_));
 NAND2x2_ASAP7_75t_R _26534_ (.A(_17957_),
    .B(net1790),
    .Y(_18022_));
 BUFx2_ASAP7_75t_R input173 (.A(net3576),
    .Y(net173));
 NAND2x2_ASAP7_75t_R _26536_ (.A(_17976_),
    .B(_17930_),
    .Y(_18024_));
 AO21x1_ASAP7_75t_R _26537_ (.A1(net1692),
    .A2(_18022_),
    .B(_18024_),
    .Y(_18025_));
 OAI21x1_ASAP7_75t_R _26538_ (.A1(_17937_),
    .A2(_18021_),
    .B(_18025_),
    .Y(_18026_));
 NAND2x2_ASAP7_75t_R _26539_ (.A(net3198),
    .B(net3196),
    .Y(_18027_));
 NAND2x2_ASAP7_75t_R _26540_ (.A(_17961_),
    .B(_17937_),
    .Y(_18028_));
 BUFx2_ASAP7_75t_R input172 (.A(net3709),
    .Y(net172));
 AO21x1_ASAP7_75t_R _26542_ (.A1(_18028_),
    .A2(_18010_),
    .B(_18024_),
    .Y(_18030_));
 OAI21x1_ASAP7_75t_R _26543_ (.A1(_17954_),
    .A2(_18027_),
    .B(_18030_),
    .Y(_18031_));
 NOR2x1_ASAP7_75t_R _26544_ (.A(_18026_),
    .B(_18031_),
    .Y(_18032_));
 NAND2x1_ASAP7_75t_R _26545_ (.A(_18018_),
    .B(_18032_),
    .Y(_18033_));
 NOR2x1_ASAP7_75t_R _26546_ (.A(_18009_),
    .B(_18033_),
    .Y(_18034_));
 BUFx2_ASAP7_75t_R input171 (.A(net3721),
    .Y(net171));
 NAND2x2_ASAP7_75t_R _26548_ (.A(net1643),
    .B(_17941_),
    .Y(_18036_));
 NOR2x2_ASAP7_75t_R _26549_ (.A(net1072),
    .B(_18036_),
    .Y(_18037_));
 NOR2x2_ASAP7_75t_R _26550_ (.A(_00641_),
    .B(_00642_),
    .Y(_18038_));
 NAND2x2_ASAP7_75t_R _26551_ (.A(_18038_),
    .B(_17930_),
    .Y(_18039_));
 INVx5_ASAP7_75t_R _26552_ (.A(net3304),
    .Y(_18040_));
 BUFx2_ASAP7_75t_R input170 (.A(net3866),
    .Y(net170));
 BUFx2_ASAP7_75t_R input169 (.A(net3751),
    .Y(net169));
 BUFx2_ASAP7_75t_R input168 (.A(net3730),
    .Y(net168));
 BUFx2_ASAP7_75t_R input167 (.A(net3664),
    .Y(net167));
 AOI211x1_ASAP7_75t_R _26557_ (.A1(net3201),
    .A2(net3124),
    .B(net3303),
    .C(net3284),
    .Y(_18045_));
 INVx4_ASAP7_75t_R _26558_ (.A(_17957_),
    .Y(_18046_));
 NOR2x2_ASAP7_75t_R _26559_ (.A(net1366),
    .B(_18046_),
    .Y(_18047_));
 NOR2x2_ASAP7_75t_R _26560_ (.A(net1365),
    .B(_17983_),
    .Y(_18048_));
 OA21x2_ASAP7_75t_R _26561_ (.A1(net3218),
    .A2(_18048_),
    .B(_18040_),
    .Y(_18049_));
 AOI211x1_ASAP7_75t_R _26562_ (.A1(_18037_),
    .A2(_18040_),
    .B(_18045_),
    .C(_18049_),
    .Y(_18050_));
 BUFx2_ASAP7_75t_R input166 (.A(net3712),
    .Y(net166));
 NAND2x2_ASAP7_75t_R _26564_ (.A(_17942_),
    .B(_17955_),
    .Y(_18052_));
 BUFx2_ASAP7_75t_R input165 (.A(net3724),
    .Y(net165));
 NAND2x2_ASAP7_75t_R _26566_ (.A(_18038_),
    .B(_17967_),
    .Y(_18054_));
 BUFx2_ASAP7_75t_R input164 (.A(net3736),
    .Y(net164));
 AO21x1_ASAP7_75t_R _26568_ (.A1(_18010_),
    .A2(net1795),
    .B(_18054_),
    .Y(_18056_));
 NAND2x2_ASAP7_75t_R _26569_ (.A(net1233),
    .B(_17942_),
    .Y(_18057_));
 BUFx2_ASAP7_75t_R input163 (.A(net3754),
    .Y(net163));
 AO21x1_ASAP7_75t_R _26571_ (.A1(net3191),
    .A2(_18057_),
    .B(_18054_),
    .Y(_18059_));
 BUFx2_ASAP7_75t_R input162 (.A(net3700),
    .Y(net162));
 NOR2x1_ASAP7_75t_R _26573_ (.A(net1367),
    .B(_18054_),
    .Y(_18061_));
 INVx1_ASAP7_75t_R _26574_ (.A(_18061_),
    .Y(_18062_));
 AND3x1_ASAP7_75t_R _26575_ (.A(_18056_),
    .B(_18059_),
    .C(_18062_),
    .Y(_18063_));
 NAND2x1_ASAP7_75t_R _26576_ (.A(_18050_),
    .B(_18063_),
    .Y(_18064_));
 NAND2x2_ASAP7_75t_R _26577_ (.A(_17975_),
    .B(_18038_),
    .Y(_18065_));
 BUFx2_ASAP7_75t_R input161 (.A(net3823),
    .Y(net161));
 AO21x1_ASAP7_75t_R _26579_ (.A1(net1532),
    .A2(_17962_),
    .B(net1909),
    .Y(_18067_));
 AO21x1_ASAP7_75t_R _26580_ (.A1(net3191),
    .A2(net1369),
    .B(net1909),
    .Y(_18068_));
 INVx4_ASAP7_75t_R _26581_ (.A(_18065_),
    .Y(_18069_));
 INVx3_ASAP7_75t_R _26582_ (.A(net3186),
    .Y(_18070_));
 NAND2x1_ASAP7_75t_R _26583_ (.A(_18069_),
    .B(_18070_),
    .Y(_18071_));
 AND3x1_ASAP7_75t_R _26584_ (.A(_18067_),
    .B(_18068_),
    .C(_18071_),
    .Y(_18072_));
 NAND2x2_ASAP7_75t_R _26585_ (.A(_17941_),
    .B(net1790),
    .Y(_18073_));
 NAND2x2_ASAP7_75t_R _26586_ (.A(_18038_),
    .B(_17996_),
    .Y(_18074_));
 BUFx2_ASAP7_75t_R input160 (.A(net3829),
    .Y(net160));
 AOI21x1_ASAP7_75t_R _26588_ (.A1(_18073_),
    .A2(_17938_),
    .B(_18074_),
    .Y(_18076_));
 INVx1_ASAP7_75t_R _26589_ (.A(_18076_),
    .Y(_18077_));
 AO21x1_ASAP7_75t_R _26590_ (.A1(_18057_),
    .A2(net1068),
    .B(_18074_),
    .Y(_18078_));
 NAND2x1_ASAP7_75t_R _26591_ (.A(_18077_),
    .B(_18078_),
    .Y(_18079_));
 BUFx2_ASAP7_75t_R input159 (.A(net3909),
    .Y(net159));
 NAND2x2_ASAP7_75t_R _26593_ (.A(net3206),
    .B(_17961_),
    .Y(_18081_));
 BUFx2_ASAP7_75t_R input158 (.A(net3784),
    .Y(net158));
 AO21x1_ASAP7_75t_R _26595_ (.A1(net3300),
    .A2(net2757),
    .B(_18074_),
    .Y(_18083_));
 OAI21x1_ASAP7_75t_R _26596_ (.A1(net2181),
    .A2(_17987_),
    .B(_18083_),
    .Y(_18084_));
 NOR2x1_ASAP7_75t_R _26597_ (.A(_18079_),
    .B(_18084_),
    .Y(_18085_));
 NAND2x1_ASAP7_75t_R _26598_ (.A(_18072_),
    .B(_18085_),
    .Y(_18086_));
 NOR2x1_ASAP7_75t_R _26599_ (.A(_18064_),
    .B(_18086_),
    .Y(_18087_));
 NAND2x2_ASAP7_75t_R _26600_ (.A(_18034_),
    .B(_18087_),
    .Y(_18088_));
 INVx1_ASAP7_75t_R _26601_ (.A(_17968_),
    .Y(_18089_));
 INVx2_ASAP7_75t_R _26602_ (.A(_17962_),
    .Y(_18090_));
 BUFx2_ASAP7_75t_R input157 (.A(net3820),
    .Y(net157));
 BUFx2_ASAP7_75t_R input156 (.A(net3760),
    .Y(net156));
 AOI21x1_ASAP7_75t_R _26605_ (.A1(net1795),
    .A2(net939),
    .B(net2364),
    .Y(_18093_));
 BUFx2_ASAP7_75t_R input155 (.A(net3851),
    .Y(net155));
 AOI21x1_ASAP7_75t_R _26607_ (.A1(_18022_),
    .A2(_17938_),
    .B(_17968_),
    .Y(_18095_));
 AOI211x1_ASAP7_75t_R _26608_ (.A1(_18089_),
    .A2(_18090_),
    .B(_18093_),
    .C(_18095_),
    .Y(_18096_));
 BUFx2_ASAP7_75t_R input154 (.A(net3886),
    .Y(net154));
 NOR2x1_ASAP7_75t_R _26610_ (.A(_17962_),
    .B(_17931_),
    .Y(_18098_));
 NOR2x1_ASAP7_75t_R _26611_ (.A(net3185),
    .B(net1746),
    .Y(_18099_));
 NOR3x1_ASAP7_75t_R _26612_ (.A(_17959_),
    .B(_18098_),
    .C(_18099_),
    .Y(_18100_));
 AO21x1_ASAP7_75t_R _26613_ (.A1(net3307),
    .A2(_18073_),
    .B(net1746),
    .Y(_18101_));
 AO21x1_ASAP7_75t_R _26614_ (.A1(net1121),
    .A2(_18057_),
    .B(net1746),
    .Y(_18102_));
 AND2x2_ASAP7_75t_R _26615_ (.A(_18101_),
    .B(_18102_),
    .Y(_18103_));
 NAND3x1_ASAP7_75t_R _26616_ (.A(_18096_),
    .B(_18100_),
    .C(_18103_),
    .Y(_18104_));
 NOR2x2_ASAP7_75t_R _26617_ (.A(_17941_),
    .B(net1070),
    .Y(_18105_));
 NAND2x2_ASAP7_75t_R _26618_ (.A(net2019),
    .B(net2751),
    .Y(_18106_));
 NOR2x2_ASAP7_75t_R _26619_ (.A(_18106_),
    .B(_18005_),
    .Y(_18107_));
 OAI21x1_ASAP7_75t_R _26620_ (.A1(_18105_),
    .A2(_18037_),
    .B(_18107_),
    .Y(_18108_));
 BUFx2_ASAP7_75t_R input153 (.A(net3763),
    .Y(net153));
 NOR2x2_ASAP7_75t_R _26622_ (.A(_17983_),
    .B(_17951_),
    .Y(_18110_));
 NAND2x1_ASAP7_75t_R _26623_ (.A(net2165),
    .B(_18110_),
    .Y(_18111_));
 BUFx2_ASAP7_75t_R input152 (.A(net3978),
    .Y(net152));
 NOR2x2_ASAP7_75t_R _26625_ (.A(_18036_),
    .B(_17951_),
    .Y(_18113_));
 NAND2x1_ASAP7_75t_R _26626_ (.A(net2165),
    .B(_18113_),
    .Y(_18114_));
 NAND3x1_ASAP7_75t_R _26627_ (.A(net3221),
    .B(_18111_),
    .C(_18114_),
    .Y(_18115_));
 OAI21x1_ASAP7_75t_R _26628_ (.A1(_17925_),
    .A2(_18048_),
    .B(_18107_),
    .Y(_18116_));
 BUFx2_ASAP7_75t_R input151 (.A(net4093),
    .Y(net151));
 NOR3x2_ASAP7_75t_R _26630_ (.B(_18005_),
    .C(_18106_),
    .Y(_18118_),
    .A(net3285));
 OAI21x1_ASAP7_75t_R _26631_ (.A1(net3201),
    .A2(net1117),
    .B(_18118_),
    .Y(_18119_));
 NAND2x1_ASAP7_75t_R _26632_ (.A(net3223),
    .B(_18119_),
    .Y(_18120_));
 NOR2x1_ASAP7_75t_R _26633_ (.A(_18115_),
    .B(_18120_),
    .Y(_18121_));
 NAND2x2_ASAP7_75t_R _26634_ (.A(_17966_),
    .B(_17995_),
    .Y(_18122_));
 NOR2x2_ASAP7_75t_R _26635_ (.A(_18106_),
    .B(_18122_),
    .Y(_18123_));
 BUFx2_ASAP7_75t_R input150 (.A(net3972),
    .Y(net150));
 NAND2x1_ASAP7_75t_R _26637_ (.A(_18113_),
    .B(_18123_),
    .Y(_18125_));
 NAND2x2_ASAP7_75t_R _26638_ (.A(_17975_),
    .B(_17928_),
    .Y(_18126_));
 NOR2x1_ASAP7_75t_R _26639_ (.A(net1075),
    .B(_18126_),
    .Y(_18127_));
 OAI21x1_ASAP7_75t_R _26640_ (.A1(net3201),
    .A2(net3308),
    .B(_18127_),
    .Y(_18128_));
 NAND2x1_ASAP7_75t_R _26641_ (.A(_18125_),
    .B(_18128_),
    .Y(_18129_));
 NOR2x2_ASAP7_75t_R _26642_ (.A(net1543),
    .B(_17947_),
    .Y(_18130_));
 NOR2x2_ASAP7_75t_R _26643_ (.A(_17983_),
    .B(_17947_),
    .Y(_18131_));
 BUFx2_ASAP7_75t_R input149 (.A(net3995),
    .Y(net149));
 OAI21x1_ASAP7_75t_R _26645_ (.A1(_18130_),
    .A2(net3207),
    .B(_18123_),
    .Y(_18133_));
 NOR2x2_ASAP7_75t_R _26646_ (.A(_17936_),
    .B(net1365),
    .Y(_18134_));
 NAND2x1_ASAP7_75t_R _26647_ (.A(_18134_),
    .B(_18123_),
    .Y(_18135_));
 NAND2x1_ASAP7_75t_R _26648_ (.A(_18123_),
    .B(_18000_),
    .Y(_18136_));
 NAND3x1_ASAP7_75t_R _26649_ (.A(_18133_),
    .B(_18135_),
    .C(_18136_),
    .Y(_18137_));
 NOR2x1_ASAP7_75t_R _26650_ (.A(_18129_),
    .B(_18137_),
    .Y(_18138_));
 NAND2x1_ASAP7_75t_R _26651_ (.A(_18121_),
    .B(_18138_),
    .Y(_18139_));
 NOR2x1_ASAP7_75t_R _26652_ (.A(_18104_),
    .B(_18139_),
    .Y(_18140_));
 BUFx2_ASAP7_75t_R input148 (.A(net3945),
    .Y(net148));
 BUFx2_ASAP7_75t_R input147 (.A(net3930),
    .Y(net147));
 NOR2x2_ASAP7_75t_R _26655_ (.A(net2750),
    .B(_17970_),
    .Y(_18143_));
 NAND2x2_ASAP7_75t_R _26656_ (.A(_17967_),
    .B(_18143_),
    .Y(_18144_));
 BUFx2_ASAP7_75t_R input146 (.A(net3802),
    .Y(net146));
 AO21x1_ASAP7_75t_R _26658_ (.A1(_17956_),
    .A2(net1622),
    .B(_18144_),
    .Y(_18146_));
 INVx6_ASAP7_75t_R _26659_ (.A(_18105_),
    .Y(_18147_));
 BUFx2_ASAP7_75t_R input145 (.A(net3781),
    .Y(net145));
 AO21x2_ASAP7_75t_R _26661_ (.A1(_18147_),
    .A2(_18081_),
    .B(net2432),
    .Y(_18149_));
 NOR2x2_ASAP7_75t_R _26662_ (.A(net1646),
    .B(net1370),
    .Y(_18150_));
 INVx4_ASAP7_75t_R _26663_ (.A(_18144_),
    .Y(_18151_));
 OAI21x1_ASAP7_75t_R _26664_ (.A1(_18000_),
    .A2(_18150_),
    .B(_18151_),
    .Y(_18152_));
 AND3x1_ASAP7_75t_R _26665_ (.A(_18146_),
    .B(_18149_),
    .C(_18152_),
    .Y(_18153_));
 NAND2x2_ASAP7_75t_R _26666_ (.A(net2019),
    .B(_17971_),
    .Y(_18154_));
 NOR2x2_ASAP7_75t_R _26667_ (.A(_18019_),
    .B(_18154_),
    .Y(_18155_));
 INVx3_ASAP7_75t_R _26668_ (.A(_18155_),
    .Y(_18156_));
 AO21x1_ASAP7_75t_R _26669_ (.A1(_18147_),
    .A2(net2908),
    .B(_18156_),
    .Y(_18157_));
 NOR2x2_ASAP7_75t_R _26670_ (.A(net2719),
    .B(_17947_),
    .Y(_18158_));
 BUFx2_ASAP7_75t_R input144 (.A(net3808),
    .Y(net144));
 OAI21x1_ASAP7_75t_R _26672_ (.A1(_18158_),
    .A2(net3207),
    .B(net2163),
    .Y(_18160_));
 OAI21x1_ASAP7_75t_R _26673_ (.A1(_18150_),
    .A2(net3367),
    .B(net2164),
    .Y(_18161_));
 AND3x1_ASAP7_75t_R _26674_ (.A(_18157_),
    .B(_18160_),
    .C(_18161_),
    .Y(_18162_));
 NAND2x1_ASAP7_75t_R _26675_ (.A(_18153_),
    .B(_18162_),
    .Y(_18163_));
 NOR2x2_ASAP7_75t_R _26676_ (.A(net2848),
    .B(net2853),
    .Y(_18164_));
 NOR2x2_ASAP7_75t_R _26677_ (.A(_18154_),
    .B(_18122_),
    .Y(_18165_));
 NAND2x2_ASAP7_75t_R _26678_ (.A(net1230),
    .B(_18165_),
    .Y(_18166_));
 NAND2x1_ASAP7_75t_R _26679_ (.A(_18165_),
    .B(_18047_),
    .Y(_18167_));
 OAI21x1_ASAP7_75t_R _26680_ (.A1(_18164_),
    .A2(_18166_),
    .B(_18167_),
    .Y(_18168_));
 NAND2x2_ASAP7_75t_R _26681_ (.A(_17975_),
    .B(_18143_),
    .Y(_18169_));
 BUFx2_ASAP7_75t_R input143 (.A(net3984),
    .Y(net143));
 AO21x1_ASAP7_75t_R _26683_ (.A1(net3188),
    .A2(net974),
    .B(_18169_),
    .Y(_18171_));
 INVx1_ASAP7_75t_R _26684_ (.A(_18171_),
    .Y(_18172_));
 AOI211x1_ASAP7_75t_R _26685_ (.A1(net3201),
    .A2(net1117),
    .B(_18169_),
    .C(net1070),
    .Y(_18173_));
 NOR3x1_ASAP7_75t_R _26686_ (.A(_18168_),
    .B(_18172_),
    .C(_18173_),
    .Y(_18174_));
 NOR2x2_ASAP7_75t_R _26687_ (.A(_18005_),
    .B(_18154_),
    .Y(_18175_));
 BUFx2_ASAP7_75t_R input142 (.A(net3585),
    .Y(net142));
 NAND2x1_ASAP7_75t_R _26689_ (.A(_17952_),
    .B(net2244),
    .Y(_18177_));
 NOR2x2_ASAP7_75t_R _26690_ (.A(_17951_),
    .B(_18046_),
    .Y(_18178_));
 BUFx2_ASAP7_75t_R input141 (.A(net3883),
    .Y(net141));
 OAI21x1_ASAP7_75t_R _26692_ (.A1(_18113_),
    .A2(_18178_),
    .B(net2246),
    .Y(_18180_));
 NAND2x1_ASAP7_75t_R _26693_ (.A(_18177_),
    .B(_18180_),
    .Y(_18181_));
 NAND2x1_ASAP7_75t_R _26694_ (.A(net2244),
    .B(_18158_),
    .Y(_18182_));
 OAI21x1_ASAP7_75t_R _26695_ (.A1(_18134_),
    .A2(_18150_),
    .B(net2244),
    .Y(_18183_));
 NAND2x1_ASAP7_75t_R _26696_ (.A(_18182_),
    .B(_18183_),
    .Y(_18184_));
 NAND2x2_ASAP7_75t_R _26697_ (.A(_17961_),
    .B(_18175_),
    .Y(_18185_));
 NOR2x1_ASAP7_75t_R _26698_ (.A(net1117),
    .B(_18185_),
    .Y(_18186_));
 NOR3x1_ASAP7_75t_R _26699_ (.A(_18181_),
    .B(_18184_),
    .C(_18186_),
    .Y(_18187_));
 NAND2x1_ASAP7_75t_R _26700_ (.A(_18174_),
    .B(_18187_),
    .Y(_18188_));
 NOR2x1_ASAP7_75t_R _26701_ (.A(_18163_),
    .B(_18188_),
    .Y(_18189_));
 NAND2x1_ASAP7_75t_R _26702_ (.A(_18140_),
    .B(_18189_),
    .Y(_18190_));
 NOR2x2_ASAP7_75t_R _26703_ (.A(_18088_),
    .B(_18190_),
    .Y(_18191_));
 NAND2x2_ASAP7_75t_R _26704_ (.A(net2557),
    .B(_18191_),
    .Y(_18192_));
 INVx2_ASAP7_75t_R _26705_ (.A(_18192_),
    .Y(_18193_));
 AO21x1_ASAP7_75t_R _26706_ (.A1(_17919_),
    .A2(_17921_),
    .B(_18193_),
    .Y(_18194_));
 NOR3x2_ASAP7_75t_R _26707_ (.B(_17682_),
    .C(net2896),
    .Y(_18195_),
    .A(net2897));
 INVx1_ASAP7_75t_R _26708_ (.A(_17698_),
    .Y(_18196_));
 NAND2x1_ASAP7_75t_R _26709_ (.A(_17710_),
    .B(_17706_),
    .Y(_18197_));
 NOR2x1_ASAP7_75t_R _26710_ (.A(_18196_),
    .B(_18197_),
    .Y(_18198_));
 INVx1_ASAP7_75t_R _26711_ (.A(_17730_),
    .Y(_18199_));
 NAND2x1_ASAP7_75t_R _26712_ (.A(_17738_),
    .B(_18199_),
    .Y(_18200_));
 NOR2x1_ASAP7_75t_R _26713_ (.A(_17722_),
    .B(_18200_),
    .Y(_18201_));
 NAND2x1_ASAP7_75t_R _26714_ (.A(_18198_),
    .B(_18201_),
    .Y(_18202_));
 NAND3x1_ASAP7_75t_R _26715_ (.A(_17766_),
    .B(_17792_),
    .C(_17776_),
    .Y(_18203_));
 NOR2x1_ASAP7_75t_R _26716_ (.A(_18202_),
    .B(_18203_),
    .Y(_18204_));
 NAND2x2_ASAP7_75t_R _26717_ (.A(_18195_),
    .B(_18204_),
    .Y(_18205_));
 NOR3x1_ASAP7_75t_R _26718_ (.A(_17837_),
    .B(_17833_),
    .C(_17829_),
    .Y(_18206_));
 NAND2x1_ASAP7_75t_R _26719_ (.A(_17850_),
    .B(_18206_),
    .Y(_18207_));
 INVx1_ASAP7_75t_R _26720_ (.A(_17800_),
    .Y(_18208_));
 NAND2x1_ASAP7_75t_R _26721_ (.A(_17807_),
    .B(_17804_),
    .Y(_18209_));
 NOR2x1_ASAP7_75t_R _26722_ (.A(_18208_),
    .B(_18209_),
    .Y(_18210_));
 INVx1_ASAP7_75t_R _26723_ (.A(_17821_),
    .Y(_18211_));
 NOR2x1_ASAP7_75t_R _26724_ (.A(_17823_),
    .B(_17822_),
    .Y(_18212_));
 NAND2x1_ASAP7_75t_R _26725_ (.A(_18211_),
    .B(_18212_),
    .Y(_18213_));
 INVx1_ASAP7_75t_R _26726_ (.A(_17819_),
    .Y(_18214_));
 NOR2x1_ASAP7_75t_R _26727_ (.A(_18213_),
    .B(_18214_),
    .Y(_18215_));
 NAND2x2_ASAP7_75t_R _26728_ (.A(_18210_),
    .B(_18215_),
    .Y(_18216_));
 NOR2x2_ASAP7_75t_R _26729_ (.A(_18207_),
    .B(_18216_),
    .Y(_18217_));
 INVx1_ASAP7_75t_R _26730_ (.A(_17882_),
    .Y(_18218_));
 NAND2x1_ASAP7_75t_R _26731_ (.A(_17885_),
    .B(_17889_),
    .Y(_18219_));
 NOR2x1_ASAP7_75t_R _26732_ (.A(_18218_),
    .B(_18219_),
    .Y(_18220_));
 INVx1_ASAP7_75t_R _26733_ (.A(_17895_),
    .Y(_18221_));
 NAND2x1_ASAP7_75t_R _26734_ (.A(_17898_),
    .B(_17901_),
    .Y(_18222_));
 NOR2x2_ASAP7_75t_R _26735_ (.A(_18221_),
    .B(_18222_),
    .Y(_18223_));
 NAND2x2_ASAP7_75t_R _26736_ (.A(_18220_),
    .B(_18223_),
    .Y(_18224_));
 INVx1_ASAP7_75t_R _26737_ (.A(_17860_),
    .Y(_18225_));
 NOR2x1_ASAP7_75t_R _26738_ (.A(_17864_),
    .B(_18225_),
    .Y(_18226_));
 NAND2x1_ASAP7_75t_R _26739_ (.A(_17875_),
    .B(_18226_),
    .Y(_18227_));
 NOR2x2_ASAP7_75t_R _26740_ (.A(_18224_),
    .B(_18227_),
    .Y(_18228_));
 NAND2x2_ASAP7_75t_R _26741_ (.A(_18217_),
    .B(_18228_),
    .Y(_18229_));
 NOR3x2_ASAP7_75t_R _26742_ (.B(_17602_),
    .C(_17545_),
    .Y(_18230_),
    .A(_17916_));
 NOR3x2_ASAP7_75t_R _26743_ (.B(_18229_),
    .C(net2143),
    .Y(_18231_),
    .A(_18205_));
 NOR2x2_ASAP7_75t_R _26744_ (.A(_18231_),
    .B(_17920_),
    .Y(_18232_));
 NAND2x1_ASAP7_75t_R _26745_ (.A(_18193_),
    .B(_18232_),
    .Y(_18233_));
 BUFx2_ASAP7_75t_R input140 (.A(net3936),
    .Y(net140));
 NOR2x2_ASAP7_75t_R _26747_ (.A(_00605_),
    .B(_00606_),
    .Y(_18235_));
 BUFx2_ASAP7_75t_R input139 (.A(net3567),
    .Y(net139));
 CKINVDCx16_ASAP7_75t_R _26749_ (.A(net1393),
    .Y(_18237_));
 NOR2x2_ASAP7_75t_R _26750_ (.A(net1680),
    .B(_18237_),
    .Y(_18238_));
 NAND2x2_ASAP7_75t_R _26751_ (.A(_18235_),
    .B(_18238_),
    .Y(_18239_));
 CKINVDCx16_ASAP7_75t_R _26752_ (.A(net1678),
    .Y(_18240_));
 NAND2x2_ASAP7_75t_R _26753_ (.A(net1397),
    .B(_18240_),
    .Y(_18241_));
 NAND2x2_ASAP7_75t_R _26754_ (.A(_18235_),
    .B(_18241_),
    .Y(_18242_));
 NAND2x1_ASAP7_75t_R _26755_ (.A(_00603_),
    .B(_00604_),
    .Y(_18243_));
 BUFx2_ASAP7_75t_R input138 (.A(net3921),
    .Y(net138));
 BUFx2_ASAP7_75t_R input137 (.A(net3832),
    .Y(net137));
 NAND2x1_ASAP7_75t_R _26758_ (.A(net2996),
    .B(_00602_),
    .Y(_18246_));
 NOR2x2_ASAP7_75t_R _26759_ (.A(_18243_),
    .B(_18246_),
    .Y(_18247_));
 INVx4_ASAP7_75t_R _26760_ (.A(_18247_),
    .Y(_18248_));
 AO21x1_ASAP7_75t_R _26761_ (.A1(_18239_),
    .A2(_18242_),
    .B(_18248_),
    .Y(_18249_));
 INVx1_ASAP7_75t_R _26762_ (.A(_18249_),
    .Y(_18250_));
 BUFx2_ASAP7_75t_R input136 (.A(net3895),
    .Y(net136));
 INVx3_ASAP7_75t_R _26764_ (.A(_00605_),
    .Y(_18252_));
 NAND2x2_ASAP7_75t_R _26765_ (.A(net2534),
    .B(_18252_),
    .Y(_18253_));
 NOR2x2_ASAP7_75t_R _26766_ (.A(net1087),
    .B(_18253_),
    .Y(_18254_));
 NAND2x1_ASAP7_75t_R _26767_ (.A(_18247_),
    .B(_18254_),
    .Y(_18255_));
 NAND2x2_ASAP7_75t_R _26768_ (.A(net1678),
    .B(net1395),
    .Y(_18256_));
 NOR2x1_ASAP7_75t_R _26769_ (.A(_18256_),
    .B(_18253_),
    .Y(_18257_));
 NAND2x2_ASAP7_75t_R _26770_ (.A(net1680),
    .B(_18237_),
    .Y(_18258_));
 NOR2x2_ASAP7_75t_R _26771_ (.A(_18253_),
    .B(_18258_),
    .Y(_18259_));
 OAI21x1_ASAP7_75t_R _26772_ (.A1(_18257_),
    .A2(_18259_),
    .B(_18247_),
    .Y(_18260_));
 NAND2x1_ASAP7_75t_R _26773_ (.A(_18255_),
    .B(_18260_),
    .Y(_18261_));
 NOR2x1_ASAP7_75t_R _26774_ (.A(_18250_),
    .B(_18261_),
    .Y(_18262_));
 INVx1_ASAP7_75t_R _26775_ (.A(_00603_),
    .Y(_18263_));
 NOR2x2_ASAP7_75t_R _26776_ (.A(_00604_),
    .B(_18263_),
    .Y(_18264_));
 AND2x4_ASAP7_75t_R _26777_ (.A(net2997),
    .B(_00602_),
    .Y(_18265_));
 NAND2x2_ASAP7_75t_R _26778_ (.A(_18264_),
    .B(_18265_),
    .Y(_18266_));
 BUFx2_ASAP7_75t_R input135 (.A(net3987),
    .Y(net135));
 NAND2x2_ASAP7_75t_R _26780_ (.A(_00605_),
    .B(_00606_),
    .Y(_18268_));
 NOR2x2_ASAP7_75t_R _26781_ (.A(net1679),
    .B(_18268_),
    .Y(_18269_));
 NOR2x2_ASAP7_75t_R _26782_ (.A(net2825),
    .B(_18258_),
    .Y(_18270_));
 OAI21x1_ASAP7_75t_R _26783_ (.A1(_18269_),
    .A2(_18270_),
    .B(_18247_),
    .Y(_18271_));
 NOR2x2_ASAP7_75t_R _26784_ (.A(_00606_),
    .B(_18252_),
    .Y(_18272_));
 NAND2x2_ASAP7_75t_R _26785_ (.A(net1864),
    .B(_18247_),
    .Y(_18273_));
 AND2x4_ASAP7_75t_R _26786_ (.A(_18271_),
    .B(_18273_),
    .Y(_18274_));
 INVx3_ASAP7_75t_R _26787_ (.A(net2996),
    .Y(_18275_));
 INVx3_ASAP7_75t_R _26788_ (.A(_00602_),
    .Y(_18276_));
 OR3x2_ASAP7_75t_R _26789_ (.A(_18275_),
    .B(_18276_),
    .C(_00603_),
    .Y(_18277_));
 AND4x2_ASAP7_75t_R _26790_ (.A(_18262_),
    .B(_18266_),
    .C(_18274_),
    .D(_18277_),
    .Y(_18278_));
 NAND3x2_ASAP7_75t_R _26791_ (.B(net2998),
    .C(_00602_),
    .Y(_18279_),
    .A(_18278_));
 INVx3_ASAP7_75t_R _26792_ (.A(_00606_),
    .Y(_18280_));
 NOR2x2_ASAP7_75t_R _26793_ (.A(_00605_),
    .B(_18280_),
    .Y(_18281_));
 NOR2x2_ASAP7_75t_R _26794_ (.A(net1395),
    .B(_18240_),
    .Y(_18282_));
 NAND2x2_ASAP7_75t_R _26795_ (.A(net2602),
    .B(_18282_),
    .Y(_18283_));
 NOR2x2_ASAP7_75t_R _26796_ (.A(net2996),
    .B(_18276_),
    .Y(_18284_));
 INVx1_ASAP7_75t_R _26797_ (.A(_00604_),
    .Y(_18285_));
 NOR2x2_ASAP7_75t_R _26798_ (.A(_00603_),
    .B(_18285_),
    .Y(_18286_));
 NAND2x2_ASAP7_75t_R _26799_ (.A(_18284_),
    .B(_18286_),
    .Y(_18287_));
 BUFx2_ASAP7_75t_R input134 (.A(net3924),
    .Y(net134));
 AO21x1_ASAP7_75t_R _26801_ (.A1(net2476),
    .A2(net2788),
    .B(_18287_),
    .Y(_18289_));
 NAND2x2_ASAP7_75t_R _26802_ (.A(net2108),
    .B(_18280_),
    .Y(_18290_));
 NOR2x2_ASAP7_75t_R _26803_ (.A(_18256_),
    .B(net2498),
    .Y(_18291_));
 INVx6_ASAP7_75t_R _26804_ (.A(_18287_),
    .Y(_18292_));
 NAND2x1_ASAP7_75t_R _26805_ (.A(_18291_),
    .B(_18292_),
    .Y(_18293_));
 AND2x2_ASAP7_75t_R _26806_ (.A(_18289_),
    .B(_18293_),
    .Y(_18294_));
 NOR2x2_ASAP7_75t_R _26807_ (.A(net2474),
    .B(net1389),
    .Y(_18295_));
 NAND2x2_ASAP7_75t_R _26808_ (.A(net3326),
    .B(_18272_),
    .Y(_18296_));
 NAND2x2_ASAP7_75t_R _26809_ (.A(net1678),
    .B(_18272_),
    .Y(_18297_));
 BUFx2_ASAP7_75t_R input133 (.A(net3960),
    .Y(net133));
 NOR2x2_ASAP7_75t_R _26811_ (.A(_00603_),
    .B(_00604_),
    .Y(_18299_));
 NAND2x2_ASAP7_75t_R _26812_ (.A(_18299_),
    .B(_18284_),
    .Y(_18300_));
 BUFx2_ASAP7_75t_R input132 (.A(net3957),
    .Y(net132));
 AO21x2_ASAP7_75t_R _26814_ (.A1(net937),
    .A2(_18297_),
    .B(_18300_),
    .Y(_18302_));
 INVx3_ASAP7_75t_R _26815_ (.A(_18300_),
    .Y(_18303_));
 AND2x6_ASAP7_75t_R _26816_ (.A(net1677),
    .B(net1391),
    .Y(_18304_));
 NAND2x2_ASAP7_75t_R _26817_ (.A(_18235_),
    .B(_18304_),
    .Y(_18305_));
 INVx5_ASAP7_75t_R _26818_ (.A(net2748),
    .Y(_18306_));
 NAND2x1_ASAP7_75t_R _26819_ (.A(_18303_),
    .B(_18306_),
    .Y(_18307_));
 BUFx2_ASAP7_75t_R input131 (.A(net3963),
    .Y(net131));
 NOR2x2_ASAP7_75t_R _26821_ (.A(_18237_),
    .B(net1579),
    .Y(_18309_));
 OAI21x1_ASAP7_75t_R _26822_ (.A1(net3281),
    .A2(_18309_),
    .B(_18303_),
    .Y(_18310_));
 AND3x1_ASAP7_75t_R _26823_ (.A(_18302_),
    .B(_18307_),
    .C(_18310_),
    .Y(_18311_));
 NAND2x1_ASAP7_75t_R _26824_ (.A(_18294_),
    .B(_18311_),
    .Y(_18312_));
 INVx8_ASAP7_75t_R _26825_ (.A(_18268_),
    .Y(_18313_));
 NAND2x2_ASAP7_75t_R _26826_ (.A(_18238_),
    .B(_18313_),
    .Y(_18314_));
 BUFx2_ASAP7_75t_R input130 (.A(net3814),
    .Y(net130));
 NAND2x2_ASAP7_75t_R _26828_ (.A(_18282_),
    .B(_18313_),
    .Y(_18316_));
 BUFx12f_ASAP7_75t_R input129 (.A(net3838),
    .Y(net129));
 NAND2x2_ASAP7_75t_R _26830_ (.A(_18284_),
    .B(_18264_),
    .Y(_18318_));
 BUFx2_ASAP7_75t_R input128 (.A(net4204),
    .Y(net128));
 AO21x1_ASAP7_75t_R _26832_ (.A1(net2043),
    .A2(net2945),
    .B(_18318_),
    .Y(_18320_));
 BUFx2_ASAP7_75t_R input127 (.A(net4198),
    .Y(net127));
 NAND2x2_ASAP7_75t_R _26834_ (.A(_18235_),
    .B(net1198),
    .Y(_18322_));
 BUFx2_ASAP7_75t_R input126 (.A(net4135),
    .Y(net126));
 AO21x1_ASAP7_75t_R _26836_ (.A1(net1254),
    .A2(net2436),
    .B(_18318_),
    .Y(_18324_));
 AND2x2_ASAP7_75t_R _26837_ (.A(_18320_),
    .B(_18324_),
    .Y(_18325_));
 BUFx2_ASAP7_75t_R input125 (.A(net4010),
    .Y(net125));
 NAND2x2_ASAP7_75t_R _26839_ (.A(net3087),
    .B(net2602),
    .Y(_18327_));
 BUFx2_ASAP7_75t_R input124 (.A(net4013),
    .Y(net124));
 AND2x4_ASAP7_75t_R _26841_ (.A(_00603_),
    .B(_00604_),
    .Y(_18329_));
 NAND2x2_ASAP7_75t_R _26842_ (.A(_18284_),
    .B(_18329_),
    .Y(_18330_));
 BUFx2_ASAP7_75t_R input123 (.A(net4033),
    .Y(net123));
 AO21x1_ASAP7_75t_R _26844_ (.A1(net2176),
    .A2(net1954),
    .B(_18330_),
    .Y(_18332_));
 NAND2x2_ASAP7_75t_R _26845_ (.A(_18235_),
    .B(_18282_),
    .Y(_18333_));
 BUFx2_ASAP7_75t_R input122 (.A(net4184),
    .Y(net122));
 NAND2x2_ASAP7_75t_R _26847_ (.A(_18240_),
    .B(_18235_),
    .Y(_18335_));
 BUFx2_ASAP7_75t_R input121 (.A(net4161),
    .Y(net121));
 AO21x1_ASAP7_75t_R _26849_ (.A1(net2050),
    .A2(_18335_),
    .B(_18330_),
    .Y(_18337_));
 AND2x2_ASAP7_75t_R _26850_ (.A(_18332_),
    .B(_18337_),
    .Y(_18338_));
 BUFx2_ASAP7_75t_R input120 (.A(net4085),
    .Y(net120));
 BUFx2_ASAP7_75t_R input119 (.A(net4079),
    .Y(net119));
 BUFx2_ASAP7_75t_R input118 (.A(net3854),
    .Y(net118));
 AOI211x1_ASAP7_75t_R _26854_ (.A1(net2999),
    .A2(net1396),
    .B(_18330_),
    .C(net2498),
    .Y(_18342_));
 NOR2x2_ASAP7_75t_R _26855_ (.A(net1580),
    .B(_18241_),
    .Y(_18343_));
 NOR2x2_ASAP7_75t_R _26856_ (.A(net2971),
    .B(net1579),
    .Y(_18344_));
 INVx5_ASAP7_75t_R _26857_ (.A(_18330_),
    .Y(_18345_));
 OA21x2_ASAP7_75t_R _26858_ (.A1(_18343_),
    .A2(_18344_),
    .B(_18345_),
    .Y(_18346_));
 NOR2x2_ASAP7_75t_R _26859_ (.A(_18342_),
    .B(_18346_),
    .Y(_18347_));
 NAND3x2_ASAP7_75t_R _26860_ (.B(_18338_),
    .C(_18347_),
    .Y(_18348_),
    .A(_18325_));
 NOR2x1_ASAP7_75t_R _26861_ (.A(_18312_),
    .B(_18348_),
    .Y(_18349_));
 INVx4_ASAP7_75t_R _26862_ (.A(net1702),
    .Y(_18350_));
 NAND2x2_ASAP7_75t_R _26863_ (.A(net2475),
    .B(net3002),
    .Y(_18351_));
 BUFx2_ASAP7_75t_R input117 (.A(net4073),
    .Y(net117));
 NOR2x2_ASAP7_75t_R _26865_ (.A(net2996),
    .B(_00602_),
    .Y(_18353_));
 NAND2x2_ASAP7_75t_R _26866_ (.A(_18353_),
    .B(_18264_),
    .Y(_18354_));
 BUFx2_ASAP7_75t_R input116 (.A(net4053),
    .Y(net116));
 AO21x1_ASAP7_75t_R _26868_ (.A1(_18350_),
    .A2(net2096),
    .B(net3178),
    .Y(_18356_));
 NAND2x2_ASAP7_75t_R _26869_ (.A(_18282_),
    .B(_18272_),
    .Y(_18357_));
 BUFx3_ASAP7_75t_R input115 (.A(net4133),
    .Y(net115));
 AO21x1_ASAP7_75t_R _26871_ (.A1(net2045),
    .A2(net2635),
    .B(net3178),
    .Y(_18359_));
 BUFx2_ASAP7_75t_R input114 (.A(net4113),
    .Y(net114));
 AO21x1_ASAP7_75t_R _26873_ (.A1(net1254),
    .A2(net2050),
    .B(net3178),
    .Y(_18361_));
 NAND3x1_ASAP7_75t_R _26874_ (.A(_18356_),
    .B(_18359_),
    .C(_18361_),
    .Y(_18362_));
 BUFx2_ASAP7_75t_R input113 (.A(net4177),
    .Y(net113));
 NAND2x2_ASAP7_75t_R _26876_ (.A(_18353_),
    .B(_18329_),
    .Y(_18364_));
 BUFx2_ASAP7_75t_R input112 (.A(net4147),
    .Y(net112));
 NAND2x2_ASAP7_75t_R _26878_ (.A(net2980),
    .B(_18280_),
    .Y(_18366_));
 BUFx2_ASAP7_75t_R input111 (.A(net4039),
    .Y(net111));
 AOI211x1_ASAP7_75t_R _26880_ (.A1(net2999),
    .A2(_18237_),
    .B(_18364_),
    .C(net2975),
    .Y(_18368_));
 INVx1_ASAP7_75t_R _26881_ (.A(_18368_),
    .Y(_18369_));
 BUFx2_ASAP7_75t_R input110 (.A(net4069),
    .Y(net110));
 INVx2_ASAP7_75t_R _26883_ (.A(_18364_),
    .Y(_18371_));
 NAND2x1_ASAP7_75t_R _26884_ (.A(_18343_),
    .B(_18371_),
    .Y(_18372_));
 AO21x1_ASAP7_75t_R _26885_ (.A1(net2473),
    .A2(net2419),
    .B(_18364_),
    .Y(_18373_));
 NAND3x1_ASAP7_75t_R _26886_ (.A(_18369_),
    .B(_18372_),
    .C(_18373_),
    .Y(_18374_));
 NOR2x1_ASAP7_75t_R _26887_ (.A(_18362_),
    .B(_18374_),
    .Y(_18375_));
 INVx1_ASAP7_75t_R _26888_ (.A(_18375_),
    .Y(_18376_));
 NAND2x2_ASAP7_75t_R _26889_ (.A(_18353_),
    .B(_18286_),
    .Y(_18377_));
 BUFx2_ASAP7_75t_R input109 (.A(net3769),
    .Y(net109));
 NOR2x1_ASAP7_75t_R _26891_ (.A(_18297_),
    .B(_18377_),
    .Y(_18379_));
 INVx1_ASAP7_75t_R _26892_ (.A(_18379_),
    .Y(_18380_));
 NAND2x2_ASAP7_75t_R _26893_ (.A(_18304_),
    .B(_18313_),
    .Y(_18381_));
 BUFx2_ASAP7_75t_R input108 (.A(net4030),
    .Y(net108));
 NAND2x2_ASAP7_75t_R _26895_ (.A(net1198),
    .B(_18313_),
    .Y(_18383_));
 BUFx2_ASAP7_75t_R input107 (.A(net4023),
    .Y(net107));
 BUFx2_ASAP7_75t_R input106 (.A(net4187),
    .Y(net106));
 AO21x1_ASAP7_75t_R _26898_ (.A1(_18381_),
    .A2(net3182),
    .B(net2981),
    .Y(_18386_));
 NAND2x1_ASAP7_75t_R _26899_ (.A(_18380_),
    .B(_18386_),
    .Y(_18387_));
 AO21x1_ASAP7_75t_R _26900_ (.A1(net2050),
    .A2(net2439),
    .B(_18377_),
    .Y(_18388_));
 BUFx2_ASAP7_75t_R input105 (.A(net4127),
    .Y(net105));
 NOR2x1_ASAP7_75t_R _26902_ (.A(net2011),
    .B(_18377_),
    .Y(_18390_));
 NAND2x1_ASAP7_75t_R _26903_ (.A(_18258_),
    .B(_18390_),
    .Y(_18391_));
 NAND2x1_ASAP7_75t_R _26904_ (.A(_18388_),
    .B(_18391_),
    .Y(_18392_));
 NOR2x1_ASAP7_75t_R _26905_ (.A(_18387_),
    .B(_18392_),
    .Y(_18393_));
 INVx3_ASAP7_75t_R _26906_ (.A(_18269_),
    .Y(_18394_));
 NAND2x2_ASAP7_75t_R _26907_ (.A(_18353_),
    .B(_18299_),
    .Y(_18395_));
 BUFx2_ASAP7_75t_R input104 (.A(net4167),
    .Y(net104));
 AO21x1_ASAP7_75t_R _26909_ (.A1(net2945),
    .A2(_18394_),
    .B(_18395_),
    .Y(_18397_));
 INVx5_ASAP7_75t_R _26910_ (.A(_18395_),
    .Y(_18398_));
 NAND2x1_ASAP7_75t_R _26911_ (.A(_18291_),
    .B(_18398_),
    .Y(_18399_));
 AND2x2_ASAP7_75t_R _26912_ (.A(_18397_),
    .B(_18399_),
    .Y(_18400_));
 NOR2x2_ASAP7_75t_R _26913_ (.A(_18241_),
    .B(_18366_),
    .Y(_18401_));
 NAND2x2_ASAP7_75t_R _26914_ (.A(net2601),
    .B(_18304_),
    .Y(_18402_));
 BUFx2_ASAP7_75t_R input103 (.A(net4067),
    .Y(net103));
 AOI21x1_ASAP7_75t_R _26916_ (.A1(_18402_),
    .A2(net2176),
    .B(_18395_),
    .Y(_18404_));
 NAND2x1_ASAP7_75t_R _26917_ (.A(net1702),
    .B(_18398_),
    .Y(_18405_));
 INVx1_ASAP7_75t_R _26918_ (.A(_18405_),
    .Y(_18406_));
 AOI211x1_ASAP7_75t_R _26919_ (.A1(_18401_),
    .A2(_18398_),
    .B(_18404_),
    .C(_18406_),
    .Y(_18407_));
 NAND3x1_ASAP7_75t_R _26920_ (.A(_18393_),
    .B(_18400_),
    .C(_18407_),
    .Y(_18408_));
 NOR2x1_ASAP7_75t_R _26921_ (.A(_18376_),
    .B(_18408_),
    .Y(_18409_));
 NAND2x1_ASAP7_75t_R _26922_ (.A(_18349_),
    .B(_18409_),
    .Y(_18410_));
 NAND2x2_ASAP7_75t_R _26923_ (.A(_18238_),
    .B(_18272_),
    .Y(_18411_));
 BUFx2_ASAP7_75t_R input102 (.A(net4125),
    .Y(net102));
 AO21x1_ASAP7_75t_R _26925_ (.A1(net2699),
    .A2(net1335),
    .B(_18266_),
    .Y(_18413_));
 BUFx2_ASAP7_75t_R input101 (.A(net4105),
    .Y(net101));
 AO21x1_ASAP7_75t_R _26927_ (.A1(_18402_),
    .A2(_18327_),
    .B(_18266_),
    .Y(_18415_));
 INVx4_ASAP7_75t_R _26928_ (.A(_18266_),
    .Y(_18416_));
 NAND2x1_ASAP7_75t_R _26929_ (.A(_18269_),
    .B(_18416_),
    .Y(_18417_));
 NAND3x1_ASAP7_75t_R _26930_ (.A(_18413_),
    .B(_18415_),
    .C(_18417_),
    .Y(_18418_));
 NAND2x2_ASAP7_75t_R _26931_ (.A(_18256_),
    .B(net2172),
    .Y(_18419_));
 AO31x2_ASAP7_75t_R _26932_ (.A1(net1254),
    .A2(net2004),
    .A3(_18419_),
    .B(_18248_),
    .Y(_18420_));
 NAND2x1_ASAP7_75t_R _26933_ (.A(_18269_),
    .B(_18247_),
    .Y(_18421_));
 INVx1_ASAP7_75t_R _26934_ (.A(_18421_),
    .Y(_18422_));
 BUFx2_ASAP7_75t_R input100 (.A(net4007),
    .Y(net100));
 AOI211x1_ASAP7_75t_R _26936_ (.A1(net1087),
    .A2(_00608_),
    .B(_18248_),
    .C(net2500),
    .Y(_18424_));
 NOR2x1_ASAP7_75t_R _26937_ (.A(_18422_),
    .B(_18424_),
    .Y(_18425_));
 NAND2x1_ASAP7_75t_R _26938_ (.A(_18420_),
    .B(_18425_),
    .Y(_18426_));
 NOR2x1_ASAP7_75t_R _26939_ (.A(_18418_),
    .B(_18426_),
    .Y(_18427_));
 NAND2x2_ASAP7_75t_R _26940_ (.A(_18299_),
    .B(_18265_),
    .Y(_18428_));
 BUFx2_ASAP7_75t_R input99 (.A(net4202),
    .Y(net99));
 NOR2x2_ASAP7_75t_R _26942_ (.A(_18428_),
    .B(_18402_),
    .Y(_18430_));
 AOI211x1_ASAP7_75t_R _26943_ (.A1(net3005),
    .A2(_00608_),
    .B(_18428_),
    .C(net2977),
    .Y(_18431_));
 NOR2x1_ASAP7_75t_R _26944_ (.A(_18430_),
    .B(_18431_),
    .Y(_18432_));
 NOR2x1_ASAP7_75t_R _26945_ (.A(_18428_),
    .B(net1755),
    .Y(_18433_));
 INVx4_ASAP7_75t_R _26946_ (.A(_18428_),
    .Y(_18434_));
 OA21x2_ASAP7_75t_R _26947_ (.A1(_18270_),
    .A2(_18269_),
    .B(_18434_),
    .Y(_18435_));
 NOR2x1_ASAP7_75t_R _26948_ (.A(_18433_),
    .B(_18435_),
    .Y(_18436_));
 NAND2x1_ASAP7_75t_R _26949_ (.A(_18432_),
    .B(_18436_),
    .Y(_18437_));
 BUFx3_ASAP7_75t_R input98 (.A(net4097),
    .Y(net98));
 NAND2x2_ASAP7_75t_R _26951_ (.A(_18286_),
    .B(_18265_),
    .Y(_18439_));
 BUFx2_ASAP7_75t_R input97 (.A(net4192),
    .Y(net97));
 AO31x2_ASAP7_75t_R _26953_ (.A1(net2747),
    .A2(_18335_),
    .A3(_18419_),
    .B(_18439_),
    .Y(_18441_));
 NAND2x2_ASAP7_75t_R _26954_ (.A(_00607_),
    .B(_18313_),
    .Y(_18442_));
 AOI21x1_ASAP7_75t_R _26955_ (.A1(_18442_),
    .A2(_18314_),
    .B(_18439_),
    .Y(_18443_));
 NOR2x2_ASAP7_75t_R _26956_ (.A(_18258_),
    .B(net2498),
    .Y(_18444_));
 NOR2x2_ASAP7_75t_R _26957_ (.A(_18241_),
    .B(net2498),
    .Y(_18445_));
 INVx1_ASAP7_75t_R _26958_ (.A(_18439_),
    .Y(_18446_));
 OA21x2_ASAP7_75t_R _26959_ (.A1(_18444_),
    .A2(_18445_),
    .B(_18446_),
    .Y(_18447_));
 NOR2x1_ASAP7_75t_R _26960_ (.A(_18443_),
    .B(_18447_),
    .Y(_18448_));
 NAND2x1_ASAP7_75t_R _26961_ (.A(_18441_),
    .B(_18448_),
    .Y(_18449_));
 NOR2x1_ASAP7_75t_R _26962_ (.A(_18437_),
    .B(_18449_),
    .Y(_18450_));
 NAND2x2_ASAP7_75t_R _26963_ (.A(_18427_),
    .B(_18450_),
    .Y(_18451_));
 INVx1_ASAP7_75t_R _26964_ (.A(_18451_),
    .Y(_18452_));
 NAND2x2_ASAP7_75t_R _26965_ (.A(net1863),
    .B(_18304_),
    .Y(_18453_));
 BUFx2_ASAP7_75t_R input96 (.A(net4194),
    .Y(net96));
 NOR2x2_ASAP7_75t_R _26967_ (.A(_00602_),
    .B(_18275_),
    .Y(_18455_));
 NAND2x2_ASAP7_75t_R _26968_ (.A(_18455_),
    .B(_18329_),
    .Y(_18456_));
 BUFx2_ASAP7_75t_R input95 (.A(net4055),
    .Y(net95));
 AO21x1_ASAP7_75t_R _26970_ (.A1(net2965),
    .A2(net3003),
    .B(_18456_),
    .Y(_18458_));
 AO21x1_ASAP7_75t_R _26971_ (.A1(net2473),
    .A2(net2106),
    .B(_18456_),
    .Y(_18459_));
 NAND2x2_ASAP7_75t_R _26972_ (.A(net1087),
    .B(_18235_),
    .Y(_18460_));
 AO21x1_ASAP7_75t_R _26973_ (.A1(_18327_),
    .A2(_18460_),
    .B(_18456_),
    .Y(_18461_));
 AND2x2_ASAP7_75t_R _26974_ (.A(_18459_),
    .B(_18461_),
    .Y(_18462_));
 NAND2x2_ASAP7_75t_R _26975_ (.A(_18458_),
    .B(_18462_),
    .Y(_18463_));
 NAND2x2_ASAP7_75t_R _26976_ (.A(_18455_),
    .B(_18264_),
    .Y(_18464_));
 BUFx2_ASAP7_75t_R input94 (.A(net4191),
    .Y(net94));
 NOR2x1_ASAP7_75t_R _26978_ (.A(net2438),
    .B(_18464_),
    .Y(_18466_));
 INVx4_ASAP7_75t_R _26979_ (.A(net1198),
    .Y(_18467_));
 NOR2x2_ASAP7_75t_R _26980_ (.A(_18253_),
    .B(_18467_),
    .Y(_18468_));
 INVx4_ASAP7_75t_R _26981_ (.A(_18464_),
    .Y(_18469_));
 OA21x2_ASAP7_75t_R _26982_ (.A1(_18259_),
    .A2(_18468_),
    .B(_18469_),
    .Y(_18470_));
 NOR2x1_ASAP7_75t_R _26983_ (.A(_18466_),
    .B(_18470_),
    .Y(_18471_));
 BUFx2_ASAP7_75t_R input93 (.A(net4199),
    .Y(net93));
 AO21x1_ASAP7_75t_R _26985_ (.A1(net2701),
    .A2(net1482),
    .B(_18464_),
    .Y(_18473_));
 AO21x1_ASAP7_75t_R _26986_ (.A1(_18383_),
    .A2(_18442_),
    .B(_18464_),
    .Y(_18474_));
 AND2x2_ASAP7_75t_R _26987_ (.A(_18473_),
    .B(_18474_),
    .Y(_18475_));
 NAND2x1_ASAP7_75t_R _26988_ (.A(_18471_),
    .B(_18475_),
    .Y(_18476_));
 NOR2x2_ASAP7_75t_R _26989_ (.A(_18463_),
    .B(_18476_),
    .Y(_18477_));
 BUFx2_ASAP7_75t_R input92 (.A(net4137),
    .Y(net92));
 NAND2x2_ASAP7_75t_R _26991_ (.A(_18455_),
    .B(_18286_),
    .Y(_18479_));
 BUFx2_ASAP7_75t_R input91 (.A(net4131),
    .Y(net91));
 AO21x1_ASAP7_75t_R _26993_ (.A1(net1335),
    .A2(net937),
    .B(_18479_),
    .Y(_18481_));
 NOR2x2_ASAP7_75t_R _26994_ (.A(net1578),
    .B(_18467_),
    .Y(_18482_));
 INVx6_ASAP7_75t_R _26995_ (.A(_18479_),
    .Y(_18483_));
 OAI21x1_ASAP7_75t_R _26996_ (.A1(_18482_),
    .A2(net2669),
    .B(_18483_),
    .Y(_18484_));
 INVx3_ASAP7_75t_R _26997_ (.A(_18297_),
    .Y(_18485_));
 NAND2x2_ASAP7_75t_R _26998_ (.A(_18485_),
    .B(_18483_),
    .Y(_18486_));
 NAND3x2_ASAP7_75t_R _26999_ (.B(_18484_),
    .C(_18486_),
    .Y(_18487_),
    .A(_18481_));
 XOR2x2_ASAP7_75t_R _27000_ (.A(net1679),
    .B(net1393),
    .Y(_18488_));
 NAND2x2_ASAP7_75t_R _27001_ (.A(net2995),
    .B(_18488_),
    .Y(_18489_));
 NAND2x2_ASAP7_75t_R _27002_ (.A(_18299_),
    .B(_18455_),
    .Y(_18490_));
 BUFx2_ASAP7_75t_R input90 (.A(net4077),
    .Y(net90));
 AO21x1_ASAP7_75t_R _27004_ (.A1(_18489_),
    .A2(_18327_),
    .B(net2595),
    .Y(_18492_));
 AOI21x1_ASAP7_75t_R _27005_ (.A1(net1483),
    .A2(net2753),
    .B(net2994),
    .Y(_18493_));
 BUFx2_ASAP7_75t_R input89 (.A(net4095),
    .Y(net89));
 AOI21x1_ASAP7_75t_R _27007_ (.A1(_18383_),
    .A2(net3003),
    .B(net2994),
    .Y(_18495_));
 NOR2x1_ASAP7_75t_R _27008_ (.A(_18493_),
    .B(_18495_),
    .Y(_18496_));
 NAND2x2_ASAP7_75t_R _27009_ (.A(_18492_),
    .B(_18496_),
    .Y(_18497_));
 NAND2x2_ASAP7_75t_R _27010_ (.A(_18401_),
    .B(_18483_),
    .Y(_18498_));
 AOI211x1_ASAP7_75t_R _27011_ (.A1(net3005),
    .A2(net1390),
    .B(_18479_),
    .C(net3246),
    .Y(_18499_));
 INVx1_ASAP7_75t_R _27012_ (.A(_18499_),
    .Y(_18500_));
 NAND2x2_ASAP7_75t_R _27013_ (.A(_18498_),
    .B(_18500_),
    .Y(_18501_));
 NOR3x2_ASAP7_75t_R _27014_ (.B(_18497_),
    .C(_18501_),
    .Y(_18502_),
    .A(_18487_));
 NAND2x2_ASAP7_75t_R _27015_ (.A(_18477_),
    .B(_18502_),
    .Y(_18503_));
 INVx1_ASAP7_75t_R _27016_ (.A(_18503_),
    .Y(_18504_));
 NAND2x1_ASAP7_75t_R _27017_ (.A(_18452_),
    .B(_18504_),
    .Y(_18505_));
 NOR2x2_ASAP7_75t_R _27018_ (.A(_18410_),
    .B(_18505_),
    .Y(_18506_));
 NAND2x2_ASAP7_75t_R _27019_ (.A(_18279_),
    .B(_18506_),
    .Y(_18507_));
 BUFx2_ASAP7_75t_R input88 (.A(net4123),
    .Y(net88));
 BUFx2_ASAP7_75t_R input87 (.A(net4183),
    .Y(net87));
 INVx2_ASAP7_75t_R _27022_ (.A(net3009),
    .Y(_18510_));
 NOR2x2_ASAP7_75t_R _27023_ (.A(net2988),
    .B(_18510_),
    .Y(_18511_));
 BUFx3_ASAP7_75t_R input86 (.A(net4149),
    .Y(net86));
 BUFx2_ASAP7_75t_R input85 (.A(net4087),
    .Y(net85));
 NAND2x2_ASAP7_75t_R _27026_ (.A(net3174),
    .B(net2984),
    .Y(_18514_));
 INVx5_ASAP7_75t_R _27027_ (.A(_18514_),
    .Y(_18515_));
 NAND2x2_ASAP7_75t_R _27028_ (.A(_18511_),
    .B(_18515_),
    .Y(_18516_));
 NOR2x2_ASAP7_75t_R _27029_ (.A(_00567_),
    .B(_00568_),
    .Y(_18517_));
 NAND2x2_ASAP7_75t_R _27030_ (.A(_18517_),
    .B(_18511_),
    .Y(_18518_));
 BUFx2_ASAP7_75t_R input84 (.A(net4043),
    .Y(net84));
 BUFx2_ASAP7_75t_R input83 (.A(net4089),
    .Y(net83));
 NAND2x2_ASAP7_75t_R _27033_ (.A(net2696),
    .B(_00562_),
    .Y(_18521_));
 BUFx2_ASAP7_75t_R input82 (.A(net3860),
    .Y(net82));
 NAND2x2_ASAP7_75t_R _27035_ (.A(_00563_),
    .B(net3211),
    .Y(_18523_));
 NOR2x2_ASAP7_75t_R _27036_ (.A(_18521_),
    .B(_18523_),
    .Y(_18524_));
 INVx3_ASAP7_75t_R _27037_ (.A(_18524_),
    .Y(_18525_));
 AO21x1_ASAP7_75t_R _27038_ (.A1(_18516_),
    .A2(net1966),
    .B(_18525_),
    .Y(_18526_));
 NOR2x2_ASAP7_75t_R _27039_ (.A(net2677),
    .B(net2988),
    .Y(_18527_));
 NAND2x2_ASAP7_75t_R _27040_ (.A(net2302),
    .B(_18515_),
    .Y(_18528_));
 BUFx2_ASAP7_75t_R input81 (.A(net4071),
    .Y(net81));
 INVx13_ASAP7_75t_R _27042_ (.A(net1471),
    .Y(_18530_));
 NOR2x2_ASAP7_75t_R _27043_ (.A(net1731),
    .B(_18530_),
    .Y(_18531_));
 NAND2x2_ASAP7_75t_R _27044_ (.A(net2387),
    .B(_18531_),
    .Y(_18532_));
 AO21x1_ASAP7_75t_R _27045_ (.A1(net3378),
    .A2(net2829),
    .B(_18525_),
    .Y(_18533_));
 BUFx2_ASAP7_75t_R input80 (.A(net4045),
    .Y(net80));
 NAND2x2_ASAP7_75t_R _27047_ (.A(net1735),
    .B(_18530_),
    .Y(_18535_));
 CKINVDCx10_ASAP7_75t_R _27048_ (.A(net1749),
    .Y(_18536_));
 NOR2x2_ASAP7_75t_R _27049_ (.A(net2308),
    .B(_18536_),
    .Y(_18537_));
 NAND2x1_ASAP7_75t_R _27050_ (.A(net2690),
    .B(_18537_),
    .Y(_18538_));
 AND3x1_ASAP7_75t_R _27051_ (.A(_18526_),
    .B(_18533_),
    .C(_18538_),
    .Y(_18539_));
 NAND2x2_ASAP7_75t_R _27052_ (.A(net2988),
    .B(_18510_),
    .Y(_18540_));
 BUFx2_ASAP7_75t_R input79 (.A(net4111),
    .Y(net79));
 INVx2_ASAP7_75t_R _27054_ (.A(_00563_),
    .Y(_18542_));
 NOR2x2_ASAP7_75t_R _27055_ (.A(net3211),
    .B(_18542_),
    .Y(_18543_));
 INVx3_ASAP7_75t_R _27056_ (.A(_18521_),
    .Y(_18544_));
 NAND2x2_ASAP7_75t_R _27057_ (.A(_18543_),
    .B(_18544_),
    .Y(_18545_));
 BUFx2_ASAP7_75t_R input78 (.A(net4195),
    .Y(net78));
 NAND2x2_ASAP7_75t_R _27059_ (.A(net1467),
    .B(net2302),
    .Y(_18547_));
 NAND2x2_ASAP7_75t_R _27060_ (.A(_18517_),
    .B(net2387),
    .Y(_18548_));
 AO21x1_ASAP7_75t_R _27061_ (.A1(_18547_),
    .A2(_18548_),
    .B(_18545_),
    .Y(_18549_));
 OAI21x1_ASAP7_75t_R _27062_ (.A1(net1567),
    .A2(net2479),
    .B(_18549_),
    .Y(_18550_));
 AO21x1_ASAP7_75t_R _27063_ (.A1(_18516_),
    .A2(net2099),
    .B(_18545_),
    .Y(_18551_));
 AND3x4_ASAP7_75t_R _27064_ (.A(net2852),
    .B(net2988),
    .C(net1474),
    .Y(_18552_));
 INVx4_ASAP7_75t_R _27065_ (.A(_18552_),
    .Y(_18553_));
 INVx11_ASAP7_75t_R _27066_ (.A(net1731),
    .Y(_18554_));
 NOR2x2_ASAP7_75t_R _27067_ (.A(net1467),
    .B(_18554_),
    .Y(_18555_));
 NAND2x2_ASAP7_75t_R _27068_ (.A(net3008),
    .B(net2988),
    .Y(_18556_));
 BUFx2_ASAP7_75t_R input77 (.A(net4081),
    .Y(net77));
 CKINVDCx8_ASAP7_75t_R _27070_ (.A(_18556_),
    .Y(_18558_));
 NAND2x2_ASAP7_75t_R _27071_ (.A(_18555_),
    .B(_18558_),
    .Y(_18559_));
 AO21x1_ASAP7_75t_R _27072_ (.A1(_18553_),
    .A2(net3376),
    .B(_18545_),
    .Y(_18560_));
 NAND2x1_ASAP7_75t_R _27073_ (.A(_18551_),
    .B(_18560_),
    .Y(_18561_));
 NOR2x1_ASAP7_75t_R _27074_ (.A(_18550_),
    .B(_18561_),
    .Y(_18562_));
 NAND2x1_ASAP7_75t_R _27075_ (.A(_18539_),
    .B(_18562_),
    .Y(_18563_));
 INVx3_ASAP7_75t_R _27076_ (.A(net2988),
    .Y(_18564_));
 NOR2x2_ASAP7_75t_R _27077_ (.A(net2676),
    .B(_18564_),
    .Y(_18565_));
 BUFx2_ASAP7_75t_R input76 (.A(net4059),
    .Y(net76));
 INVx3_ASAP7_75t_R _27079_ (.A(_00564_),
    .Y(_18567_));
 NOR2x2_ASAP7_75t_R _27080_ (.A(_00563_),
    .B(_18567_),
    .Y(_18568_));
 NAND2x2_ASAP7_75t_R _27081_ (.A(_18568_),
    .B(_18544_),
    .Y(_18569_));
 INVx4_ASAP7_75t_R _27082_ (.A(_18569_),
    .Y(_18570_));
 NAND2x1_ASAP7_75t_R _27083_ (.A(net2555),
    .B(_18570_),
    .Y(_18571_));
 INVx2_ASAP7_75t_R _27084_ (.A(net2829),
    .Y(_18572_));
 NAND2x1_ASAP7_75t_R _27085_ (.A(_18572_),
    .B(_18570_),
    .Y(_18573_));
 OAI21x1_ASAP7_75t_R _27086_ (.A1(_18515_),
    .A2(_18571_),
    .B(_18573_),
    .Y(_18574_));
 NAND2x2_ASAP7_75t_R _27087_ (.A(_18555_),
    .B(_18511_),
    .Y(_18575_));
 AO21x2_ASAP7_75t_R _27088_ (.A1(_18575_),
    .A2(_18518_),
    .B(_18569_),
    .Y(_18576_));
 AO21x2_ASAP7_75t_R _27089_ (.A1(_18553_),
    .A2(net3377),
    .B(_18569_),
    .Y(_18577_));
 NAND2x1_ASAP7_75t_R _27090_ (.A(_18576_),
    .B(_18577_),
    .Y(_18578_));
 NOR2x1_ASAP7_75t_R _27091_ (.A(_18574_),
    .B(_18578_),
    .Y(_18579_));
 BUFx2_ASAP7_75t_R input75 (.A(net3939),
    .Y(net75));
 NAND2x2_ASAP7_75t_R _27093_ (.A(net2678),
    .B(_18564_),
    .Y(_18581_));
 BUFx2_ASAP7_75t_R input74 (.A(net3650),
    .Y(net74));
 NOR2x2_ASAP7_75t_R _27095_ (.A(net1731),
    .B(net2527),
    .Y(_18583_));
 INVx3_ASAP7_75t_R _27096_ (.A(_18583_),
    .Y(_18584_));
 NOR2x2_ASAP7_75t_R _27097_ (.A(net1737),
    .B(net1728),
    .Y(_18585_));
 INVx1_ASAP7_75t_R _27098_ (.A(_18585_),
    .Y(_18586_));
 NOR2x2_ASAP7_75t_R _27099_ (.A(_00563_),
    .B(net3211),
    .Y(_18587_));
 NAND2x2_ASAP7_75t_R _27100_ (.A(_18587_),
    .B(_18544_),
    .Y(_18588_));
 AO21x1_ASAP7_75t_R _27101_ (.A1(_18584_),
    .A2(_18586_),
    .B(_18588_),
    .Y(_18589_));
 NOR2x2_ASAP7_75t_R _27102_ (.A(net1471),
    .B(net1563),
    .Y(_18590_));
 NAND2x1_ASAP7_75t_R _27103_ (.A(_18542_),
    .B(_18567_),
    .Y(_18591_));
 NOR2x2_ASAP7_75t_R _27104_ (.A(_18521_),
    .B(_18591_),
    .Y(_18592_));
 NAND2x1_ASAP7_75t_R _27105_ (.A(_18590_),
    .B(_18592_),
    .Y(_18593_));
 NAND2x2_ASAP7_75t_R _27106_ (.A(net2388),
    .B(_18555_),
    .Y(_18594_));
 AO21x1_ASAP7_75t_R _27107_ (.A1(_18528_),
    .A2(net2386),
    .B(_18588_),
    .Y(_18595_));
 AND3x1_ASAP7_75t_R _27108_ (.A(_18589_),
    .B(_18593_),
    .C(_18595_),
    .Y(_18596_));
 NAND2x1_ASAP7_75t_R _27109_ (.A(_18579_),
    .B(_18596_),
    .Y(_18597_));
 NOR2x2_ASAP7_75t_R _27110_ (.A(_18563_),
    .B(_18597_),
    .Y(_18598_));
 INVx1_ASAP7_75t_R _27111_ (.A(_18598_),
    .Y(_18599_));
 NAND2x2_ASAP7_75t_R _27112_ (.A(_18565_),
    .B(_18531_),
    .Y(_18600_));
 NAND2x2_ASAP7_75t_R _27113_ (.A(_18530_),
    .B(net2387),
    .Y(_18601_));
 INVx2_ASAP7_75t_R _27114_ (.A(net2696),
    .Y(_18602_));
 NOR2x2_ASAP7_75t_R _27115_ (.A(_00562_),
    .B(_18602_),
    .Y(_18603_));
 NAND2x2_ASAP7_75t_R _27116_ (.A(_18603_),
    .B(_18568_),
    .Y(_18604_));
 AO21x1_ASAP7_75t_R _27117_ (.A1(_18600_),
    .A2(_18601_),
    .B(_18604_),
    .Y(_18605_));
 AO21x1_ASAP7_75t_R _27118_ (.A1(net1966),
    .A2(net1730),
    .B(_18604_),
    .Y(_18606_));
 AND2x2_ASAP7_75t_R _27119_ (.A(_18605_),
    .B(_18606_),
    .Y(_18607_));
 NOR2x2_ASAP7_75t_R _27120_ (.A(net1565),
    .B(net3208),
    .Y(_18608_));
 BUFx2_ASAP7_75t_R input73 (.A(net4186),
    .Y(net73));
 AND2x2_ASAP7_75t_R _27122_ (.A(net1748),
    .B(net1069),
    .Y(_18610_));
 NAND2x2_ASAP7_75t_R _27123_ (.A(_18587_),
    .B(_18603_),
    .Y(_18611_));
 INVx4_ASAP7_75t_R _27124_ (.A(_18611_),
    .Y(_18612_));
 OAI21x1_ASAP7_75t_R _27125_ (.A1(_18608_),
    .A2(_18610_),
    .B(_18612_),
    .Y(_18613_));
 NOR2x2_ASAP7_75t_R _27126_ (.A(_18530_),
    .B(net1571),
    .Y(_18614_));
 NAND2x1_ASAP7_75t_R _27127_ (.A(_18614_),
    .B(_18612_),
    .Y(_18615_));
 AND2x2_ASAP7_75t_R _27128_ (.A(_18613_),
    .B(_18615_),
    .Y(_18616_));
 NAND2x2_ASAP7_75t_R _27129_ (.A(_18535_),
    .B(net2101),
    .Y(_18617_));
 AO21x1_ASAP7_75t_R _27130_ (.A1(_18586_),
    .A2(_18617_),
    .B(net2414),
    .Y(_18618_));
 AND3x4_ASAP7_75t_R _27131_ (.A(_18607_),
    .B(_18616_),
    .C(_18618_),
    .Y(_18619_));
 NOR2x1_ASAP7_75t_R _27132_ (.A(net1738),
    .B(_18536_),
    .Y(_18620_));
 INVx2_ASAP7_75t_R _27133_ (.A(_18620_),
    .Y(_18621_));
 BUFx2_ASAP7_75t_R input72 (.A(net4037),
    .Y(net72));
 NAND2x2_ASAP7_75t_R _27135_ (.A(_18530_),
    .B(_18565_),
    .Y(_18623_));
 INVx3_ASAP7_75t_R _27136_ (.A(_18523_),
    .Y(_18624_));
 NAND2x2_ASAP7_75t_R _27137_ (.A(_18603_),
    .B(_18624_),
    .Y(_18625_));
 AO21x1_ASAP7_75t_R _27138_ (.A1(_18621_),
    .A2(_18623_),
    .B(_18625_),
    .Y(_18626_));
 NAND2x2_ASAP7_75t_R _27139_ (.A(_18531_),
    .B(_18558_),
    .Y(_18627_));
 BUFx2_ASAP7_75t_R input71 (.A(net4018),
    .Y(net71));
 AO21x1_ASAP7_75t_R _27141_ (.A1(_18627_),
    .A2(net1965),
    .B(_18625_),
    .Y(_18629_));
 AND2x2_ASAP7_75t_R _27142_ (.A(_18626_),
    .B(_18629_),
    .Y(_18630_));
 INVx1_ASAP7_75t_R _27143_ (.A(_18630_),
    .Y(_18631_));
 NAND2x2_ASAP7_75t_R _27144_ (.A(net2886),
    .B(_18567_),
    .Y(_18632_));
 INVx3_ASAP7_75t_R _27145_ (.A(_00562_),
    .Y(_18633_));
 NAND2x2_ASAP7_75t_R _27146_ (.A(net2696),
    .B(_18633_),
    .Y(_18634_));
 NOR2x2_ASAP7_75t_R _27147_ (.A(_18632_),
    .B(_18634_),
    .Y(_18635_));
 NOR2x2_ASAP7_75t_R _27148_ (.A(_18535_),
    .B(_18581_),
    .Y(_18636_));
 NAND2x2_ASAP7_75t_R _27149_ (.A(net1469),
    .B(_18554_),
    .Y(_18637_));
 NOR2x2_ASAP7_75t_R _27150_ (.A(_18637_),
    .B(_18581_),
    .Y(_18638_));
 OA21x2_ASAP7_75t_R _27151_ (.A1(_18636_),
    .A2(_18638_),
    .B(_18635_),
    .Y(_18639_));
 AO21x1_ASAP7_75t_R _27152_ (.A1(_18635_),
    .A2(_18585_),
    .B(_18639_),
    .Y(_18640_));
 NAND2x2_ASAP7_75t_R _27153_ (.A(_18543_),
    .B(_18603_),
    .Y(_18641_));
 NOR2x1_ASAP7_75t_R _27154_ (.A(_18600_),
    .B(_18641_),
    .Y(_18642_));
 NAND2x2_ASAP7_75t_R _27155_ (.A(_18565_),
    .B(_18555_),
    .Y(_18643_));
 NOR2x1_ASAP7_75t_R _27156_ (.A(_18643_),
    .B(_18641_),
    .Y(_18644_));
 NOR2x1_ASAP7_75t_R _27157_ (.A(_18548_),
    .B(_18641_),
    .Y(_18645_));
 OR3x2_ASAP7_75t_R _27158_ (.A(_18642_),
    .B(_18644_),
    .C(_18645_),
    .Y(_18646_));
 NOR3x1_ASAP7_75t_R _27159_ (.A(_18631_),
    .B(_18640_),
    .C(_18646_),
    .Y(_18647_));
 NAND2x1_ASAP7_75t_R _27160_ (.A(_18619_),
    .B(_18647_),
    .Y(_18648_));
 NOR2x1_ASAP7_75t_R _27161_ (.A(_18599_),
    .B(_18648_),
    .Y(_18649_));
 NOR2x2_ASAP7_75t_R _27162_ (.A(_18514_),
    .B(_18556_),
    .Y(_18650_));
 CKINVDCx5p33_ASAP7_75t_R _27163_ (.A(_18650_),
    .Y(_18651_));
 BUFx2_ASAP7_75t_R input70 (.A(net3981),
    .Y(net70));
 NAND2x2_ASAP7_75t_R _27165_ (.A(net1011),
    .B(net2102),
    .Y(_18653_));
 NOR2x2_ASAP7_75t_R _27166_ (.A(net2696),
    .B(_00562_),
    .Y(_18654_));
 NAND2x2_ASAP7_75t_R _27167_ (.A(_18654_),
    .B(_18624_),
    .Y(_18655_));
 AO21x1_ASAP7_75t_R _27168_ (.A1(_18651_),
    .A2(_18653_),
    .B(_18655_),
    .Y(_18656_));
 NAND2x2_ASAP7_75t_R _27169_ (.A(net1469),
    .B(_18565_),
    .Y(_18657_));
 NOR2x1_ASAP7_75t_R _27170_ (.A(_18657_),
    .B(_18655_),
    .Y(_18658_));
 INVx1_ASAP7_75t_R _27171_ (.A(_18658_),
    .Y(_18659_));
 BUFx2_ASAP7_75t_R input69 (.A(net4049),
    .Y(net69));
 AO21x1_ASAP7_75t_R _27173_ (.A1(net2398),
    .A2(_18601_),
    .B(_18655_),
    .Y(_18661_));
 AND3x2_ASAP7_75t_R _27174_ (.A(_18656_),
    .B(_18659_),
    .C(_18661_),
    .Y(_18662_));
 INVx1_ASAP7_75t_R _27175_ (.A(_18662_),
    .Y(_18663_));
 BUFx2_ASAP7_75t_R input68 (.A(net4063),
    .Y(net68));
 BUFx2_ASAP7_75t_R input67 (.A(net3889),
    .Y(net67));
 NAND2x2_ASAP7_75t_R _27178_ (.A(_18654_),
    .B(_18543_),
    .Y(_18666_));
 BUFx2_ASAP7_75t_R input66 (.A(net3998),
    .Y(net66));
 AO21x1_ASAP7_75t_R _27180_ (.A1(net1404),
    .A2(net2421),
    .B(_18666_),
    .Y(_18668_));
 AO21x1_ASAP7_75t_R _27181_ (.A1(_18528_),
    .A2(net2398),
    .B(_18666_),
    .Y(_18669_));
 INVx2_ASAP7_75t_R _27182_ (.A(_18654_),
    .Y(_18670_));
 NOR2x2_ASAP7_75t_R _27183_ (.A(_18632_),
    .B(_18670_),
    .Y(_18671_));
 INVx3_ASAP7_75t_R _27184_ (.A(_18548_),
    .Y(_18672_));
 NAND2x1_ASAP7_75t_R _27185_ (.A(_18671_),
    .B(_18672_),
    .Y(_18673_));
 INVx3_ASAP7_75t_R _27186_ (.A(_18517_),
    .Y(_18674_));
 NOR2x2_ASAP7_75t_R _27187_ (.A(_18674_),
    .B(_18540_),
    .Y(_18675_));
 NAND2x2_ASAP7_75t_R _27188_ (.A(_18675_),
    .B(_18671_),
    .Y(_18676_));
 AND3x2_ASAP7_75t_R _27189_ (.A(_18669_),
    .B(_18673_),
    .C(_18676_),
    .Y(_18677_));
 NAND2x1_ASAP7_75t_R _27190_ (.A(_18668_),
    .B(_18677_),
    .Y(_18678_));
 NOR2x1_ASAP7_75t_R _27191_ (.A(_18663_),
    .B(_18678_),
    .Y(_18679_));
 NAND2x2_ASAP7_75t_R _27192_ (.A(net1748),
    .B(_18535_),
    .Y(_18680_));
 INVx1_ASAP7_75t_R _27193_ (.A(_18680_),
    .Y(_18681_));
 NAND2x2_ASAP7_75t_R _27194_ (.A(_18654_),
    .B(_18568_),
    .Y(_18682_));
 INVx5_ASAP7_75t_R _27195_ (.A(_18682_),
    .Y(_18683_));
 OA211x2_ASAP7_75t_R _27196_ (.A1(net2555),
    .A2(_18681_),
    .B(_18683_),
    .C(_18637_),
    .Y(_18684_));
 NAND2x2_ASAP7_75t_R _27197_ (.A(_18531_),
    .B(_18511_),
    .Y(_18685_));
 BUFx2_ASAP7_75t_R input65 (.A(net4099),
    .Y(net65));
 NAND2x2_ASAP7_75t_R _27199_ (.A(_18530_),
    .B(net2101),
    .Y(_18687_));
 AO21x1_ASAP7_75t_R _27200_ (.A1(_18685_),
    .A2(_18687_),
    .B(net2545),
    .Y(_18688_));
 NAND2x1_ASAP7_75t_R _27201_ (.A(_18552_),
    .B(_18683_),
    .Y(_18689_));
 NOR2x2_ASAP7_75t_R _27202_ (.A(net1728),
    .B(net3210),
    .Y(_18690_));
 NAND2x1_ASAP7_75t_R _27203_ (.A(_18690_),
    .B(_18683_),
    .Y(_18691_));
 NAND3x1_ASAP7_75t_R _27204_ (.A(_18688_),
    .B(_18689_),
    .C(_18691_),
    .Y(_18692_));
 NOR2x1_ASAP7_75t_R _27205_ (.A(_18684_),
    .B(_18692_),
    .Y(_18693_));
 NOR2x2_ASAP7_75t_R _27206_ (.A(net1563),
    .B(_18637_),
    .Y(_18694_));
 NAND2x2_ASAP7_75t_R _27207_ (.A(_18654_),
    .B(_18587_),
    .Y(_18695_));
 INVx4_ASAP7_75t_R _27208_ (.A(_18695_),
    .Y(_18696_));
 NAND2x1_ASAP7_75t_R _27209_ (.A(_18694_),
    .B(_18696_),
    .Y(_18697_));
 AO21x1_ASAP7_75t_R _27210_ (.A1(_18528_),
    .A2(_18594_),
    .B(_18695_),
    .Y(_18698_));
 NAND2x1_ASAP7_75t_R _27211_ (.A(_18697_),
    .B(_18698_),
    .Y(_18699_));
 BUFx2_ASAP7_75t_R input64 (.A(net4057),
    .Y(net64));
 BUFx2_ASAP7_75t_R input63 (.A(net4041),
    .Y(net63));
 NAND2x2_ASAP7_75t_R _27214_ (.A(net1467),
    .B(_18511_),
    .Y(_18702_));
 NOR2x2_ASAP7_75t_R _27215_ (.A(net2182),
    .B(_18702_),
    .Y(_18703_));
 OA21x2_ASAP7_75t_R _27216_ (.A1(_18690_),
    .A2(_18552_),
    .B(_18696_),
    .Y(_18704_));
 NOR3x1_ASAP7_75t_R _27217_ (.A(_18699_),
    .B(_18703_),
    .C(_18704_),
    .Y(_18705_));
 NAND2x1_ASAP7_75t_R _27218_ (.A(_18693_),
    .B(_18705_),
    .Y(_18706_));
 INVx1_ASAP7_75t_R _27219_ (.A(_18706_),
    .Y(_18707_));
 NAND2x1_ASAP7_75t_R _27220_ (.A(_18679_),
    .B(_18707_),
    .Y(_18708_));
 BUFx2_ASAP7_75t_R input62 (.A(net4129),
    .Y(net62));
 BUFx2_ASAP7_75t_R input61 (.A(net4115),
    .Y(net61));
 NOR2x2_ASAP7_75t_R _27223_ (.A(net2696),
    .B(_18633_),
    .Y(_18711_));
 NAND2x2_ASAP7_75t_R _27224_ (.A(_18711_),
    .B(_18568_),
    .Y(_18712_));
 AO221x2_ASAP7_75t_R _27225_ (.A1(net3090),
    .A2(_18554_),
    .B1(net1570),
    .B2(_18536_),
    .C(net3324),
    .Y(_18713_));
 NAND2x2_ASAP7_75t_R _27226_ (.A(_18587_),
    .B(_18711_),
    .Y(_18714_));
 AO21x1_ASAP7_75t_R _27227_ (.A1(_18553_),
    .A2(_18617_),
    .B(_18714_),
    .Y(_18715_));
 AO21x1_ASAP7_75t_R _27228_ (.A1(_18623_),
    .A2(net2433),
    .B(_18714_),
    .Y(_18716_));
 AND2x2_ASAP7_75t_R _27229_ (.A(_18715_),
    .B(_18716_),
    .Y(_18717_));
 INVx3_ASAP7_75t_R _27230_ (.A(_18712_),
    .Y(_18718_));
 NAND2x2_ASAP7_75t_R _27231_ (.A(net2979),
    .B(_18718_),
    .Y(_18719_));
 NAND3x2_ASAP7_75t_R _27232_ (.B(_18717_),
    .C(_18719_),
    .Y(_18720_),
    .A(_18713_));
 NAND2x2_ASAP7_75t_R _27233_ (.A(net3004),
    .B(_18558_),
    .Y(_18721_));
 BUFx2_ASAP7_75t_R input60 (.A(net4200),
    .Y(net60));
 NAND2x2_ASAP7_75t_R _27235_ (.A(_18711_),
    .B(_18624_),
    .Y(_18723_));
 AO21x1_ASAP7_75t_R _27236_ (.A1(_18651_),
    .A2(_18721_),
    .B(_18723_),
    .Y(_18724_));
 INVx4_ASAP7_75t_R _27237_ (.A(_18723_),
    .Y(_18725_));
 NAND2x1_ASAP7_75t_R _27238_ (.A(_18614_),
    .B(_18725_),
    .Y(_18726_));
 NAND2x1_ASAP7_75t_R _27239_ (.A(_18638_),
    .B(_18725_),
    .Y(_18727_));
 NAND3x1_ASAP7_75t_R _27240_ (.A(_18724_),
    .B(_18726_),
    .C(_18727_),
    .Y(_18728_));
 NAND2x2_ASAP7_75t_R _27241_ (.A(_18711_),
    .B(_18543_),
    .Y(_18729_));
 AO21x1_ASAP7_75t_R _27242_ (.A1(_18575_),
    .A2(_18518_),
    .B(net2694),
    .Y(_18730_));
 AO21x1_ASAP7_75t_R _27243_ (.A1(_18627_),
    .A2(_18721_),
    .B(net2694),
    .Y(_18731_));
 AND2x2_ASAP7_75t_R _27244_ (.A(_18730_),
    .B(_18731_),
    .Y(_18732_));
 AO21x1_ASAP7_75t_R _27245_ (.A1(_18600_),
    .A2(_18643_),
    .B(_18729_),
    .Y(_18733_));
 AO21x1_ASAP7_75t_R _27246_ (.A1(_18528_),
    .A2(_18548_),
    .B(_18729_),
    .Y(_18734_));
 AND2x2_ASAP7_75t_R _27247_ (.A(_18733_),
    .B(_18734_),
    .Y(_18735_));
 NAND2x1_ASAP7_75t_R _27248_ (.A(_18732_),
    .B(_18735_),
    .Y(_18736_));
 NOR2x1_ASAP7_75t_R _27249_ (.A(_18728_),
    .B(_18736_),
    .Y(_18737_));
 INVx1_ASAP7_75t_R _27250_ (.A(_18737_),
    .Y(_18738_));
 NOR2x2_ASAP7_75t_R _27251_ (.A(_18720_),
    .B(_18738_),
    .Y(_18739_));
 INVx1_ASAP7_75t_R _27252_ (.A(_18739_),
    .Y(_18740_));
 NOR2x2_ASAP7_75t_R _27253_ (.A(_18708_),
    .B(_18740_),
    .Y(_18741_));
 NAND2x2_ASAP7_75t_R _27254_ (.A(_18649_),
    .B(_18741_),
    .Y(_18742_));
 XOR2x1_ASAP7_75t_R _27255_ (.A(_18507_),
    .Y(_18743_),
    .B(_18742_));
 AOI21x1_ASAP7_75t_R _27256_ (.A1(_18194_),
    .A2(_18233_),
    .B(_18743_),
    .Y(_18744_));
 AO21x1_ASAP7_75t_R _27257_ (.A1(_17919_),
    .A2(_17921_),
    .B(_18192_),
    .Y(_18745_));
 NAND2x1_ASAP7_75t_R _27258_ (.A(_18192_),
    .B(_18232_),
    .Y(_18746_));
 INVx1_ASAP7_75t_R _27259_ (.A(_18743_),
    .Y(_18747_));
 AOI21x1_ASAP7_75t_R _27260_ (.A1(_18745_),
    .A2(_18746_),
    .B(_18747_),
    .Y(_18748_));
 BUFx2_ASAP7_75t_R input59 (.A(net4109),
    .Y(net59));
 BUFx2_ASAP7_75t_R input58 (.A(net4091),
    .Y(net58));
 OAI21x1_ASAP7_75t_R _27263_ (.A1(_18744_),
    .A2(_18748_),
    .B(net397),
    .Y(_18751_));
 NAND2x1_ASAP7_75t_R _27264_ (.A(_17528_),
    .B(_18751_),
    .Y(_18752_));
 XOR2x2_ASAP7_75t_R _27265_ (.A(_18752_),
    .B(_14672_),
    .Y(_00121_));
 CKINVDCx20_ASAP7_75t_R _27266_ (.A(net395),
    .Y(_18753_));
 BUFx2_ASAP7_75t_R input57 (.A(net4083),
    .Y(net57));
 BUFx2_ASAP7_75t_R input56 (.A(net4065),
    .Y(net56));
 AND2x2_ASAP7_75t_R _27269_ (.A(net390),
    .B(_00914_),
    .Y(_18756_));
 INVx2_ASAP7_75t_R _27270_ (.A(_18232_),
    .Y(_18757_));
 BUFx2_ASAP7_75t_R input55 (.A(net4101),
    .Y(net55));
 AOI21x1_ASAP7_75t_R _27272_ (.A1(net2015),
    .A2(net1081),
    .B(_17566_),
    .Y(_18759_));
 AOI21x1_ASAP7_75t_R _27273_ (.A1(net1082),
    .A2(net1098),
    .B(_17566_),
    .Y(_18760_));
 NOR2x1_ASAP7_75t_R _27274_ (.A(_18759_),
    .B(_18760_),
    .Y(_18761_));
 BUFx2_ASAP7_75t_R input54 (.A(net4103),
    .Y(net54));
 AO31x2_ASAP7_75t_R _27276_ (.A1(net936),
    .A2(_17626_),
    .A3(_17665_),
    .B(_17566_),
    .Y(_18763_));
 NAND2x1_ASAP7_75t_R _27277_ (.A(_18761_),
    .B(_18763_),
    .Y(_18764_));
 AO21x1_ASAP7_75t_R _27278_ (.A1(_17845_),
    .A2(_17695_),
    .B(_17547_),
    .Y(_18765_));
 AO21x1_ASAP7_75t_R _27279_ (.A1(_17834_),
    .A2(net1816),
    .B(_17547_),
    .Y(_18766_));
 NAND2x1_ASAP7_75t_R _27280_ (.A(net1901),
    .B(_17548_),
    .Y(_18767_));
 NAND3x1_ASAP7_75t_R _27281_ (.A(_18765_),
    .B(_18766_),
    .C(_18767_),
    .Y(_18768_));
 NOR2x1_ASAP7_75t_R _27282_ (.A(_18764_),
    .B(_18768_),
    .Y(_18769_));
 BUFx2_ASAP7_75t_R input53 (.A(net4196),
    .Y(net53));
 AO21x1_ASAP7_75t_R _27284_ (.A1(net2202),
    .A2(_17756_),
    .B(_17614_),
    .Y(_18771_));
 BUFx2_ASAP7_75t_R input52 (.A(net4151),
    .Y(net52));
 AO21x1_ASAP7_75t_R _27286_ (.A1(_17834_),
    .A2(_17575_),
    .B(_17614_),
    .Y(_18773_));
 NAND2x1_ASAP7_75t_R _27287_ (.A(_17609_),
    .B(_17618_),
    .Y(_18774_));
 NAND3x1_ASAP7_75t_R _27288_ (.A(_18771_),
    .B(_18773_),
    .C(_18774_),
    .Y(_18775_));
 BUFx2_ASAP7_75t_R input51 (.A(net4163),
    .Y(net51));
 AO31x2_ASAP7_75t_R _27290_ (.A1(net2630),
    .A2(net2893),
    .A3(net1097),
    .B(_17589_),
    .Y(_18777_));
 NAND2x1_ASAP7_75t_R _27291_ (.A(_17604_),
    .B(_17609_),
    .Y(_18778_));
 OA21x2_ASAP7_75t_R _27292_ (.A1(_17605_),
    .A2(net1832),
    .B(_18778_),
    .Y(_18779_));
 NAND2x1_ASAP7_75t_R _27293_ (.A(_18777_),
    .B(_18779_),
    .Y(_18780_));
 NOR2x1_ASAP7_75t_R _27294_ (.A(_18775_),
    .B(_18780_),
    .Y(_18781_));
 NAND2x1_ASAP7_75t_R _27295_ (.A(_18769_),
    .B(_18781_),
    .Y(_18782_));
 AO21x1_ASAP7_75t_R _27296_ (.A1(net936),
    .A2(_17562_),
    .B(net2484),
    .Y(_18783_));
 AO21x1_ASAP7_75t_R _27297_ (.A1(_17645_),
    .A2(_17551_),
    .B(_17641_),
    .Y(_18784_));
 NAND2x1_ASAP7_75t_R _27298_ (.A(_17661_),
    .B(_17650_),
    .Y(_18785_));
 NAND3x1_ASAP7_75t_R _27299_ (.A(_18783_),
    .B(_18784_),
    .C(_18785_),
    .Y(_18786_));
 AO21x1_ASAP7_75t_R _27300_ (.A1(net1097),
    .A2(_17834_),
    .B(_17629_),
    .Y(_18787_));
 NOR2x2_ASAP7_75t_R _27301_ (.A(_17608_),
    .B(net1973),
    .Y(_18788_));
 INVx3_ASAP7_75t_R _27302_ (.A(_17629_),
    .Y(_18789_));
 NAND2x1_ASAP7_75t_R _27303_ (.A(_18788_),
    .B(_18789_),
    .Y(_18790_));
 NAND3x1_ASAP7_75t_R _27304_ (.A(_18787_),
    .B(_17900_),
    .C(_18790_),
    .Y(_18791_));
 NOR2x1_ASAP7_75t_R _27305_ (.A(_18786_),
    .B(_18791_),
    .Y(_18792_));
 BUFx2_ASAP7_75t_R input50 (.A(net3880),
    .Y(net50));
 AO31x2_ASAP7_75t_R _27307_ (.A1(net2630),
    .A2(_17813_),
    .A3(net1097),
    .B(net3313),
    .Y(_18794_));
 AOI211x1_ASAP7_75t_R _27308_ (.A1(net1123),
    .A2(net1186),
    .B(net3313),
    .C(net1974),
    .Y(_18795_));
 OA21x2_ASAP7_75t_R _27309_ (.A1(_17788_),
    .A2(net2640),
    .B(_17671_),
    .Y(_18796_));
 NOR2x1_ASAP7_75t_R _27310_ (.A(_18795_),
    .B(_18796_),
    .Y(_18797_));
 NAND2x1_ASAP7_75t_R _27311_ (.A(_18794_),
    .B(_18797_),
    .Y(_18798_));
 NOR2x2_ASAP7_75t_R _27312_ (.A(net1816),
    .B(_17657_),
    .Y(_18799_));
 AOI21x1_ASAP7_75t_R _27313_ (.A1(_17586_),
    .A2(_17813_),
    .B(net2847),
    .Y(_18800_));
 NOR2x1_ASAP7_75t_R _27314_ (.A(_18799_),
    .B(_18800_),
    .Y(_18801_));
 AO21x1_ASAP7_75t_R _27315_ (.A1(_17626_),
    .A2(net2899),
    .B(net2847),
    .Y(_18802_));
 BUFx2_ASAP7_75t_R input49 (.A(net4193),
    .Y(net49));
 AO21x1_ASAP7_75t_R _27317_ (.A1(net2202),
    .A2(net941),
    .B(net2847),
    .Y(_18804_));
 NAND3x1_ASAP7_75t_R _27318_ (.A(_18801_),
    .B(_18802_),
    .C(_18804_),
    .Y(_18805_));
 NOR2x1_ASAP7_75t_R _27319_ (.A(_18798_),
    .B(_18805_),
    .Y(_18806_));
 NAND2x2_ASAP7_75t_R _27320_ (.A(_18792_),
    .B(_18806_),
    .Y(_18807_));
 NOR2x2_ASAP7_75t_R _27321_ (.A(_18807_),
    .B(_18782_),
    .Y(_18808_));
 AO21x1_ASAP7_75t_R _27322_ (.A1(net1098),
    .A2(net1097),
    .B(net2909),
    .Y(_18809_));
 AO21x1_ASAP7_75t_R _27323_ (.A1(_17831_),
    .A2(_17756_),
    .B(net2909),
    .Y(_18810_));
 NAND3x1_ASAP7_75t_R _27324_ (.A(_17836_),
    .B(_18809_),
    .C(_18810_),
    .Y(_18811_));
 NAND2x1_ASAP7_75t_R _27325_ (.A(_17571_),
    .B(_17782_),
    .Y(_18812_));
 INVx1_ASAP7_75t_R _27326_ (.A(_18812_),
    .Y(_18813_));
 AOI21x1_ASAP7_75t_R _27327_ (.A1(net936),
    .A2(_17756_),
    .B(_17777_),
    .Y(_18814_));
 AOI21x1_ASAP7_75t_R _27328_ (.A1(_17555_),
    .A2(_18813_),
    .B(_18814_),
    .Y(_18815_));
 OA21x2_ASAP7_75t_R _27329_ (.A1(_17661_),
    .A2(_17673_),
    .B(_17782_),
    .Y(_18816_));
 NOR2x1_ASAP7_75t_R _27330_ (.A(_17779_),
    .B(_18816_),
    .Y(_18817_));
 NAND2x1_ASAP7_75t_R _27331_ (.A(_18815_),
    .B(_18817_),
    .Y(_18818_));
 NOR2x1_ASAP7_75t_R _27332_ (.A(_18811_),
    .B(_18818_),
    .Y(_18819_));
 AO21x1_ASAP7_75t_R _27333_ (.A1(_17626_),
    .A2(net941),
    .B(_17744_),
    .Y(_18820_));
 AO21x1_ASAP7_75t_R _27334_ (.A1(net1097),
    .A2(_17834_),
    .B(_17744_),
    .Y(_18821_));
 AO21x1_ASAP7_75t_R _27335_ (.A1(_17813_),
    .A2(net2630),
    .B(_17744_),
    .Y(_18822_));
 NAND3x1_ASAP7_75t_R _27336_ (.A(_18820_),
    .B(_18821_),
    .C(_18822_),
    .Y(_18823_));
 AO31x2_ASAP7_75t_R _27337_ (.A1(net2903),
    .A2(net3193),
    .A3(net1081),
    .B(_17759_),
    .Y(_18824_));
 NOR2x2_ASAP7_75t_R _27338_ (.A(_17601_),
    .B(_17781_),
    .Y(_18825_));
 OA21x2_ASAP7_75t_R _27339_ (.A1(_17788_),
    .A2(net2640),
    .B(_18825_),
    .Y(_18826_));
 AOI211x1_ASAP7_75t_R _27340_ (.A1(net2907),
    .A2(_17533_),
    .B(_17759_),
    .C(_17557_),
    .Y(_18827_));
 NOR2x1_ASAP7_75t_R _27341_ (.A(_18826_),
    .B(_18827_),
    .Y(_18828_));
 NAND2x1_ASAP7_75t_R _27342_ (.A(_18824_),
    .B(_18828_),
    .Y(_18829_));
 NOR2x1_ASAP7_75t_R _27343_ (.A(_18823_),
    .B(_18829_),
    .Y(_18830_));
 NAND2x1_ASAP7_75t_R _27344_ (.A(_18819_),
    .B(_18830_),
    .Y(_18831_));
 AO21x1_ASAP7_75t_R _27345_ (.A1(net936),
    .A2(_17756_),
    .B(_17691_),
    .Y(_18832_));
 OAI21x1_ASAP7_75t_R _27346_ (.A1(_17758_),
    .A2(_17691_),
    .B(_18832_),
    .Y(_18833_));
 NOR2x2_ASAP7_75t_R _27347_ (.A(net2880),
    .B(net1975),
    .Y(_18834_));
 OAI21x1_ASAP7_75t_R _27348_ (.A1(_17694_),
    .A2(_18834_),
    .B(net3086),
    .Y(_18835_));
 NAND3x1_ASAP7_75t_R _27349_ (.A(_18835_),
    .B(_17907_),
    .C(_17908_),
    .Y(_18836_));
 OA21x2_ASAP7_75t_R _27350_ (.A1(_17679_),
    .A2(_17731_),
    .B(_17801_),
    .Y(_18837_));
 NOR3x1_ASAP7_75t_R _27351_ (.A(_18833_),
    .B(_18836_),
    .C(_18837_),
    .Y(_18838_));
 NAND2x1_ASAP7_75t_R _27352_ (.A(_17733_),
    .B(_18834_),
    .Y(_18839_));
 AO21x1_ASAP7_75t_R _27353_ (.A1(_17626_),
    .A2(_17695_),
    .B(_17725_),
    .Y(_18840_));
 NAND2x1_ASAP7_75t_R _27354_ (.A(_18839_),
    .B(_18840_),
    .Y(_18841_));
 BUFx2_ASAP7_75t_R input48 (.A(net4185),
    .Y(net48));
 AOI211x1_ASAP7_75t_R _27356_ (.A1(net2862),
    .A2(net2879),
    .B(_17712_),
    .C(_17575_),
    .Y(_18843_));
 OA21x2_ASAP7_75t_R _27357_ (.A1(_17780_),
    .A2(_17661_),
    .B(_17714_),
    .Y(_18844_));
 NOR2x1_ASAP7_75t_R _27358_ (.A(_18843_),
    .B(_18844_),
    .Y(_18845_));
 AND2x2_ASAP7_75t_R _27359_ (.A(_17811_),
    .B(_17715_),
    .Y(_18846_));
 NAND2x1_ASAP7_75t_R _27360_ (.A(_18845_),
    .B(_18846_),
    .Y(_18847_));
 NOR2x1_ASAP7_75t_R _27361_ (.A(_18841_),
    .B(_18847_),
    .Y(_18848_));
 NAND2x1_ASAP7_75t_R _27362_ (.A(_18838_),
    .B(_18848_),
    .Y(_18849_));
 NOR2x1_ASAP7_75t_R _27363_ (.A(_18831_),
    .B(_18849_),
    .Y(_18850_));
 NAND2x2_ASAP7_75t_R _27364_ (.A(_18808_),
    .B(_18850_),
    .Y(_18851_));
 NOR2x2_ASAP7_75t_R _27365_ (.A(_18230_),
    .B(_18851_),
    .Y(_18852_));
 AO21x1_ASAP7_75t_R _27366_ (.A1(net3302),
    .A2(_17963_),
    .B(net2364),
    .Y(_18853_));
 AO21x1_ASAP7_75t_R _27367_ (.A1(net2908),
    .A2(net1839),
    .B(_17968_),
    .Y(_18854_));
 BUFx2_ASAP7_75t_R input47 (.A(net3863),
    .Y(net47));
 AO21x1_ASAP7_75t_R _27369_ (.A1(_18073_),
    .A2(net3190),
    .B(net2364),
    .Y(_18856_));
 AND3x1_ASAP7_75t_R _27370_ (.A(_18853_),
    .B(_18854_),
    .C(_18856_),
    .Y(_18857_));
 AO21x1_ASAP7_75t_R _27371_ (.A1(_18073_),
    .A2(net3284),
    .B(net1746),
    .Y(_18858_));
 INVx1_ASAP7_75t_R _27372_ (.A(_18098_),
    .Y(_18859_));
 NOR2x2_ASAP7_75t_R _27373_ (.A(net2823),
    .B(net2059),
    .Y(_18860_));
 NAND2x1_ASAP7_75t_R _27374_ (.A(_18860_),
    .B(_17932_),
    .Y(_18861_));
 AND3x1_ASAP7_75t_R _27375_ (.A(_18858_),
    .B(_18859_),
    .C(_18861_),
    .Y(_18862_));
 AND2x2_ASAP7_75t_R _27376_ (.A(_18857_),
    .B(_18862_),
    .Y(_18863_));
 NAND2x2_ASAP7_75t_R _27377_ (.A(_17996_),
    .B(_17928_),
    .Y(_18864_));
 AO21x1_ASAP7_75t_R _27378_ (.A1(net3302),
    .A2(_17962_),
    .B(_18864_),
    .Y(_18865_));
 AOI211x1_ASAP7_75t_R _27379_ (.A1(net3201),
    .A2(net3308),
    .B(net2060),
    .C(_18864_),
    .Y(_18866_));
 INVx2_ASAP7_75t_R _27380_ (.A(_18866_),
    .Y(_18867_));
 NAND2x1_ASAP7_75t_R _27381_ (.A(_18865_),
    .B(_18867_),
    .Y(_18868_));
 NOR2x2_ASAP7_75t_R _27382_ (.A(net3366),
    .B(net1365),
    .Y(_18869_));
 OA21x2_ASAP7_75t_R _27383_ (.A1(net3218),
    .A2(_18869_),
    .B(_18123_),
    .Y(_18870_));
 BUFx2_ASAP7_75t_R input46 (.A(net4159),
    .Y(net46));
 OAI21x1_ASAP7_75t_R _27385_ (.A1(net1121),
    .A2(_18126_),
    .B(_18133_),
    .Y(_18872_));
 NOR2x1_ASAP7_75t_R _27386_ (.A(_18870_),
    .B(_18872_),
    .Y(_18873_));
 OA21x2_ASAP7_75t_R _27387_ (.A1(_18178_),
    .A2(_18110_),
    .B(_18123_),
    .Y(_18874_));
 INVx1_ASAP7_75t_R _27388_ (.A(_18874_),
    .Y(_18875_));
 AND2x2_ASAP7_75t_R _27389_ (.A(_18875_),
    .B(_18128_),
    .Y(_18876_));
 NAND2x1_ASAP7_75t_R _27390_ (.A(_18873_),
    .B(_18876_),
    .Y(_18877_));
 NOR2x1_ASAP7_75t_R _27391_ (.A(_18868_),
    .B(_18877_),
    .Y(_18878_));
 NAND2x1_ASAP7_75t_R _27392_ (.A(_18863_),
    .B(_18878_),
    .Y(_18879_));
 AO21x1_ASAP7_75t_R _27393_ (.A1(_18028_),
    .A2(net1622),
    .B(net2446),
    .Y(_18880_));
 NAND2x2_ASAP7_75t_R _27394_ (.A(_17954_),
    .B(net1790),
    .Y(_18881_));
 BUFx2_ASAP7_75t_R input45 (.A(net4141),
    .Y(net45));
 NAND2x2_ASAP7_75t_R _27396_ (.A(net3204),
    .B(net1790),
    .Y(_18883_));
 BUFx2_ASAP7_75t_R input44 (.A(net4121),
    .Y(net44));
 AO21x1_ASAP7_75t_R _27398_ (.A1(net3212),
    .A2(_18883_),
    .B(net2446),
    .Y(_18885_));
 AO21x1_ASAP7_75t_R _27399_ (.A1(net3306),
    .A2(net1068),
    .B(net2446),
    .Y(_18886_));
 AND3x1_ASAP7_75t_R _27400_ (.A(_18880_),
    .B(_18885_),
    .C(_18886_),
    .Y(_18887_));
 NAND2x1_ASAP7_75t_R _27401_ (.A(net3343),
    .B(net2163),
    .Y(_18888_));
 NAND2x1_ASAP7_75t_R _27402_ (.A(_18888_),
    .B(_18160_),
    .Y(_18889_));
 NAND2x1_ASAP7_75t_R _27403_ (.A(net3192),
    .B(_18860_),
    .Y(_18890_));
 BUFx2_ASAP7_75t_R input43 (.A(net3969),
    .Y(net43));
 AO21x1_ASAP7_75t_R _27405_ (.A1(net2757),
    .A2(net1529),
    .B(_18156_),
    .Y(_18892_));
 NAND2x1_ASAP7_75t_R _27406_ (.A(_18890_),
    .B(_18892_),
    .Y(_18893_));
 NOR2x1_ASAP7_75t_R _27407_ (.A(_18889_),
    .B(_18893_),
    .Y(_18894_));
 AND2x2_ASAP7_75t_R _27408_ (.A(_18887_),
    .B(_18894_),
    .Y(_18895_));
 OA21x2_ASAP7_75t_R _27409_ (.A1(_18070_),
    .A2(_18113_),
    .B(_18175_),
    .Y(_18896_));
 NOR2x1_ASAP7_75t_R _27410_ (.A(_17937_),
    .B(_18185_),
    .Y(_18897_));
 OA21x2_ASAP7_75t_R _27411_ (.A1(_18158_),
    .A2(_17925_),
    .B(_18175_),
    .Y(_18898_));
 OR3x1_ASAP7_75t_R _27412_ (.A(_18896_),
    .B(_18897_),
    .C(_18898_),
    .Y(_18899_));
 NOR2x2_ASAP7_75t_R _27413_ (.A(net1070),
    .B(_18046_),
    .Y(_18900_));
 NOR2x2_ASAP7_75t_R _27414_ (.A(net1072),
    .B(_17983_),
    .Y(_18901_));
 OA21x2_ASAP7_75t_R _27415_ (.A1(_18900_),
    .A2(_18901_),
    .B(_18165_),
    .Y(_18902_));
 AOI21x1_ASAP7_75t_R _27416_ (.A1(_18070_),
    .A2(_18165_),
    .B(_18902_),
    .Y(_18903_));
 INVx1_ASAP7_75t_R _27417_ (.A(_18166_),
    .Y(_18904_));
 NAND2x1_ASAP7_75t_R _27418_ (.A(net1542),
    .B(_18904_),
    .Y(_18905_));
 BUFx2_ASAP7_75t_R input42 (.A(net3658),
    .Y(net42));
 AO21x1_ASAP7_75t_R _27420_ (.A1(net3212),
    .A2(net1693),
    .B(_18169_),
    .Y(_18907_));
 AND2x2_ASAP7_75t_R _27421_ (.A(_18905_),
    .B(_18907_),
    .Y(_18908_));
 NAND2x1_ASAP7_75t_R _27422_ (.A(_18903_),
    .B(_18908_),
    .Y(_18909_));
 NOR2x1_ASAP7_75t_R _27423_ (.A(_18899_),
    .B(_18909_),
    .Y(_18910_));
 NAND2x2_ASAP7_75t_R _27424_ (.A(_18895_),
    .B(_18910_),
    .Y(_18911_));
 NOR2x2_ASAP7_75t_R _27425_ (.A(_18879_),
    .B(_18911_),
    .Y(_18912_));
 AO21x2_ASAP7_75t_R _27426_ (.A1(net1795),
    .A2(net2908),
    .B(_18012_),
    .Y(_18913_));
 BUFx2_ASAP7_75t_R input41 (.A(net3872),
    .Y(net41));
 AO21x1_ASAP7_75t_R _27428_ (.A1(_18883_),
    .A2(net3284),
    .B(net3216),
    .Y(_18915_));
 INVx3_ASAP7_75t_R _27429_ (.A(_18012_),
    .Y(_18916_));
 NAND2x2_ASAP7_75t_R _27430_ (.A(_18037_),
    .B(_18916_),
    .Y(_18917_));
 NAND3x2_ASAP7_75t_R _27431_ (.B(_18915_),
    .C(_18917_),
    .Y(_18918_),
    .A(_18913_));
 BUFx2_ASAP7_75t_R input40 (.A(net4016),
    .Y(net40));
 NAND2x1_ASAP7_75t_R _27433_ (.A(_18037_),
    .B(net3092),
    .Y(_18920_));
 OA21x2_ASAP7_75t_R _27434_ (.A1(_18027_),
    .A2(_17954_),
    .B(_18920_),
    .Y(_18921_));
 NOR2x1_ASAP7_75t_R _27435_ (.A(net1050),
    .B(_18024_),
    .Y(_18922_));
 NOR2x2_ASAP7_75t_R _27436_ (.A(_18036_),
    .B(net1365),
    .Y(_18923_));
 OA21x2_ASAP7_75t_R _27437_ (.A1(_18923_),
    .A2(net2844),
    .B(net3092),
    .Y(_18924_));
 NOR2x1_ASAP7_75t_R _27438_ (.A(_18922_),
    .B(_18924_),
    .Y(_18925_));
 NAND2x1_ASAP7_75t_R _27439_ (.A(_18921_),
    .B(_18925_),
    .Y(_18926_));
 NOR2x2_ASAP7_75t_R _27440_ (.A(_18918_),
    .B(_18926_),
    .Y(_18927_));
 AO21x1_ASAP7_75t_R _27441_ (.A1(_18010_),
    .A2(net2757),
    .B(_17997_),
    .Y(_18928_));
 NAND2x1_ASAP7_75t_R _27442_ (.A(_18110_),
    .B(_18006_),
    .Y(_18929_));
 NAND2x1_ASAP7_75t_R _27443_ (.A(_18901_),
    .B(_18006_),
    .Y(_18930_));
 NAND2x1_ASAP7_75t_R _27444_ (.A(net2718),
    .B(net1791),
    .Y(_18931_));
 NOR2x1_ASAP7_75t_R _27445_ (.A(_18931_),
    .B(_17997_),
    .Y(_18932_));
 INVx1_ASAP7_75t_R _27446_ (.A(_18932_),
    .Y(_18933_));
 AND4x2_ASAP7_75t_R _27447_ (.A(_18928_),
    .B(_18929_),
    .C(_18930_),
    .D(_18933_),
    .Y(_18934_));
 NAND2x1_ASAP7_75t_R _27448_ (.A(net1644),
    .B(_17961_),
    .Y(_18935_));
 AO21x1_ASAP7_75t_R _27449_ (.A1(net939),
    .A2(_18935_),
    .B(net1955),
    .Y(_18936_));
 AO21x1_ASAP7_75t_R _27450_ (.A1(net1689),
    .A2(_18022_),
    .B(net1955),
    .Y(_18937_));
 AO21x1_ASAP7_75t_R _27451_ (.A1(net1121),
    .A2(_18057_),
    .B(net1955),
    .Y(_18938_));
 AND3x2_ASAP7_75t_R _27452_ (.A(_18936_),
    .B(_18937_),
    .C(_18938_),
    .Y(_18939_));
 NAND3x2_ASAP7_75t_R _27453_ (.B(_18934_),
    .C(_18939_),
    .Y(_18940_),
    .A(_18927_));
 INVx2_ASAP7_75t_R _27454_ (.A(net3200),
    .Y(_18941_));
 AOI21x1_ASAP7_75t_R _27455_ (.A1(net1145),
    .A2(_17980_),
    .B(_18074_),
    .Y(_18942_));
 OA21x2_ASAP7_75t_R _27456_ (.A1(_18923_),
    .A2(_18869_),
    .B(_18941_),
    .Y(_18943_));
 AOI211x1_ASAP7_75t_R _27457_ (.A1(_18941_),
    .A2(_18113_),
    .B(_18942_),
    .C(_18943_),
    .Y(_18944_));
 AO21x1_ASAP7_75t_R _27458_ (.A1(net1349),
    .A2(_17987_),
    .B(net1908),
    .Y(_18945_));
 AO21x1_ASAP7_75t_R _27459_ (.A1(net3191),
    .A2(net1068),
    .B(net1907),
    .Y(_18946_));
 NAND2x1_ASAP7_75t_R _27460_ (.A(net3220),
    .B(_18069_),
    .Y(_18947_));
 AND3x1_ASAP7_75t_R _27461_ (.A(_18945_),
    .B(_18946_),
    .C(_18947_),
    .Y(_18948_));
 AND2x2_ASAP7_75t_R _27462_ (.A(_18944_),
    .B(_18948_),
    .Y(_18949_));
 BUFx2_ASAP7_75t_R input39 (.A(net4153),
    .Y(net39));
 AOI211x1_ASAP7_75t_R _27464_ (.A1(net1061),
    .A2(net1644),
    .B(net2057),
    .C(net2303),
    .Y(_18951_));
 INVx4_ASAP7_75t_R _27465_ (.A(_18054_),
    .Y(_18952_));
 OA21x2_ASAP7_75t_R _27466_ (.A1(net3091),
    .A2(_18901_),
    .B(_18952_),
    .Y(_18953_));
 NOR2x1_ASAP7_75t_R _27467_ (.A(_18951_),
    .B(_18953_),
    .Y(_18954_));
 AO21x1_ASAP7_75t_R _27468_ (.A1(net3306),
    .A2(net1068),
    .B(net2303),
    .Y(_18955_));
 OA21x2_ASAP7_75t_R _27469_ (.A1(net3213),
    .A2(net2303),
    .B(_18955_),
    .Y(_18956_));
 NAND2x1_ASAP7_75t_R _27470_ (.A(_18954_),
    .B(_18956_),
    .Y(_18957_));
 NAND2x2_ASAP7_75t_R _27471_ (.A(net3366),
    .B(net1231),
    .Y(_18958_));
 AO21x1_ASAP7_75t_R _27472_ (.A1(net3306),
    .A2(_18958_),
    .B(net3303),
    .Y(_18959_));
 OA21x2_ASAP7_75t_R _27473_ (.A1(_18022_),
    .A2(net3303),
    .B(_18959_),
    .Y(_18960_));
 NOR2x1_ASAP7_75t_R _27474_ (.A(net1074),
    .B(_18039_),
    .Y(_18961_));
 NOR2x2_ASAP7_75t_R _27475_ (.A(_18039_),
    .B(net3199),
    .Y(_18962_));
 AOI221x1_ASAP7_75t_R _27476_ (.A1(_18040_),
    .A2(net1858),
    .B1(_18164_),
    .B2(_18961_),
    .C(_18962_),
    .Y(_18963_));
 NAND2x1_ASAP7_75t_R _27477_ (.A(_18960_),
    .B(_18963_),
    .Y(_18964_));
 NOR2x1_ASAP7_75t_R _27478_ (.A(_18957_),
    .B(_18964_),
    .Y(_18965_));
 NAND2x1_ASAP7_75t_R _27479_ (.A(_18949_),
    .B(_18965_),
    .Y(_18966_));
 NOR2x2_ASAP7_75t_R _27480_ (.A(_18966_),
    .B(_18940_),
    .Y(_18967_));
 NAND3x2_ASAP7_75t_R _27481_ (.B(_18912_),
    .C(_18967_),
    .Y(_18968_),
    .A(_17974_));
 XNOR2x2_ASAP7_75t_R _27482_ (.A(_18852_),
    .B(_18968_),
    .Y(_18969_));
 NOR2x2_ASAP7_75t_R _27483_ (.A(_18969_),
    .B(_18757_),
    .Y(_18970_));
 XOR2x2_ASAP7_75t_R _27484_ (.A(_18968_),
    .B(_18852_),
    .Y(_18971_));
 NOR2x1_ASAP7_75t_R _27485_ (.A(_18232_),
    .B(_18971_),
    .Y(_18972_));
 BUFx2_ASAP7_75t_R input38 (.A(net4143),
    .Y(net38));
 BUFx2_ASAP7_75t_R input37 (.A(net3793),
    .Y(net37));
 NAND2x2_ASAP7_75t_R _27488_ (.A(_18637_),
    .B(_18558_),
    .Y(_18975_));
 AO21x1_ASAP7_75t_R _27489_ (.A1(_18617_),
    .A2(_18975_),
    .B(net2394),
    .Y(_18976_));
 OA21x2_ASAP7_75t_R _27490_ (.A1(net2394),
    .A2(net3379),
    .B(_18976_),
    .Y(_18977_));
 BUFx2_ASAP7_75t_R input36 (.A(net3966),
    .Y(net36));
 BUFx2_ASAP7_75t_R input35 (.A(net4155),
    .Y(net35));
 BUFx2_ASAP7_75t_R input34 (.A(net4169),
    .Y(net34));
 AO21x1_ASAP7_75t_R _27494_ (.A1(net2089),
    .A2(_18680_),
    .B(net3324),
    .Y(_18981_));
 OA21x2_ASAP7_75t_R _27495_ (.A1(net1823),
    .A2(net3324),
    .B(_18981_),
    .Y(_18982_));
 NAND2x1_ASAP7_75t_R _27496_ (.A(_18977_),
    .B(_18982_),
    .Y(_18983_));
 BUFx2_ASAP7_75t_R input33 (.A(net4035),
    .Y(net33));
 BUFx2_ASAP7_75t_R input32 (.A(net4051),
    .Y(net32));
 BUFx2_ASAP7_75t_R input31 (.A(net4021),
    .Y(net31));
 AO21x1_ASAP7_75t_R _27500_ (.A1(net1388),
    .A2(_18548_),
    .B(net2693),
    .Y(_18987_));
 AO21x1_ASAP7_75t_R _27501_ (.A1(_18627_),
    .A2(net2421),
    .B(net2693),
    .Y(_18988_));
 NAND2x1_ASAP7_75t_R _27502_ (.A(_18987_),
    .B(_18988_),
    .Y(_18989_));
 INVx1_ASAP7_75t_R _27503_ (.A(_18989_),
    .Y(_18990_));
 NAND2x1_ASAP7_75t_R _27504_ (.A(_18610_),
    .B(_18725_),
    .Y(_18991_));
 NAND2x2_ASAP7_75t_R _27505_ (.A(_18565_),
    .B(net3004),
    .Y(_18992_));
 BUFx2_ASAP7_75t_R input30 (.A(net4145),
    .Y(net30));
 BUFx2_ASAP7_75t_R input29 (.A(net4165),
    .Y(net29));
 AO21x1_ASAP7_75t_R _27508_ (.A1(net2177),
    .A2(_18992_),
    .B(net2317),
    .Y(_18995_));
 NAND2x1_ASAP7_75t_R _27509_ (.A(_18991_),
    .B(_18995_),
    .Y(_18996_));
 INVx1_ASAP7_75t_R _27510_ (.A(_18617_),
    .Y(_18997_));
 NAND2x1_ASAP7_75t_R _27511_ (.A(_18997_),
    .B(_18725_),
    .Y(_18998_));
 AO21x1_ASAP7_75t_R _27512_ (.A1(_18651_),
    .A2(net2421),
    .B(net2317),
    .Y(_18999_));
 NAND2x1_ASAP7_75t_R _27513_ (.A(_18998_),
    .B(_18999_),
    .Y(_19000_));
 NOR2x1_ASAP7_75t_R _27514_ (.A(_18996_),
    .B(_19000_),
    .Y(_19001_));
 NAND2x1_ASAP7_75t_R _27515_ (.A(_18990_),
    .B(_19001_),
    .Y(_19002_));
 NOR2x2_ASAP7_75t_R _27516_ (.A(_18983_),
    .B(_19002_),
    .Y(_19003_));
 NAND2x1_ASAP7_75t_R _27517_ (.A(_18637_),
    .B(net2555),
    .Y(_19004_));
 BUFx2_ASAP7_75t_R input28 (.A(net3907),
    .Y(net28));
 AO21x1_ASAP7_75t_R _27519_ (.A1(_18621_),
    .A2(_19004_),
    .B(net2546),
    .Y(_19006_));
 NOR2x1_ASAP7_75t_R _27520_ (.A(_18530_),
    .B(net2631),
    .Y(_19007_));
 NAND2x1_ASAP7_75t_R _27521_ (.A(_19007_),
    .B(_18683_),
    .Y(_19008_));
 BUFx2_ASAP7_75t_R input27 (.A(net3990),
    .Y(net27));
 AO21x1_ASAP7_75t_R _27523_ (.A1(_18651_),
    .A2(net2405),
    .B(net2546),
    .Y(_19010_));
 AND3x1_ASAP7_75t_R _27524_ (.A(_19006_),
    .B(_19008_),
    .C(_19010_),
    .Y(_19011_));
 NOR2x2_ASAP7_75t_R _27525_ (.A(net1472),
    .B(net1729),
    .Y(_19012_));
 INVx2_ASAP7_75t_R _27526_ (.A(_19012_),
    .Y(_19013_));
 AO21x1_ASAP7_75t_R _27527_ (.A1(_18627_),
    .A2(_19013_),
    .B(net2304),
    .Y(_19014_));
 AO21x1_ASAP7_75t_R _27528_ (.A1(net1388),
    .A2(net1569),
    .B(net2304),
    .Y(_19015_));
 NOR2x1_ASAP7_75t_R _27529_ (.A(_18695_),
    .B(_18516_),
    .Y(_19016_));
 INVx1_ASAP7_75t_R _27530_ (.A(_19016_),
    .Y(_19017_));
 AND3x1_ASAP7_75t_R _27531_ (.A(_19014_),
    .B(_19015_),
    .C(_19017_),
    .Y(_19018_));
 AND2x2_ASAP7_75t_R _27532_ (.A(_19011_),
    .B(_19018_),
    .Y(_19019_));
 BUFx2_ASAP7_75t_R input26 (.A(net3875),
    .Y(net26));
 AO21x1_ASAP7_75t_R _27534_ (.A1(net2633),
    .A2(net2421),
    .B(_18666_),
    .Y(_19021_));
 BUFx2_ASAP7_75t_R input25 (.A(net4047),
    .Y(net25));
 AO21x1_ASAP7_75t_R _27536_ (.A1(net1307),
    .A2(net1388),
    .B(_18666_),
    .Y(_19023_));
 NOR2x1_ASAP7_75t_R _27537_ (.A(net1569),
    .B(_18666_),
    .Y(_19024_));
 INVx1_ASAP7_75t_R _27538_ (.A(_19024_),
    .Y(_19025_));
 NAND3x2_ASAP7_75t_R _27539_ (.B(_19023_),
    .C(_19025_),
    .Y(_19026_),
    .A(_19021_));
 BUFx2_ASAP7_75t_R input24 (.A(net4179),
    .Y(net24));
 AOI211x1_ASAP7_75t_R _27541_ (.A1(net3090),
    .A2(net3380),
    .B(_18655_),
    .C(_18536_),
    .Y(_19028_));
 INVx1_ASAP7_75t_R _27542_ (.A(_19028_),
    .Y(_19029_));
 AO21x1_ASAP7_75t_R _27543_ (.A1(net2177),
    .A2(_18992_),
    .B(_18655_),
    .Y(_19030_));
 NOR2x2_ASAP7_75t_R _27544_ (.A(net2993),
    .B(_18670_),
    .Y(_19031_));
 NAND2x2_ASAP7_75t_R _27545_ (.A(net2992),
    .B(_19031_),
    .Y(_19032_));
 NAND3x2_ASAP7_75t_R _27546_ (.B(_19030_),
    .C(_19032_),
    .Y(_19033_),
    .A(_19029_));
 NOR2x2_ASAP7_75t_R _27547_ (.A(_19026_),
    .B(_19033_),
    .Y(_19034_));
 NAND3x2_ASAP7_75t_R _27548_ (.B(_19019_),
    .C(_19034_),
    .Y(_19035_),
    .A(_19003_));
 NAND2x2_ASAP7_75t_R _27549_ (.A(net2309),
    .B(_18558_),
    .Y(_19036_));
 BUFx2_ASAP7_75t_R input23 (.A(net4119),
    .Y(net23));
 AO21x1_ASAP7_75t_R _27551_ (.A1(_18584_),
    .A2(_19036_),
    .B(net2414),
    .Y(_19038_));
 BUFx2_ASAP7_75t_R input22 (.A(net4117),
    .Y(net22));
 AO21x2_ASAP7_75t_R _27553_ (.A1(net2760),
    .A2(net2433),
    .B(net2414),
    .Y(_19040_));
 NAND2x2_ASAP7_75t_R _27554_ (.A(_18675_),
    .B(_18612_),
    .Y(_19041_));
 NAND3x2_ASAP7_75t_R _27555_ (.B(_19040_),
    .C(_19041_),
    .Y(_19042_),
    .A(_19038_));
 BUFx2_ASAP7_75t_R input21 (.A(net4189),
    .Y(net21));
 OR3x4_ASAP7_75t_R _27557_ (.A(net2615),
    .B(net1565),
    .C(_18555_),
    .Y(_19044_));
 AO21x1_ASAP7_75t_R _27558_ (.A1(_18586_),
    .A2(net2631),
    .B(net2615),
    .Y(_19045_));
 INVx2_ASAP7_75t_R _27559_ (.A(_18604_),
    .Y(_19046_));
 NAND2x2_ASAP7_75t_R _27560_ (.A(_18537_),
    .B(_19046_),
    .Y(_19047_));
 NAND3x2_ASAP7_75t_R _27561_ (.B(_19045_),
    .C(_19047_),
    .Y(_19048_),
    .A(_19044_));
 NOR2x2_ASAP7_75t_R _27562_ (.A(_19042_),
    .B(_19048_),
    .Y(_19049_));
 INVx1_ASAP7_75t_R _27563_ (.A(_19049_),
    .Y(_19050_));
 BUFx2_ASAP7_75t_R input20 (.A(net4139),
    .Y(net20));
 AO21x1_ASAP7_75t_R _27565_ (.A1(_18553_),
    .A2(net2405),
    .B(net2620),
    .Y(_19052_));
 OAI21x1_ASAP7_75t_R _27566_ (.A1(net2620),
    .A2(_18687_),
    .B(_19052_),
    .Y(_19053_));
 NOR2x1_ASAP7_75t_R _27567_ (.A(_18992_),
    .B(_18641_),
    .Y(_19054_));
 OR3x1_ASAP7_75t_R _27568_ (.A(_18642_),
    .B(_18645_),
    .C(_19054_),
    .Y(_19055_));
 NOR2x2_ASAP7_75t_R _27569_ (.A(_19053_),
    .B(_19055_),
    .Y(_19056_));
 NOR2x2_ASAP7_75t_R _27570_ (.A(net1726),
    .B(_18637_),
    .Y(_19057_));
 NOR2x2_ASAP7_75t_R _27571_ (.A(_18523_),
    .B(_18634_),
    .Y(_19058_));
 NAND2x1_ASAP7_75t_R _27572_ (.A(net2735),
    .B(_19058_),
    .Y(_19059_));
 NOR2x2_ASAP7_75t_R _27573_ (.A(_18514_),
    .B(_18581_),
    .Y(_19060_));
 NAND2x1_ASAP7_75t_R _27574_ (.A(_19060_),
    .B(_19058_),
    .Y(_19061_));
 NAND2x1_ASAP7_75t_R _27575_ (.A(_18650_),
    .B(_19058_),
    .Y(_19062_));
 AND3x1_ASAP7_75t_R _27576_ (.A(_19059_),
    .B(_19061_),
    .C(_19062_),
    .Y(_19063_));
 AO21x1_ASAP7_75t_R _27577_ (.A1(net3090),
    .A2(_18554_),
    .B(_18536_),
    .Y(_19064_));
 NAND2x1_ASAP7_75t_R _27578_ (.A(_18554_),
    .B(net2555),
    .Y(_19065_));
 BUFx2_ASAP7_75t_R input19 (.A(net4173),
    .Y(net19));
 AO21x1_ASAP7_75t_R _27580_ (.A1(_19064_),
    .A2(_19065_),
    .B(_18625_),
    .Y(_19067_));
 AND2x2_ASAP7_75t_R _27581_ (.A(_19063_),
    .B(_19067_),
    .Y(_19068_));
 NAND2x1_ASAP7_75t_R _27582_ (.A(_19056_),
    .B(_19068_),
    .Y(_19069_));
 NOR2x1_ASAP7_75t_R _27583_ (.A(_19050_),
    .B(_19069_),
    .Y(_19070_));
 AO21x1_ASAP7_75t_R _27584_ (.A1(net1404),
    .A2(net3215),
    .B(net2479),
    .Y(_19071_));
 INVx1_ASAP7_75t_R _27585_ (.A(_19071_),
    .Y(_19072_));
 NAND2x2_ASAP7_75t_R _27586_ (.A(_18565_),
    .B(_18515_),
    .Y(_19073_));
 BUFx2_ASAP7_75t_R input18 (.A(net4061),
    .Y(net18));
 AO21x1_ASAP7_75t_R _27588_ (.A1(_19073_),
    .A2(_18992_),
    .B(_18545_),
    .Y(_19075_));
 INVx1_ASAP7_75t_R _27589_ (.A(_19075_),
    .Y(_19076_));
 BUFx2_ASAP7_75t_R input17 (.A(net4208),
    .Y(net17));
 NOR2x2_ASAP7_75t_R _27591_ (.A(_19013_),
    .B(net2479),
    .Y(_19078_));
 NOR3x2_ASAP7_75t_R _27592_ (.B(_19076_),
    .C(_19078_),
    .Y(_19079_),
    .A(_19072_));
 AO21x1_ASAP7_75t_R _27593_ (.A1(net2177),
    .A2(_18623_),
    .B(_18525_),
    .Y(_19080_));
 AO21x1_ASAP7_75t_R _27594_ (.A1(net1307),
    .A2(net1388),
    .B(_18525_),
    .Y(_19081_));
 AND2x2_ASAP7_75t_R _27595_ (.A(_19080_),
    .B(_19081_),
    .Y(_19082_));
 NOR2x2_ASAP7_75t_R _27596_ (.A(_18581_),
    .B(_18674_),
    .Y(_19083_));
 OAI21x1_ASAP7_75t_R _27597_ (.A1(_18636_),
    .A2(_19083_),
    .B(_18524_),
    .Y(_19084_));
 NAND2x1_ASAP7_75t_R _27598_ (.A(net2690),
    .B(_18638_),
    .Y(_19085_));
 NAND2x1_ASAP7_75t_R _27599_ (.A(_19012_),
    .B(net2690),
    .Y(_19086_));
 AND3x2_ASAP7_75t_R _27600_ (.A(_19084_),
    .B(_19085_),
    .C(_19086_),
    .Y(_19087_));
 NAND3x1_ASAP7_75t_R _27601_ (.A(_19079_),
    .B(_19082_),
    .C(_19087_),
    .Y(_19088_));
 BUFx2_ASAP7_75t_R input16 (.A(net3915),
    .Y(net16));
 OAI21x1_ASAP7_75t_R _27603_ (.A1(_18585_),
    .A2(net2991),
    .B(_18592_),
    .Y(_19090_));
 OAI21x1_ASAP7_75t_R _27604_ (.A1(net1404),
    .A2(_18588_),
    .B(_19090_),
    .Y(_19091_));
 NOR2x2_ASAP7_75t_R _27605_ (.A(_18588_),
    .B(_19073_),
    .Y(_19092_));
 INVx1_ASAP7_75t_R _27606_ (.A(_18547_),
    .Y(_19093_));
 OA21x2_ASAP7_75t_R _27607_ (.A1(_18672_),
    .A2(_19093_),
    .B(_18592_),
    .Y(_19094_));
 NOR3x2_ASAP7_75t_R _27608_ (.B(_19092_),
    .C(_19094_),
    .Y(_19095_),
    .A(_19091_));
 BUFx2_ASAP7_75t_R input15 (.A(net3892),
    .Y(net15));
 AO21x1_ASAP7_75t_R _27610_ (.A1(net1404),
    .A2(net2633),
    .B(_18569_),
    .Y(_19097_));
 AND2x2_ASAP7_75t_R _27611_ (.A(_18577_),
    .B(_19097_),
    .Y(_19098_));
 AOI211x1_ASAP7_75t_R _27612_ (.A1(net1473),
    .A2(net3380),
    .B(_18569_),
    .C(_18536_),
    .Y(_19099_));
 NOR2x1_ASAP7_75t_R _27613_ (.A(_18515_),
    .B(_18571_),
    .Y(_19100_));
 NOR2x1_ASAP7_75t_R _27614_ (.A(_19099_),
    .B(_19100_),
    .Y(_19101_));
 NAND3x1_ASAP7_75t_R _27615_ (.A(_19095_),
    .B(_19098_),
    .C(_19101_),
    .Y(_19102_));
 NOR2x1_ASAP7_75t_R _27616_ (.A(_19088_),
    .B(_19102_),
    .Y(_19103_));
 NAND2x1_ASAP7_75t_R _27617_ (.A(_19070_),
    .B(_19103_),
    .Y(_19104_));
 NOR2x2_ASAP7_75t_R _27618_ (.A(_19035_),
    .B(_19104_),
    .Y(_19105_));
 NAND2x1_ASAP7_75t_R _27619_ (.A(_19105_),
    .B(_18742_),
    .Y(_19106_));
 OA21x2_ASAP7_75t_R _27620_ (.A1(_18690_),
    .A2(_18585_),
    .B(_18524_),
    .Y(_19107_));
 OAI21x1_ASAP7_75t_R _27621_ (.A1(_19060_),
    .A2(_18638_),
    .B(_18524_),
    .Y(_19108_));
 NAND2x1_ASAP7_75t_R _27622_ (.A(_19108_),
    .B(_19084_),
    .Y(_19109_));
 NOR2x1_ASAP7_75t_R _27623_ (.A(_19107_),
    .B(_19109_),
    .Y(_19110_));
 AO21x1_ASAP7_75t_R _27624_ (.A1(_18594_),
    .A2(_18680_),
    .B(_18525_),
    .Y(_19111_));
 INVx1_ASAP7_75t_R _27625_ (.A(_19111_),
    .Y(_19112_));
 NAND2x1_ASAP7_75t_R _27626_ (.A(_18524_),
    .B(_18590_),
    .Y(_19113_));
 NOR2x2_ASAP7_75t_R _27627_ (.A(net1009),
    .B(net1563),
    .Y(_19114_));
 OAI21x1_ASAP7_75t_R _27628_ (.A1(_19114_),
    .A2(_18694_),
    .B(_18524_),
    .Y(_19115_));
 NAND2x1_ASAP7_75t_R _27629_ (.A(_19113_),
    .B(_19115_),
    .Y(_19116_));
 NOR2x1_ASAP7_75t_R _27630_ (.A(_19112_),
    .B(_19116_),
    .Y(_19117_));
 OR3x1_ASAP7_75t_R _27631_ (.A(_18602_),
    .B(_18633_),
    .C(net2887),
    .Y(_19118_));
 AND4x2_ASAP7_75t_R _27632_ (.A(_19110_),
    .B(_19117_),
    .C(net2479),
    .D(_19118_),
    .Y(_19119_));
 NAND3x2_ASAP7_75t_R _27633_ (.B(net2697),
    .C(net2869),
    .Y(_19120_),
    .A(_19119_));
 INVx3_ASAP7_75t_R _27634_ (.A(_19120_),
    .Y(_19121_));
 INVx1_ASAP7_75t_R _27635_ (.A(_19003_),
    .Y(_19122_));
 NAND2x1_ASAP7_75t_R _27636_ (.A(_19034_),
    .B(_19019_),
    .Y(_19123_));
 NOR2x2_ASAP7_75t_R _27637_ (.A(_19122_),
    .B(_19123_),
    .Y(_19124_));
 INVx1_ASAP7_75t_R _27638_ (.A(_19079_),
    .Y(_19125_));
 NAND2x1_ASAP7_75t_R _27639_ (.A(_19082_),
    .B(_19087_),
    .Y(_19126_));
 NOR2x1_ASAP7_75t_R _27640_ (.A(_19125_),
    .B(_19126_),
    .Y(_19127_));
 NAND2x1_ASAP7_75t_R _27641_ (.A(_19098_),
    .B(_19101_),
    .Y(_19128_));
 INVx1_ASAP7_75t_R _27642_ (.A(_19095_),
    .Y(_19129_));
 NOR2x1_ASAP7_75t_R _27643_ (.A(_19128_),
    .B(_19129_),
    .Y(_19130_));
 NAND2x1_ASAP7_75t_R _27644_ (.A(_19127_),
    .B(_19130_),
    .Y(_19131_));
 NAND3x1_ASAP7_75t_R _27645_ (.A(_19049_),
    .B(_19068_),
    .C(_19056_),
    .Y(_19132_));
 NOR2x1_ASAP7_75t_R _27646_ (.A(_19131_),
    .B(_19132_),
    .Y(_19133_));
 NAND2x2_ASAP7_75t_R _27647_ (.A(_19124_),
    .B(_19133_),
    .Y(_19134_));
 NOR2x1_ASAP7_75t_R _27648_ (.A(_18646_),
    .B(_18640_),
    .Y(_19135_));
 NAND2x1_ASAP7_75t_R _27649_ (.A(_18630_),
    .B(_19135_),
    .Y(_19136_));
 INVx1_ASAP7_75t_R _27650_ (.A(_18619_),
    .Y(_19137_));
 NOR2x1_ASAP7_75t_R _27651_ (.A(_19136_),
    .B(_19137_),
    .Y(_19138_));
 NAND2x1_ASAP7_75t_R _27652_ (.A(_18598_),
    .B(_19138_),
    .Y(_19139_));
 NAND3x1_ASAP7_75t_R _27653_ (.A(_18662_),
    .B(_18677_),
    .C(_18668_),
    .Y(_19140_));
 NOR2x1_ASAP7_75t_R _27654_ (.A(_19140_),
    .B(_18706_),
    .Y(_19141_));
 NAND2x2_ASAP7_75t_R _27655_ (.A(_18739_),
    .B(_19141_),
    .Y(_19142_));
 NOR2x2_ASAP7_75t_R _27656_ (.A(_19139_),
    .B(_19142_),
    .Y(_19143_));
 OAI21x1_ASAP7_75t_R _27657_ (.A1(_19121_),
    .A2(_19134_),
    .B(_19143_),
    .Y(_19144_));
 NAND2x2_ASAP7_75t_R _27658_ (.A(_19106_),
    .B(_19144_),
    .Y(_19145_));
 OAI21x1_ASAP7_75t_R _27659_ (.A1(net1199),
    .A2(_18273_),
    .B(_18421_),
    .Y(_19146_));
 NAND2x1_ASAP7_75t_R _27660_ (.A(_18255_),
    .B(_18249_),
    .Y(_19147_));
 NOR2x1_ASAP7_75t_R _27661_ (.A(_19146_),
    .B(_19147_),
    .Y(_19148_));
 OA21x2_ASAP7_75t_R _27662_ (.A1(_18254_),
    .A2(_18401_),
    .B(_18416_),
    .Y(_19149_));
 INVx3_ASAP7_75t_R _27663_ (.A(_18442_),
    .Y(_19150_));
 NAND2x1_ASAP7_75t_R _27664_ (.A(_19150_),
    .B(_18416_),
    .Y(_19151_));
 AO21x1_ASAP7_75t_R _27665_ (.A1(net1755),
    .A2(_18453_),
    .B(_18266_),
    .Y(_19152_));
 NAND2x1_ASAP7_75t_R _27666_ (.A(_19151_),
    .B(_19152_),
    .Y(_19153_));
 NOR2x1_ASAP7_75t_R _27667_ (.A(_19149_),
    .B(_19153_),
    .Y(_19154_));
 NAND2x1_ASAP7_75t_R _27668_ (.A(_19148_),
    .B(_19154_),
    .Y(_19155_));
 NOR2x2_ASAP7_75t_R _27669_ (.A(net2498),
    .B(_18467_),
    .Y(_19156_));
 OA21x2_ASAP7_75t_R _27670_ (.A1(_19156_),
    .A2(_18444_),
    .B(_18434_),
    .Y(_19157_));
 NOR2x1_ASAP7_75t_R _27671_ (.A(_19157_),
    .B(_18435_),
    .Y(_19158_));
 AOI211x1_ASAP7_75t_R _27672_ (.A1(net2999),
    .A2(_18237_),
    .B(_18428_),
    .C(net2977),
    .Y(_19159_));
 NOR2x2_ASAP7_75t_R _27673_ (.A(_18240_),
    .B(net2009),
    .Y(_19160_));
 OA21x2_ASAP7_75t_R _27674_ (.A1(_19160_),
    .A2(_18468_),
    .B(_18434_),
    .Y(_19161_));
 NOR2x1_ASAP7_75t_R _27675_ (.A(_19159_),
    .B(_19161_),
    .Y(_19162_));
 NOR2x1_ASAP7_75t_R _27676_ (.A(net3326),
    .B(net2498),
    .Y(_19163_));
 INVx1_ASAP7_75t_R _27677_ (.A(_19163_),
    .Y(_19164_));
 NOR2x1_ASAP7_75t_R _27678_ (.A(_18439_),
    .B(_19164_),
    .Y(_19165_));
 AOI21x1_ASAP7_75t_R _27679_ (.A1(_18394_),
    .A2(_18381_),
    .B(_18439_),
    .Y(_19166_));
 NOR2x1_ASAP7_75t_R _27680_ (.A(_19165_),
    .B(_19166_),
    .Y(_19167_));
 NAND3x1_ASAP7_75t_R _27681_ (.A(_19158_),
    .B(_19162_),
    .C(_19167_),
    .Y(_19168_));
 NOR2x1_ASAP7_75t_R _27682_ (.A(_19155_),
    .B(_19168_),
    .Y(_19169_));
 NOR2x2_ASAP7_75t_R _27683_ (.A(net2973),
    .B(_18490_),
    .Y(_19170_));
 NAND2x2_ASAP7_75t_R _27684_ (.A(net2602),
    .B(_18238_),
    .Y(_19171_));
 BUFx2_ASAP7_75t_R input14 (.A(net4181),
    .Y(net14));
 AOI21x1_ASAP7_75t_R _27686_ (.A1(net2176),
    .A2(net1606),
    .B(net2595),
    .Y(_19173_));
 NAND2x2_ASAP7_75t_R _27687_ (.A(_18237_),
    .B(_18313_),
    .Y(_19174_));
 AOI21x1_ASAP7_75t_R _27688_ (.A1(_19174_),
    .A2(net2965),
    .B(net2994),
    .Y(_19175_));
 AOI211x1_ASAP7_75t_R _27689_ (.A1(_19170_),
    .A2(net2972),
    .B(_19173_),
    .C(_19175_),
    .Y(_19176_));
 AO21x1_ASAP7_75t_R _27690_ (.A1(net2347),
    .A2(_18327_),
    .B(_18479_),
    .Y(_19177_));
 NAND2x1_ASAP7_75t_R _27691_ (.A(_18498_),
    .B(_19177_),
    .Y(_19178_));
 BUFx2_ASAP7_75t_R input13 (.A(net4157),
    .Y(net13));
 AO21x2_ASAP7_75t_R _27693_ (.A1(_18316_),
    .A2(_18394_),
    .B(_18479_),
    .Y(_19180_));
 AO21x1_ASAP7_75t_R _27694_ (.A1(net2251),
    .A2(net2965),
    .B(_18479_),
    .Y(_19181_));
 NAND2x1_ASAP7_75t_R _27695_ (.A(_19180_),
    .B(_19181_),
    .Y(_19182_));
 NOR2x1_ASAP7_75t_R _27696_ (.A(_19178_),
    .B(_19182_),
    .Y(_19183_));
 NAND2x1_ASAP7_75t_R _27697_ (.A(_19176_),
    .B(_19183_),
    .Y(_19184_));
 INVx4_ASAP7_75t_R _27698_ (.A(_18456_),
    .Y(_19185_));
 NAND2x1_ASAP7_75t_R _27699_ (.A(net2533),
    .B(_19185_),
    .Y(_19186_));
 AO21x1_ASAP7_75t_R _27700_ (.A1(net2106),
    .A2(net3181),
    .B(_18456_),
    .Y(_19187_));
 NAND2x1_ASAP7_75t_R _27701_ (.A(_19186_),
    .B(_19187_),
    .Y(_19188_));
 NAND2x1_ASAP7_75t_R _27702_ (.A(_19163_),
    .B(_19185_),
    .Y(_19189_));
 AO21x1_ASAP7_75t_R _27703_ (.A1(net2964),
    .A2(_18383_),
    .B(_18456_),
    .Y(_19190_));
 NAND2x1_ASAP7_75t_R _27704_ (.A(_19189_),
    .B(_19190_),
    .Y(_19191_));
 NOR2x1_ASAP7_75t_R _27705_ (.A(_19188_),
    .B(_19191_),
    .Y(_19192_));
 AO21x1_ASAP7_75t_R _27706_ (.A1(_18381_),
    .A2(net1483),
    .B(net3312),
    .Y(_19193_));
 BUFx2_ASAP7_75t_R input12 (.A(net4203),
    .Y(net12));
 AO21x1_ASAP7_75t_R _27708_ (.A1(net2250),
    .A2(_18351_),
    .B(net3312),
    .Y(_19195_));
 AO21x1_ASAP7_75t_R _27709_ (.A1(_18305_),
    .A2(net2438),
    .B(net3312),
    .Y(_19196_));
 AND3x1_ASAP7_75t_R _27710_ (.A(_19193_),
    .B(_19195_),
    .C(_19196_),
    .Y(_19197_));
 NAND2x1_ASAP7_75t_R _27711_ (.A(_19192_),
    .B(_19197_),
    .Y(_19198_));
 NOR2x2_ASAP7_75t_R _27712_ (.A(_19184_),
    .B(_19198_),
    .Y(_19199_));
 NAND2x2_ASAP7_75t_R _27713_ (.A(_19169_),
    .B(_19199_),
    .Y(_19200_));
 AO21x1_ASAP7_75t_R _27714_ (.A1(net2473),
    .A2(net2250),
    .B(_18330_),
    .Y(_19201_));
 INVx3_ASAP7_75t_R _27715_ (.A(net2439),
    .Y(_19202_));
 NAND2x1_ASAP7_75t_R _27716_ (.A(_19202_),
    .B(_18345_),
    .Y(_19203_));
 AND2x2_ASAP7_75t_R _27717_ (.A(_19201_),
    .B(_19203_),
    .Y(_19204_));
 NOR2x2_ASAP7_75t_R _27718_ (.A(net2498),
    .B(net2968),
    .Y(_19205_));
 OAI21x1_ASAP7_75t_R _27719_ (.A1(_18343_),
    .A2(_19205_),
    .B(_18345_),
    .Y(_19206_));
 AOI21x1_ASAP7_75t_R _27720_ (.A1(net3248),
    .A2(net2043),
    .B(_18318_),
    .Y(_19207_));
 AOI21x1_ASAP7_75t_R _27721_ (.A1(net2974),
    .A2(net2095),
    .B(_18318_),
    .Y(_19208_));
 NOR2x1_ASAP7_75t_R _27722_ (.A(_19207_),
    .B(_19208_),
    .Y(_19209_));
 NAND3x1_ASAP7_75t_R _27723_ (.A(_19204_),
    .B(_19206_),
    .C(_19209_),
    .Y(_19210_));
 AO21x1_ASAP7_75t_R _27724_ (.A1(net2095),
    .A2(_18327_),
    .B(net2982),
    .Y(_19211_));
 OAI21x1_ASAP7_75t_R _27725_ (.A1(net3281),
    .A2(net2669),
    .B(_18292_),
    .Y(_19212_));
 NAND2x1_ASAP7_75t_R _27726_ (.A(_18444_),
    .B(_18292_),
    .Y(_19213_));
 AND3x1_ASAP7_75t_R _27727_ (.A(_19211_),
    .B(_19212_),
    .C(_19213_),
    .Y(_19214_));
 AO21x1_ASAP7_75t_R _27728_ (.A1(net2176),
    .A2(_18327_),
    .B(_18300_),
    .Y(_19215_));
 BUFx2_ASAP7_75t_R input11 (.A(net4004),
    .Y(net11));
 AO21x1_ASAP7_75t_R _27730_ (.A1(net2671),
    .A2(net2050),
    .B(_18300_),
    .Y(_19217_));
 OAI21x1_ASAP7_75t_R _27731_ (.A1(_18309_),
    .A2(net3283),
    .B(_18303_),
    .Y(_19218_));
 AND3x1_ASAP7_75t_R _27732_ (.A(_19215_),
    .B(_19217_),
    .C(_19218_),
    .Y(_19219_));
 NAND2x1_ASAP7_75t_R _27733_ (.A(_19214_),
    .B(_19219_),
    .Y(_19220_));
 NOR2x1_ASAP7_75t_R _27734_ (.A(_19210_),
    .B(_19220_),
    .Y(_19221_));
 AO21x1_ASAP7_75t_R _27735_ (.A1(net2969),
    .A2(net2440),
    .B(_18377_),
    .Y(_19222_));
 INVx2_ASAP7_75t_R _27736_ (.A(net2250),
    .Y(_19223_));
 INVx3_ASAP7_75t_R _27737_ (.A(_18377_),
    .Y(_19224_));
 OAI21x1_ASAP7_75t_R _27738_ (.A1(_19160_),
    .A2(_19223_),
    .B(_19224_),
    .Y(_19225_));
 NAND2x1_ASAP7_75t_R _27739_ (.A(_18445_),
    .B(_19224_),
    .Y(_19226_));
 AND3x1_ASAP7_75t_R _27740_ (.A(_19222_),
    .B(_19225_),
    .C(_19226_),
    .Y(_19227_));
 BUFx2_ASAP7_75t_R input10 (.A(net4175),
    .Y(net10));
 AO21x1_ASAP7_75t_R _27742_ (.A1(net1753),
    .A2(net1821),
    .B(_18395_),
    .Y(_19229_));
 AO21x1_ASAP7_75t_R _27743_ (.A1(net2671),
    .A2(net2439),
    .B(_18395_),
    .Y(_19230_));
 NAND2x1_ASAP7_75t_R _27744_ (.A(_18468_),
    .B(_18398_),
    .Y(_19231_));
 AND3x1_ASAP7_75t_R _27745_ (.A(_19229_),
    .B(_19230_),
    .C(_19231_),
    .Y(_19232_));
 NAND2x1_ASAP7_75t_R _27746_ (.A(_19227_),
    .B(_19232_),
    .Y(_19233_));
 AO21x1_ASAP7_75t_R _27747_ (.A1(_18467_),
    .A2(net2971),
    .B(_18366_),
    .Y(_19234_));
 BUFx2_ASAP7_75t_R input9 (.A(net4107),
    .Y(net9));
 AOI21x1_ASAP7_75t_R _27749_ (.A1(net1606),
    .A2(_19234_),
    .B(_18354_),
    .Y(_19236_));
 INVx2_ASAP7_75t_R _27750_ (.A(_18354_),
    .Y(_19237_));
 OA21x2_ASAP7_75t_R _27751_ (.A1(_18482_),
    .A2(_18270_),
    .B(_19237_),
    .Y(_19238_));
 AOI211x1_ASAP7_75t_R _27752_ (.A1(net1087),
    .A2(net2990),
    .B(_18354_),
    .C(net2499),
    .Y(_19239_));
 NOR3x1_ASAP7_75t_R _27753_ (.A(_19236_),
    .B(_19238_),
    .C(_19239_),
    .Y(_19240_));
 BUFx2_ASAP7_75t_R input8 (.A(net4205),
    .Y(net8));
 AO21x1_ASAP7_75t_R _27755_ (.A1(net2635),
    .A2(net1484),
    .B(_18364_),
    .Y(_19242_));
 AO21x1_ASAP7_75t_R _27756_ (.A1(_18381_),
    .A2(net3183),
    .B(_18364_),
    .Y(_19243_));
 NAND2x1_ASAP7_75t_R _27757_ (.A(_19242_),
    .B(_19243_),
    .Y(_19244_));
 AO21x1_ASAP7_75t_R _27758_ (.A1(net2747),
    .A2(_18335_),
    .B(_18364_),
    .Y(_19245_));
 OAI21x1_ASAP7_75t_R _27759_ (.A1(_18364_),
    .A2(net1954),
    .B(_19245_),
    .Y(_19246_));
 NOR2x1_ASAP7_75t_R _27760_ (.A(_19244_),
    .B(_19246_),
    .Y(_19247_));
 NAND2x1_ASAP7_75t_R _27761_ (.A(_19240_),
    .B(_19247_),
    .Y(_19248_));
 NOR2x1_ASAP7_75t_R _27762_ (.A(_19233_),
    .B(_19248_),
    .Y(_19249_));
 NAND2x1_ASAP7_75t_R _27763_ (.A(_19221_),
    .B(_19249_),
    .Y(_19250_));
 NOR2x2_ASAP7_75t_R _27764_ (.A(_19200_),
    .B(_19250_),
    .Y(_19251_));
 NAND2x2_ASAP7_75t_R _27765_ (.A(_18279_),
    .B(_19251_),
    .Y(_19252_));
 XOR2x2_ASAP7_75t_R _27766_ (.A(_19145_),
    .B(_19252_),
    .Y(_19253_));
 OAI21x1_ASAP7_75t_R _27767_ (.A1(_18970_),
    .A2(_18972_),
    .B(_19253_),
    .Y(_19254_));
 NOR2x2_ASAP7_75t_R _27768_ (.A(_18971_),
    .B(_18757_),
    .Y(_19255_));
 NOR2x1_ASAP7_75t_R _27769_ (.A(_18232_),
    .B(_18969_),
    .Y(_19256_));
 INVx2_ASAP7_75t_R _27770_ (.A(_19252_),
    .Y(_19257_));
 XOR2x2_ASAP7_75t_R _27771_ (.A(_19145_),
    .B(_19257_),
    .Y(_19258_));
 OAI21x1_ASAP7_75t_R _27772_ (.A1(_19255_),
    .A2(_19256_),
    .B(_19258_),
    .Y(_19259_));
 BUFx2_ASAP7_75t_R input7 (.A(net4171),
    .Y(net7));
 BUFx2_ASAP7_75t_R input6 (.A(net4206),
    .Y(net6));
 AOI21x1_ASAP7_75t_R _27775_ (.A1(_19254_),
    .A2(_19259_),
    .B(net390),
    .Y(_19262_));
 OAI21x1_ASAP7_75t_R _27776_ (.A1(_18756_),
    .A2(_19262_),
    .B(_14620_),
    .Y(_19263_));
 BUFx2_ASAP7_75t_R input5 (.A(net4190),
    .Y(net5));
 NOR2x1_ASAP7_75t_R _27778_ (.A(net397),
    .B(_00914_),
    .Y(_19265_));
 OAI21x1_ASAP7_75t_R _27779_ (.A1(_19256_),
    .A2(_19255_),
    .B(_19253_),
    .Y(_19266_));
 OAI21x1_ASAP7_75t_R _27780_ (.A1(_18970_),
    .A2(_18972_),
    .B(_19258_),
    .Y(_19267_));
 BUFx2_ASAP7_75t_R input4 (.A(net4201),
    .Y(net4));
 AOI21x1_ASAP7_75t_R _27782_ (.A1(_19266_),
    .A2(_19267_),
    .B(net390),
    .Y(_19269_));
 OAI21x1_ASAP7_75t_R _27783_ (.A1(_19265_),
    .A2(_19269_),
    .B(net2198),
    .Y(_19270_));
 NAND2x2_ASAP7_75t_R _27784_ (.A(_19263_),
    .B(_19270_),
    .Y(_00122_));
 BUFx2_ASAP7_75t_R input3 (.A(net4075),
    .Y(net3));
 BUFx2_ASAP7_75t_R input2 (.A(net4197),
    .Y(net2));
 AO21x1_ASAP7_75t_R _27787_ (.A1(net1097),
    .A2(_17586_),
    .B(_17759_),
    .Y(_19273_));
 AO21x1_ASAP7_75t_R _27788_ (.A1(net2202),
    .A2(net2451),
    .B(_17759_),
    .Y(_19274_));
 NAND2x1_ASAP7_75t_R _27789_ (.A(_19273_),
    .B(_19274_),
    .Y(_19275_));
 AO21x1_ASAP7_75t_R _27790_ (.A1(net2202),
    .A2(net2899),
    .B(_17744_),
    .Y(_19276_));
 AO21x1_ASAP7_75t_R _27791_ (.A1(net2014),
    .A2(net3195),
    .B(_17744_),
    .Y(_19277_));
 OA21x2_ASAP7_75t_R _27792_ (.A1(_17744_),
    .A2(net1097),
    .B(_19277_),
    .Y(_19278_));
 NAND2x1_ASAP7_75t_R _27793_ (.A(_19276_),
    .B(_19278_),
    .Y(_19279_));
 NOR2x1_ASAP7_75t_R _27794_ (.A(_19275_),
    .B(_19279_),
    .Y(_19280_));
 AO21x1_ASAP7_75t_R _27795_ (.A1(_17834_),
    .A2(net3193),
    .B(net2758),
    .Y(_19281_));
 NOR2x1_ASAP7_75t_R _27796_ (.A(net1901),
    .B(_17788_),
    .Y(_19282_));
 AO21x1_ASAP7_75t_R _27797_ (.A1(_19282_),
    .A2(net941),
    .B(net2758),
    .Y(_19283_));
 NAND2x1_ASAP7_75t_R _27798_ (.A(_19281_),
    .B(_19283_),
    .Y(_19284_));
 NAND2x1_ASAP7_75t_R _27799_ (.A(net2642),
    .B(_17782_),
    .Y(_19285_));
 AO21x1_ASAP7_75t_R _27800_ (.A1(net2202),
    .A2(net941),
    .B(_17777_),
    .Y(_19286_));
 NAND2x1_ASAP7_75t_R _27801_ (.A(_19285_),
    .B(_19286_),
    .Y(_19287_));
 AO21x1_ASAP7_75t_R _27802_ (.A1(net1030),
    .A2(net1081),
    .B(_17777_),
    .Y(_19288_));
 AO21x1_ASAP7_75t_R _27803_ (.A1(_17639_),
    .A2(net1082),
    .B(_17777_),
    .Y(_19289_));
 NAND2x1_ASAP7_75t_R _27804_ (.A(_19288_),
    .B(_19289_),
    .Y(_19290_));
 NOR3x1_ASAP7_75t_R _27805_ (.A(_19284_),
    .B(_19287_),
    .C(_19290_),
    .Y(_19291_));
 NAND2x1_ASAP7_75t_R _27806_ (.A(_19280_),
    .B(_19291_),
    .Y(_19292_));
 AO21x1_ASAP7_75t_R _27807_ (.A1(_17845_),
    .A2(_17665_),
    .B(_17701_),
    .Y(_19293_));
 NAND2x2_ASAP7_75t_R _27808_ (.A(net1003),
    .B(_17608_),
    .Y(_19294_));
 AO21x1_ASAP7_75t_R _27809_ (.A1(net2236),
    .A2(_19294_),
    .B(_17701_),
    .Y(_19295_));
 NAND3x1_ASAP7_75t_R _27810_ (.A(_17910_),
    .B(_19293_),
    .C(_19295_),
    .Y(_19296_));
 OA21x2_ASAP7_75t_R _27811_ (.A1(_17678_),
    .A2(_17576_),
    .B(_17801_),
    .Y(_19297_));
 OA21x2_ASAP7_75t_R _27812_ (.A1(_17788_),
    .A2(_18788_),
    .B(_17801_),
    .Y(_19298_));
 OA21x2_ASAP7_75t_R _27813_ (.A1(_17661_),
    .A2(_17780_),
    .B(_17801_),
    .Y(_19299_));
 OR3x1_ASAP7_75t_R _27814_ (.A(_19297_),
    .B(_19298_),
    .C(_19299_),
    .Y(_19300_));
 NOR2x1_ASAP7_75t_R _27815_ (.A(_19296_),
    .B(_19300_),
    .Y(_19301_));
 AO21x1_ASAP7_75t_R _27816_ (.A1(_17746_),
    .A2(net1973),
    .B(_17725_),
    .Y(_19302_));
 NAND2x2_ASAP7_75t_R _27817_ (.A(_17733_),
    .B(_17553_),
    .Y(_19303_));
 AO21x1_ASAP7_75t_R _27818_ (.A1(net1097),
    .A2(_17834_),
    .B(_17725_),
    .Y(_19304_));
 NAND3x2_ASAP7_75t_R _27819_ (.B(_19303_),
    .C(_19304_),
    .Y(_19305_),
    .A(_19302_));
 AO21x1_ASAP7_75t_R _27820_ (.A1(net936),
    .A2(net2202),
    .B(_17712_),
    .Y(_19306_));
 OAI21x1_ASAP7_75t_R _27821_ (.A1(_17758_),
    .A2(net2881),
    .B(_19306_),
    .Y(_19307_));
 AO21x1_ASAP7_75t_R _27822_ (.A1(net3193),
    .A2(net2630),
    .B(net2881),
    .Y(_19308_));
 OAI21x1_ASAP7_75t_R _27823_ (.A1(_17639_),
    .A2(net2881),
    .B(_19308_),
    .Y(_19309_));
 NOR3x2_ASAP7_75t_R _27824_ (.B(_19307_),
    .C(_19309_),
    .Y(_19310_),
    .A(_19305_));
 NAND2x2_ASAP7_75t_R _27825_ (.A(_19301_),
    .B(_19310_),
    .Y(_19311_));
 NOR2x2_ASAP7_75t_R _27826_ (.A(_19311_),
    .B(_19292_),
    .Y(_19312_));
 OA21x2_ASAP7_75t_R _27827_ (.A1(_17661_),
    .A2(_17780_),
    .B(_17618_),
    .Y(_19313_));
 AO21x1_ASAP7_75t_R _27828_ (.A1(_17618_),
    .A2(_17539_),
    .B(_19313_),
    .Y(_19314_));
 AO21x1_ASAP7_75t_R _27829_ (.A1(net2902),
    .A2(_17538_),
    .B(_17589_),
    .Y(_19315_));
 AO21x1_ASAP7_75t_R _27830_ (.A1(_17746_),
    .A2(_17557_),
    .B(_17589_),
    .Y(_19316_));
 NAND2x1_ASAP7_75t_R _27831_ (.A(_19315_),
    .B(_19316_),
    .Y(_19317_));
 AOI211x1_ASAP7_75t_R _27832_ (.A1(_17618_),
    .A2(_17694_),
    .B(_19314_),
    .C(_19317_),
    .Y(_19318_));
 AOI211x1_ASAP7_75t_R _27833_ (.A1(net2862),
    .A2(net2891),
    .B(_17566_),
    .C(net2902),
    .Y(_19319_));
 OA21x2_ASAP7_75t_R _27834_ (.A1(_17576_),
    .A2(_17679_),
    .B(_17569_),
    .Y(_19320_));
 NOR2x1_ASAP7_75t_R _27835_ (.A(_19319_),
    .B(_19320_),
    .Y(_19321_));
 AO21x1_ASAP7_75t_R _27836_ (.A1(net936),
    .A2(_17562_),
    .B(_17566_),
    .Y(_19322_));
 NAND3x1_ASAP7_75t_R _27837_ (.A(_19321_),
    .B(_17574_),
    .C(_19322_),
    .Y(_19323_));
 AO21x1_ASAP7_75t_R _27838_ (.A1(net1030),
    .A2(net1081),
    .B(_17547_),
    .Y(_19324_));
 OA21x2_ASAP7_75t_R _27839_ (.A1(_17547_),
    .A2(net1097),
    .B(_19324_),
    .Y(_19325_));
 OA211x2_ASAP7_75t_R _27840_ (.A1(net2862),
    .A2(net2879),
    .B(_17548_),
    .C(_17561_),
    .Y(_19326_));
 INVx1_ASAP7_75t_R _27841_ (.A(_19326_),
    .Y(_19327_));
 NAND2x1_ASAP7_75t_R _27842_ (.A(_19325_),
    .B(_19327_),
    .Y(_19328_));
 NOR2x1_ASAP7_75t_R _27843_ (.A(_19323_),
    .B(_19328_),
    .Y(_19329_));
 NAND2x1_ASAP7_75t_R _27844_ (.A(_19318_),
    .B(_19329_),
    .Y(_19330_));
 OA21x2_ASAP7_75t_R _27845_ (.A1(_17788_),
    .A2(_17607_),
    .B(_17650_),
    .Y(_19331_));
 AOI21x1_ASAP7_75t_R _27846_ (.A1(_17632_),
    .A2(_17647_),
    .B(net2484),
    .Y(_19332_));
 OR3x1_ASAP7_75t_R _27847_ (.A(_19331_),
    .B(_17894_),
    .C(_19332_),
    .Y(_19333_));
 OA21x2_ASAP7_75t_R _27848_ (.A1(_18788_),
    .A2(_17774_),
    .B(_18789_),
    .Y(_19334_));
 OA21x2_ASAP7_75t_R _27849_ (.A1(net2906),
    .A2(_17673_),
    .B(_18789_),
    .Y(_19335_));
 NOR2x1_ASAP7_75t_R _27850_ (.A(_19294_),
    .B(_17629_),
    .Y(_19336_));
 OR3x1_ASAP7_75t_R _27851_ (.A(_19334_),
    .B(_19335_),
    .C(_19336_),
    .Y(_19337_));
 NOR2x1_ASAP7_75t_R _27852_ (.A(_19333_),
    .B(_19337_),
    .Y(_19338_));
 AO21x1_ASAP7_75t_R _27853_ (.A1(_17845_),
    .A2(_17695_),
    .B(net2889),
    .Y(_19339_));
 AO21x1_ASAP7_75t_R _27854_ (.A1(net997),
    .A2(net1380),
    .B(net2889),
    .Y(_19340_));
 AND2x2_ASAP7_75t_R _27855_ (.A(_19339_),
    .B(_19340_),
    .Y(_19341_));
 AO21x1_ASAP7_75t_R _27856_ (.A1(net2893),
    .A2(net1097),
    .B(net2889),
    .Y(_19342_));
 AO21x1_ASAP7_75t_R _27857_ (.A1(_17813_),
    .A2(_17586_),
    .B(net2889),
    .Y(_19343_));
 NAND3x2_ASAP7_75t_R _27858_ (.B(_19342_),
    .C(_19343_),
    .Y(_19344_),
    .A(_19341_));
 AO21x1_ASAP7_75t_R _27859_ (.A1(net2532),
    .A2(_17647_),
    .B(_17657_),
    .Y(_19345_));
 INVx1_ASAP7_75t_R _27860_ (.A(_17888_),
    .Y(_19346_));
 AND2x2_ASAP7_75t_R _27861_ (.A(_19345_),
    .B(_19346_),
    .Y(_19347_));
 AO21x1_ASAP7_75t_R _27862_ (.A1(net997),
    .A2(net2597),
    .B(_17657_),
    .Y(_19348_));
 AO21x1_ASAP7_75t_R _27863_ (.A1(_17756_),
    .A2(net1380),
    .B(_17657_),
    .Y(_19349_));
 NAND2x1_ASAP7_75t_R _27864_ (.A(_17694_),
    .B(_17662_),
    .Y(_19350_));
 AND3x1_ASAP7_75t_R _27865_ (.A(_19348_),
    .B(_19349_),
    .C(_19350_),
    .Y(_19351_));
 NAND2x1_ASAP7_75t_R _27866_ (.A(_19351_),
    .B(_19347_),
    .Y(_19352_));
 NOR2x2_ASAP7_75t_R _27867_ (.A(_19344_),
    .B(_19352_),
    .Y(_19353_));
 NAND2x2_ASAP7_75t_R _27868_ (.A(_19353_),
    .B(_19338_),
    .Y(_19354_));
 NOR2x2_ASAP7_75t_R _27869_ (.A(_19330_),
    .B(_19354_),
    .Y(_19355_));
 NAND2x2_ASAP7_75t_R _27870_ (.A(_19312_),
    .B(_19355_),
    .Y(_19356_));
 AO21x1_ASAP7_75t_R _27871_ (.A1(net3306),
    .A2(_18057_),
    .B(net3216),
    .Y(_19357_));
 AO21x1_ASAP7_75t_R _27872_ (.A1(_18883_),
    .A2(_18022_),
    .B(net3216),
    .Y(_19358_));
 NAND2x2_ASAP7_75t_R _27873_ (.A(_18090_),
    .B(_18916_),
    .Y(_19359_));
 NAND3x2_ASAP7_75t_R _27874_ (.B(_19358_),
    .C(_19359_),
    .Y(_19360_),
    .A(_19357_));
 NAND2x1_ASAP7_75t_R _27875_ (.A(net2718),
    .B(_17961_),
    .Y(_19361_));
 AO21x1_ASAP7_75t_R _27876_ (.A1(_19361_),
    .A2(net2058),
    .B(_18024_),
    .Y(_19362_));
 AO21x2_ASAP7_75t_R _27877_ (.A1(_17980_),
    .A2(_18057_),
    .B(_18024_),
    .Y(_19363_));
 NAND2x2_ASAP7_75t_R _27878_ (.A(net3343),
    .B(net2730),
    .Y(_19364_));
 NAND3x2_ASAP7_75t_R _27879_ (.B(_19363_),
    .C(_19364_),
    .Y(_19365_),
    .A(_19362_));
 NOR2x2_ASAP7_75t_R _27880_ (.A(_19360_),
    .B(_19365_),
    .Y(_19366_));
 AO21x1_ASAP7_75t_R _27881_ (.A1(net1121),
    .A2(_18057_),
    .B(_17997_),
    .Y(_19367_));
 OA21x2_ASAP7_75t_R _27882_ (.A1(net3213),
    .A2(_17997_),
    .B(_19367_),
    .Y(_19368_));
 OA211x2_ASAP7_75t_R _27883_ (.A1(net3201),
    .A2(net3124),
    .B(_18006_),
    .C(_17955_),
    .Y(_19369_));
 INVx1_ASAP7_75t_R _27884_ (.A(_19369_),
    .Y(_19370_));
 NAND2x2_ASAP7_75t_R _27885_ (.A(_19368_),
    .B(_19370_),
    .Y(_19371_));
 AO21x1_ASAP7_75t_R _27886_ (.A1(net939),
    .A2(_17987_),
    .B(net1955),
    .Y(_19372_));
 AND2x2_ASAP7_75t_R _27887_ (.A(_19372_),
    .B(_17986_),
    .Y(_19373_));
 AO21x1_ASAP7_75t_R _27888_ (.A1(_17938_),
    .A2(net1690),
    .B(net1955),
    .Y(_19374_));
 AO21x1_ASAP7_75t_R _27889_ (.A1(net3224),
    .A2(net3191),
    .B(net3205),
    .Y(_19375_));
 INVx2_ASAP7_75t_R _27890_ (.A(_17977_),
    .Y(_19376_));
 NAND2x1_ASAP7_75t_R _27891_ (.A(_18923_),
    .B(_19376_),
    .Y(_19377_));
 AND3x1_ASAP7_75t_R _27892_ (.A(_19374_),
    .B(_19375_),
    .C(_19377_),
    .Y(_19378_));
 NAND2x2_ASAP7_75t_R _27893_ (.A(_19373_),
    .B(_19378_),
    .Y(_19379_));
 NOR2x1_ASAP7_75t_R _27894_ (.A(_19371_),
    .B(_19379_),
    .Y(_19380_));
 NAND2x1_ASAP7_75t_R _27895_ (.A(_19366_),
    .B(_19380_),
    .Y(_19381_));
 AOI21x1_ASAP7_75t_R _27896_ (.A1(net1624),
    .A2(net1348),
    .B(_18039_),
    .Y(_19382_));
 AOI21x1_ASAP7_75t_R _27897_ (.A1(_18040_),
    .A2(_17952_),
    .B(_19382_),
    .Y(_19383_));
 AO21x1_ASAP7_75t_R _27898_ (.A1(_18010_),
    .A2(net2757),
    .B(_18039_),
    .Y(_19384_));
 NAND2x1_ASAP7_75t_R _27899_ (.A(_17923_),
    .B(_17942_),
    .Y(_19385_));
 AO21x2_ASAP7_75t_R _27900_ (.A1(_18073_),
    .A2(_19385_),
    .B(_18039_),
    .Y(_19386_));
 NAND3x2_ASAP7_75t_R _27901_ (.B(_19384_),
    .C(_19386_),
    .Y(_19387_),
    .A(_19383_));
 AO21x1_ASAP7_75t_R _27902_ (.A1(net939),
    .A2(net974),
    .B(net2303),
    .Y(_19388_));
 AO21x1_ASAP7_75t_R _27903_ (.A1(net1532),
    .A2(_17962_),
    .B(net2303),
    .Y(_19389_));
 AND2x2_ASAP7_75t_R _27904_ (.A(_19388_),
    .B(_19389_),
    .Y(_19390_));
 AO21x1_ASAP7_75t_R _27905_ (.A1(net3213),
    .A2(net1689),
    .B(_18054_),
    .Y(_19391_));
 AO21x1_ASAP7_75t_R _27906_ (.A1(net3306),
    .A2(_18958_),
    .B(_18054_),
    .Y(_19392_));
 NAND3x1_ASAP7_75t_R _27907_ (.A(_19390_),
    .B(_19391_),
    .C(_19392_),
    .Y(_19393_));
 NOR2x1_ASAP7_75t_R _27908_ (.A(_19387_),
    .B(_19393_),
    .Y(_19394_));
 AOI211x1_ASAP7_75t_R _27909_ (.A1(net3201),
    .A2(net1117),
    .B(_18074_),
    .C(net3285),
    .Y(_19395_));
 INVx1_ASAP7_75t_R _27910_ (.A(_19395_),
    .Y(_19396_));
 AO21x1_ASAP7_75t_R _27911_ (.A1(net3214),
    .A2(net1689),
    .B(net2181),
    .Y(_19397_));
 AO21x1_ASAP7_75t_R _27912_ (.A1(net939),
    .A2(net974),
    .B(net2181),
    .Y(_19398_));
 AND3x1_ASAP7_75t_R _27913_ (.A(_19396_),
    .B(_19397_),
    .C(_19398_),
    .Y(_19399_));
 AO21x1_ASAP7_75t_R _27914_ (.A1(_18028_),
    .A2(net2757),
    .B(net1912),
    .Y(_19400_));
 NAND2x1_ASAP7_75t_R _27915_ (.A(_17952_),
    .B(_18069_),
    .Y(_19401_));
 AND2x2_ASAP7_75t_R _27916_ (.A(_19400_),
    .B(_19401_),
    .Y(_19402_));
 NOR2x2_ASAP7_75t_R _27917_ (.A(_17947_),
    .B(net1910),
    .Y(_19403_));
 AOI22x1_ASAP7_75t_R _27918_ (.A1(_19403_),
    .A2(net3124),
    .B1(_17925_),
    .B2(_18069_),
    .Y(_19404_));
 AND2x2_ASAP7_75t_R _27919_ (.A(_19402_),
    .B(_19404_),
    .Y(_19405_));
 NAND2x1_ASAP7_75t_R _27920_ (.A(_19399_),
    .B(_19405_),
    .Y(_19406_));
 INVx1_ASAP7_75t_R _27921_ (.A(_19406_),
    .Y(_19407_));
 NAND2x1_ASAP7_75t_R _27922_ (.A(_19394_),
    .B(_19407_),
    .Y(_19408_));
 NOR2x1_ASAP7_75t_R _27923_ (.A(_19381_),
    .B(_19408_),
    .Y(_19409_));
 AO21x1_ASAP7_75t_R _27924_ (.A1(_18010_),
    .A2(net1795),
    .B(_18156_),
    .Y(_19410_));
 AO21x1_ASAP7_75t_R _27925_ (.A1(net1121),
    .A2(net1050),
    .B(_18156_),
    .Y(_19411_));
 NAND2x1_ASAP7_75t_R _27926_ (.A(net3192),
    .B(_18923_),
    .Y(_19412_));
 AND3x1_ASAP7_75t_R _27927_ (.A(_19410_),
    .B(_19411_),
    .C(_19412_),
    .Y(_19413_));
 AO21x1_ASAP7_75t_R _27928_ (.A1(_18057_),
    .A2(net1068),
    .B(net2446),
    .Y(_19414_));
 NAND2x1_ASAP7_75t_R _27929_ (.A(_18923_),
    .B(_18151_),
    .Y(_19415_));
 NAND2x1_ASAP7_75t_R _27930_ (.A(_18900_),
    .B(_18151_),
    .Y(_19416_));
 NAND2x1_ASAP7_75t_R _27931_ (.A(_18110_),
    .B(_18151_),
    .Y(_19417_));
 AND4x1_ASAP7_75t_R _27932_ (.A(_19414_),
    .B(_19415_),
    .C(_19416_),
    .D(_19417_),
    .Y(_19418_));
 NAND2x2_ASAP7_75t_R _27933_ (.A(_19413_),
    .B(_19418_),
    .Y(_19419_));
 AO21x1_ASAP7_75t_R _27934_ (.A1(_18883_),
    .A2(_18057_),
    .B(_18169_),
    .Y(_19420_));
 NAND2x1_ASAP7_75t_R _27935_ (.A(net3299),
    .B(_18900_),
    .Y(_19421_));
 AND3x2_ASAP7_75t_R _27936_ (.A(_18171_),
    .B(_19420_),
    .C(_19421_),
    .Y(_19422_));
 NAND2x2_ASAP7_75t_R _27937_ (.A(_17996_),
    .B(_18143_),
    .Y(_19423_));
 AO31x2_ASAP7_75t_R _27938_ (.A1(net1529),
    .A2(net1795),
    .A3(net974),
    .B(_19423_),
    .Y(_19424_));
 AO21x1_ASAP7_75t_R _27939_ (.A1(net1675),
    .A2(_18022_),
    .B(_19423_),
    .Y(_19425_));
 AO21x1_ASAP7_75t_R _27940_ (.A1(net1121),
    .A2(_18057_),
    .B(_19423_),
    .Y(_19426_));
 AND2x2_ASAP7_75t_R _27941_ (.A(_19425_),
    .B(_19426_),
    .Y(_19427_));
 NAND3x2_ASAP7_75t_R _27942_ (.B(_19424_),
    .C(_19427_),
    .Y(_19428_),
    .A(_19422_));
 NOR2x2_ASAP7_75t_R _27943_ (.A(_19419_),
    .B(_19428_),
    .Y(_19429_));
 INVx1_ASAP7_75t_R _27944_ (.A(_19429_),
    .Y(_19430_));
 AOI211x1_ASAP7_75t_R _27945_ (.A1(net3201),
    .A2(net1117),
    .B(net1371),
    .C(net2364),
    .Y(_19431_));
 INVx1_ASAP7_75t_R _27946_ (.A(_19431_),
    .Y(_19432_));
 AO21x1_ASAP7_75t_R _27947_ (.A1(net3306),
    .A2(_18057_),
    .B(net2364),
    .Y(_19433_));
 AO21x1_ASAP7_75t_R _27948_ (.A1(net939),
    .A2(net2757),
    .B(net2364),
    .Y(_19434_));
 AND3x1_ASAP7_75t_R _27949_ (.A(_19432_),
    .B(_19433_),
    .C(_19434_),
    .Y(_19435_));
 INVx1_ASAP7_75t_R _27950_ (.A(_17959_),
    .Y(_19436_));
 AO21x1_ASAP7_75t_R _27951_ (.A1(_18010_),
    .A2(_17963_),
    .B(net1746),
    .Y(_19437_));
 NAND2x1_ASAP7_75t_R _27952_ (.A(_19436_),
    .B(_19437_),
    .Y(_19438_));
 AO22x1_ASAP7_75t_R _27953_ (.A1(_18923_),
    .A2(_17932_),
    .B1(_17948_),
    .B2(net2720),
    .Y(_19439_));
 NOR2x1_ASAP7_75t_R _27954_ (.A(_19438_),
    .B(_19439_),
    .Y(_19440_));
 NAND2x1_ASAP7_75t_R _27955_ (.A(_19435_),
    .B(_19440_),
    .Y(_19441_));
 INVx1_ASAP7_75t_R _27956_ (.A(_19441_),
    .Y(_19442_));
 NAND2x1_ASAP7_75t_R _27957_ (.A(net2166),
    .B(_18000_),
    .Y(_19443_));
 OA211x2_ASAP7_75t_R _27958_ (.A1(net1057),
    .A2(net1117),
    .B(net2680),
    .C(_17934_),
    .Y(_19444_));
 INVx1_ASAP7_75t_R _27959_ (.A(_19444_),
    .Y(_19445_));
 NAND2x2_ASAP7_75t_R _27960_ (.A(_19443_),
    .B(_19445_),
    .Y(_19446_));
 AO21x1_ASAP7_75t_R _27961_ (.A1(net1795),
    .A2(net939),
    .B(_18126_),
    .Y(_19447_));
 NAND2x1_ASAP7_75t_R _27962_ (.A(net3308),
    .B(net1815),
    .Y(_19448_));
 AO21x1_ASAP7_75t_R _27963_ (.A1(net1676),
    .A2(_19448_),
    .B(_18126_),
    .Y(_19449_));
 NAND2x2_ASAP7_75t_R _27964_ (.A(_18105_),
    .B(_18123_),
    .Y(_19450_));
 NAND3x2_ASAP7_75t_R _27965_ (.B(_19449_),
    .C(_19450_),
    .Y(_19451_),
    .A(_19447_));
 AO21x1_ASAP7_75t_R _27966_ (.A1(_18147_),
    .A2(_18081_),
    .B(_18864_),
    .Y(_19452_));
 OAI21x1_ASAP7_75t_R _27967_ (.A1(_18864_),
    .A2(net2060),
    .B(_19452_),
    .Y(_19453_));
 NOR3x2_ASAP7_75t_R _27968_ (.B(net3342),
    .C(_19453_),
    .Y(_19454_),
    .A(_19446_));
 NAND2x1_ASAP7_75t_R _27969_ (.A(_19442_),
    .B(_19454_),
    .Y(_19455_));
 NOR2x2_ASAP7_75t_R _27970_ (.A(_19430_),
    .B(_19455_),
    .Y(_19456_));
 NAND2x2_ASAP7_75t_R _27971_ (.A(_19409_),
    .B(_19456_),
    .Y(_19457_));
 NAND2x1_ASAP7_75t_R _27972_ (.A(net3346),
    .B(_19457_),
    .Y(_19458_));
 NOR2x1_ASAP7_75t_R _27973_ (.A(net3346),
    .B(_19457_),
    .Y(_19459_));
 INVx1_ASAP7_75t_R _27974_ (.A(_19459_),
    .Y(_19460_));
 AO21x1_ASAP7_75t_R _27975_ (.A1(net2043),
    .A2(net2634),
    .B(_18456_),
    .Y(_19461_));
 AO21x1_ASAP7_75t_R _27976_ (.A1(net1606),
    .A2(_18335_),
    .B(_18456_),
    .Y(_19462_));
 AND2x2_ASAP7_75t_R _27977_ (.A(_19461_),
    .B(_19462_),
    .Y(_19463_));
 NOR2x1_ASAP7_75t_R _27978_ (.A(net2250),
    .B(_18464_),
    .Y(_19464_));
 NOR2x2_ASAP7_75t_R _27979_ (.A(_18258_),
    .B(_18366_),
    .Y(_19465_));
 OA21x2_ASAP7_75t_R _27980_ (.A1(_19202_),
    .A2(_19465_),
    .B(_18469_),
    .Y(_19466_));
 NOR2x1_ASAP7_75t_R _27981_ (.A(_19464_),
    .B(_19466_),
    .Y(_19467_));
 AO21x1_ASAP7_75t_R _27982_ (.A1(net2634),
    .A2(net2638),
    .B(net3312),
    .Y(_19468_));
 AND3x1_ASAP7_75t_R _27983_ (.A(_19463_),
    .B(_19467_),
    .C(_19468_),
    .Y(_19469_));
 INVx1_ASAP7_75t_R _27984_ (.A(_18493_),
    .Y(_19470_));
 AO21x1_ASAP7_75t_R _27985_ (.A1(_18351_),
    .A2(net2004),
    .B(net2595),
    .Y(_19471_));
 INVx3_ASAP7_75t_R _27986_ (.A(_18490_),
    .Y(_19472_));
 NAND2x1_ASAP7_75t_R _27987_ (.A(_18482_),
    .B(_19472_),
    .Y(_19473_));
 NAND3x1_ASAP7_75t_R _27988_ (.A(_19470_),
    .B(_19471_),
    .C(_19473_),
    .Y(_19474_));
 AO21x1_ASAP7_75t_R _27989_ (.A1(_18467_),
    .A2(net2971),
    .B(net3246),
    .Y(_19475_));
 AO21x1_ASAP7_75t_R _27990_ (.A1(_19475_),
    .A2(_18489_),
    .B(net3282),
    .Y(_19476_));
 AO21x1_ASAP7_75t_R _27991_ (.A1(net2699),
    .A2(net937),
    .B(net3282),
    .Y(_19477_));
 OA21x2_ASAP7_75t_R _27992_ (.A1(net2452),
    .A2(net3282),
    .B(_19477_),
    .Y(_19478_));
 NAND2x1_ASAP7_75t_R _27993_ (.A(_19476_),
    .B(_19478_),
    .Y(_19479_));
 NOR2x1_ASAP7_75t_R _27994_ (.A(_19474_),
    .B(_19479_),
    .Y(_19480_));
 NAND2x1_ASAP7_75t_R _27995_ (.A(_19469_),
    .B(_19480_),
    .Y(_19481_));
 NOR2x1_ASAP7_75t_R _27996_ (.A(net1087),
    .B(_18273_),
    .Y(_19482_));
 INVx1_ASAP7_75t_R _27997_ (.A(_19482_),
    .Y(_19483_));
 AO21x1_ASAP7_75t_R _27998_ (.A1(net1606),
    .A2(_18242_),
    .B(_18248_),
    .Y(_19484_));
 AO21x1_ASAP7_75t_R _27999_ (.A1(_18314_),
    .A2(net2452),
    .B(_18248_),
    .Y(_19485_));
 NAND3x1_ASAP7_75t_R _28000_ (.A(_19483_),
    .B(_19484_),
    .C(_19485_),
    .Y(_19486_));
 OA21x2_ASAP7_75t_R _28001_ (.A1(_18482_),
    .A2(_18445_),
    .B(_18416_),
    .Y(_19487_));
 OA21x2_ASAP7_75t_R _28002_ (.A1(_19160_),
    .A2(_18468_),
    .B(_18416_),
    .Y(_19488_));
 NOR2x1_ASAP7_75t_R _28003_ (.A(_18460_),
    .B(_18266_),
    .Y(_19489_));
 OR3x1_ASAP7_75t_R _28004_ (.A(_19487_),
    .B(_19488_),
    .C(_19489_),
    .Y(_19490_));
 NOR2x1_ASAP7_75t_R _28005_ (.A(_19486_),
    .B(_19490_),
    .Y(_19491_));
 AO21x1_ASAP7_75t_R _28006_ (.A1(net1606),
    .A2(_18351_),
    .B(net2989),
    .Y(_19492_));
 NAND2x2_ASAP7_75t_R _28007_ (.A(_18241_),
    .B(_18313_),
    .Y(_19493_));
 AO21x1_ASAP7_75t_R _28008_ (.A1(_19493_),
    .A2(net2498),
    .B(net2989),
    .Y(_19494_));
 NAND2x1_ASAP7_75t_R _28009_ (.A(_19202_),
    .B(_18446_),
    .Y(_19495_));
 NAND3x1_ASAP7_75t_R _28010_ (.A(_19492_),
    .B(_19494_),
    .C(_19495_),
    .Y(_19496_));
 OA21x2_ASAP7_75t_R _28011_ (.A1(_19202_),
    .A2(_19465_),
    .B(_18434_),
    .Y(_19497_));
 NOR2x1_ASAP7_75t_R _28012_ (.A(_18430_),
    .B(_19497_),
    .Y(_19498_));
 AO21x1_ASAP7_75t_R _28013_ (.A1(_18381_),
    .A2(net2452),
    .B(_18428_),
    .Y(_19499_));
 AO21x1_ASAP7_75t_R _28014_ (.A1(net2634),
    .A2(net1335),
    .B(_18428_),
    .Y(_19500_));
 NAND3x1_ASAP7_75t_R _28015_ (.A(_19498_),
    .B(_19499_),
    .C(_19500_),
    .Y(_19501_));
 NOR2x1_ASAP7_75t_R _28016_ (.A(_19496_),
    .B(_19501_),
    .Y(_19502_));
 NAND2x1_ASAP7_75t_R _28017_ (.A(_19491_),
    .B(_19502_),
    .Y(_19503_));
 NOR2x2_ASAP7_75t_R _28018_ (.A(_19481_),
    .B(_19503_),
    .Y(_19504_));
 AO21x1_ASAP7_75t_R _28019_ (.A1(net1254),
    .A2(net2004),
    .B(net2985),
    .Y(_19505_));
 OA21x2_ASAP7_75t_R _28020_ (.A1(net1606),
    .A2(net2985),
    .B(_19505_),
    .Y(_19506_));
 OA211x2_ASAP7_75t_R _28021_ (.A1(net2999),
    .A2(_18237_),
    .B(_18292_),
    .C(_18272_),
    .Y(_19507_));
 INVx1_ASAP7_75t_R _28022_ (.A(_19507_),
    .Y(_19508_));
 NAND2x1_ASAP7_75t_R _28023_ (.A(_19506_),
    .B(_19508_),
    .Y(_19509_));
 AO21x1_ASAP7_75t_R _28024_ (.A1(net1335),
    .A2(net1821),
    .B(net2970),
    .Y(_19510_));
 AND2x2_ASAP7_75t_R _28025_ (.A(_19510_),
    .B(_18310_),
    .Y(_19511_));
 BUFx2_ASAP7_75t_R input1 (.A(net4188),
    .Y(net1));
 AOI211x1_ASAP7_75t_R _28027_ (.A1(net2999),
    .A2(_18237_),
    .B(net2970),
    .C(net2010),
    .Y(_19513_));
 INVx1_ASAP7_75t_R _28028_ (.A(_19513_),
    .Y(_19514_));
 AO21x1_ASAP7_75t_R _28029_ (.A1(net2748),
    .A2(net1254),
    .B(net2970),
    .Y(_19515_));
 NAND3x1_ASAP7_75t_R _28030_ (.A(_19511_),
    .B(_19514_),
    .C(_19515_),
    .Y(_19516_));
 NOR2x1_ASAP7_75t_R _28031_ (.A(_19509_),
    .B(_19516_),
    .Y(_19517_));
 AO21x1_ASAP7_75t_R _28032_ (.A1(net2095),
    .A2(net1954),
    .B(_18318_),
    .Y(_19518_));
 INVx1_ASAP7_75t_R _28033_ (.A(_18460_),
    .Y(_19519_));
 INVx2_ASAP7_75t_R _28034_ (.A(_18318_),
    .Y(_19520_));
 NAND2x2_ASAP7_75t_R _28035_ (.A(_19519_),
    .B(_19520_),
    .Y(_19521_));
 NAND2x1_ASAP7_75t_R _28036_ (.A(net3281),
    .B(_19520_),
    .Y(_19522_));
 NAND3x1_ASAP7_75t_R _28037_ (.A(_19518_),
    .B(_19521_),
    .C(_19522_),
    .Y(_19523_));
 AO21x1_ASAP7_75t_R _28038_ (.A1(_18350_),
    .A2(_19493_),
    .B(_18330_),
    .Y(_19524_));
 AO21x1_ASAP7_75t_R _28039_ (.A1(net1335),
    .A2(_18460_),
    .B(_18330_),
    .Y(_19525_));
 NAND2x1_ASAP7_75t_R _28040_ (.A(_19160_),
    .B(_18345_),
    .Y(_19526_));
 NAND2x1_ASAP7_75t_R _28041_ (.A(_19205_),
    .B(_18345_),
    .Y(_19527_));
 AND3x1_ASAP7_75t_R _28042_ (.A(_19525_),
    .B(_19526_),
    .C(_19527_),
    .Y(_19528_));
 NAND2x1_ASAP7_75t_R _28043_ (.A(_19524_),
    .B(_19528_),
    .Y(_19529_));
 NOR2x1_ASAP7_75t_R _28044_ (.A(_19523_),
    .B(_19529_),
    .Y(_19530_));
 NAND2x1_ASAP7_75t_R _28045_ (.A(_19517_),
    .B(_19530_),
    .Y(_19531_));
 AO21x1_ASAP7_75t_R _28046_ (.A1(net2176),
    .A2(net1606),
    .B(net2981),
    .Y(_19532_));
 AO21x1_ASAP7_75t_R _28047_ (.A1(net1335),
    .A2(net937),
    .B(net2981),
    .Y(_19533_));
 OR2x2_ASAP7_75t_R _28048_ (.A(net2788),
    .B(net2981),
    .Y(_19534_));
 NAND3x1_ASAP7_75t_R _28049_ (.A(_19532_),
    .B(_19533_),
    .C(_19534_),
    .Y(_19535_));
 AO21x1_ASAP7_75t_R _28050_ (.A1(net2050),
    .A2(net2437),
    .B(_18395_),
    .Y(_19536_));
 AND2x2_ASAP7_75t_R _28051_ (.A(_19536_),
    .B(_18405_),
    .Y(_19537_));
 AO21x1_ASAP7_75t_R _28052_ (.A1(_18381_),
    .A2(net2638),
    .B(_18395_),
    .Y(_19538_));
 NAND2x2_ASAP7_75t_R _28053_ (.A(_18398_),
    .B(_18485_),
    .Y(_19539_));
 AND2x2_ASAP7_75t_R _28054_ (.A(_19538_),
    .B(_19539_),
    .Y(_19540_));
 NAND2x1_ASAP7_75t_R _28055_ (.A(_19537_),
    .B(_19540_),
    .Y(_19541_));
 NOR2x1_ASAP7_75t_R _28056_ (.A(_19535_),
    .B(_19541_),
    .Y(_19542_));
 NAND2x2_ASAP7_75t_R _28057_ (.A(_18488_),
    .B(net3001),
    .Y(_19543_));
 AOI21x1_ASAP7_75t_R _28058_ (.A1(net1483),
    .A2(_19543_),
    .B(_18364_),
    .Y(_19544_));
 INVx1_ASAP7_75t_R _28059_ (.A(_19544_),
    .Y(_19545_));
 AO21x1_ASAP7_75t_R _28060_ (.A1(net2045),
    .A2(net2638),
    .B(_18364_),
    .Y(_19546_));
 NAND2x1_ASAP7_75t_R _28061_ (.A(_18291_),
    .B(_18371_),
    .Y(_19547_));
 AO21x1_ASAP7_75t_R _28062_ (.A1(_18419_),
    .A2(net2004),
    .B(_18364_),
    .Y(_19548_));
 AND4x1_ASAP7_75t_R _28063_ (.A(_19545_),
    .B(_19546_),
    .C(_19547_),
    .D(_19548_),
    .Y(_19549_));
 AOI21x1_ASAP7_75t_R _28064_ (.A1(net2638),
    .A2(net2045),
    .B(_18354_),
    .Y(_19550_));
 AO21x1_ASAP7_75t_R _28065_ (.A1(net2668),
    .A2(_19237_),
    .B(_19550_),
    .Y(_19551_));
 AO21x1_ASAP7_75t_R _28066_ (.A1(net1335),
    .A2(net937),
    .B(net3178),
    .Y(_19552_));
 INVx1_ASAP7_75t_R _28067_ (.A(_19552_),
    .Y(_19553_));
 AO21x1_ASAP7_75t_R _28068_ (.A1(net2963),
    .A2(_18335_),
    .B(net3178),
    .Y(_19554_));
 AO21x1_ASAP7_75t_R _28069_ (.A1(net2176),
    .A2(net1606),
    .B(net3178),
    .Y(_19555_));
 NAND2x1_ASAP7_75t_R _28070_ (.A(_19554_),
    .B(_19555_),
    .Y(_19556_));
 NOR3x1_ASAP7_75t_R _28071_ (.A(_19551_),
    .B(_19553_),
    .C(_19556_),
    .Y(_19557_));
 NAND3x1_ASAP7_75t_R _28072_ (.A(_19542_),
    .B(_19549_),
    .C(_19557_),
    .Y(_19558_));
 NOR2x1_ASAP7_75t_R _28073_ (.A(_19531_),
    .B(_19558_),
    .Y(_19559_));
 NAND2x2_ASAP7_75t_R _28074_ (.A(_19504_),
    .B(_19559_),
    .Y(_19560_));
 AOI21x1_ASAP7_75t_R _28075_ (.A1(_19458_),
    .A2(_19460_),
    .B(_19560_),
    .Y(_19561_));
 INVx1_ASAP7_75t_R _28076_ (.A(_19387_),
    .Y(_19562_));
 AND4x1_ASAP7_75t_R _28077_ (.A(_19388_),
    .B(_19391_),
    .C(_19389_),
    .D(_19392_),
    .Y(_19563_));
 NAND2x1_ASAP7_75t_R _28078_ (.A(_19562_),
    .B(_19563_),
    .Y(_19564_));
 NOR2x1_ASAP7_75t_R _28079_ (.A(_19406_),
    .B(_19564_),
    .Y(_19565_));
 INVx1_ASAP7_75t_R _28080_ (.A(_19366_),
    .Y(_19566_));
 NOR3x2_ASAP7_75t_R _28081_ (.B(_19379_),
    .C(_19371_),
    .Y(_19567_),
    .A(_19566_));
 NAND2x2_ASAP7_75t_R _28082_ (.A(_19565_),
    .B(_19567_),
    .Y(_19568_));
 INVx1_ASAP7_75t_R _28083_ (.A(_19451_),
    .Y(_19569_));
 AOI211x1_ASAP7_75t_R _28084_ (.A1(_18000_),
    .A2(net2166),
    .B(_19444_),
    .C(_19453_),
    .Y(_19570_));
 NAND2x1_ASAP7_75t_R _28085_ (.A(_19569_),
    .B(_19570_),
    .Y(_19571_));
 NOR2x1_ASAP7_75t_R _28086_ (.A(_19441_),
    .B(_19571_),
    .Y(_19572_));
 NAND2x1_ASAP7_75t_R _28087_ (.A(_19429_),
    .B(_19572_),
    .Y(_19573_));
 NOR2x2_ASAP7_75t_R _28088_ (.A(_19568_),
    .B(_19573_),
    .Y(_19574_));
 NAND2x1_ASAP7_75t_R _28089_ (.A(net3346),
    .B(_19574_),
    .Y(_19575_));
 NOR2x2_ASAP7_75t_R _28090_ (.A(net3346),
    .B(_19574_),
    .Y(_19576_));
 INVx1_ASAP7_75t_R _28091_ (.A(_19576_),
    .Y(_19577_));
 INVx1_ASAP7_75t_R _28092_ (.A(_19560_),
    .Y(_19578_));
 AOI21x1_ASAP7_75t_R _28093_ (.A1(_19575_),
    .A2(_19577_),
    .B(_19578_),
    .Y(_19579_));
 INVx1_ASAP7_75t_R _28094_ (.A(_18714_),
    .Y(_19580_));
 OA21x2_ASAP7_75t_R _28095_ (.A1(_18694_),
    .A2(_18675_),
    .B(_19580_),
    .Y(_19581_));
 NAND2x2_ASAP7_75t_R _28096_ (.A(net1735),
    .B(_18558_),
    .Y(_19582_));
 TAPCELL_ASAP7_75t_R TAP_829 ();
 TAPCELL_ASAP7_75t_R TAP_828 ();
 AOI21x1_ASAP7_75t_R _28099_ (.A1(_19582_),
    .A2(net1404),
    .B(net2394),
    .Y(_19585_));
 AOI21x1_ASAP7_75t_R _28100_ (.A1(net1307),
    .A2(net1388),
    .B(net2394),
    .Y(_19586_));
 NOR3x1_ASAP7_75t_R _28101_ (.A(_19581_),
    .B(_19585_),
    .C(_19586_),
    .Y(_19587_));
 AOI211x1_ASAP7_75t_R _28102_ (.A1(net1469),
    .A2(net1733),
    .B(_18712_),
    .C(net1727),
    .Y(_19588_));
 NOR2x1_ASAP7_75t_R _28103_ (.A(net2633),
    .B(_18712_),
    .Y(_19589_));
 TAPCELL_ASAP7_75t_R TAP_827 ();
 AOI21x1_ASAP7_75t_R _28105_ (.A1(_18992_),
    .A2(net2029),
    .B(net3325),
    .Y(_19591_));
 NOR3x1_ASAP7_75t_R _28106_ (.A(_19588_),
    .B(_19589_),
    .C(_19591_),
    .Y(_19592_));
 NAND2x1_ASAP7_75t_R _28107_ (.A(_19587_),
    .B(_19592_),
    .Y(_19593_));
 AO21x1_ASAP7_75t_R _28108_ (.A1(net2089),
    .A2(net2142),
    .B(net2317),
    .Y(_19594_));
 NAND2x1_ASAP7_75t_R _28109_ (.A(_18672_),
    .B(_18725_),
    .Y(_19595_));
 AND2x2_ASAP7_75t_R _28110_ (.A(_19594_),
    .B(_19595_),
    .Y(_19596_));
 AOI21x1_ASAP7_75t_R _28111_ (.A1(_18536_),
    .A2(net2029),
    .B(_18729_),
    .Y(_19597_));
 INVx1_ASAP7_75t_R _28112_ (.A(_18729_),
    .Y(_19598_));
 OA21x2_ASAP7_75t_R _28113_ (.A1(_19007_),
    .A2(_18690_),
    .B(_19598_),
    .Y(_19599_));
 NOR2x1_ASAP7_75t_R _28114_ (.A(_19597_),
    .B(_19599_),
    .Y(_19600_));
 AO21x1_ASAP7_75t_R _28115_ (.A1(net3376),
    .A2(_18617_),
    .B(net2317),
    .Y(_19601_));
 NAND3x1_ASAP7_75t_R _28116_ (.A(_19596_),
    .B(_19600_),
    .C(_19601_),
    .Y(_19602_));
 NOR2x1_ASAP7_75t_R _28117_ (.A(_19593_),
    .B(_19602_),
    .Y(_19603_));
 NAND2x2_ASAP7_75t_R _28118_ (.A(_18608_),
    .B(_18671_),
    .Y(_19604_));
 AO21x1_ASAP7_75t_R _28119_ (.A1(_18528_),
    .A2(_18548_),
    .B(_18666_),
    .Y(_19605_));
 NAND2x1_ASAP7_75t_R _28120_ (.A(_19604_),
    .B(_19605_),
    .Y(_19606_));
 OR2x2_ASAP7_75t_R _28121_ (.A(_18666_),
    .B(_18653_),
    .Y(_19607_));
 AO21x1_ASAP7_75t_R _28122_ (.A1(_18627_),
    .A2(net3381),
    .B(_18666_),
    .Y(_19608_));
 NAND2x1_ASAP7_75t_R _28123_ (.A(_19607_),
    .B(_19608_),
    .Y(_19609_));
 NOR2x1_ASAP7_75t_R _28124_ (.A(_19606_),
    .B(_19609_),
    .Y(_19610_));
 NAND2x1_ASAP7_75t_R _28125_ (.A(_18675_),
    .B(_19031_),
    .Y(_19611_));
 AO21x1_ASAP7_75t_R _28126_ (.A1(_18528_),
    .A2(_18601_),
    .B(_18655_),
    .Y(_19612_));
 NAND2x1_ASAP7_75t_R _28127_ (.A(_19611_),
    .B(_19612_),
    .Y(_19613_));
 NOR2x2_ASAP7_75t_R _28128_ (.A(_18556_),
    .B(_18674_),
    .Y(_19614_));
 OA31x2_ASAP7_75t_R _28129_ (.A1(_18583_),
    .A2(_19614_),
    .A3(net2979),
    .B1(_19031_),
    .Y(_19615_));
 NOR2x1_ASAP7_75t_R _28130_ (.A(_19613_),
    .B(_19615_),
    .Y(_19616_));
 NAND2x1_ASAP7_75t_R _28131_ (.A(_19610_),
    .B(_19616_),
    .Y(_19617_));
 AO21x1_ASAP7_75t_R _28132_ (.A1(net1404),
    .A2(_18702_),
    .B(net2304),
    .Y(_19618_));
 AO21x1_ASAP7_75t_R _28133_ (.A1(net1388),
    .A2(_18548_),
    .B(net2304),
    .Y(_19619_));
 NAND2x1_ASAP7_75t_R _28134_ (.A(_18675_),
    .B(_18696_),
    .Y(_19620_));
 AND3x1_ASAP7_75t_R _28135_ (.A(_19618_),
    .B(_19619_),
    .C(_19620_),
    .Y(_19621_));
 NOR2x1_ASAP7_75t_R _28136_ (.A(_18531_),
    .B(_18680_),
    .Y(_19622_));
 OA21x2_ASAP7_75t_R _28137_ (.A1(_18614_),
    .A2(_18608_),
    .B(_18683_),
    .Y(_19623_));
 NOR2x1_ASAP7_75t_R _28138_ (.A(_18682_),
    .B(net1404),
    .Y(_19624_));
 AOI211x1_ASAP7_75t_R _28139_ (.A1(_18683_),
    .A2(_19622_),
    .B(_19623_),
    .C(_19624_),
    .Y(_19625_));
 NAND2x1_ASAP7_75t_R _28140_ (.A(_19621_),
    .B(_19625_),
    .Y(_19626_));
 NOR2x1_ASAP7_75t_R _28141_ (.A(_19617_),
    .B(_19626_),
    .Y(_19627_));
 NAND2x1_ASAP7_75t_R _28142_ (.A(_19603_),
    .B(_19627_),
    .Y(_19628_));
 OA21x2_ASAP7_75t_R _28143_ (.A1(_18608_),
    .A2(_18614_),
    .B(_18635_),
    .Y(_19629_));
 OA21x2_ASAP7_75t_R _28144_ (.A1(_19083_),
    .A2(net2979),
    .B(_18635_),
    .Y(_19630_));
 AOI211x1_ASAP7_75t_R _28145_ (.A1(_18635_),
    .A2(_19622_),
    .B(_19629_),
    .C(_19630_),
    .Y(_19631_));
 NAND2x1_ASAP7_75t_R _28146_ (.A(net2555),
    .B(_19058_),
    .Y(_19632_));
 AO21x1_ASAP7_75t_R _28147_ (.A1(net1307),
    .A2(net2386),
    .B(_18625_),
    .Y(_19633_));
 NAND2x1_ASAP7_75t_R _28148_ (.A(_19632_),
    .B(_19633_),
    .Y(_19634_));
 NAND2x2_ASAP7_75t_R _28149_ (.A(_19058_),
    .B(_19614_),
    .Y(_19635_));
 NOR2x1_ASAP7_75t_R _28150_ (.A(_18517_),
    .B(_18581_),
    .Y(_19636_));
 NAND2x1_ASAP7_75t_R _28151_ (.A(_19058_),
    .B(_19636_),
    .Y(_19637_));
 NAND3x1_ASAP7_75t_R _28152_ (.A(_19059_),
    .B(_19635_),
    .C(_19637_),
    .Y(_19638_));
 NOR2x1_ASAP7_75t_R _28153_ (.A(_19634_),
    .B(_19638_),
    .Y(_19639_));
 NAND2x1_ASAP7_75t_R _28154_ (.A(_19631_),
    .B(_19639_),
    .Y(_19640_));
 OA21x2_ASAP7_75t_R _28155_ (.A1(_19060_),
    .A2(_18585_),
    .B(_18612_),
    .Y(_19641_));
 OA21x2_ASAP7_75t_R _28156_ (.A1(_18694_),
    .A2(_18608_),
    .B(_18612_),
    .Y(_19642_));
 AOI211x1_ASAP7_75t_R _28157_ (.A1(net1468),
    .A2(net1735),
    .B(_18611_),
    .C(_18536_),
    .Y(_19643_));
 NOR3x1_ASAP7_75t_R _28158_ (.A(_19641_),
    .B(_19642_),
    .C(_19643_),
    .Y(_19644_));
 OA21x2_ASAP7_75t_R _28159_ (.A1(_18590_),
    .A2(_18537_),
    .B(_19046_),
    .Y(_19645_));
 AO21x1_ASAP7_75t_R _28160_ (.A1(net1404),
    .A2(_18516_),
    .B(_18604_),
    .Y(_19646_));
 NOR2x2_ASAP7_75t_R _28161_ (.A(net1730),
    .B(net2578),
    .Y(_19647_));
 NAND2x1_ASAP7_75t_R _28162_ (.A(net1069),
    .B(_19647_),
    .Y(_19648_));
 NAND2x1_ASAP7_75t_R _28163_ (.A(_19646_),
    .B(_19648_),
    .Y(_19649_));
 NOR2x1_ASAP7_75t_R _28164_ (.A(_19645_),
    .B(_19649_),
    .Y(_19650_));
 NAND2x1_ASAP7_75t_R _28165_ (.A(_19644_),
    .B(_19650_),
    .Y(_19651_));
 NOR2x1_ASAP7_75t_R _28166_ (.A(_19640_),
    .B(_19651_),
    .Y(_19652_));
 AO21x1_ASAP7_75t_R _28167_ (.A1(_18657_),
    .A2(_18992_),
    .B(_18588_),
    .Y(_19653_));
 AO21x1_ASAP7_75t_R _28168_ (.A1(net1388),
    .A2(_18547_),
    .B(_18588_),
    .Y(_19654_));
 AND2x2_ASAP7_75t_R _28169_ (.A(_19653_),
    .B(_19654_),
    .Y(_19655_));
 INVx1_ASAP7_75t_R _28170_ (.A(_19636_),
    .Y(_19656_));
 NOR2x1_ASAP7_75t_R _28171_ (.A(_18569_),
    .B(_19656_),
    .Y(_19657_));
 OA21x2_ASAP7_75t_R _28172_ (.A1(net2979),
    .A2(_19012_),
    .B(_18570_),
    .Y(_19658_));
 NOR2x1_ASAP7_75t_R _28173_ (.A(_19657_),
    .B(_19658_),
    .Y(_19659_));
 OA21x2_ASAP7_75t_R _28174_ (.A1(_18584_),
    .A2(_18588_),
    .B(_19090_),
    .Y(_19660_));
 NAND3x1_ASAP7_75t_R _28175_ (.A(_19655_),
    .B(_19659_),
    .C(_19660_),
    .Y(_19661_));
 AO21x1_ASAP7_75t_R _28176_ (.A1(net1404),
    .A2(net2052),
    .B(net2479),
    .Y(_19662_));
 AO21x1_ASAP7_75t_R _28177_ (.A1(_18623_),
    .A2(net1388),
    .B(_18545_),
    .Y(_19663_));
 INVx3_ASAP7_75t_R _28178_ (.A(_18545_),
    .Y(_19664_));
 NAND2x1_ASAP7_75t_R _28179_ (.A(_18552_),
    .B(_19664_),
    .Y(_19665_));
 AND3x1_ASAP7_75t_R _28180_ (.A(_19662_),
    .B(_19663_),
    .C(_19665_),
    .Y(_19666_));
 NAND2x1_ASAP7_75t_R _28181_ (.A(_19113_),
    .B(_19111_),
    .Y(_19667_));
 NAND2x1_ASAP7_75t_R _28182_ (.A(_18524_),
    .B(_18636_),
    .Y(_19668_));
 NAND3x1_ASAP7_75t_R _28183_ (.A(net2776),
    .B(_19668_),
    .C(_19086_),
    .Y(_19669_));
 NOR2x1_ASAP7_75t_R _28184_ (.A(_19667_),
    .B(_19669_),
    .Y(_19670_));
 NAND2x1_ASAP7_75t_R _28185_ (.A(_19666_),
    .B(_19670_),
    .Y(_19671_));
 NOR2x1_ASAP7_75t_R _28186_ (.A(_19661_),
    .B(_19671_),
    .Y(_19672_));
 NAND2x1_ASAP7_75t_R _28187_ (.A(_19652_),
    .B(_19672_),
    .Y(_19673_));
 NOR2x2_ASAP7_75t_R _28188_ (.A(_19628_),
    .B(_19673_),
    .Y(_19674_));
 NAND2x2_ASAP7_75t_R _28189_ (.A(_19120_),
    .B(_19674_),
    .Y(_19675_));
 XOR2x2_ASAP7_75t_R _28190_ (.A(_18852_),
    .B(_19675_),
    .Y(_19676_));
 OA21x2_ASAP7_75t_R _28191_ (.A1(_19561_),
    .A2(_19579_),
    .B(_19676_),
    .Y(_19677_));
 NAND2x1_ASAP7_75t_R _28192_ (.A(_19675_),
    .B(_18852_),
    .Y(_19678_));
 INVx1_ASAP7_75t_R _28193_ (.A(_19675_),
    .Y(_19679_));
 OAI21x1_ASAP7_75t_R _28194_ (.A1(net2143),
    .A2(_18851_),
    .B(_19679_),
    .Y(_19680_));
 AOI211x1_ASAP7_75t_R _28195_ (.A1(_19678_),
    .A2(_19680_),
    .B(_19579_),
    .C(_19561_),
    .Y(_19681_));
 NOR2x2_ASAP7_75t_R _28196_ (.A(_19681_),
    .B(_19677_),
    .Y(_19682_));
 TAPCELL_ASAP7_75t_R TAP_826 ();
 NOR2x1_ASAP7_75t_R _28198_ (.A(net397),
    .B(_00913_),
    .Y(_19684_));
 AOI21x1_ASAP7_75t_R _28199_ (.A1(net397),
    .A2(_19682_),
    .B(_19684_),
    .Y(_19685_));
 XOR2x1_ASAP7_75t_R _28200_ (.A(_19685_),
    .Y(_00123_),
    .B(net3527));
 NOR2x1_ASAP7_75t_R _28201_ (.A(net397),
    .B(_00912_),
    .Y(_19686_));
 INVx1_ASAP7_75t_R _28202_ (.A(_19686_),
    .Y(_19687_));
 XOR2x2_ASAP7_75t_R _28203_ (.A(net3346),
    .B(_18229_),
    .Y(_19688_));
 AOI211x1_ASAP7_75t_R _28204_ (.A1(net3090),
    .A2(_18554_),
    .B(net2632),
    .C(net1565),
    .Y(_19689_));
 AOI21x1_ASAP7_75t_R _28205_ (.A1(net2631),
    .A2(_19036_),
    .B(net2632),
    .Y(_19690_));
 AOI211x1_ASAP7_75t_R _28206_ (.A1(_18570_),
    .A2(_18672_),
    .B(_19689_),
    .C(_19690_),
    .Y(_19691_));
 AO21x1_ASAP7_75t_R _28207_ (.A1(_18621_),
    .A2(_19073_),
    .B(_18588_),
    .Y(_19692_));
 NAND2x1_ASAP7_75t_R _28208_ (.A(_18552_),
    .B(_18592_),
    .Y(_19693_));
 AO21x1_ASAP7_75t_R _28209_ (.A1(net2067),
    .A2(_18685_),
    .B(_18588_),
    .Y(_19694_));
 AND3x1_ASAP7_75t_R _28210_ (.A(_19692_),
    .B(_19693_),
    .C(_19694_),
    .Y(_19695_));
 NAND2x1_ASAP7_75t_R _28211_ (.A(_19695_),
    .B(_19691_),
    .Y(_19696_));
 AO21x1_ASAP7_75t_R _28212_ (.A1(_18627_),
    .A2(net3377),
    .B(_18525_),
    .Y(_19697_));
 AO21x1_ASAP7_75t_R _28213_ (.A1(_18643_),
    .A2(_18680_),
    .B(_18525_),
    .Y(_19698_));
 AND3x1_ASAP7_75t_R _28214_ (.A(_19697_),
    .B(_19698_),
    .C(_19084_),
    .Y(_19699_));
 AOI211x1_ASAP7_75t_R _28215_ (.A1(net3090),
    .A2(net1736),
    .B(_18545_),
    .C(net1565),
    .Y(_19700_));
 NOR2x1_ASAP7_75t_R _28216_ (.A(_18721_),
    .B(_18545_),
    .Y(_19701_));
 AO21x1_ASAP7_75t_R _28217_ (.A1(_18636_),
    .A2(_19664_),
    .B(_19701_),
    .Y(_19702_));
 AOI211x1_ASAP7_75t_R _28218_ (.A1(_19664_),
    .A2(_19093_),
    .B(_19700_),
    .C(_19702_),
    .Y(_19703_));
 NAND2x1_ASAP7_75t_R _28219_ (.A(_19699_),
    .B(_19703_),
    .Y(_19704_));
 NOR2x1_ASAP7_75t_R _28220_ (.A(_19696_),
    .B(_19704_),
    .Y(_19705_));
 AO21x1_ASAP7_75t_R _28221_ (.A1(_18685_),
    .A2(net1966),
    .B(net2580),
    .Y(_19706_));
 OA21x2_ASAP7_75t_R _28222_ (.A1(_18627_),
    .A2(net2615),
    .B(_19706_),
    .Y(_19707_));
 AO21x1_ASAP7_75t_R _28223_ (.A1(_18584_),
    .A2(net3381),
    .B(net2414),
    .Y(_19708_));
 AO21x1_ASAP7_75t_R _28224_ (.A1(net2028),
    .A2(net2829),
    .B(net2414),
    .Y(_19709_));
 AND2x2_ASAP7_75t_R _28225_ (.A(_19708_),
    .B(_19709_),
    .Y(_19710_));
 AO21x1_ASAP7_75t_R _28226_ (.A1(_19073_),
    .A2(_18992_),
    .B(net2580),
    .Y(_19711_));
 AO21x1_ASAP7_75t_R _28227_ (.A1(net2760),
    .A2(_18594_),
    .B(net2580),
    .Y(_19712_));
 AND2x2_ASAP7_75t_R _28228_ (.A(_19711_),
    .B(_19712_),
    .Y(_19713_));
 NAND3x2_ASAP7_75t_R _28229_ (.B(_19710_),
    .C(_19713_),
    .Y(_19714_),
    .A(_19707_));
 AO21x1_ASAP7_75t_R _28230_ (.A1(_18685_),
    .A2(net3377),
    .B(_18625_),
    .Y(_19715_));
 AO21x1_ASAP7_75t_R _28231_ (.A1(net2433),
    .A2(_18548_),
    .B(_18625_),
    .Y(_19716_));
 NAND2x1_ASAP7_75t_R _28232_ (.A(_19058_),
    .B(_18608_),
    .Y(_19717_));
 AND3x1_ASAP7_75t_R _28233_ (.A(_19715_),
    .B(_19716_),
    .C(_19717_),
    .Y(_19718_));
 TAPCELL_ASAP7_75t_R TAP_825 ();
 AO21x1_ASAP7_75t_R _28235_ (.A1(_18685_),
    .A2(net3381),
    .B(_18641_),
    .Y(_19720_));
 AO21x1_ASAP7_75t_R _28236_ (.A1(net2760),
    .A2(_18548_),
    .B(_18641_),
    .Y(_19721_));
 OA211x2_ASAP7_75t_R _28237_ (.A1(net2142),
    .A2(_18641_),
    .B(_19720_),
    .C(_19721_),
    .Y(_19722_));
 NAND2x2_ASAP7_75t_R _28238_ (.A(_19718_),
    .B(_19722_),
    .Y(_19723_));
 NOR2x2_ASAP7_75t_R _28239_ (.A(_19714_),
    .B(_19723_),
    .Y(_19724_));
 NAND2x2_ASAP7_75t_R _28240_ (.A(_19705_),
    .B(_19724_),
    .Y(_19725_));
 OA21x2_ASAP7_75t_R _28241_ (.A1(_18620_),
    .A2(_18590_),
    .B(_18696_),
    .Y(_19726_));
 OA21x2_ASAP7_75t_R _28242_ (.A1(_19614_),
    .A2(_18650_),
    .B(_18696_),
    .Y(_19727_));
 NOR3x1_ASAP7_75t_R _28243_ (.A(_19726_),
    .B(_19727_),
    .C(_18703_),
    .Y(_19728_));
 AO21x1_ASAP7_75t_R _28244_ (.A1(_18637_),
    .A2(_18535_),
    .B(net1568),
    .Y(_19729_));
 AO21x1_ASAP7_75t_R _28245_ (.A1(_19729_),
    .A2(_18680_),
    .B(net2545),
    .Y(_19730_));
 OA21x2_ASAP7_75t_R _28246_ (.A1(net2545),
    .A2(_18687_),
    .B(_19730_),
    .Y(_19731_));
 NAND2x1_ASAP7_75t_R _28247_ (.A(_19728_),
    .B(_19731_),
    .Y(_19732_));
 AO21x1_ASAP7_75t_R _28248_ (.A1(_18528_),
    .A2(_18601_),
    .B(_18666_),
    .Y(_19733_));
 NAND2x1_ASAP7_75t_R _28249_ (.A(_18694_),
    .B(_18671_),
    .Y(_19734_));
 AND3x1_ASAP7_75t_R _28250_ (.A(_19733_),
    .B(_19604_),
    .C(_19734_),
    .Y(_19735_));
 AO21x1_ASAP7_75t_R _28251_ (.A1(net2012),
    .A2(_18518_),
    .B(_18666_),
    .Y(_19736_));
 AO21x1_ASAP7_75t_R _28252_ (.A1(_18559_),
    .A2(_18721_),
    .B(_18666_),
    .Y(_19737_));
 NAND2x1_ASAP7_75t_R _28253_ (.A(_19057_),
    .B(_18671_),
    .Y(_19738_));
 AND3x1_ASAP7_75t_R _28254_ (.A(_19736_),
    .B(_19737_),
    .C(_19738_),
    .Y(_19739_));
 NAND2x1_ASAP7_75t_R _28255_ (.A(_19739_),
    .B(_19735_),
    .Y(_19740_));
 AO21x1_ASAP7_75t_R _28256_ (.A1(_18536_),
    .A2(net1564),
    .B(_18637_),
    .Y(_19741_));
 AO21x1_ASAP7_75t_R _28257_ (.A1(_19741_),
    .A2(_18623_),
    .B(_18655_),
    .Y(_19742_));
 AO21x1_ASAP7_75t_R _28258_ (.A1(net3376),
    .A2(net3381),
    .B(_18655_),
    .Y(_19743_));
 AO21x1_ASAP7_75t_R _28259_ (.A1(net1825),
    .A2(_18653_),
    .B(_18655_),
    .Y(_19744_));
 NAND3x1_ASAP7_75t_R _28260_ (.A(_19742_),
    .B(_19743_),
    .C(_19744_),
    .Y(_19745_));
 NOR3x1_ASAP7_75t_R _28261_ (.A(_19732_),
    .B(_19740_),
    .C(_19745_),
    .Y(_19746_));
 AO21x1_ASAP7_75t_R _28262_ (.A1(net1307),
    .A2(net2386),
    .B(_18712_),
    .Y(_19747_));
 NAND2x1_ASAP7_75t_R _28263_ (.A(_18608_),
    .B(_18718_),
    .Y(_19748_));
 OA211x2_ASAP7_75t_R _28264_ (.A1(_18712_),
    .A2(_18653_),
    .B(_19747_),
    .C(_19748_),
    .Y(_19749_));
 AO21x1_ASAP7_75t_R _28265_ (.A1(net2067),
    .A2(_18702_),
    .B(_18714_),
    .Y(_19750_));
 AO21x1_ASAP7_75t_R _28266_ (.A1(_18643_),
    .A2(net2029),
    .B(_18714_),
    .Y(_19751_));
 AO21x1_ASAP7_75t_R _28267_ (.A1(_18528_),
    .A2(net2433),
    .B(_18714_),
    .Y(_19752_));
 OR2x2_ASAP7_75t_R _28268_ (.A(_18714_),
    .B(_18975_),
    .Y(_19753_));
 AND4x1_ASAP7_75t_R _28269_ (.A(_19750_),
    .B(_19751_),
    .C(_19752_),
    .D(_19753_),
    .Y(_19754_));
 AO21x1_ASAP7_75t_R _28270_ (.A1(net2029),
    .A2(_18992_),
    .B(_18729_),
    .Y(_19755_));
 OAI21x1_ASAP7_75t_R _28271_ (.A1(net2694),
    .A2(_18547_),
    .B(_19755_),
    .Y(_19756_));
 AND3x1_ASAP7_75t_R _28272_ (.A(_18725_),
    .B(_18559_),
    .C(_18601_),
    .Y(_19757_));
 AO21x2_ASAP7_75t_R _28273_ (.A1(_18559_),
    .A2(_18721_),
    .B(net2694),
    .Y(_19758_));
 INVx1_ASAP7_75t_R _28274_ (.A(_19758_),
    .Y(_19759_));
 NOR3x1_ASAP7_75t_R _28275_ (.A(_19756_),
    .B(_19757_),
    .C(_19759_),
    .Y(_19760_));
 AND3x1_ASAP7_75t_R _28276_ (.A(_19749_),
    .B(_19754_),
    .C(_19760_),
    .Y(_19761_));
 NAND2x1_ASAP7_75t_R _28277_ (.A(_19761_),
    .B(_19746_),
    .Y(_19762_));
 NOR2x2_ASAP7_75t_R _28278_ (.A(_19725_),
    .B(_19762_),
    .Y(_19763_));
 XOR2x2_ASAP7_75t_R _28279_ (.A(_19763_),
    .B(_19143_),
    .Y(_19764_));
 NOR2x1_ASAP7_75t_R _28280_ (.A(_19688_),
    .B(_19764_),
    .Y(_19765_));
 AND2x2_ASAP7_75t_R _28281_ (.A(_19764_),
    .B(_19688_),
    .Y(_19766_));
 NAND2x1_ASAP7_75t_R _28282_ (.A(_18107_),
    .B(_18901_),
    .Y(_19767_));
 NAND2x1_ASAP7_75t_R _28283_ (.A(net2680),
    .B(net1857),
    .Y(_19768_));
 NAND2x1_ASAP7_75t_R _28284_ (.A(_18107_),
    .B(_18131_),
    .Y(_19769_));
 AND4x1_ASAP7_75t_R _28285_ (.A(_19767_),
    .B(_19768_),
    .C(_19769_),
    .D(_18111_),
    .Y(_19770_));
 AO21x1_ASAP7_75t_R _28286_ (.A1(net2908),
    .A2(net974),
    .B(_18126_),
    .Y(_19771_));
 OA21x2_ASAP7_75t_R _28287_ (.A1(net3306),
    .A2(_18126_),
    .B(_19771_),
    .Y(_19772_));
 AND2x2_ASAP7_75t_R _28288_ (.A(_19770_),
    .B(_19772_),
    .Y(_19773_));
 AO21x1_ASAP7_75t_R _28289_ (.A1(_17984_),
    .A2(_17987_),
    .B(_17968_),
    .Y(_19774_));
 INVx1_ASAP7_75t_R _28290_ (.A(_18095_),
    .Y(_19775_));
 NAND2x1_ASAP7_75t_R _28291_ (.A(net3367),
    .B(_18089_),
    .Y(_19776_));
 NAND3x1_ASAP7_75t_R _28292_ (.A(_19774_),
    .B(_19775_),
    .C(_19776_),
    .Y(_19777_));
 INVx1_ASAP7_75t_R _28293_ (.A(_19777_),
    .Y(_19778_));
 AO21x1_ASAP7_75t_R _28294_ (.A1(net1795),
    .A2(net939),
    .B(net1746),
    .Y(_19779_));
 AO21x1_ASAP7_75t_R _28295_ (.A1(_17963_),
    .A2(net2757),
    .B(net1746),
    .Y(_19780_));
 AND2x2_ASAP7_75t_R _28296_ (.A(_19779_),
    .B(_19780_),
    .Y(_19781_));
 AO21x1_ASAP7_75t_R _28297_ (.A1(net3306),
    .A2(net3189),
    .B(net1746),
    .Y(_19782_));
 NAND2x1_ASAP7_75t_R _28298_ (.A(net3219),
    .B(_17932_),
    .Y(_19783_));
 AND2x2_ASAP7_75t_R _28299_ (.A(_19782_),
    .B(_19783_),
    .Y(_19784_));
 NAND3x1_ASAP7_75t_R _28300_ (.A(_19778_),
    .B(_19781_),
    .C(_19784_),
    .Y(_19785_));
 INVx1_ASAP7_75t_R _28301_ (.A(_19785_),
    .Y(_19786_));
 NAND2x1_ASAP7_75t_R _28302_ (.A(_19773_),
    .B(_19786_),
    .Y(_19787_));
 AO21x1_ASAP7_75t_R _28303_ (.A1(_18014_),
    .A2(_17999_),
    .B(_19423_),
    .Y(_19788_));
 NAND2x1_ASAP7_75t_R _28304_ (.A(_18175_),
    .B(net3207),
    .Y(_19789_));
 AND2x2_ASAP7_75t_R _28305_ (.A(_18175_),
    .B(_18150_),
    .Y(_19790_));
 INVx1_ASAP7_75t_R _28306_ (.A(_19790_),
    .Y(_19791_));
 AND3x2_ASAP7_75t_R _28307_ (.A(_19788_),
    .B(_19789_),
    .C(_19791_),
    .Y(_19792_));
 AO21x1_ASAP7_75t_R _28308_ (.A1(net3188),
    .A2(net1839),
    .B(_18169_),
    .Y(_19793_));
 NAND2x1_ASAP7_75t_R _28309_ (.A(_19421_),
    .B(_19793_),
    .Y(_19794_));
 OA31x2_ASAP7_75t_R _28310_ (.A1(_18134_),
    .A2(_18923_),
    .A3(_18131_),
    .B1(net3299),
    .Y(_19795_));
 NOR2x2_ASAP7_75t_R _28311_ (.A(_19794_),
    .B(_19795_),
    .Y(_19796_));
 OAI22x1_ASAP7_75t_R _28312_ (.A1(_18185_),
    .A2(_17937_),
    .B1(_19423_),
    .B2(net1795),
    .Y(_19797_));
 INVx1_ASAP7_75t_R _28313_ (.A(_19797_),
    .Y(_19798_));
 NAND3x2_ASAP7_75t_R _28314_ (.B(_19796_),
    .C(_19798_),
    .Y(_19799_),
    .A(_19792_));
 INVx1_ASAP7_75t_R _28315_ (.A(_19799_),
    .Y(_19800_));
 AO21x1_ASAP7_75t_R _28316_ (.A1(_18010_),
    .A2(_18081_),
    .B(_18156_),
    .Y(_19801_));
 NOR2x2_ASAP7_75t_R _28317_ (.A(net1071),
    .B(net1543),
    .Y(_19802_));
 NAND2x1_ASAP7_75t_R _28318_ (.A(_19802_),
    .B(net3192),
    .Y(_19803_));
 AND3x2_ASAP7_75t_R _28319_ (.A(_19801_),
    .B(_19803_),
    .C(_18890_),
    .Y(_19804_));
 AO21x2_ASAP7_75t_R _28320_ (.A1(_18052_),
    .A2(net1622),
    .B(net2946),
    .Y(_19805_));
 NAND2x2_ASAP7_75t_R _28321_ (.A(_19416_),
    .B(_19805_),
    .Y(_19806_));
 AO21x1_ASAP7_75t_R _28322_ (.A1(_18883_),
    .A2(_18073_),
    .B(net2446),
    .Y(_19807_));
 OAI21x1_ASAP7_75t_R _28323_ (.A1(net3284),
    .A2(net2446),
    .B(_19807_),
    .Y(_19808_));
 NOR2x2_ASAP7_75t_R _28324_ (.A(_19808_),
    .B(_19806_),
    .Y(_19809_));
 AO21x1_ASAP7_75t_R _28325_ (.A1(net1121),
    .A2(_17980_),
    .B(_18156_),
    .Y(_19810_));
 OA21x2_ASAP7_75t_R _28326_ (.A1(_18156_),
    .A2(net1693),
    .B(_19810_),
    .Y(_19811_));
 NAND3x2_ASAP7_75t_R _28327_ (.B(_19809_),
    .C(_19811_),
    .Y(_19812_),
    .A(_19804_));
 INVx1_ASAP7_75t_R _28328_ (.A(_19812_),
    .Y(_19813_));
 NAND2x1_ASAP7_75t_R _28329_ (.A(_19800_),
    .B(_19813_),
    .Y(_19814_));
 NOR2x2_ASAP7_75t_R _28330_ (.A(_19787_),
    .B(_19814_),
    .Y(_19815_));
 AO21x1_ASAP7_75t_R _28331_ (.A1(net2821),
    .A2(net974),
    .B(net2303),
    .Y(_19816_));
 AO21x1_ASAP7_75t_R _28332_ (.A1(_18022_),
    .A2(_18958_),
    .B(net2303),
    .Y(_19817_));
 NAND2x2_ASAP7_75t_R _28333_ (.A(net2878),
    .B(_18952_),
    .Y(_19818_));
 NAND3x2_ASAP7_75t_R _28334_ (.B(_19817_),
    .C(_19818_),
    .Y(_19819_),
    .A(_19816_));
 NAND2x1_ASAP7_75t_R _28335_ (.A(_18040_),
    .B(_18070_),
    .Y(_19820_));
 AO21x1_ASAP7_75t_R _28336_ (.A1(_18147_),
    .A2(net2757),
    .B(net3305),
    .Y(_19821_));
 NAND2x2_ASAP7_75t_R _28337_ (.A(_19820_),
    .B(_19821_),
    .Y(_19822_));
 NOR2x1_ASAP7_75t_R _28338_ (.A(net3285),
    .B(net3304),
    .Y(_19823_));
 INVx2_ASAP7_75t_R _28339_ (.A(_19823_),
    .Y(_19824_));
 AO21x1_ASAP7_75t_R _28340_ (.A1(_18883_),
    .A2(_18022_),
    .B(net3305),
    .Y(_19825_));
 NAND2x2_ASAP7_75t_R _28341_ (.A(_19824_),
    .B(_19825_),
    .Y(_19826_));
 NOR3x2_ASAP7_75t_R _28342_ (.B(_19822_),
    .C(_19826_),
    .Y(_19827_),
    .A(_19819_));
 AO21x1_ASAP7_75t_R _28343_ (.A1(_18010_),
    .A2(net1532),
    .B(net2181),
    .Y(_19828_));
 AO21x1_ASAP7_75t_R _28344_ (.A1(net939),
    .A2(_17987_),
    .B(net2181),
    .Y(_19829_));
 AND2x2_ASAP7_75t_R _28345_ (.A(_19828_),
    .B(_19829_),
    .Y(_19830_));
 AOI211x1_ASAP7_75t_R _28346_ (.A1(net1062),
    .A2(net3124),
    .B(net2181),
    .C(net3284),
    .Y(_19831_));
 NOR2x1_ASAP7_75t_R _28347_ (.A(_18022_),
    .B(_18074_),
    .Y(_19832_));
 AOI211x1_ASAP7_75t_R _28348_ (.A1(_18869_),
    .A2(_18941_),
    .B(_19831_),
    .C(_19832_),
    .Y(_19833_));
 NAND2x1_ASAP7_75t_R _28349_ (.A(_19830_),
    .B(_19833_),
    .Y(_19834_));
 AO21x1_ASAP7_75t_R _28350_ (.A1(net1691),
    .A2(_18073_),
    .B(net1907),
    .Y(_19835_));
 OA21x2_ASAP7_75t_R _28351_ (.A1(net1121),
    .A2(net1907),
    .B(_19835_),
    .Y(_19836_));
 AO21x1_ASAP7_75t_R _28352_ (.A1(net3301),
    .A2(_17962_),
    .B(net1907),
    .Y(_19837_));
 NAND2x1_ASAP7_75t_R _28353_ (.A(net1857),
    .B(_18069_),
    .Y(_19838_));
 AND3x1_ASAP7_75t_R _28354_ (.A(_19837_),
    .B(_18071_),
    .C(_19838_),
    .Y(_19839_));
 NAND2x1_ASAP7_75t_R _28355_ (.A(_19836_),
    .B(_19839_),
    .Y(_19840_));
 NOR2x2_ASAP7_75t_R _28356_ (.A(_19834_),
    .B(_19840_),
    .Y(_19841_));
 NAND2x2_ASAP7_75t_R _28357_ (.A(_19827_),
    .B(_19841_),
    .Y(_19842_));
 AO21x1_ASAP7_75t_R _28358_ (.A1(net1532),
    .A2(net3217),
    .B(net3205),
    .Y(_19843_));
 AO21x1_ASAP7_75t_R _28359_ (.A1(net939),
    .A2(net974),
    .B(net3205),
    .Y(_19844_));
 NAND2x1_ASAP7_75t_R _28360_ (.A(_19376_),
    .B(_18070_),
    .Y(_19845_));
 AND3x1_ASAP7_75t_R _28361_ (.A(_19843_),
    .B(_19844_),
    .C(_19845_),
    .Y(_19846_));
 AO21x1_ASAP7_75t_R _28362_ (.A1(_17938_),
    .A2(_18022_),
    .B(net1955),
    .Y(_19847_));
 AO21x1_ASAP7_75t_R _28363_ (.A1(_18057_),
    .A2(_18958_),
    .B(net1955),
    .Y(_19848_));
 AND2x2_ASAP7_75t_R _28364_ (.A(_19847_),
    .B(_19848_),
    .Y(_19849_));
 AND2x2_ASAP7_75t_R _28365_ (.A(_19846_),
    .B(_19849_),
    .Y(_19850_));
 AO21x1_ASAP7_75t_R _28366_ (.A1(net2908),
    .A2(_19361_),
    .B(_18024_),
    .Y(_19851_));
 NAND2x1_ASAP7_75t_R _28367_ (.A(net3196),
    .B(_17925_),
    .Y(_19852_));
 OA21x2_ASAP7_75t_R _28368_ (.A1(_18021_),
    .A2(_18164_),
    .B(_19852_),
    .Y(_19853_));
 NAND2x1_ASAP7_75t_R _28369_ (.A(_19851_),
    .B(_19853_),
    .Y(_19854_));
 AO21x2_ASAP7_75t_R _28370_ (.A1(_18036_),
    .A2(_17983_),
    .B(net1365),
    .Y(_19855_));
 AO21x1_ASAP7_75t_R _28371_ (.A1(_19855_),
    .A2(net3284),
    .B(net3123),
    .Y(_19856_));
 AO21x1_ASAP7_75t_R _28372_ (.A1(net1795),
    .A2(net974),
    .B(net3123),
    .Y(_19857_));
 NAND3x2_ASAP7_75t_R _28373_ (.B(_19359_),
    .C(_19857_),
    .Y(_19858_),
    .A(_19856_));
 NOR2x2_ASAP7_75t_R _28374_ (.A(_19854_),
    .B(_19858_),
    .Y(_19859_));
 AO21x1_ASAP7_75t_R _28375_ (.A1(_18881_),
    .A2(net1068),
    .B(_17997_),
    .Y(_19860_));
 AO21x1_ASAP7_75t_R _28376_ (.A1(net3187),
    .A2(net1623),
    .B(_17997_),
    .Y(_19861_));
 AND3x4_ASAP7_75t_R _28377_ (.A(_18928_),
    .B(_19860_),
    .C(_19861_),
    .Y(_19862_));
 NAND3x2_ASAP7_75t_R _28378_ (.B(_19859_),
    .C(_19862_),
    .Y(_19863_),
    .A(_19850_));
 NOR2x2_ASAP7_75t_R _28379_ (.A(_19863_),
    .B(_19842_),
    .Y(_19864_));
 AO21x1_ASAP7_75t_R _28380_ (.A1(_17572_),
    .A2(_17562_),
    .B(_17691_),
    .Y(_19865_));
 INVx1_ASAP7_75t_R _28381_ (.A(_17693_),
    .Y(_19866_));
 NAND2x1_ASAP7_75t_R _28382_ (.A(_17801_),
    .B(_17576_),
    .Y(_19867_));
 NAND3x1_ASAP7_75t_R _28383_ (.A(_19865_),
    .B(_19866_),
    .C(_19867_),
    .Y(_19868_));
 AO21x1_ASAP7_75t_R _28384_ (.A1(_17845_),
    .A2(_17624_),
    .B(_17701_),
    .Y(_19869_));
 AO21x1_ASAP7_75t_R _28385_ (.A1(_17685_),
    .A2(net2597),
    .B(_17701_),
    .Y(_19870_));
 NAND2x1_ASAP7_75t_R _28386_ (.A(_19869_),
    .B(_19870_),
    .Y(_19871_));
 AO21x1_ASAP7_75t_R _28387_ (.A1(_17813_),
    .A2(net2385),
    .B(_17701_),
    .Y(_19872_));
 OAI21x1_ASAP7_75t_R _28388_ (.A1(_17701_),
    .A2(net1082),
    .B(_19872_),
    .Y(_19873_));
 NOR3x1_ASAP7_75t_R _28389_ (.A(_19868_),
    .B(_19871_),
    .C(_19873_),
    .Y(_19874_));
 AO21x1_ASAP7_75t_R _28390_ (.A1(net2598),
    .A2(net1381),
    .B(_17725_),
    .Y(_19875_));
 NAND2x2_ASAP7_75t_R _28391_ (.A(_17616_),
    .B(_17733_),
    .Y(_19876_));
 AND3x1_ASAP7_75t_R _28392_ (.A(_19875_),
    .B(_17820_),
    .C(_19876_),
    .Y(_19877_));
 AO21x1_ASAP7_75t_R _28393_ (.A1(_17756_),
    .A2(net1381),
    .B(net2881),
    .Y(_19878_));
 OA21x2_ASAP7_75t_R _28394_ (.A1(_17813_),
    .A2(net2881),
    .B(_19878_),
    .Y(_19879_));
 AND2x2_ASAP7_75t_R _28395_ (.A(_19879_),
    .B(_19877_),
    .Y(_19880_));
 AND2x4_ASAP7_75t_R _28396_ (.A(_19880_),
    .B(_19874_),
    .Y(_19881_));
 AO21x1_ASAP7_75t_R _28397_ (.A1(_17813_),
    .A2(net2385),
    .B(_17759_),
    .Y(_19882_));
 OAI21x1_ASAP7_75t_R _28398_ (.A1(net1098),
    .A2(_17759_),
    .B(_19882_),
    .Y(_19883_));
 AO21x1_ASAP7_75t_R _28399_ (.A1(_17626_),
    .A2(_17695_),
    .B(_17759_),
    .Y(_19884_));
 INVx1_ASAP7_75t_R _28400_ (.A(_18827_),
    .Y(_19885_));
 NAND2x1_ASAP7_75t_R _28401_ (.A(_19884_),
    .B(_19885_),
    .Y(_19886_));
 NOR2x1_ASAP7_75t_R _28402_ (.A(_19883_),
    .B(_19886_),
    .Y(_19887_));
 AO21x2_ASAP7_75t_R _28403_ (.A1(net2598),
    .A2(net1381),
    .B(_17744_),
    .Y(_19888_));
 AO21x1_ASAP7_75t_R _28404_ (.A1(_17834_),
    .A2(_17647_),
    .B(_17744_),
    .Y(_19889_));
 NOR2x2_ASAP7_75t_R _28405_ (.A(_17617_),
    .B(_17781_),
    .Y(_19890_));
 NAND2x1_ASAP7_75t_R _28406_ (.A(_19890_),
    .B(_17788_),
    .Y(_19891_));
 NAND2x1_ASAP7_75t_R _28407_ (.A(net1007),
    .B(_19890_),
    .Y(_19892_));
 AND4x1_ASAP7_75t_R _28408_ (.A(_19888_),
    .B(_19889_),
    .C(_19891_),
    .D(_19892_),
    .Y(_19893_));
 NAND2x1_ASAP7_75t_R _28409_ (.A(_19887_),
    .B(_19893_),
    .Y(_19894_));
 AOI22x1_ASAP7_75t_R _28410_ (.A1(_18813_),
    .A2(_17555_),
    .B1(net1901),
    .B2(_17782_),
    .Y(_19895_));
 AO21x1_ASAP7_75t_R _28411_ (.A1(_17593_),
    .A2(_17596_),
    .B(_17777_),
    .Y(_19896_));
 AO21x1_ASAP7_75t_R _28412_ (.A1(net2013),
    .A2(_17586_),
    .B(_17777_),
    .Y(_19897_));
 AND2x2_ASAP7_75t_R _28413_ (.A(_19896_),
    .B(_19897_),
    .Y(_19898_));
 AND2x2_ASAP7_75t_R _28414_ (.A(_19895_),
    .B(_19898_),
    .Y(_19899_));
 AO21x1_ASAP7_75t_R _28415_ (.A1(_17685_),
    .A2(net2599),
    .B(net2758),
    .Y(_19900_));
 AO21x1_ASAP7_75t_R _28416_ (.A1(_17639_),
    .A2(net2236),
    .B(net2758),
    .Y(_19901_));
 NAND2x1_ASAP7_75t_R _28417_ (.A(_17788_),
    .B(_17771_),
    .Y(_19902_));
 NAND2x1_ASAP7_75t_R _28418_ (.A(_17678_),
    .B(_17771_),
    .Y(_19903_));
 AND4x1_ASAP7_75t_R _28419_ (.A(_19900_),
    .B(_19901_),
    .C(_19902_),
    .D(_19903_),
    .Y(_19904_));
 NAND2x1_ASAP7_75t_R _28420_ (.A(_19904_),
    .B(_19899_),
    .Y(_19905_));
 NOR2x1_ASAP7_75t_R _28421_ (.A(_19894_),
    .B(_19905_),
    .Y(_19906_));
 NAND2x2_ASAP7_75t_R _28422_ (.A(_19881_),
    .B(_19906_),
    .Y(_19907_));
 INVx2_ASAP7_75t_R _28423_ (.A(_19907_),
    .Y(_19908_));
 AO21x1_ASAP7_75t_R _28424_ (.A1(_17756_),
    .A2(net941),
    .B(net3313),
    .Y(_19909_));
 AO21x1_ASAP7_75t_R _28425_ (.A1(net1082),
    .A2(_17586_),
    .B(net3313),
    .Y(_19910_));
 NAND2x1_ASAP7_75t_R _28426_ (.A(net2640),
    .B(_17671_),
    .Y(_19911_));
 NAND3x1_ASAP7_75t_R _28427_ (.A(_19909_),
    .B(_19910_),
    .C(_19911_),
    .Y(_19912_));
 NOR3x1_ASAP7_75t_R _28428_ (.A(_17887_),
    .B(_18799_),
    .C(_17659_),
    .Y(_19913_));
 NOR2x1_ASAP7_75t_R _28429_ (.A(_17657_),
    .B(_17756_),
    .Y(_19914_));
 INVx1_ASAP7_75t_R _28430_ (.A(_19914_),
    .Y(_19915_));
 AO21x1_ASAP7_75t_R _28431_ (.A1(_17758_),
    .A2(net2899),
    .B(net2847),
    .Y(_19916_));
 NAND3x1_ASAP7_75t_R _28432_ (.A(_19913_),
    .B(_19915_),
    .C(_19916_),
    .Y(_19917_));
 NOR2x1_ASAP7_75t_R _28433_ (.A(_19912_),
    .B(_19917_),
    .Y(_19918_));
 AO21x1_ASAP7_75t_R _28434_ (.A1(_17756_),
    .A2(net1380),
    .B(_17641_),
    .Y(_19919_));
 AOI211x1_ASAP7_75t_R _28435_ (.A1(net1123),
    .A2(net2891),
    .B(_17641_),
    .C(net1103),
    .Y(_19920_));
 INVx1_ASAP7_75t_R _28436_ (.A(_19920_),
    .Y(_19921_));
 NAND2x1_ASAP7_75t_R _28437_ (.A(_19919_),
    .B(_19921_),
    .Y(_19922_));
 NOR2x1_ASAP7_75t_R _28438_ (.A(_17641_),
    .B(net2894),
    .Y(_19923_));
 NOR3x1_ASAP7_75t_R _28439_ (.A(_19923_),
    .B(_17646_),
    .C(_17648_),
    .Y(_19924_));
 INVx1_ASAP7_75t_R _28440_ (.A(_19924_),
    .Y(_19925_));
 NOR2x1_ASAP7_75t_R _28441_ (.A(_19922_),
    .B(_19925_),
    .Y(_19926_));
 INVx1_ASAP7_75t_R _28442_ (.A(_19926_),
    .Y(_19927_));
 AO21x1_ASAP7_75t_R _28443_ (.A1(_17845_),
    .A2(_17665_),
    .B(_17629_),
    .Y(_19928_));
 AO21x1_ASAP7_75t_R _28444_ (.A1(net997),
    .A2(_17562_),
    .B(_17629_),
    .Y(_19929_));
 AND2x2_ASAP7_75t_R _28445_ (.A(_19928_),
    .B(_19929_),
    .Y(_19930_));
 AO21x1_ASAP7_75t_R _28446_ (.A1(_17834_),
    .A2(net1816),
    .B(_17629_),
    .Y(_19931_));
 AOI211x1_ASAP7_75t_R _28447_ (.A1(net1123),
    .A2(net2879),
    .B(_17629_),
    .C(_17575_),
    .Y(_19932_));
 INVx1_ASAP7_75t_R _28448_ (.A(_19932_),
    .Y(_19933_));
 NAND3x2_ASAP7_75t_R _28449_ (.B(_19931_),
    .C(_19933_),
    .Y(_19934_),
    .A(_19930_));
 NOR2x2_ASAP7_75t_R _28450_ (.A(_19927_),
    .B(_19934_),
    .Y(_19935_));
 NAND2x2_ASAP7_75t_R _28451_ (.A(_19918_),
    .B(_19935_),
    .Y(_19936_));
 AO21x1_ASAP7_75t_R _28452_ (.A1(_17845_),
    .A2(net2901),
    .B(_17566_),
    .Y(_19937_));
 AO21x1_ASAP7_75t_R _28453_ (.A1(net997),
    .A2(net1380),
    .B(_17566_),
    .Y(_19938_));
 NAND2x1_ASAP7_75t_R _28454_ (.A(_17558_),
    .B(_17569_),
    .Y(_19939_));
 AND3x1_ASAP7_75t_R _28455_ (.A(_19937_),
    .B(_19938_),
    .C(_19939_),
    .Y(_19940_));
 AO21x1_ASAP7_75t_R _28456_ (.A1(_17639_),
    .A2(net1816),
    .B(_17566_),
    .Y(_19941_));
 AO21x1_ASAP7_75t_R _28457_ (.A1(net2015),
    .A2(_17586_),
    .B(_17566_),
    .Y(_19942_));
 AND2x2_ASAP7_75t_R _28458_ (.A(_19941_),
    .B(_19942_),
    .Y(_19943_));
 AND2x2_ASAP7_75t_R _28459_ (.A(_19940_),
    .B(_19943_),
    .Y(_19944_));
 AO21x1_ASAP7_75t_R _28460_ (.A1(_17746_),
    .A2(_17756_),
    .B(_17589_),
    .Y(_19945_));
 AO21x1_ASAP7_75t_R _28461_ (.A1(net2013),
    .A2(net1081),
    .B(_17589_),
    .Y(_19946_));
 AO21x2_ASAP7_75t_R _28462_ (.A1(_17815_),
    .A2(net2892),
    .B(_17589_),
    .Y(_19947_));
 NAND3x2_ASAP7_75t_R _28463_ (.B(_19946_),
    .C(_19947_),
    .Y(_19948_),
    .A(_19945_));
 AO31x2_ASAP7_75t_R _28464_ (.A1(net2202),
    .A2(net941),
    .A3(_17695_),
    .B(_17614_),
    .Y(_19949_));
 NAND2x1_ASAP7_75t_R _28465_ (.A(net1002),
    .B(_17618_),
    .Y(_19950_));
 AND2x2_ASAP7_75t_R _28466_ (.A(_17855_),
    .B(_19950_),
    .Y(_19951_));
 NAND2x1_ASAP7_75t_R _28467_ (.A(_19949_),
    .B(_19951_),
    .Y(_19952_));
 NOR2x2_ASAP7_75t_R _28468_ (.A(_19948_),
    .B(_19952_),
    .Y(_19953_));
 AO21x1_ASAP7_75t_R _28469_ (.A1(_17756_),
    .A2(net1380),
    .B(_17547_),
    .Y(_19954_));
 AO21x1_ASAP7_75t_R _28470_ (.A1(net1788),
    .A2(net2630),
    .B(_17547_),
    .Y(_19955_));
 NAND2x1_ASAP7_75t_R _28471_ (.A(_17694_),
    .B(_17548_),
    .Y(_19956_));
 AND3x2_ASAP7_75t_R _28472_ (.A(_19954_),
    .B(_19955_),
    .C(_19956_),
    .Y(_19957_));
 NAND3x2_ASAP7_75t_R _28473_ (.B(_19953_),
    .C(_19957_),
    .Y(_19958_),
    .A(_19944_));
 NOR2x2_ASAP7_75t_R _28474_ (.A(_19936_),
    .B(_19958_),
    .Y(_19959_));
 AOI22x1_ASAP7_75t_R _28475_ (.A1(_19815_),
    .A2(_19864_),
    .B1(_19908_),
    .B2(_19959_),
    .Y(_19960_));
 NAND2x2_ASAP7_75t_R _28476_ (.A(_19959_),
    .B(_19908_),
    .Y(_19961_));
 NAND2x2_ASAP7_75t_R _28477_ (.A(_19864_),
    .B(_19815_),
    .Y(_19962_));
 NOR2x2_ASAP7_75t_R _28478_ (.A(_19961_),
    .B(_19962_),
    .Y(_19963_));
 AO21x2_ASAP7_75t_R _28479_ (.A1(net2753),
    .A2(net1482),
    .B(_18464_),
    .Y(_19964_));
 NAND2x2_ASAP7_75t_R _28480_ (.A(_18482_),
    .B(_18469_),
    .Y(_19965_));
 NOR2x1_ASAP7_75t_R _28481_ (.A(net2109),
    .B(net3312),
    .Y(_19966_));
 INVx1_ASAP7_75t_R _28482_ (.A(_19966_),
    .Y(_19967_));
 NAND3x2_ASAP7_75t_R _28483_ (.B(_19965_),
    .C(_19967_),
    .Y(_19968_),
    .A(_19964_));
 AO21x2_ASAP7_75t_R _28484_ (.A1(net1087),
    .A2(_18237_),
    .B(net2093),
    .Y(_19969_));
 AO21x1_ASAP7_75t_R _28485_ (.A1(_19969_),
    .A2(_19164_),
    .B(_18456_),
    .Y(_19970_));
 NAND2x2_ASAP7_75t_R _28486_ (.A(_18259_),
    .B(_19185_),
    .Y(_19971_));
 AO21x1_ASAP7_75t_R _28487_ (.A1(net2963),
    .A2(net1254),
    .B(_18456_),
    .Y(_19972_));
 NAND3x2_ASAP7_75t_R _28488_ (.B(_19971_),
    .C(_19972_),
    .Y(_19973_),
    .A(_19970_));
 NOR2x2_ASAP7_75t_R _28489_ (.A(_19968_),
    .B(_19973_),
    .Y(_19974_));
 AO21x1_ASAP7_75t_R _28490_ (.A1(net2176),
    .A2(net1954),
    .B(net3282),
    .Y(_19975_));
 AO21x1_ASAP7_75t_R _28491_ (.A1(net2004),
    .A2(_18335_),
    .B(net3282),
    .Y(_19976_));
 NAND2x1_ASAP7_75t_R _28492_ (.A(_18444_),
    .B(_18483_),
    .Y(_19977_));
 AND4x2_ASAP7_75t_R _28493_ (.A(_19180_),
    .B(_19975_),
    .C(_19976_),
    .D(_19977_),
    .Y(_19978_));
 AO21x1_ASAP7_75t_R _28494_ (.A1(net2634),
    .A2(net1335),
    .B(net2595),
    .Y(_19979_));
 NAND2x1_ASAP7_75t_R _28495_ (.A(net1390),
    .B(net2533),
    .Y(_19980_));
 AO21x1_ASAP7_75t_R _28496_ (.A1(_19980_),
    .A2(net2004),
    .B(net2595),
    .Y(_19981_));
 AND3x2_ASAP7_75t_R _28497_ (.A(_19979_),
    .B(_19981_),
    .C(_19473_),
    .Y(_19982_));
 NAND3x2_ASAP7_75t_R _28498_ (.B(_19978_),
    .C(_19982_),
    .Y(_19983_),
    .A(_19974_));
 AO21x1_ASAP7_75t_R _28499_ (.A1(_19969_),
    .A2(net1821),
    .B(_18266_),
    .Y(_19984_));
 NAND2x1_ASAP7_75t_R _28500_ (.A(_18306_),
    .B(_18416_),
    .Y(_19985_));
 NAND3x1_ASAP7_75t_R _28501_ (.A(_19984_),
    .B(_19985_),
    .C(_18415_),
    .Y(_19986_));
 AO21x1_ASAP7_75t_R _28502_ (.A1(net2452),
    .A2(net2638),
    .B(_18248_),
    .Y(_19987_));
 OA21x2_ASAP7_75t_R _28503_ (.A1(_18444_),
    .A2(_18445_),
    .B(_18247_),
    .Y(_19988_));
 INVx1_ASAP7_75t_R _28504_ (.A(_19988_),
    .Y(_19989_));
 NAND2x1_ASAP7_75t_R _28505_ (.A(_19987_),
    .B(_19989_),
    .Y(_19990_));
 OA31x2_ASAP7_75t_R _28506_ (.A1(_18401_),
    .A2(_18306_),
    .A3(_18468_),
    .B1(_18247_),
    .Y(_19991_));
 NOR3x1_ASAP7_75t_R _28507_ (.A(_19986_),
    .B(_19990_),
    .C(_19991_),
    .Y(_19992_));
 OA21x2_ASAP7_75t_R _28508_ (.A1(_19156_),
    .A2(_18291_),
    .B(_18434_),
    .Y(_19993_));
 AO21x1_ASAP7_75t_R _28509_ (.A1(_18306_),
    .A2(_18434_),
    .B(_19993_),
    .Y(_19994_));
 NOR2x1_ASAP7_75t_R _28510_ (.A(net2989),
    .B(net2452),
    .Y(_19995_));
 NOR2x1_ASAP7_75t_R _28511_ (.A(net2989),
    .B(net2634),
    .Y(_19996_));
 NOR2x1_ASAP7_75t_R _28512_ (.A(net1482),
    .B(net2989),
    .Y(_19997_));
 OR3x1_ASAP7_75t_R _28513_ (.A(_19995_),
    .B(_19996_),
    .C(_19997_),
    .Y(_19998_));
 AOI211x1_ASAP7_75t_R _28514_ (.A1(_19465_),
    .A2(_18446_),
    .B(_19994_),
    .C(_19998_),
    .Y(_19999_));
 NAND2x1_ASAP7_75t_R _28515_ (.A(_19992_),
    .B(_19999_),
    .Y(_20000_));
 NOR2x2_ASAP7_75t_R _28516_ (.A(_19983_),
    .B(_20000_),
    .Y(_20001_));
 AO21x1_ASAP7_75t_R _28517_ (.A1(net2965),
    .A2(net937),
    .B(net3178),
    .Y(_20002_));
 AO21x1_ASAP7_75t_R _28518_ (.A1(net2419),
    .A2(_18335_),
    .B(net3178),
    .Y(_20003_));
 NAND2x1_ASAP7_75t_R _28519_ (.A(net2668),
    .B(_19237_),
    .Y(_20004_));
 NAND3x1_ASAP7_75t_R _28520_ (.A(_20002_),
    .B(_20003_),
    .C(_20004_),
    .Y(_20005_));
 AO31x2_ASAP7_75t_R _28521_ (.A1(net2095),
    .A2(net2976),
    .A3(net1954),
    .B(_18364_),
    .Y(_20006_));
 AO21x1_ASAP7_75t_R _28522_ (.A1(net3183),
    .A2(net3003),
    .B(_18364_),
    .Y(_20007_));
 NAND3x1_ASAP7_75t_R _28523_ (.A(_20006_),
    .B(_19547_),
    .C(_20007_),
    .Y(_20008_));
 NOR2x1_ASAP7_75t_R _28524_ (.A(_20005_),
    .B(_20008_),
    .Y(_20009_));
 AO21x1_ASAP7_75t_R _28525_ (.A1(_18381_),
    .A2(_18394_),
    .B(_18395_),
    .Y(_20010_));
 AO21x1_ASAP7_75t_R _28526_ (.A1(net2965),
    .A2(net937),
    .B(_18395_),
    .Y(_20011_));
 AO21x1_ASAP7_75t_R _28527_ (.A1(_18419_),
    .A2(net1254),
    .B(_18395_),
    .Y(_20012_));
 NAND3x1_ASAP7_75t_R _28528_ (.A(_20010_),
    .B(_20011_),
    .C(_20012_),
    .Y(_20013_));
 AO21x1_ASAP7_75t_R _28529_ (.A1(net2096),
    .A2(net2419),
    .B(_18377_),
    .Y(_20014_));
 AO21x1_ASAP7_75t_R _28530_ (.A1(net2671),
    .A2(net2437),
    .B(_18377_),
    .Y(_20015_));
 NAND2x1_ASAP7_75t_R _28531_ (.A(_19224_),
    .B(_18306_),
    .Y(_20016_));
 AND3x1_ASAP7_75t_R _28532_ (.A(_20014_),
    .B(_20015_),
    .C(_20016_),
    .Y(_20017_));
 AO21x1_ASAP7_75t_R _28533_ (.A1(net2045),
    .A2(net2452),
    .B(net2981),
    .Y(_20018_));
 AND3x1_ASAP7_75t_R _28534_ (.A(_20018_),
    .B(_18380_),
    .C(_19226_),
    .Y(_20019_));
 NAND2x1_ASAP7_75t_R _28535_ (.A(_20017_),
    .B(_20019_),
    .Y(_20020_));
 NOR2x1_ASAP7_75t_R _28536_ (.A(_20013_),
    .B(_20020_),
    .Y(_20021_));
 NAND2x1_ASAP7_75t_R _28537_ (.A(_20009_),
    .B(_20021_),
    .Y(_20022_));
 AO21x1_ASAP7_75t_R _28538_ (.A1(net2965),
    .A2(_19493_),
    .B(_18330_),
    .Y(_20023_));
 AO21x1_ASAP7_75t_R _28539_ (.A1(_18489_),
    .A2(_18350_),
    .B(_18330_),
    .Y(_20024_));
 NAND2x1_ASAP7_75t_R _28540_ (.A(_20023_),
    .B(_20024_),
    .Y(_20025_));
 AO21x1_ASAP7_75t_R _28541_ (.A1(net2699),
    .A2(net937),
    .B(_18318_),
    .Y(_20026_));
 NAND2x1_ASAP7_75t_R _28542_ (.A(_19522_),
    .B(_20026_),
    .Y(_20027_));
 AO21x2_ASAP7_75t_R _28543_ (.A1(net2476),
    .A2(net2505),
    .B(_18318_),
    .Y(_20028_));
 NAND3x1_ASAP7_75t_R _28544_ (.A(_20028_),
    .B(_18324_),
    .C(_19521_),
    .Y(_20029_));
 NOR3x1_ASAP7_75t_R _28545_ (.A(_20025_),
    .B(_20027_),
    .C(_20029_),
    .Y(_20030_));
 NOR2x1_ASAP7_75t_R _28546_ (.A(net1483),
    .B(_18287_),
    .Y(_20031_));
 INVx1_ASAP7_75t_R _28547_ (.A(_20031_),
    .Y(_20032_));
 NAND2x1_ASAP7_75t_R _28548_ (.A(_18293_),
    .B(_20032_),
    .Y(_20033_));
 NOR2x1_ASAP7_75t_R _28549_ (.A(_18394_),
    .B(net2985),
    .Y(_20034_));
 OA21x2_ASAP7_75t_R _28550_ (.A1(_19223_),
    .A2(_19202_),
    .B(_18292_),
    .Y(_20035_));
 OR3x1_ASAP7_75t_R _28551_ (.A(_20033_),
    .B(_20034_),
    .C(_20035_),
    .Y(_20036_));
 AO21x1_ASAP7_75t_R _28552_ (.A1(_18402_),
    .A2(net1954),
    .B(_18300_),
    .Y(_20037_));
 AO21x1_ASAP7_75t_R _28553_ (.A1(net2107),
    .A2(net2437),
    .B(_18300_),
    .Y(_20038_));
 NAND2x1_ASAP7_75t_R _28554_ (.A(_19465_),
    .B(_18303_),
    .Y(_20039_));
 AND3x1_ASAP7_75t_R _28555_ (.A(_20037_),
    .B(_20038_),
    .C(_20039_),
    .Y(_20040_));
 AO21x1_ASAP7_75t_R _28556_ (.A1(net1754),
    .A2(net1483),
    .B(_18300_),
    .Y(_20041_));
 AO21x1_ASAP7_75t_R _28557_ (.A1(net2452),
    .A2(net2638),
    .B(_18300_),
    .Y(_20042_));
 NAND2x1_ASAP7_75t_R _28558_ (.A(_18291_),
    .B(_18303_),
    .Y(_20043_));
 AND3x1_ASAP7_75t_R _28559_ (.A(_20041_),
    .B(_20042_),
    .C(_20043_),
    .Y(_20044_));
 NAND2x1_ASAP7_75t_R _28560_ (.A(_20040_),
    .B(_20044_),
    .Y(_20045_));
 NOR2x1_ASAP7_75t_R _28561_ (.A(_20036_),
    .B(_20045_),
    .Y(_20046_));
 NAND2x1_ASAP7_75t_R _28562_ (.A(_20030_),
    .B(_20046_),
    .Y(_20047_));
 NOR2x1_ASAP7_75t_R _28563_ (.A(_20022_),
    .B(_20047_),
    .Y(_20048_));
 NAND2x2_ASAP7_75t_R _28564_ (.A(_20001_),
    .B(_20048_),
    .Y(_20049_));
 OAI21x1_ASAP7_75t_R _28565_ (.A1(_19960_),
    .A2(_19963_),
    .B(net2986),
    .Y(_20050_));
 INVx1_ASAP7_75t_R _28566_ (.A(_19953_),
    .Y(_20051_));
 NAND3x1_ASAP7_75t_R _28567_ (.A(_19957_),
    .B(_19940_),
    .C(_19943_),
    .Y(_20052_));
 NOR2x1_ASAP7_75t_R _28568_ (.A(_20051_),
    .B(_20052_),
    .Y(_20053_));
 INVx1_ASAP7_75t_R _28569_ (.A(_19936_),
    .Y(_20054_));
 NAND2x1_ASAP7_75t_R _28570_ (.A(_20053_),
    .B(_20054_),
    .Y(_20055_));
 NOR2x2_ASAP7_75t_R _28571_ (.A(_19907_),
    .B(_20055_),
    .Y(_20056_));
 NOR2x1_ASAP7_75t_R _28572_ (.A(_19962_),
    .B(_20056_),
    .Y(_20057_));
 INVx1_ASAP7_75t_R _28573_ (.A(_19773_),
    .Y(_20058_));
 NOR2x1_ASAP7_75t_R _28574_ (.A(_19785_),
    .B(_20058_),
    .Y(_20059_));
 NOR2x1_ASAP7_75t_R _28575_ (.A(_19799_),
    .B(_19812_),
    .Y(_20060_));
 NAND2x2_ASAP7_75t_R _28576_ (.A(_20059_),
    .B(_20060_),
    .Y(_20061_));
 INVx1_ASAP7_75t_R _28577_ (.A(_19859_),
    .Y(_20062_));
 NAND3x1_ASAP7_75t_R _28578_ (.A(_19862_),
    .B(net3180),
    .C(_19849_),
    .Y(_20063_));
 NOR2x1_ASAP7_75t_R _28579_ (.A(_20062_),
    .B(_20063_),
    .Y(_20064_));
 INVx1_ASAP7_75t_R _28580_ (.A(_19842_),
    .Y(_20065_));
 NAND2x1_ASAP7_75t_R _28581_ (.A(_20064_),
    .B(_20065_),
    .Y(_20066_));
 NOR2x2_ASAP7_75t_R _28582_ (.A(_20061_),
    .B(_20066_),
    .Y(_20067_));
 NOR2x1_ASAP7_75t_R _28583_ (.A(_19961_),
    .B(_20067_),
    .Y(_20068_));
 INVx1_ASAP7_75t_R _28584_ (.A(net2986),
    .Y(_20069_));
 OAI21x1_ASAP7_75t_R _28585_ (.A1(_20057_),
    .A2(_20068_),
    .B(_20069_),
    .Y(_20070_));
 NAND2x1_ASAP7_75t_R _28586_ (.A(_20050_),
    .B(_20070_),
    .Y(_20071_));
 OAI21x1_ASAP7_75t_R _28587_ (.A1(_19765_),
    .A2(_19766_),
    .B(_20071_),
    .Y(_20072_));
 NAND2x1_ASAP7_75t_R _28588_ (.A(_19961_),
    .B(_19962_),
    .Y(_20073_));
 NAND2x1_ASAP7_75t_R _28589_ (.A(_20056_),
    .B(_20067_),
    .Y(_20074_));
 AOI21x1_ASAP7_75t_R _28590_ (.A1(_20073_),
    .A2(_20074_),
    .B(_20069_),
    .Y(_20075_));
 NAND2x1_ASAP7_75t_R _28591_ (.A(_19962_),
    .B(_20056_),
    .Y(_20076_));
 NAND2x1_ASAP7_75t_R _28592_ (.A(_19961_),
    .B(_20067_),
    .Y(_20077_));
 AOI21x1_ASAP7_75t_R _28593_ (.A1(_20076_),
    .A2(_20077_),
    .B(net2987),
    .Y(_20078_));
 NOR2x1_ASAP7_75t_R _28594_ (.A(_20075_),
    .B(_20078_),
    .Y(_20079_));
 XOR2x1_ASAP7_75t_R _28595_ (.A(_19764_),
    .Y(_20080_),
    .B(_19688_));
 NAND2x1_ASAP7_75t_R _28596_ (.A(_20080_),
    .B(_20079_),
    .Y(_20081_));
 TAPCELL_ASAP7_75t_R TAP_824 ();
 AOI21x1_ASAP7_75t_R _28598_ (.A1(_20072_),
    .A2(_20081_),
    .B(net390),
    .Y(_20083_));
 INVx1_ASAP7_75t_R _28599_ (.A(_20083_),
    .Y(_20084_));
 AOI21x1_ASAP7_75t_R _28600_ (.A1(_19687_),
    .A2(_20084_),
    .B(net3533),
    .Y(_20085_));
 NOR3x1_ASAP7_75t_R _28601_ (.A(_20083_),
    .B(_14629_),
    .C(_19686_),
    .Y(_20086_));
 NOR2x1_ASAP7_75t_R _28602_ (.A(_20086_),
    .B(_20085_),
    .Y(_00124_));
 AND2x2_ASAP7_75t_R _28603_ (.A(net390),
    .B(_00911_),
    .Y(_20087_));
 XOR2x2_ASAP7_75t_R _28604_ (.A(_19961_),
    .B(_17905_),
    .Y(_20088_));
 AO21x1_ASAP7_75t_R _28605_ (.A1(net2407),
    .A2(net2438),
    .B(_18428_),
    .Y(_20089_));
 OAI21x1_ASAP7_75t_R _28606_ (.A1(net2051),
    .A2(_18428_),
    .B(_20089_),
    .Y(_20090_));
 OA211x2_ASAP7_75t_R _28607_ (.A1(net1087),
    .A2(_18237_),
    .B(_18434_),
    .C(net1864),
    .Y(_20091_));
 NOR2x1_ASAP7_75t_R _28608_ (.A(_20090_),
    .B(_20091_),
    .Y(_20092_));
 NOR2x1_ASAP7_75t_R _28609_ (.A(_19165_),
    .B(_18443_),
    .Y(_20093_));
 AO21x1_ASAP7_75t_R _28610_ (.A1(_18460_),
    .A2(_18335_),
    .B(net2989),
    .Y(_20094_));
 AO21x1_ASAP7_75t_R _28611_ (.A1(_18402_),
    .A2(_18327_),
    .B(net2989),
    .Y(_20095_));
 AND3x1_ASAP7_75t_R _28612_ (.A(_20093_),
    .B(_20094_),
    .C(_20095_),
    .Y(_20096_));
 NAND2x1_ASAP7_75t_R _28613_ (.A(_20092_),
    .B(_20096_),
    .Y(_20097_));
 AO21x1_ASAP7_75t_R _28614_ (.A1(_18402_),
    .A2(_18242_),
    .B(_18248_),
    .Y(_20098_));
 NAND2x1_ASAP7_75t_R _28615_ (.A(_18247_),
    .B(_18291_),
    .Y(_20099_));
 AND3x2_ASAP7_75t_R _28616_ (.A(_20098_),
    .B(_18271_),
    .C(_20099_),
    .Y(_20100_));
 AO21x1_ASAP7_75t_R _28617_ (.A1(net937),
    .A2(net3247),
    .B(_18266_),
    .Y(_20101_));
 NAND2x1_ASAP7_75t_R _28618_ (.A(_18482_),
    .B(_18416_),
    .Y(_20102_));
 AND2x2_ASAP7_75t_R _28619_ (.A(_20101_),
    .B(_20102_),
    .Y(_20103_));
 AO21x1_ASAP7_75t_R _28620_ (.A1(net2747),
    .A2(net2407),
    .B(_18266_),
    .Y(_20104_));
 OA21x2_ASAP7_75t_R _28621_ (.A1(net2051),
    .A2(_18266_),
    .B(_20104_),
    .Y(_20105_));
 NAND3x2_ASAP7_75t_R _28622_ (.B(_20103_),
    .C(_20105_),
    .Y(_20106_),
    .A(_20100_));
 NOR2x2_ASAP7_75t_R _28623_ (.A(_20097_),
    .B(_20106_),
    .Y(_20107_));
 INVx1_ASAP7_75t_R _28624_ (.A(_20107_),
    .Y(_20108_));
 AOI211x1_ASAP7_75t_R _28625_ (.A1(net2999),
    .A2(_18237_),
    .B(net3282),
    .C(net2974),
    .Y(_20109_));
 OA21x2_ASAP7_75t_R _28626_ (.A1(_18259_),
    .A2(_18468_),
    .B(_18483_),
    .Y(_20110_));
 NOR2x2_ASAP7_75t_R _28627_ (.A(_20109_),
    .B(_20110_),
    .Y(_20111_));
 NAND2x2_ASAP7_75t_R _28628_ (.A(_18445_),
    .B(_18483_),
    .Y(_20112_));
 AO21x1_ASAP7_75t_R _28629_ (.A1(_18381_),
    .A2(net2638),
    .B(net3282),
    .Y(_20113_));
 NAND3x2_ASAP7_75t_R _28630_ (.B(net3286),
    .C(_20113_),
    .Y(_20114_),
    .A(_20111_));
 AO21x2_ASAP7_75t_R _28631_ (.A1(_19171_),
    .A2(_18351_),
    .B(_18490_),
    .Y(_20115_));
 OA21x2_ASAP7_75t_R _28632_ (.A1(net2974),
    .A2(net2595),
    .B(_20115_),
    .Y(_20116_));
 AO21x1_ASAP7_75t_R _28633_ (.A1(net1753),
    .A2(net1483),
    .B(net2994),
    .Y(_20117_));
 NAND2x1_ASAP7_75t_R _28634_ (.A(_18344_),
    .B(_19472_),
    .Y(_20118_));
 NAND2x1_ASAP7_75t_R _28635_ (.A(_18485_),
    .B(_19472_),
    .Y(_20119_));
 AND3x1_ASAP7_75t_R _28636_ (.A(_20117_),
    .B(_20118_),
    .C(_20119_),
    .Y(_20120_));
 NAND2x1_ASAP7_75t_R _28637_ (.A(_20116_),
    .B(_20120_),
    .Y(_20121_));
 NOR2x2_ASAP7_75t_R _28638_ (.A(_20114_),
    .B(_20121_),
    .Y(_20122_));
 AO21x1_ASAP7_75t_R _28639_ (.A1(net2251),
    .A2(net2965),
    .B(_18456_),
    .Y(_20123_));
 NAND2x1_ASAP7_75t_R _28640_ (.A(_18482_),
    .B(_19185_),
    .Y(_20124_));
 AND3x2_ASAP7_75t_R _28641_ (.A(_20123_),
    .B(_19186_),
    .C(_20124_),
    .Y(_20125_));
 NAND2x1_ASAP7_75t_R _28642_ (.A(_19150_),
    .B(_18469_),
    .Y(_20126_));
 NAND2x1_ASAP7_75t_R _28643_ (.A(_18444_),
    .B(_18469_),
    .Y(_20127_));
 AND3x2_ASAP7_75t_R _28644_ (.A(_18473_),
    .B(_20126_),
    .C(_20127_),
    .Y(_20128_));
 AO21x1_ASAP7_75t_R _28645_ (.A1(_18350_),
    .A2(net1254),
    .B(net3312),
    .Y(_20129_));
 NAND3x2_ASAP7_75t_R _28646_ (.B(_20128_),
    .C(_20129_),
    .Y(_20130_),
    .A(_20125_));
 INVx1_ASAP7_75t_R _28647_ (.A(_20130_),
    .Y(_20131_));
 NAND2x1_ASAP7_75t_R _28648_ (.A(_20122_),
    .B(_20131_),
    .Y(_20132_));
 NOR2x2_ASAP7_75t_R _28649_ (.A(_20108_),
    .B(_20132_),
    .Y(_20133_));
 AO21x1_ASAP7_75t_R _28650_ (.A1(_18350_),
    .A2(net2788),
    .B(_18318_),
    .Y(_20134_));
 AO21x1_ASAP7_75t_R _28651_ (.A1(net1335),
    .A2(net2638),
    .B(_18318_),
    .Y(_20135_));
 AND2x2_ASAP7_75t_R _28652_ (.A(_20134_),
    .B(_20135_),
    .Y(_20136_));
 NAND2x1_ASAP7_75t_R _28653_ (.A(net1702),
    .B(_18345_),
    .Y(_20137_));
 AND3x1_ASAP7_75t_R _28654_ (.A(_18337_),
    .B(_20137_),
    .C(_19206_),
    .Y(_20138_));
 NAND2x1_ASAP7_75t_R _28655_ (.A(_20136_),
    .B(_20138_),
    .Y(_20139_));
 AO21x1_ASAP7_75t_R _28656_ (.A1(net2043),
    .A2(net2945),
    .B(net2985),
    .Y(_20140_));
 NAND3x1_ASAP7_75t_R _28657_ (.A(_20140_),
    .B(_18289_),
    .C(_20032_),
    .Y(_20141_));
 AO21x1_ASAP7_75t_R _28658_ (.A1(net2043),
    .A2(net2634),
    .B(net2970),
    .Y(_20142_));
 AO21x1_ASAP7_75t_R _28659_ (.A1(net2473),
    .A2(net2250),
    .B(net2970),
    .Y(_20143_));
 NAND3x1_ASAP7_75t_R _28660_ (.A(_20142_),
    .B(_20143_),
    .C(_20039_),
    .Y(_20144_));
 NOR2x1_ASAP7_75t_R _28661_ (.A(_20141_),
    .B(_20144_),
    .Y(_20145_));
 INVx1_ASAP7_75t_R _28662_ (.A(_20145_),
    .Y(_20146_));
 NOR2x2_ASAP7_75t_R _28663_ (.A(_20139_),
    .B(_20146_),
    .Y(_20147_));
 INVx1_ASAP7_75t_R _28664_ (.A(_20147_),
    .Y(_20148_));
 AO21x1_ASAP7_75t_R _28665_ (.A1(net1753),
    .A2(net2965),
    .B(_18364_),
    .Y(_20149_));
 NAND2x1_ASAP7_75t_R _28666_ (.A(_18371_),
    .B(_19150_),
    .Y(_20150_));
 AND3x1_ASAP7_75t_R _28667_ (.A(_20149_),
    .B(_19548_),
    .C(_20150_),
    .Y(_20151_));
 AO21x1_ASAP7_75t_R _28668_ (.A1(net2045),
    .A2(_18442_),
    .B(_18354_),
    .Y(_20152_));
 NOR2x1_ASAP7_75t_R _28669_ (.A(_18354_),
    .B(net1753),
    .Y(_20153_));
 INVx1_ASAP7_75t_R _28670_ (.A(_20153_),
    .Y(_20154_));
 AND2x2_ASAP7_75t_R _28671_ (.A(_20152_),
    .B(_20154_),
    .Y(_20155_));
 INVx1_ASAP7_75t_R _28672_ (.A(_18335_),
    .Y(_20156_));
 OA21x2_ASAP7_75t_R _28673_ (.A1(net1702),
    .A2(net2849),
    .B(_19237_),
    .Y(_20157_));
 AOI21x1_ASAP7_75t_R _28674_ (.A1(_20156_),
    .A2(_19237_),
    .B(_20157_),
    .Y(_20158_));
 AND3x2_ASAP7_75t_R _28675_ (.A(_20151_),
    .B(_20155_),
    .C(_20158_),
    .Y(_20159_));
 AO21x1_ASAP7_75t_R _28676_ (.A1(net2045),
    .A2(net2638),
    .B(_18377_),
    .Y(_20160_));
 AO21x1_ASAP7_75t_R _28677_ (.A1(net2634),
    .A2(net1483),
    .B(_18377_),
    .Y(_20161_));
 NAND2x1_ASAP7_75t_R _28678_ (.A(net2669),
    .B(_19224_),
    .Y(_20162_));
 AND3x1_ASAP7_75t_R _28679_ (.A(_20160_),
    .B(_20161_),
    .C(_20162_),
    .Y(_20163_));
 AO21x1_ASAP7_75t_R _28680_ (.A1(net2176),
    .A2(_18366_),
    .B(_18395_),
    .Y(_20164_));
 AND2x2_ASAP7_75t_R _28681_ (.A(_20164_),
    .B(_18399_),
    .Y(_20165_));
 OA21x2_ASAP7_75t_R _28682_ (.A1(net2096),
    .A2(net2981),
    .B(_18388_),
    .Y(_20166_));
 AND3x2_ASAP7_75t_R _28683_ (.A(_20163_),
    .B(_20165_),
    .C(_20166_),
    .Y(_20167_));
 NAND2x1_ASAP7_75t_R _28684_ (.A(_20159_),
    .B(_20167_),
    .Y(_20168_));
 NOR2x2_ASAP7_75t_R _28685_ (.A(_20148_),
    .B(_20168_),
    .Y(_20169_));
 NAND2x2_ASAP7_75t_R _28686_ (.A(_20133_),
    .B(_20169_),
    .Y(_20170_));
 XOR2x1_ASAP7_75t_R _28687_ (.A(_20088_),
    .Y(_20171_),
    .B(net2537));
 AO21x1_ASAP7_75t_R _28688_ (.A1(_18584_),
    .A2(net2405),
    .B(_18641_),
    .Y(_20172_));
 AO21x1_ASAP7_75t_R _28689_ (.A1(net3378),
    .A2(net2760),
    .B(net2620),
    .Y(_20173_));
 AO21x1_ASAP7_75t_R _28690_ (.A1(net2028),
    .A2(_18623_),
    .B(net2620),
    .Y(_20174_));
 AO21x1_ASAP7_75t_R _28691_ (.A1(net1388),
    .A2(_18548_),
    .B(net2620),
    .Y(_20175_));
 AND3x1_ASAP7_75t_R _28692_ (.A(_20173_),
    .B(_20174_),
    .C(_20175_),
    .Y(_20176_));
 NAND2x1_ASAP7_75t_R _28693_ (.A(_20172_),
    .B(_20176_),
    .Y(_20177_));
 AO21x1_ASAP7_75t_R _28694_ (.A1(net3378),
    .A2(net1388),
    .B(_18625_),
    .Y(_20178_));
 OA21x2_ASAP7_75t_R _28695_ (.A1(net2177),
    .A2(_18625_),
    .B(_20178_),
    .Y(_20179_));
 NAND2x1_ASAP7_75t_R _28696_ (.A(_18690_),
    .B(_19058_),
    .Y(_20180_));
 AND4x1_ASAP7_75t_R _28697_ (.A(_19635_),
    .B(_19637_),
    .C(_20180_),
    .D(_19062_),
    .Y(_20181_));
 NAND2x1_ASAP7_75t_R _28698_ (.A(_20179_),
    .B(_20181_),
    .Y(_20182_));
 NOR2x2_ASAP7_75t_R _28699_ (.A(_20177_),
    .B(_20182_),
    .Y(_20183_));
 TAPCELL_ASAP7_75t_R TAP_823 ();
 AO21x1_ASAP7_75t_R _28701_ (.A1(_18516_),
    .A2(net1965),
    .B(_18588_),
    .Y(_20185_));
 OA21x2_ASAP7_75t_R _28702_ (.A1(_18528_),
    .A2(_18588_),
    .B(_20185_),
    .Y(_20186_));
 AO21x1_ASAP7_75t_R _28703_ (.A1(net3215),
    .A2(net1965),
    .B(_18569_),
    .Y(_20187_));
 NAND2x2_ASAP7_75t_R _28704_ (.A(net2735),
    .B(_18570_),
    .Y(_20188_));
 AND3x1_ASAP7_75t_R _28705_ (.A(_20187_),
    .B(_20188_),
    .C(_18573_),
    .Y(_20189_));
 NAND2x1_ASAP7_75t_R _28706_ (.A(_20186_),
    .B(_20189_),
    .Y(_20190_));
 OA31x2_ASAP7_75t_R _28707_ (.A1(_18585_),
    .A2(_18636_),
    .A3(_18638_),
    .B1(net2690),
    .Y(_20191_));
 NOR2x2_ASAP7_75t_R _28708_ (.A(net1069),
    .B(_18536_),
    .Y(_20192_));
 OA31x2_ASAP7_75t_R _28709_ (.A1(_18675_),
    .A2(_20192_),
    .A3(_18537_),
    .B1(net2690),
    .Y(_20193_));
 NOR2x1_ASAP7_75t_R _28710_ (.A(_20191_),
    .B(_20193_),
    .Y(_20194_));
 AO21x1_ASAP7_75t_R _28711_ (.A1(_18975_),
    .A2(_18702_),
    .B(_18545_),
    .Y(_20195_));
 NAND2x1_ASAP7_75t_R _28712_ (.A(_20192_),
    .B(_19664_),
    .Y(_20196_));
 AND3x1_ASAP7_75t_R _28713_ (.A(_19075_),
    .B(_20195_),
    .C(_20196_),
    .Y(_20197_));
 NAND2x1_ASAP7_75t_R _28714_ (.A(_20194_),
    .B(_20197_),
    .Y(_20198_));
 NOR2x2_ASAP7_75t_R _28715_ (.A(_20190_),
    .B(_20198_),
    .Y(_20199_));
 AO21x1_ASAP7_75t_R _28716_ (.A1(_19073_),
    .A2(net2142),
    .B(net2414),
    .Y(_20200_));
 OA21x2_ASAP7_75t_R _28717_ (.A1(net1307),
    .A2(net2414),
    .B(_20200_),
    .Y(_20201_));
 AO21x1_ASAP7_75t_R _28718_ (.A1(net1404),
    .A2(net3215),
    .B(net2414),
    .Y(_20202_));
 OA21x2_ASAP7_75t_R _28719_ (.A1(net2405),
    .A2(net2414),
    .B(_20202_),
    .Y(_20203_));
 NAND2x1_ASAP7_75t_R _28720_ (.A(_20201_),
    .B(_20203_),
    .Y(_20204_));
 AOI22x1_ASAP7_75t_R _28721_ (.A1(_19647_),
    .A2(net1010),
    .B1(_18638_),
    .B2(_19046_),
    .Y(_20205_));
 OR3x4_ASAP7_75t_R _28722_ (.A(_18604_),
    .B(net1736),
    .C(net1566),
    .Y(_20206_));
 AO21x1_ASAP7_75t_R _28723_ (.A1(net1307),
    .A2(_18601_),
    .B(net2578),
    .Y(_20207_));
 NAND3x2_ASAP7_75t_R _28724_ (.B(_20206_),
    .C(_20207_),
    .Y(_20208_),
    .A(_20205_));
 NOR2x2_ASAP7_75t_R _28725_ (.A(_20204_),
    .B(_20208_),
    .Y(_20209_));
 NAND3x2_ASAP7_75t_R _28726_ (.B(_20199_),
    .C(_20209_),
    .Y(_20210_),
    .A(_20183_));
 AO21x1_ASAP7_75t_R _28727_ (.A1(_18516_),
    .A2(_19036_),
    .B(net2317),
    .Y(_20211_));
 AO21x1_ASAP7_75t_R _28728_ (.A1(net1307),
    .A2(net2386),
    .B(net2317),
    .Y(_20212_));
 NAND2x2_ASAP7_75t_R _28729_ (.A(_18590_),
    .B(_18725_),
    .Y(_20213_));
 NAND3x2_ASAP7_75t_R _28730_ (.B(_20212_),
    .C(_20213_),
    .Y(_20214_),
    .A(_20211_));
 AO21x1_ASAP7_75t_R _28731_ (.A1(net3215),
    .A2(_18518_),
    .B(net2694),
    .Y(_20215_));
 NAND2x2_ASAP7_75t_R _28732_ (.A(_19758_),
    .B(_20215_),
    .Y(_20216_));
 AO21x1_ASAP7_75t_R _28733_ (.A1(_19729_),
    .A2(_18536_),
    .B(net2693),
    .Y(_20217_));
 INVx1_ASAP7_75t_R _28734_ (.A(_20217_),
    .Y(_20218_));
 NOR3x2_ASAP7_75t_R _28735_ (.B(_20216_),
    .C(_20218_),
    .Y(_20219_),
    .A(_20214_));
 INVx1_ASAP7_75t_R _28736_ (.A(_20219_),
    .Y(_20220_));
 AO21x1_ASAP7_75t_R _28737_ (.A1(net3376),
    .A2(net3381),
    .B(net3324),
    .Y(_20221_));
 AO21x1_ASAP7_75t_R _28738_ (.A1(net1823),
    .A2(_18518_),
    .B(net3324),
    .Y(_20222_));
 AO21x1_ASAP7_75t_R _28739_ (.A1(net2504),
    .A2(_18548_),
    .B(net3324),
    .Y(_20223_));
 AND3x2_ASAP7_75t_R _28740_ (.A(_20221_),
    .B(_20222_),
    .C(_20223_),
    .Y(_20224_));
 AO21x1_ASAP7_75t_R _28741_ (.A1(_19073_),
    .A2(_18992_),
    .B(net2394),
    .Y(_20225_));
 AO21x1_ASAP7_75t_R _28742_ (.A1(net1388),
    .A2(_18548_),
    .B(_18714_),
    .Y(_20226_));
 NOR2x1_ASAP7_75t_R _28743_ (.A(net2398),
    .B(_18714_),
    .Y(_20227_));
 INVx1_ASAP7_75t_R _28744_ (.A(_20227_),
    .Y(_20228_));
 AND3x2_ASAP7_75t_R _28745_ (.A(_20225_),
    .B(_20226_),
    .C(_20228_),
    .Y(_20229_));
 AOI211x1_ASAP7_75t_R _28746_ (.A1(net1470),
    .A2(_18554_),
    .B(net2394),
    .C(net2631),
    .Y(_20230_));
 NOR2x1_ASAP7_75t_R _28747_ (.A(_18714_),
    .B(net2405),
    .Y(_20231_));
 AOI211x1_ASAP7_75t_R _28748_ (.A1(_19057_),
    .A2(_19580_),
    .B(_20230_),
    .C(_20231_),
    .Y(_20232_));
 NAND3x2_ASAP7_75t_R _28749_ (.B(_20229_),
    .C(_20232_),
    .Y(_20233_),
    .A(_20224_));
 NOR2x1_ASAP7_75t_R _28750_ (.A(_20220_),
    .B(_20233_),
    .Y(_20234_));
 AO21x1_ASAP7_75t_R _28751_ (.A1(net2067),
    .A2(_18702_),
    .B(net2413),
    .Y(_20235_));
 NAND2x1_ASAP7_75t_R _28752_ (.A(_19057_),
    .B(_18683_),
    .Y(_20236_));
 AND3x1_ASAP7_75t_R _28753_ (.A(_20235_),
    .B(_20236_),
    .C(_18691_),
    .Y(_20237_));
 AO21x1_ASAP7_75t_R _28754_ (.A1(net2028),
    .A2(_18992_),
    .B(net2413),
    .Y(_20238_));
 AO21x1_ASAP7_75t_R _28755_ (.A1(net1388),
    .A2(_18548_),
    .B(net2413),
    .Y(_20239_));
 NAND2x1_ASAP7_75t_R _28756_ (.A(_20192_),
    .B(_18683_),
    .Y(_20240_));
 AND3x1_ASAP7_75t_R _28757_ (.A(_20238_),
    .B(_20239_),
    .C(_20240_),
    .Y(_20241_));
 NAND2x1_ASAP7_75t_R _28758_ (.A(_18537_),
    .B(_18696_),
    .Y(_20242_));
 AO21x1_ASAP7_75t_R _28759_ (.A1(_18600_),
    .A2(_18623_),
    .B(_18695_),
    .Y(_20243_));
 NAND2x1_ASAP7_75t_R _28760_ (.A(_20242_),
    .B(_20243_),
    .Y(_20244_));
 AO21x1_ASAP7_75t_R _28761_ (.A1(_18516_),
    .A2(net1966),
    .B(net2292),
    .Y(_20245_));
 AO21x1_ASAP7_75t_R _28762_ (.A1(_18651_),
    .A2(_19013_),
    .B(_18695_),
    .Y(_20246_));
 NAND2x1_ASAP7_75t_R _28763_ (.A(_20245_),
    .B(_20246_),
    .Y(_20247_));
 NOR2x1_ASAP7_75t_R _28764_ (.A(_20244_),
    .B(_20247_),
    .Y(_20248_));
 NAND3x1_ASAP7_75t_R _28765_ (.A(_20237_),
    .B(_20241_),
    .C(_20248_),
    .Y(_20249_));
 OAI21x1_ASAP7_75t_R _28766_ (.A1(_18650_),
    .A2(_19057_),
    .B(_19031_),
    .Y(_20250_));
 NAND2x1_ASAP7_75t_R _28767_ (.A(_19614_),
    .B(_19031_),
    .Y(_20251_));
 NAND2x1_ASAP7_75t_R _28768_ (.A(_19060_),
    .B(_19031_),
    .Y(_20252_));
 AND3x1_ASAP7_75t_R _28769_ (.A(_20250_),
    .B(_20251_),
    .C(_20252_),
    .Y(_20253_));
 NAND2x1_ASAP7_75t_R _28770_ (.A(net1750),
    .B(_19031_),
    .Y(_20254_));
 AND3x1_ASAP7_75t_R _28771_ (.A(_18659_),
    .B(_19611_),
    .C(_20254_),
    .Y(_20255_));
 NAND2x1_ASAP7_75t_R _28772_ (.A(_20253_),
    .B(_20255_),
    .Y(_20256_));
 INVx1_ASAP7_75t_R _28773_ (.A(_18601_),
    .Y(_20257_));
 NAND2x1_ASAP7_75t_R _28774_ (.A(_20257_),
    .B(_18671_),
    .Y(_20258_));
 NAND2x1_ASAP7_75t_R _28775_ (.A(_20258_),
    .B(_18676_),
    .Y(_20259_));
 INVx1_ASAP7_75t_R _28776_ (.A(_19738_),
    .Y(_20260_));
 OA21x2_ASAP7_75t_R _28777_ (.A1(_19083_),
    .A2(_19060_),
    .B(_18671_),
    .Y(_20261_));
 OR3x2_ASAP7_75t_R _28778_ (.A(_20259_),
    .B(_20260_),
    .C(_20261_),
    .Y(_20262_));
 NOR2x2_ASAP7_75t_R _28779_ (.A(_20256_),
    .B(_20262_),
    .Y(_20263_));
 INVx1_ASAP7_75t_R _28780_ (.A(_20263_),
    .Y(_20264_));
 NOR2x1_ASAP7_75t_R _28781_ (.A(_20249_),
    .B(_20264_),
    .Y(_20265_));
 NAND2x2_ASAP7_75t_R _28782_ (.A(_20234_),
    .B(_20265_),
    .Y(_20266_));
 NOR2x2_ASAP7_75t_R _28783_ (.A(_20210_),
    .B(_20266_),
    .Y(_20267_));
 NOR2x2_ASAP7_75t_R _28784_ (.A(_20267_),
    .B(_18742_),
    .Y(_20268_));
 AND3x1_ASAP7_75t_R _28785_ (.A(_20237_),
    .B(_20241_),
    .C(_20248_),
    .Y(_20269_));
 NAND2x1_ASAP7_75t_R _28786_ (.A(_20263_),
    .B(_20269_),
    .Y(_20270_));
 INVx1_ASAP7_75t_R _28787_ (.A(_20233_),
    .Y(_20271_));
 NAND2x1_ASAP7_75t_R _28788_ (.A(_20219_),
    .B(_20271_),
    .Y(_20272_));
 NOR2x2_ASAP7_75t_R _28789_ (.A(_20270_),
    .B(_20272_),
    .Y(_20273_));
 INVx1_ASAP7_75t_R _28790_ (.A(_20210_),
    .Y(_20274_));
 NAND2x2_ASAP7_75t_R _28791_ (.A(_20273_),
    .B(_20274_),
    .Y(_20275_));
 NOR2x2_ASAP7_75t_R _28792_ (.A(_19143_),
    .B(_20275_),
    .Y(_20276_));
 NOR2x2_ASAP7_75t_R _28793_ (.A(_20268_),
    .B(_20276_),
    .Y(_20277_));
 AO21x1_ASAP7_75t_R _28794_ (.A1(net1081),
    .A2(_17538_),
    .B(_17777_),
    .Y(_20278_));
 AND2x2_ASAP7_75t_R _28795_ (.A(_19896_),
    .B(_20278_),
    .Y(_20279_));
 NAND2x1_ASAP7_75t_R _28796_ (.A(_18788_),
    .B(_17782_),
    .Y(_20280_));
 AO21x1_ASAP7_75t_R _28797_ (.A1(_17626_),
    .A2(net2899),
    .B(_17777_),
    .Y(_20281_));
 NAND3x1_ASAP7_75t_R _28798_ (.A(_20279_),
    .B(_20280_),
    .C(_20281_),
    .Y(_20282_));
 OA21x2_ASAP7_75t_R _28799_ (.A1(_17575_),
    .A2(net2909),
    .B(_17835_),
    .Y(_20283_));
 OA21x2_ASAP7_75t_R _28800_ (.A1(_18788_),
    .A2(_17774_),
    .B(_17771_),
    .Y(_20284_));
 NOR2x1_ASAP7_75t_R _28801_ (.A(_17770_),
    .B(_17626_),
    .Y(_20285_));
 AOI211x1_ASAP7_75t_R _28802_ (.A1(_17771_),
    .A2(_17786_),
    .B(_20284_),
    .C(_20285_),
    .Y(_20286_));
 NAND2x1_ASAP7_75t_R _28803_ (.A(_20283_),
    .B(_20286_),
    .Y(_20287_));
 NOR2x1_ASAP7_75t_R _28804_ (.A(_20282_),
    .B(_20287_),
    .Y(_20288_));
 OA21x2_ASAP7_75t_R _28805_ (.A1(_18788_),
    .A2(_17558_),
    .B(_18825_),
    .Y(_20289_));
 NOR2x1_ASAP7_75t_R _28806_ (.A(net2902),
    .B(_17759_),
    .Y(_20290_));
 NOR2x1_ASAP7_75t_R _28807_ (.A(net2901),
    .B(_17759_),
    .Y(_20291_));
 OR3x1_ASAP7_75t_R _28808_ (.A(_20289_),
    .B(_20290_),
    .C(_20291_),
    .Y(_20292_));
 OA21x2_ASAP7_75t_R _28809_ (.A1(_17679_),
    .A2(_17731_),
    .B(_19890_),
    .Y(_20293_));
 NOR2x1_ASAP7_75t_R _28810_ (.A(_17744_),
    .B(net2600),
    .Y(_20294_));
 NOR2x1_ASAP7_75t_R _28811_ (.A(_17758_),
    .B(_17744_),
    .Y(_20295_));
 OR4x1_ASAP7_75t_R _28812_ (.A(_20293_),
    .B(_20294_),
    .C(_17749_),
    .D(_20295_),
    .Y(_20296_));
 NOR2x1_ASAP7_75t_R _28813_ (.A(_20292_),
    .B(_20296_),
    .Y(_20297_));
 NAND2x1_ASAP7_75t_R _28814_ (.A(_20288_),
    .B(_20297_),
    .Y(_20298_));
 AO21x1_ASAP7_75t_R _28815_ (.A1(net2893),
    .A2(_17892_),
    .B(_17691_),
    .Y(_20299_));
 AO21x1_ASAP7_75t_R _28816_ (.A1(_17562_),
    .A2(net1380),
    .B(_17691_),
    .Y(_20300_));
 NAND2x1_ASAP7_75t_R _28817_ (.A(_17801_),
    .B(_17788_),
    .Y(_20301_));
 AND3x1_ASAP7_75t_R _28818_ (.A(_20299_),
    .B(_20300_),
    .C(_20301_),
    .Y(_20302_));
 OA21x2_ASAP7_75t_R _28819_ (.A1(_17701_),
    .A2(_17756_),
    .B(_17912_),
    .Y(_20303_));
 AO21x1_ASAP7_75t_R _28820_ (.A1(_17639_),
    .A2(_19294_),
    .B(_17701_),
    .Y(_20304_));
 AND3x1_ASAP7_75t_R _28821_ (.A(_20302_),
    .B(_20303_),
    .C(_20304_),
    .Y(_20305_));
 AO21x1_ASAP7_75t_R _28822_ (.A1(net2598),
    .A2(_17756_),
    .B(net2882),
    .Y(_20306_));
 AO21x1_ASAP7_75t_R _28823_ (.A1(net2532),
    .A2(_17586_),
    .B(net2882),
    .Y(_20307_));
 NAND2x1_ASAP7_75t_R _28824_ (.A(_17774_),
    .B(_17714_),
    .Y(_20308_));
 AND3x1_ASAP7_75t_R _28825_ (.A(_20306_),
    .B(_20307_),
    .C(_20308_),
    .Y(_20309_));
 NAND2x1_ASAP7_75t_R _28826_ (.A(_18839_),
    .B(_17729_),
    .Y(_20310_));
 INVx1_ASAP7_75t_R _28827_ (.A(_20310_),
    .Y(_20311_));
 AO21x1_ASAP7_75t_R _28828_ (.A1(_17639_),
    .A2(net2892),
    .B(_17725_),
    .Y(_20312_));
 OA21x2_ASAP7_75t_R _28829_ (.A1(_17575_),
    .A2(_17725_),
    .B(_20312_),
    .Y(_20313_));
 AND3x1_ASAP7_75t_R _28830_ (.A(_20309_),
    .B(_20311_),
    .C(_20313_),
    .Y(_20314_));
 NAND2x1_ASAP7_75t_R _28831_ (.A(_20305_),
    .B(_20314_),
    .Y(_20315_));
 NOR2x1_ASAP7_75t_R _28832_ (.A(_20298_),
    .B(_20315_),
    .Y(_20316_));
 AO21x1_ASAP7_75t_R _28833_ (.A1(net936),
    .A2(_17756_),
    .B(net2847),
    .Y(_20317_));
 OA21x2_ASAP7_75t_R _28834_ (.A1(_17758_),
    .A2(net2847),
    .B(_20317_),
    .Y(_20318_));
 NAND2x1_ASAP7_75t_R _28835_ (.A(_19347_),
    .B(_20318_),
    .Y(_20319_));
 NOR2x2_ASAP7_75t_R _28836_ (.A(_17670_),
    .B(net997),
    .Y(_20320_));
 OA21x2_ASAP7_75t_R _28837_ (.A1(_17757_),
    .A2(_17609_),
    .B(_17671_),
    .Y(_20321_));
 NOR2x1_ASAP7_75t_R _28838_ (.A(_20320_),
    .B(_20321_),
    .Y(_20322_));
 NAND2x1_ASAP7_75t_R _28839_ (.A(net2906),
    .B(_17671_),
    .Y(_20323_));
 NAND2x1_ASAP7_75t_R _28840_ (.A(_20323_),
    .B(_17674_),
    .Y(_20324_));
 AOI21x1_ASAP7_75t_R _28841_ (.A1(_17886_),
    .A2(_17671_),
    .B(_20324_),
    .Y(_20325_));
 NAND2x1_ASAP7_75t_R _28842_ (.A(_20322_),
    .B(_20325_),
    .Y(_20326_));
 NOR2x1_ASAP7_75t_R _28843_ (.A(_20319_),
    .B(_20326_),
    .Y(_20327_));
 OA21x2_ASAP7_75t_R _28844_ (.A1(_17676_),
    .A2(_17774_),
    .B(_18789_),
    .Y(_20328_));
 AOI211x1_ASAP7_75t_R _28845_ (.A1(net1123),
    .A2(net1187),
    .B(net1103),
    .C(_17629_),
    .Y(_20329_));
 AOI21x1_ASAP7_75t_R _28846_ (.A1(_17632_),
    .A2(_17834_),
    .B(_17629_),
    .Y(_20330_));
 OR3x1_ASAP7_75t_R _28847_ (.A(_20328_),
    .B(_20329_),
    .C(_20330_),
    .Y(_20331_));
 AO21x1_ASAP7_75t_R _28848_ (.A1(_17813_),
    .A2(_17582_),
    .B(_17641_),
    .Y(_20332_));
 INVx1_ASAP7_75t_R _28849_ (.A(_19923_),
    .Y(_20333_));
 AND3x1_ASAP7_75t_R _28850_ (.A(_20332_),
    .B(_18784_),
    .C(_20333_),
    .Y(_20334_));
 OAI21x1_ASAP7_75t_R _28851_ (.A1(_17756_),
    .A2(net2484),
    .B(_20334_),
    .Y(_20335_));
 NOR2x1_ASAP7_75t_R _28852_ (.A(_20331_),
    .B(_20335_),
    .Y(_20336_));
 NAND2x1_ASAP7_75t_R _28853_ (.A(_20327_),
    .B(_20336_),
    .Y(_20337_));
 OA21x2_ASAP7_75t_R _28854_ (.A1(net2906),
    .A2(_17673_),
    .B(_17569_),
    .Y(_20338_));
 AOI21x1_ASAP7_75t_R _28855_ (.A1(_17678_),
    .A2(_17569_),
    .B(_20338_),
    .Y(_20339_));
 AND2x2_ASAP7_75t_R _28856_ (.A(_17549_),
    .B(_17554_),
    .Y(_20340_));
 AO21x1_ASAP7_75t_R _28857_ (.A1(net1089),
    .A2(_17608_),
    .B(net1103),
    .Y(_20341_));
 AO21x1_ASAP7_75t_R _28858_ (.A1(_20341_),
    .A2(net941),
    .B(_17547_),
    .Y(_20342_));
 AO21x1_ASAP7_75t_R _28859_ (.A1(net2202),
    .A2(net2451),
    .B(_17566_),
    .Y(_20343_));
 AND4x1_ASAP7_75t_R _28860_ (.A(_20339_),
    .B(_20340_),
    .C(_20342_),
    .D(_20343_),
    .Y(_20344_));
 AO21x1_ASAP7_75t_R _28861_ (.A1(net936),
    .A2(net2901),
    .B(_17614_),
    .Y(_20345_));
 AO21x1_ASAP7_75t_R _28862_ (.A1(net1788),
    .A2(net1082),
    .B(_17614_),
    .Y(_20346_));
 OA211x2_ASAP7_75t_R _28863_ (.A1(net1832),
    .A2(_19950_),
    .B(_20345_),
    .C(_20346_),
    .Y(_20347_));
 AND3x1_ASAP7_75t_R _28864_ (.A(_18779_),
    .B(_19947_),
    .C(_17591_),
    .Y(_20348_));
 AND2x2_ASAP7_75t_R _28865_ (.A(_20347_),
    .B(_20348_),
    .Y(_20349_));
 NAND2x1_ASAP7_75t_R _28866_ (.A(_20344_),
    .B(_20349_),
    .Y(_20350_));
 NOR2x1_ASAP7_75t_R _28867_ (.A(_20337_),
    .B(_20350_),
    .Y(_20351_));
 NAND2x2_ASAP7_75t_R _28868_ (.A(_20316_),
    .B(_20351_),
    .Y(_20352_));
 AO21x1_ASAP7_75t_R _28869_ (.A1(net939),
    .A2(_18081_),
    .B(net3123),
    .Y(_20353_));
 AO21x1_ASAP7_75t_R _28870_ (.A1(_18881_),
    .A2(_18022_),
    .B(net3123),
    .Y(_20354_));
 AO21x1_ASAP7_75t_R _28871_ (.A1(net1068),
    .A2(_18002_),
    .B(net3123),
    .Y(_20355_));
 AND3x1_ASAP7_75t_R _28872_ (.A(_20353_),
    .B(_20354_),
    .C(_20355_),
    .Y(_20356_));
 OA21x2_ASAP7_75t_R _28873_ (.A1(_18021_),
    .A2(_17937_),
    .B(_19852_),
    .Y(_20357_));
 AND2x2_ASAP7_75t_R _28874_ (.A(_18921_),
    .B(_20357_),
    .Y(_20358_));
 NAND2x1_ASAP7_75t_R _28875_ (.A(_20356_),
    .B(_20358_),
    .Y(_20359_));
 AO21x1_ASAP7_75t_R _28876_ (.A1(_18010_),
    .A2(net3184),
    .B(net3205),
    .Y(_20360_));
 AO21x1_ASAP7_75t_R _28877_ (.A1(_18881_),
    .A2(net1690),
    .B(net3205),
    .Y(_20361_));
 NAND2x1_ASAP7_75t_R _28878_ (.A(net2792),
    .B(_19376_),
    .Y(_20362_));
 AND3x1_ASAP7_75t_R _28879_ (.A(_20360_),
    .B(_20361_),
    .C(_20362_),
    .Y(_20363_));
 NAND2x1_ASAP7_75t_R _28880_ (.A(_18006_),
    .B(net1857),
    .Y(_20364_));
 AO21x1_ASAP7_75t_R _28881_ (.A1(_18010_),
    .A2(net1530),
    .B(_17997_),
    .Y(_20365_));
 AND3x1_ASAP7_75t_R _28882_ (.A(_18007_),
    .B(_20364_),
    .C(_20365_),
    .Y(_20366_));
 NAND2x1_ASAP7_75t_R _28883_ (.A(_20363_),
    .B(_20366_),
    .Y(_20367_));
 NOR2x2_ASAP7_75t_R _28884_ (.A(_20359_),
    .B(_20367_),
    .Y(_20368_));
 INVx1_ASAP7_75t_R _28885_ (.A(_20368_),
    .Y(_20369_));
 INVx1_ASAP7_75t_R _28886_ (.A(_18958_),
    .Y(_20370_));
 AOI211x1_ASAP7_75t_R _28887_ (.A1(net1062),
    .A2(net1117),
    .B(_18054_),
    .C(net1369),
    .Y(_20371_));
 AO21x1_ASAP7_75t_R _28888_ (.A1(_20370_),
    .A2(_18952_),
    .B(_20371_),
    .Y(_20372_));
 AO21x1_ASAP7_75t_R _28889_ (.A1(net2821),
    .A2(net939),
    .B(net3304),
    .Y(_20373_));
 NAND2x2_ASAP7_75t_R _28890_ (.A(_18105_),
    .B(_18040_),
    .Y(_20374_));
 NAND3x2_ASAP7_75t_R _28891_ (.B(_19386_),
    .C(_20374_),
    .Y(_20375_),
    .A(_20373_));
 NAND2x2_ASAP7_75t_R _28892_ (.A(_18113_),
    .B(_18952_),
    .Y(_20376_));
 AO21x1_ASAP7_75t_R _28893_ (.A1(_18010_),
    .A2(_18147_),
    .B(net2303),
    .Y(_20377_));
 NAND2x2_ASAP7_75t_R _28894_ (.A(_20376_),
    .B(_20377_),
    .Y(_20378_));
 NOR3x2_ASAP7_75t_R _28895_ (.B(_20375_),
    .C(_20378_),
    .Y(_20379_),
    .A(_20372_));
 AO21x1_ASAP7_75t_R _28896_ (.A1(_18010_),
    .A2(net3217),
    .B(net3200),
    .Y(_20380_));
 AO21x1_ASAP7_75t_R _28897_ (.A1(net3184),
    .A2(net974),
    .B(net3200),
    .Y(_20381_));
 NAND2x1_ASAP7_75t_R _28898_ (.A(net2877),
    .B(_18941_),
    .Y(_20382_));
 AND3x2_ASAP7_75t_R _28899_ (.A(_20380_),
    .B(_20381_),
    .C(_20382_),
    .Y(_20383_));
 AO21x1_ASAP7_75t_R _28900_ (.A1(net1690),
    .A2(net3285),
    .B(net1907),
    .Y(_20384_));
 AND2x2_ASAP7_75t_R _28901_ (.A(_20384_),
    .B(_18071_),
    .Y(_20385_));
 OA21x2_ASAP7_75t_R _28902_ (.A1(_18883_),
    .A2(net2181),
    .B(_18078_),
    .Y(_20386_));
 NAND3x2_ASAP7_75t_R _28903_ (.B(_20385_),
    .C(_20386_),
    .Y(_20387_),
    .A(_20383_));
 INVx1_ASAP7_75t_R _28904_ (.A(_20387_),
    .Y(_20388_));
 NAND2x1_ASAP7_75t_R _28905_ (.A(_20379_),
    .B(_20388_),
    .Y(_20389_));
 NOR2x2_ASAP7_75t_R _28906_ (.A(_20369_),
    .B(_20389_),
    .Y(_20390_));
 AO21x1_ASAP7_75t_R _28907_ (.A1(net1795),
    .A2(net2908),
    .B(_18126_),
    .Y(_20391_));
 AO21x1_ASAP7_75t_R _28908_ (.A1(net3307),
    .A2(_18958_),
    .B(_18126_),
    .Y(_20392_));
 NAND2x2_ASAP7_75t_R _28909_ (.A(_18123_),
    .B(net1859),
    .Y(_20393_));
 NAND3x2_ASAP7_75t_R _28910_ (.B(_20392_),
    .C(_20393_),
    .Y(_20394_),
    .A(_20391_));
 OA21x2_ASAP7_75t_R _28911_ (.A1(net3218),
    .A2(_18134_),
    .B(_18107_),
    .Y(_20395_));
 AO21x1_ASAP7_75t_R _28912_ (.A1(net1815),
    .A2(net2680),
    .B(_20395_),
    .Y(_20396_));
 NAND2x2_ASAP7_75t_R _28913_ (.A(net3222),
    .B(_18867_),
    .Y(_20397_));
 NOR3x2_ASAP7_75t_R _28914_ (.B(_20396_),
    .C(_20397_),
    .Y(_20398_),
    .A(_20394_));
 NOR2x1_ASAP7_75t_R _28915_ (.A(net3186),
    .B(_17931_),
    .Y(_20399_));
 NOR2x1_ASAP7_75t_R _28916_ (.A(_20399_),
    .B(_17964_),
    .Y(_20400_));
 NOR2x1_ASAP7_75t_R _28917_ (.A(_17938_),
    .B(_17931_),
    .Y(_20401_));
 INVx1_ASAP7_75t_R _28918_ (.A(_20401_),
    .Y(_20402_));
 NAND2x1_ASAP7_75t_R _28919_ (.A(net2720),
    .B(_17948_),
    .Y(_20403_));
 AND3x1_ASAP7_75t_R _28920_ (.A(_20400_),
    .B(_20402_),
    .C(_20403_),
    .Y(_20404_));
 AO21x1_ASAP7_75t_R _28921_ (.A1(_17980_),
    .A2(net3189),
    .B(_17968_),
    .Y(_20405_));
 AO21x1_ASAP7_75t_R _28922_ (.A1(_17987_),
    .A2(net1624),
    .B(_17968_),
    .Y(_20406_));
 NOR2x1_ASAP7_75t_R _28923_ (.A(_18081_),
    .B(_17968_),
    .Y(_20407_));
 INVx1_ASAP7_75t_R _28924_ (.A(_20407_),
    .Y(_20408_));
 NAND2x1_ASAP7_75t_R _28925_ (.A(net2842),
    .B(_18089_),
    .Y(_20409_));
 AND4x1_ASAP7_75t_R _28926_ (.A(_20405_),
    .B(_20406_),
    .C(_20408_),
    .D(_20409_),
    .Y(_20410_));
 NAND2x1_ASAP7_75t_R _28927_ (.A(_20404_),
    .B(_20410_),
    .Y(_20411_));
 INVx1_ASAP7_75t_R _28928_ (.A(_20411_),
    .Y(_20412_));
 NAND2x1_ASAP7_75t_R _28929_ (.A(_20398_),
    .B(_20412_),
    .Y(_20413_));
 AO21x1_ASAP7_75t_R _28930_ (.A1(net3186),
    .A2(net1839),
    .B(_18156_),
    .Y(_20414_));
 NAND2x1_ASAP7_75t_R _28931_ (.A(net2163),
    .B(net3091),
    .Y(_20415_));
 AND3x1_ASAP7_75t_R _28932_ (.A(_20414_),
    .B(_18888_),
    .C(_20415_),
    .Y(_20416_));
 AO21x1_ASAP7_75t_R _28933_ (.A1(_18073_),
    .A2(net3191),
    .B(_18144_),
    .Y(_20417_));
 NAND2x1_ASAP7_75t_R _28934_ (.A(_18105_),
    .B(_18151_),
    .Y(_20418_));
 AND4x1_ASAP7_75t_R _28935_ (.A(_18146_),
    .B(_20417_),
    .C(_20418_),
    .D(_19417_),
    .Y(_20419_));
 NAND2x1_ASAP7_75t_R _28936_ (.A(_20416_),
    .B(_20419_),
    .Y(_20420_));
 OA21x2_ASAP7_75t_R _28937_ (.A1(_18178_),
    .A2(_18113_),
    .B(net3299),
    .Y(_20421_));
 NOR2x1_ASAP7_75t_R _28938_ (.A(_18169_),
    .B(_18028_),
    .Y(_20422_));
 AOI211x1_ASAP7_75t_R _28939_ (.A1(_17952_),
    .A2(net3299),
    .B(_20421_),
    .C(_20422_),
    .Y(_20423_));
 AO21x1_ASAP7_75t_R _28940_ (.A1(_18014_),
    .A2(_18002_),
    .B(_19423_),
    .Y(_20424_));
 NAND2x1_ASAP7_75t_R _28941_ (.A(_20424_),
    .B(_19791_),
    .Y(_20425_));
 NAND2x2_ASAP7_75t_R _28942_ (.A(net2245),
    .B(_18113_),
    .Y(_20426_));
 AO21x1_ASAP7_75t_R _28943_ (.A1(_18028_),
    .A2(_18081_),
    .B(_19423_),
    .Y(_20427_));
 NAND2x1_ASAP7_75t_R _28944_ (.A(_20426_),
    .B(_20427_),
    .Y(_20428_));
 NOR2x2_ASAP7_75t_R _28945_ (.A(_20425_),
    .B(_20428_),
    .Y(_20429_));
 NAND2x1_ASAP7_75t_R _28946_ (.A(net3343),
    .B(_18046_),
    .Y(_20430_));
 AO21x1_ASAP7_75t_R _28947_ (.A1(_20430_),
    .A2(net3284),
    .B(_18169_),
    .Y(_20431_));
 NAND3x2_ASAP7_75t_R _28948_ (.B(_20429_),
    .C(_20431_),
    .Y(_20432_),
    .A(_20423_));
 NOR2x2_ASAP7_75t_R _28949_ (.A(_20420_),
    .B(_20432_),
    .Y(_20433_));
 INVx1_ASAP7_75t_R _28950_ (.A(_20433_),
    .Y(_20434_));
 NOR2x2_ASAP7_75t_R _28951_ (.A(_20413_),
    .B(_20434_),
    .Y(_20435_));
 NAND2x2_ASAP7_75t_R _28952_ (.A(_20390_),
    .B(_20435_),
    .Y(_20436_));
 XOR2x2_ASAP7_75t_R _28953_ (.A(_20352_),
    .B(_20436_),
    .Y(_20437_));
 XOR2x1_ASAP7_75t_R _28954_ (.A(_20277_),
    .Y(_20438_),
    .B(_20437_));
 NAND2x1_ASAP7_75t_R _28955_ (.A(_20438_),
    .B(_20171_),
    .Y(_20439_));
 XOR2x2_ASAP7_75t_R _28956_ (.A(_19961_),
    .B(_18229_),
    .Y(_20440_));
 XOR2x1_ASAP7_75t_R _28957_ (.A(_20440_),
    .Y(_20441_),
    .B(net2537));
 INVx1_ASAP7_75t_R _28958_ (.A(_20379_),
    .Y(_20442_));
 NOR2x1_ASAP7_75t_R _28959_ (.A(_20387_),
    .B(_20442_),
    .Y(_20443_));
 NAND2x1_ASAP7_75t_R _28960_ (.A(_20368_),
    .B(_20443_),
    .Y(_20444_));
 INVx1_ASAP7_75t_R _28961_ (.A(_20398_),
    .Y(_20445_));
 NOR2x1_ASAP7_75t_R _28962_ (.A(_20411_),
    .B(_20445_),
    .Y(_20446_));
 NAND2x2_ASAP7_75t_R _28963_ (.A(_20433_),
    .B(_20446_),
    .Y(_20447_));
 NOR2x2_ASAP7_75t_R _28964_ (.A(_20444_),
    .B(_20447_),
    .Y(_20448_));
 XOR2x2_ASAP7_75t_R _28965_ (.A(_20352_),
    .B(_20448_),
    .Y(_20449_));
 XOR2x1_ASAP7_75t_R _28966_ (.A(_20277_),
    .Y(_20450_),
    .B(_20449_));
 NAND2x1_ASAP7_75t_R _28967_ (.A(_20441_),
    .B(_20450_),
    .Y(_20451_));
 TAPCELL_ASAP7_75t_R TAP_822 ();
 TAPCELL_ASAP7_75t_R TAP_821 ();
 AOI21x1_ASAP7_75t_R _28970_ (.A1(_20439_),
    .A2(_20451_),
    .B(net390),
    .Y(_20454_));
 OAI21x1_ASAP7_75t_R _28971_ (.A1(_20087_),
    .A2(_20454_),
    .B(_14682_),
    .Y(_20455_));
 NOR2x1_ASAP7_75t_R _28972_ (.A(net397),
    .B(_00911_),
    .Y(_20456_));
 NAND2x1_ASAP7_75t_R _28973_ (.A(_20441_),
    .B(_20438_),
    .Y(_20457_));
 NAND2x1_ASAP7_75t_R _28974_ (.A(_20450_),
    .B(_20171_),
    .Y(_20458_));
 AOI21x1_ASAP7_75t_R _28975_ (.A1(_20457_),
    .A2(_20458_),
    .B(net390),
    .Y(_20459_));
 OAI21x1_ASAP7_75t_R _28976_ (.A1(_20456_),
    .A2(_20459_),
    .B(_00448_),
    .Y(_20460_));
 NAND2x2_ASAP7_75t_R _28977_ (.A(_20455_),
    .B(_20460_),
    .Y(_00125_));
 NOR2x1_ASAP7_75t_R _28978_ (.A(net397),
    .B(_00910_),
    .Y(_20461_));
 INVx1_ASAP7_75t_R _28979_ (.A(_20461_),
    .Y(_20462_));
 NAND2x2_ASAP7_75t_R _28980_ (.A(_17764_),
    .B(_17762_),
    .Y(_20463_));
 OA31x2_ASAP7_75t_R _28981_ (.A1(_17609_),
    .A2(_17774_),
    .A3(net1901),
    .B1(_18825_),
    .Y(_20464_));
 OAI21x1_ASAP7_75t_R _28982_ (.A1(_18834_),
    .A2(_17788_),
    .B(_19890_),
    .Y(_20465_));
 AO21x1_ASAP7_75t_R _28983_ (.A1(_17639_),
    .A2(_17647_),
    .B(_17744_),
    .Y(_20466_));
 NAND2x2_ASAP7_75t_R _28984_ (.A(_20465_),
    .B(_20466_),
    .Y(_20467_));
 NOR3x2_ASAP7_75t_R _28985_ (.B(_20464_),
    .C(_20467_),
    .Y(_20468_),
    .A(_20463_));
 OA21x2_ASAP7_75t_R _28986_ (.A1(_18812_),
    .A2(_17638_),
    .B(_20280_),
    .Y(_20469_));
 AO21x1_ASAP7_75t_R _28987_ (.A1(net1030),
    .A2(net2630),
    .B(_17777_),
    .Y(_20470_));
 NAND2x1_ASAP7_75t_R _28988_ (.A(_19896_),
    .B(_20470_),
    .Y(_20471_));
 INVx1_ASAP7_75t_R _28989_ (.A(_20471_),
    .Y(_20472_));
 NAND2x1_ASAP7_75t_R _28990_ (.A(_20469_),
    .B(_20472_),
    .Y(_20473_));
 NOR2x1_ASAP7_75t_R _28991_ (.A(net2759),
    .B(_17845_),
    .Y(_20474_));
 NOR2x1_ASAP7_75t_R _28992_ (.A(_20474_),
    .B(_20284_),
    .Y(_20475_));
 AO21x1_ASAP7_75t_R _28993_ (.A1(net1030),
    .A2(net1081),
    .B(net2758),
    .Y(_20476_));
 AO21x1_ASAP7_75t_R _28994_ (.A1(_17834_),
    .A2(net1082),
    .B(net2758),
    .Y(_20477_));
 NAND2x1_ASAP7_75t_R _28995_ (.A(_20476_),
    .B(_20477_),
    .Y(_20478_));
 INVx1_ASAP7_75t_R _28996_ (.A(_20478_),
    .Y(_20479_));
 NAND2x1_ASAP7_75t_R _28997_ (.A(_20475_),
    .B(_20479_),
    .Y(_20480_));
 NOR2x1_ASAP7_75t_R _28998_ (.A(_20473_),
    .B(_20480_),
    .Y(_20481_));
 NAND2x1_ASAP7_75t_R _28999_ (.A(_20468_),
    .B(_20481_),
    .Y(_20482_));
 AO21x1_ASAP7_75t_R _29000_ (.A1(net1082),
    .A2(_17575_),
    .B(net2883),
    .Y(_20483_));
 OAI21x1_ASAP7_75t_R _29001_ (.A1(net2883),
    .A2(net2451),
    .B(_20483_),
    .Y(_20484_));
 AO21x1_ASAP7_75t_R _29002_ (.A1(_17813_),
    .A2(net1081),
    .B(_17725_),
    .Y(_20485_));
 NAND2x2_ASAP7_75t_R _29003_ (.A(net2087),
    .B(_17733_),
    .Y(_20486_));
 OAI21x1_ASAP7_75t_R _29004_ (.A1(_18834_),
    .A2(_17745_),
    .B(_17733_),
    .Y(_20487_));
 NAND3x2_ASAP7_75t_R _29005_ (.B(_20486_),
    .C(_20487_),
    .Y(_20488_),
    .A(_20485_));
 NOR2x2_ASAP7_75t_R _29006_ (.A(_20484_),
    .B(_20488_),
    .Y(_20489_));
 AOI221x1_ASAP7_75t_R _29007_ (.A1(net1123),
    .A2(net2879),
    .B1(_17575_),
    .B2(net2902),
    .C(_17701_),
    .Y(_20490_));
 INVx1_ASAP7_75t_R _29008_ (.A(_17912_),
    .Y(_20491_));
 AO21x1_ASAP7_75t_R _29009_ (.A1(net3086),
    .A2(_18834_),
    .B(_20491_),
    .Y(_20492_));
 NOR2x2_ASAP7_75t_R _29010_ (.A(_20490_),
    .B(_20492_),
    .Y(_20493_));
 AO21x1_ASAP7_75t_R _29011_ (.A1(_17756_),
    .A2(net941),
    .B(_17691_),
    .Y(_20494_));
 NAND2x1_ASAP7_75t_R _29012_ (.A(_20301_),
    .B(_20494_),
    .Y(_20495_));
 AO21x1_ASAP7_75t_R _29013_ (.A1(net1030),
    .A2(net1081),
    .B(_17691_),
    .Y(_20496_));
 AO21x1_ASAP7_75t_R _29014_ (.A1(_17639_),
    .A2(_17647_),
    .B(net3088),
    .Y(_20497_));
 NAND2x1_ASAP7_75t_R _29015_ (.A(_20496_),
    .B(_20497_),
    .Y(_20498_));
 NOR2x2_ASAP7_75t_R _29016_ (.A(_20495_),
    .B(_20498_),
    .Y(_20499_));
 NAND3x2_ASAP7_75t_R _29017_ (.B(_20493_),
    .C(_20499_),
    .Y(_20500_),
    .A(_20489_));
 NOR2x1_ASAP7_75t_R _29018_ (.A(_20500_),
    .B(_20482_),
    .Y(_20501_));
 NAND2x1_ASAP7_75t_R _29019_ (.A(_17607_),
    .B(_17618_),
    .Y(_20502_));
 NAND3x1_ASAP7_75t_R _29020_ (.A(_17855_),
    .B(_18771_),
    .C(_20502_),
    .Y(_20503_));
 NOR2x1_ASAP7_75t_R _29021_ (.A(net2904),
    .B(_17589_),
    .Y(_20504_));
 OAI21x1_ASAP7_75t_R _29022_ (.A1(net2862),
    .A2(net2879),
    .B(_20504_),
    .Y(_20505_));
 NAND2x1_ASAP7_75t_R _29023_ (.A(_17604_),
    .B(_17788_),
    .Y(_20506_));
 AO21x1_ASAP7_75t_R _29024_ (.A1(_17813_),
    .A2(net2630),
    .B(_17589_),
    .Y(_20507_));
 NAND3x1_ASAP7_75t_R _29025_ (.A(_20505_),
    .B(_20506_),
    .C(_20507_),
    .Y(_20508_));
 NOR2x1_ASAP7_75t_R _29026_ (.A(_20503_),
    .B(_20508_),
    .Y(_20509_));
 AOI211x1_ASAP7_75t_R _29027_ (.A1(net2862),
    .A2(net2879),
    .B(_17566_),
    .C(_17575_),
    .Y(_20510_));
 INVx1_ASAP7_75t_R _29028_ (.A(_20510_),
    .Y(_20511_));
 AO21x1_ASAP7_75t_R _29029_ (.A1(_17572_),
    .A2(net941),
    .B(_17566_),
    .Y(_20512_));
 AO21x1_ASAP7_75t_R _29030_ (.A1(_17639_),
    .A2(_17647_),
    .B(_17566_),
    .Y(_20513_));
 NAND3x1_ASAP7_75t_R _29031_ (.A(_20511_),
    .B(_20512_),
    .C(_20513_),
    .Y(_20514_));
 NOR2x1_ASAP7_75t_R _29032_ (.A(net936),
    .B(_17547_),
    .Y(_20515_));
 AOI211x1_ASAP7_75t_R _29033_ (.A1(net2862),
    .A2(net2879),
    .B(_17547_),
    .C(net1103),
    .Y(_20516_));
 NOR2x1_ASAP7_75t_R _29034_ (.A(_20515_),
    .B(_20516_),
    .Y(_20517_));
 AO21x1_ASAP7_75t_R _29035_ (.A1(net1097),
    .A2(net1082),
    .B(_17547_),
    .Y(_20518_));
 AO21x1_ASAP7_75t_R _29036_ (.A1(_17645_),
    .A2(net3194),
    .B(_17547_),
    .Y(_20519_));
 AND2x2_ASAP7_75t_R _29037_ (.A(_20518_),
    .B(_20519_),
    .Y(_20520_));
 NAND2x1_ASAP7_75t_R _29038_ (.A(_20517_),
    .B(_20520_),
    .Y(_20521_));
 NOR2x1_ASAP7_75t_R _29039_ (.A(_20514_),
    .B(_20521_),
    .Y(_20522_));
 NAND2x2_ASAP7_75t_R _29040_ (.A(_20509_),
    .B(_20522_),
    .Y(_20523_));
 AO21x2_ASAP7_75t_R _29041_ (.A1(_17626_),
    .A2(_17845_),
    .B(_17629_),
    .Y(_20524_));
 AO21x1_ASAP7_75t_R _29042_ (.A1(net1081),
    .A2(net1082),
    .B(_17629_),
    .Y(_20525_));
 NAND2x2_ASAP7_75t_R _29043_ (.A(_17558_),
    .B(_18789_),
    .Y(_20526_));
 NAND3x2_ASAP7_75t_R _29044_ (.B(_20525_),
    .C(_20526_),
    .Y(_20527_),
    .A(_20524_));
 AO21x1_ASAP7_75t_R _29045_ (.A1(net1097),
    .A2(_17892_),
    .B(net2484),
    .Y(_20528_));
 AO21x1_ASAP7_75t_R _29046_ (.A1(_17562_),
    .A2(net941),
    .B(net2484),
    .Y(_20529_));
 NAND2x2_ASAP7_75t_R _29047_ (.A(net2640),
    .B(_17650_),
    .Y(_20530_));
 NAND3x2_ASAP7_75t_R _29048_ (.B(_20529_),
    .C(_20530_),
    .Y(_20531_),
    .A(_20528_));
 NOR2x2_ASAP7_75t_R _29049_ (.A(_20527_),
    .B(_20531_),
    .Y(_20532_));
 AO21x1_ASAP7_75t_R _29050_ (.A1(_17639_),
    .A2(net1097),
    .B(net2847),
    .Y(_20533_));
 NAND2x1_ASAP7_75t_R _29051_ (.A(_19346_),
    .B(_20533_),
    .Y(_20534_));
 AO21x1_ASAP7_75t_R _29052_ (.A1(_17758_),
    .A2(_17695_),
    .B(net2847),
    .Y(_20535_));
 NAND2x1_ASAP7_75t_R _29053_ (.A(_20535_),
    .B(_19348_),
    .Y(_20536_));
 NOR2x2_ASAP7_75t_R _29054_ (.A(_20534_),
    .B(_20536_),
    .Y(_20537_));
 OAI21x1_ASAP7_75t_R _29055_ (.A1(net1082),
    .A2(_17670_),
    .B(_17672_),
    .Y(_20538_));
 OA21x2_ASAP7_75t_R _29056_ (.A1(_17757_),
    .A2(_17694_),
    .B(_17671_),
    .Y(_20539_));
 NOR3x2_ASAP7_75t_R _29057_ (.B(_20539_),
    .C(_20320_),
    .Y(_20540_),
    .A(_20538_));
 NAND3x2_ASAP7_75t_R _29058_ (.B(_20537_),
    .C(_20540_),
    .Y(_20541_),
    .A(_20532_));
 NOR2x2_ASAP7_75t_R _29059_ (.A(_20523_),
    .B(_20541_),
    .Y(_20542_));
 NAND2x2_ASAP7_75t_R _29060_ (.A(_20501_),
    .B(_20542_),
    .Y(_20543_));
 NOR2x2_ASAP7_75t_R _29061_ (.A(net2143),
    .B(_20543_),
    .Y(_20544_));
 OAI21x1_ASAP7_75t_R _29062_ (.A1(net3367),
    .A2(_18000_),
    .B(net3092),
    .Y(_20545_));
 OAI21x1_ASAP7_75t_R _29063_ (.A1(_17925_),
    .A2(net2843),
    .B(net3092),
    .Y(_20546_));
 NAND2x2_ASAP7_75t_R _29064_ (.A(net3092),
    .B(net3091),
    .Y(_20547_));
 NAND3x2_ASAP7_75t_R _29065_ (.B(_20546_),
    .C(_20547_),
    .Y(_20548_),
    .A(_20545_));
 NOR2x2_ASAP7_75t_R _29066_ (.A(net3216),
    .B(_19855_),
    .Y(_20549_));
 NAND2x2_ASAP7_75t_R _29067_ (.A(_19802_),
    .B(_18916_),
    .Y(_20550_));
 NAND2x2_ASAP7_75t_R _29068_ (.A(_20550_),
    .B(_18913_),
    .Y(_20551_));
 NOR3x2_ASAP7_75t_R _29069_ (.B(_20549_),
    .C(_20551_),
    .Y(_20552_),
    .A(_20548_));
 INVx1_ASAP7_75t_R _29070_ (.A(_20552_),
    .Y(_20553_));
 AOI211x1_ASAP7_75t_R _29071_ (.A1(net3201),
    .A2(net3124),
    .B(_17997_),
    .C(net1073),
    .Y(_20554_));
 AND3x1_ASAP7_75t_R _29072_ (.A(_18006_),
    .B(_17923_),
    .C(net3201),
    .Y(_20555_));
 AOI211x1_ASAP7_75t_R _29073_ (.A1(_18113_),
    .A2(_18006_),
    .B(_20554_),
    .C(_20555_),
    .Y(_20556_));
 AOI211x1_ASAP7_75t_R _29074_ (.A1(net1059),
    .A2(net3308),
    .B(net1369),
    .C(net1955),
    .Y(_20557_));
 INVx1_ASAP7_75t_R _29075_ (.A(_20557_),
    .Y(_20558_));
 AO21x1_ASAP7_75t_R _29076_ (.A1(_17984_),
    .A2(net974),
    .B(net1955),
    .Y(_20559_));
 AO21x1_ASAP7_75t_R _29077_ (.A1(net1121),
    .A2(_18002_),
    .B(net1955),
    .Y(_20560_));
 AND3x2_ASAP7_75t_R _29078_ (.A(_20558_),
    .B(_20559_),
    .C(_20560_),
    .Y(_20561_));
 NAND2x1_ASAP7_75t_R _29079_ (.A(_20556_),
    .B(_20561_),
    .Y(_20562_));
 NOR2x1_ASAP7_75t_R _29080_ (.A(_20553_),
    .B(_20562_),
    .Y(_20563_));
 AO21x1_ASAP7_75t_R _29081_ (.A1(_17987_),
    .A2(net974),
    .B(net1911),
    .Y(_20564_));
 OAI21x1_ASAP7_75t_R _29082_ (.A1(_17963_),
    .A2(net1911),
    .B(_20564_),
    .Y(_20565_));
 AO21x1_ASAP7_75t_R _29083_ (.A1(net1121),
    .A2(_18022_),
    .B(net2181),
    .Y(_20566_));
 AO21x1_ASAP7_75t_R _29084_ (.A1(net2796),
    .A2(_18147_),
    .B(net2181),
    .Y(_20567_));
 NAND2x2_ASAP7_75t_R _29085_ (.A(_20566_),
    .B(_20567_),
    .Y(_20568_));
 NOR2x1_ASAP7_75t_R _29086_ (.A(net1911),
    .B(net3213),
    .Y(_20569_));
 AO21x1_ASAP7_75t_R _29087_ (.A1(net1117),
    .A2(_19403_),
    .B(_20569_),
    .Y(_20570_));
 NOR3x2_ASAP7_75t_R _29088_ (.B(_20568_),
    .C(_20570_),
    .Y(_20571_),
    .A(_20565_));
 INVx2_ASAP7_75t_R _29089_ (.A(_20571_),
    .Y(_20572_));
 AO21x1_ASAP7_75t_R _29090_ (.A1(_18147_),
    .A2(_17962_),
    .B(net2303),
    .Y(_20573_));
 AO21x1_ASAP7_75t_R _29091_ (.A1(_18883_),
    .A2(_18022_),
    .B(net2303),
    .Y(_20574_));
 AND3x1_ASAP7_75t_R _29092_ (.A(_20573_),
    .B(_20574_),
    .C(_20376_),
    .Y(_20575_));
 AO21x1_ASAP7_75t_R _29093_ (.A1(_17938_),
    .A2(net3213),
    .B(_18039_),
    .Y(_20576_));
 OAI21x1_ASAP7_75t_R _29094_ (.A1(_17983_),
    .A2(_19824_),
    .B(_20576_),
    .Y(_20577_));
 NOR2x1_ASAP7_75t_R _29095_ (.A(_18039_),
    .B(net1350),
    .Y(_20578_));
 OR3x2_ASAP7_75t_R _29096_ (.A(_20578_),
    .B(_18962_),
    .C(_18961_),
    .Y(_20579_));
 NOR2x2_ASAP7_75t_R _29097_ (.A(_20577_),
    .B(_20579_),
    .Y(_20580_));
 NAND2x1_ASAP7_75t_R _29098_ (.A(_20575_),
    .B(_20580_),
    .Y(_20581_));
 NOR2x1_ASAP7_75t_R _29099_ (.A(_20572_),
    .B(_20581_),
    .Y(_20582_));
 NAND2x1_ASAP7_75t_R _29100_ (.A(_20563_),
    .B(_20582_),
    .Y(_20583_));
 OA21x2_ASAP7_75t_R _29101_ (.A1(net3091),
    .A2(_18860_),
    .B(_18151_),
    .Y(_20584_));
 AND3x1_ASAP7_75t_R _29102_ (.A(_18151_),
    .B(net3343),
    .C(_17983_),
    .Y(_20585_));
 NOR2x2_ASAP7_75t_R _29103_ (.A(_20584_),
    .B(_20585_),
    .Y(_20586_));
 AND2x2_ASAP7_75t_R _29104_ (.A(_18160_),
    .B(_18161_),
    .Y(_20587_));
 OA21x2_ASAP7_75t_R _29105_ (.A1(_18178_),
    .A2(_18110_),
    .B(net3192),
    .Y(_20588_));
 AOI21x1_ASAP7_75t_R _29106_ (.A1(_18037_),
    .A2(net3192),
    .B(_20588_),
    .Y(_20589_));
 NAND3x2_ASAP7_75t_R _29107_ (.B(_20587_),
    .C(_20589_),
    .Y(_20590_),
    .A(_20586_));
 OAI21x1_ASAP7_75t_R _29108_ (.A1(_17937_),
    .A2(_18185_),
    .B(_20426_),
    .Y(_20591_));
 OA21x2_ASAP7_75t_R _29109_ (.A1(_18000_),
    .A2(net3207),
    .B(net2245),
    .Y(_20592_));
 NOR3x1_ASAP7_75t_R _29110_ (.A(_20591_),
    .B(_19790_),
    .C(_20592_),
    .Y(_20593_));
 OA21x2_ASAP7_75t_R _29111_ (.A1(_18047_),
    .A2(_18869_),
    .B(_18165_),
    .Y(_20594_));
 NOR2x1_ASAP7_75t_R _29112_ (.A(_18164_),
    .B(_18166_),
    .Y(_20595_));
 NOR2x1_ASAP7_75t_R _29113_ (.A(_20594_),
    .B(_20595_),
    .Y(_20596_));
 NOR2x1_ASAP7_75t_R _29114_ (.A(_18169_),
    .B(net1529),
    .Y(_20597_));
 NOR2x1_ASAP7_75t_R _29115_ (.A(_20597_),
    .B(_20421_),
    .Y(_20598_));
 AND2x2_ASAP7_75t_R _29116_ (.A(_20598_),
    .B(_20596_),
    .Y(_20599_));
 NAND2x2_ASAP7_75t_R _29117_ (.A(_20593_),
    .B(_20599_),
    .Y(_20600_));
 NOR2x2_ASAP7_75t_R _29118_ (.A(_20590_),
    .B(_20600_),
    .Y(_20601_));
 AOI221x1_ASAP7_75t_R _29119_ (.A1(net1057),
    .A2(net3124),
    .B1(net3284),
    .B2(net1371),
    .C(net1746),
    .Y(_20602_));
 AO21x1_ASAP7_75t_R _29120_ (.A1(_17932_),
    .A2(_18860_),
    .B(_17964_),
    .Y(_20603_));
 NOR2x1_ASAP7_75t_R _29121_ (.A(_20602_),
    .B(_20603_),
    .Y(_20604_));
 AOI21x1_ASAP7_75t_R _29122_ (.A1(_17958_),
    .A2(net3186),
    .B(_17968_),
    .Y(_20605_));
 NOR2x1_ASAP7_75t_R _29123_ (.A(_20407_),
    .B(_20605_),
    .Y(_20606_));
 AO21x1_ASAP7_75t_R _29124_ (.A1(net1675),
    .A2(_18073_),
    .B(net2364),
    .Y(_20607_));
 AO21x1_ASAP7_75t_R _29125_ (.A1(net1121),
    .A2(_18057_),
    .B(net2364),
    .Y(_20608_));
 NAND3x1_ASAP7_75t_R _29126_ (.A(_20606_),
    .B(_20607_),
    .C(_20608_),
    .Y(_20609_));
 INVx1_ASAP7_75t_R _29127_ (.A(_20609_),
    .Y(_20610_));
 NAND2x1_ASAP7_75t_R _29128_ (.A(_20610_),
    .B(_20604_),
    .Y(_20611_));
 AO21x1_ASAP7_75t_R _29129_ (.A1(_18022_),
    .A2(net3284),
    .B(_18126_),
    .Y(_20612_));
 OAI21x1_ASAP7_75t_R _29130_ (.A1(_18010_),
    .A2(_18126_),
    .B(_20612_),
    .Y(_20613_));
 INVx1_ASAP7_75t_R _29131_ (.A(_20613_),
    .Y(_20614_));
 NAND2x1_ASAP7_75t_R _29132_ (.A(_19452_),
    .B(_18867_),
    .Y(_20615_));
 AO21x1_ASAP7_75t_R _29133_ (.A1(_17980_),
    .A2(net3189),
    .B(_18864_),
    .Y(_20616_));
 NAND2x2_ASAP7_75t_R _29134_ (.A(net2680),
    .B(_18134_),
    .Y(_20617_));
 NAND3x2_ASAP7_75t_R _29135_ (.B(_20617_),
    .C(net3223),
    .Y(_20618_),
    .A(_20616_));
 NOR2x1_ASAP7_75t_R _29136_ (.A(_20615_),
    .B(_20618_),
    .Y(_20619_));
 NAND2x1_ASAP7_75t_R _29137_ (.A(_20614_),
    .B(_20619_),
    .Y(_20620_));
 NOR2x1_ASAP7_75t_R _29138_ (.A(_20620_),
    .B(_20611_),
    .Y(_20621_));
 NAND2x2_ASAP7_75t_R _29139_ (.A(_20601_),
    .B(_20621_),
    .Y(_20622_));
 NOR2x2_ASAP7_75t_R _29140_ (.A(_20583_),
    .B(_20622_),
    .Y(_20623_));
 NAND2x2_ASAP7_75t_R _29141_ (.A(_17974_),
    .B(_20623_),
    .Y(_20624_));
 NOR2x1_ASAP7_75t_R _29142_ (.A(_20544_),
    .B(_20624_),
    .Y(_20625_));
 INVx1_ASAP7_75t_R _29143_ (.A(_20532_),
    .Y(_20626_));
 NAND2x1_ASAP7_75t_R _29144_ (.A(_20537_),
    .B(_20540_),
    .Y(_20627_));
 NOR2x1_ASAP7_75t_R _29145_ (.A(_20626_),
    .B(_20627_),
    .Y(_20628_));
 INVx1_ASAP7_75t_R _29146_ (.A(_20523_),
    .Y(_20629_));
 NAND2x1_ASAP7_75t_R _29147_ (.A(_20628_),
    .B(_20629_),
    .Y(_20630_));
 INVx1_ASAP7_75t_R _29148_ (.A(_20468_),
    .Y(_20631_));
 INVx1_ASAP7_75t_R _29149_ (.A(_20469_),
    .Y(_20632_));
 NOR2x1_ASAP7_75t_R _29150_ (.A(_20471_),
    .B(_20632_),
    .Y(_20633_));
 INVx1_ASAP7_75t_R _29151_ (.A(_20475_),
    .Y(_20634_));
 NOR2x1_ASAP7_75t_R _29152_ (.A(_20478_),
    .B(_20634_),
    .Y(_20635_));
 NAND2x1_ASAP7_75t_R _29153_ (.A(_20633_),
    .B(_20635_),
    .Y(_20636_));
 NOR2x1_ASAP7_75t_R _29154_ (.A(_20631_),
    .B(_20636_),
    .Y(_20637_));
 INVx1_ASAP7_75t_R _29155_ (.A(_20500_),
    .Y(_20638_));
 NAND2x1_ASAP7_75t_R _29156_ (.A(_20637_),
    .B(_20638_),
    .Y(_20639_));
 NOR2x1_ASAP7_75t_R _29157_ (.A(_20630_),
    .B(_20639_),
    .Y(_20640_));
 NAND2x1_ASAP7_75t_R _29158_ (.A(_17918_),
    .B(_20640_),
    .Y(_20641_));
 INVx4_ASAP7_75t_R _29159_ (.A(_17974_),
    .Y(_20642_));
 NAND3x1_ASAP7_75t_R _29160_ (.A(_20571_),
    .B(_20580_),
    .C(_20575_),
    .Y(_20643_));
 NAND3x1_ASAP7_75t_R _29161_ (.A(_20552_),
    .B(_20556_),
    .C(_20561_),
    .Y(_20644_));
 NOR2x1_ASAP7_75t_R _29162_ (.A(_20643_),
    .B(_20644_),
    .Y(_20645_));
 NOR3x1_ASAP7_75t_R _29163_ (.A(_20618_),
    .B(_20615_),
    .C(_20613_),
    .Y(_20646_));
 INVx1_ASAP7_75t_R _29164_ (.A(_20604_),
    .Y(_20647_));
 NOR2x1_ASAP7_75t_R _29165_ (.A(_20609_),
    .B(_20647_),
    .Y(_20648_));
 NAND2x1_ASAP7_75t_R _29166_ (.A(_20646_),
    .B(_20648_),
    .Y(_20649_));
 INVx1_ASAP7_75t_R _29167_ (.A(_20601_),
    .Y(_20650_));
 NOR2x2_ASAP7_75t_R _29168_ (.A(_20649_),
    .B(_20650_),
    .Y(_20651_));
 NAND2x2_ASAP7_75t_R _29169_ (.A(_20645_),
    .B(_20651_),
    .Y(_20652_));
 NOR2x2_ASAP7_75t_R _29170_ (.A(_20642_),
    .B(_20652_),
    .Y(_20653_));
 NOR2x1_ASAP7_75t_R _29171_ (.A(_20641_),
    .B(_20653_),
    .Y(_20654_));
 AND3x1_ASAP7_75t_R _29172_ (.A(_18262_),
    .B(_18266_),
    .C(_18274_),
    .Y(_20655_));
 NAND2x2_ASAP7_75t_R _29173_ (.A(_18277_),
    .B(_20655_),
    .Y(_20656_));
 NOR3x2_ASAP7_75t_R _29174_ (.B(_18275_),
    .C(_18276_),
    .Y(_20657_),
    .A(_20656_));
 AO21x1_ASAP7_75t_R _29175_ (.A1(_18453_),
    .A2(net1482),
    .B(_18266_),
    .Y(_20658_));
 NAND2x1_ASAP7_75t_R _29176_ (.A(_20102_),
    .B(_20658_),
    .Y(_20659_));
 AO21x1_ASAP7_75t_R _29177_ (.A1(net1254),
    .A2(net2004),
    .B(_18266_),
    .Y(_20660_));
 AO21x1_ASAP7_75t_R _29178_ (.A1(_18350_),
    .A2(_18402_),
    .B(_18266_),
    .Y(_20661_));
 NAND2x1_ASAP7_75t_R _29179_ (.A(_20660_),
    .B(_20661_),
    .Y(_20662_));
 NOR2x2_ASAP7_75t_R _29180_ (.A(_20659_),
    .B(_20662_),
    .Y(_20663_));
 AO21x1_ASAP7_75t_R _29181_ (.A1(net1954),
    .A2(net2978),
    .B(_18428_),
    .Y(_20664_));
 OAI21x1_ASAP7_75t_R _29182_ (.A1(_18314_),
    .A2(_18428_),
    .B(_20664_),
    .Y(_20665_));
 NAND2x1_ASAP7_75t_R _29183_ (.A(net1392),
    .B(_18235_),
    .Y(_20666_));
 AO21x1_ASAP7_75t_R _29184_ (.A1(_20666_),
    .A2(net2008),
    .B(_18439_),
    .Y(_20667_));
 AO21x1_ASAP7_75t_R _29185_ (.A1(_19164_),
    .A2(_19493_),
    .B(_18439_),
    .Y(_20668_));
 NAND2x2_ASAP7_75t_R _29186_ (.A(_20667_),
    .B(_20668_),
    .Y(_20669_));
 NOR2x2_ASAP7_75t_R _29187_ (.A(_20665_),
    .B(_20669_),
    .Y(_20670_));
 OAI21x1_ASAP7_75t_R _29188_ (.A1(net1199),
    .A2(_18273_),
    .B(_18271_),
    .Y(_20671_));
 AOI221x1_ASAP7_75t_R _29189_ (.A1(net1087),
    .A2(_18237_),
    .B1(net2008),
    .B2(net2977),
    .C(_18248_),
    .Y(_20672_));
 NOR2x2_ASAP7_75t_R _29190_ (.A(_20671_),
    .B(_20672_),
    .Y(_20673_));
 NAND3x2_ASAP7_75t_R _29191_ (.B(_20670_),
    .C(_20673_),
    .Y(_20674_),
    .A(_20663_));
 AOI211x1_ASAP7_75t_R _29192_ (.A1(net2999),
    .A2(_18237_),
    .B(net3312),
    .C(_18290_),
    .Y(_20675_));
 INVx1_ASAP7_75t_R _29193_ (.A(_20675_),
    .Y(_20676_));
 AO21x1_ASAP7_75t_R _29194_ (.A1(_18350_),
    .A2(_18402_),
    .B(net3312),
    .Y(_20677_));
 NAND3x1_ASAP7_75t_R _29195_ (.A(_20676_),
    .B(_19965_),
    .C(_20677_),
    .Y(_20678_));
 AO31x2_ASAP7_75t_R _29196_ (.A1(net937),
    .A2(net2044),
    .A3(net2634),
    .B(_18456_),
    .Y(_20679_));
 NAND2x1_ASAP7_75t_R _29197_ (.A(_20679_),
    .B(_18462_),
    .Y(_20680_));
 NOR2x1_ASAP7_75t_R _29198_ (.A(_20678_),
    .B(_20680_),
    .Y(_20681_));
 AO31x2_ASAP7_75t_R _29199_ (.A1(_18489_),
    .A2(_18351_),
    .A3(net1954),
    .B(net2595),
    .Y(_20682_));
 NAND2x1_ASAP7_75t_R _29200_ (.A(net2669),
    .B(_19472_),
    .Y(_20683_));
 AND2x2_ASAP7_75t_R _29201_ (.A(_20117_),
    .B(_20683_),
    .Y(_20684_));
 NAND2x1_ASAP7_75t_R _29202_ (.A(_20682_),
    .B(_20684_),
    .Y(_20685_));
 OA21x2_ASAP7_75t_R _29203_ (.A1(_19202_),
    .A2(_19465_),
    .B(_18483_),
    .Y(_20686_));
 NOR2x1_ASAP7_75t_R _29204_ (.A(_20110_),
    .B(_20686_),
    .Y(_20687_));
 AND2x2_ASAP7_75t_R _29205_ (.A(_19180_),
    .B(_20112_),
    .Y(_20688_));
 NAND2x1_ASAP7_75t_R _29206_ (.A(_20687_),
    .B(_20688_),
    .Y(_20689_));
 NOR2x2_ASAP7_75t_R _29207_ (.A(_20685_),
    .B(_20689_),
    .Y(_20690_));
 NAND2x2_ASAP7_75t_R _29208_ (.A(_20681_),
    .B(_20690_),
    .Y(_20691_));
 NOR2x2_ASAP7_75t_R _29209_ (.A(_20674_),
    .B(_20691_),
    .Y(_20692_));
 AO21x1_ASAP7_75t_R _29210_ (.A1(net1254),
    .A2(net2435),
    .B(net2982),
    .Y(_20693_));
 AO21x1_ASAP7_75t_R _29211_ (.A1(net1606),
    .A2(net1954),
    .B(net2983),
    .Y(_20694_));
 NAND2x1_ASAP7_75t_R _29212_ (.A(_20693_),
    .B(_20694_),
    .Y(_20695_));
 AO21x1_ASAP7_75t_R _29213_ (.A1(_18381_),
    .A2(net2945),
    .B(net2985),
    .Y(_20696_));
 NAND2x2_ASAP7_75t_R _29214_ (.A(_18343_),
    .B(_18292_),
    .Y(_20697_));
 NAND2x2_ASAP7_75t_R _29215_ (.A(net3283),
    .B(_18292_),
    .Y(_20698_));
 NAND3x2_ASAP7_75t_R _29216_ (.B(_20697_),
    .C(_20698_),
    .Y(_20699_),
    .A(_20696_));
 NOR2x2_ASAP7_75t_R _29217_ (.A(_20695_),
    .B(_20699_),
    .Y(_20700_));
 AO21x1_ASAP7_75t_R _29218_ (.A1(_18381_),
    .A2(net1821),
    .B(_18318_),
    .Y(_20701_));
 NAND2x1_ASAP7_75t_R _29219_ (.A(_20701_),
    .B(_20028_),
    .Y(_20702_));
 AO21x1_ASAP7_75t_R _29220_ (.A1(net2963),
    .A2(net2437),
    .B(_18330_),
    .Y(_20703_));
 OAI21x1_ASAP7_75t_R _29221_ (.A1(net2849),
    .A2(net1702),
    .B(_18345_),
    .Y(_20704_));
 NAND2x1_ASAP7_75t_R _29222_ (.A(_18482_),
    .B(_18345_),
    .Y(_20705_));
 NAND3x1_ASAP7_75t_R _29223_ (.A(_20703_),
    .B(_20704_),
    .C(_20705_),
    .Y(_20706_));
 NOR2x1_ASAP7_75t_R _29224_ (.A(_20702_),
    .B(_20706_),
    .Y(_20707_));
 AOI211x1_ASAP7_75t_R _29225_ (.A1(net1087),
    .A2(_18237_),
    .B(net2970),
    .C(net3246),
    .Y(_20708_));
 INVx1_ASAP7_75t_R _29226_ (.A(_20708_),
    .Y(_20709_));
 AO21x1_ASAP7_75t_R _29227_ (.A1(_19969_),
    .A2(net937),
    .B(net2970),
    .Y(_20710_));
 AO21x1_ASAP7_75t_R _29228_ (.A1(net1254),
    .A2(_18460_),
    .B(net2970),
    .Y(_20711_));
 AND3x2_ASAP7_75t_R _29229_ (.A(_20709_),
    .B(_20710_),
    .C(_20711_),
    .Y(_20712_));
 NAND3x1_ASAP7_75t_R _29230_ (.A(_20700_),
    .B(_20707_),
    .C(_20712_),
    .Y(_20713_));
 AO21x1_ASAP7_75t_R _29231_ (.A1(_18381_),
    .A2(net2452),
    .B(net2981),
    .Y(_20714_));
 AO21x1_ASAP7_75t_R _29232_ (.A1(net1254),
    .A2(net1954),
    .B(net2981),
    .Y(_20715_));
 NAND2x1_ASAP7_75t_R _29233_ (.A(_18291_),
    .B(_19224_),
    .Y(_20716_));
 NAND3x1_ASAP7_75t_R _29234_ (.A(_20714_),
    .B(_20715_),
    .C(_20716_),
    .Y(_20717_));
 AO31x2_ASAP7_75t_R _29235_ (.A1(net2452),
    .A2(net937),
    .A3(net1821),
    .B(_18395_),
    .Y(_20718_));
 AOI21x1_ASAP7_75t_R _29236_ (.A1(net2671),
    .A2(net2969),
    .B(_18395_),
    .Y(_20719_));
 AOI21x1_ASAP7_75t_R _29237_ (.A1(_19223_),
    .A2(_18398_),
    .B(_20719_),
    .Y(_20720_));
 NAND2x1_ASAP7_75t_R _29238_ (.A(_20718_),
    .B(_20720_),
    .Y(_20721_));
 NOR2x1_ASAP7_75t_R _29239_ (.A(_20717_),
    .B(_20721_),
    .Y(_20722_));
 NOR2x1_ASAP7_75t_R _29240_ (.A(_18354_),
    .B(net3003),
    .Y(_20723_));
 NOR3x1_ASAP7_75t_R _29241_ (.A(_19550_),
    .B(_20153_),
    .C(_20723_),
    .Y(_20724_));
 AO21x1_ASAP7_75t_R _29242_ (.A1(net2097),
    .A2(net1954),
    .B(net3178),
    .Y(_20725_));
 AND2x2_ASAP7_75t_R _29243_ (.A(_20724_),
    .B(_20725_),
    .Y(_20726_));
 NOR2x1_ASAP7_75t_R _29244_ (.A(net2011),
    .B(_18364_),
    .Y(_20727_));
 AOI21x1_ASAP7_75t_R _29245_ (.A1(net1959),
    .A2(_19543_),
    .B(_18364_),
    .Y(_20728_));
 NOR2x1_ASAP7_75t_R _29246_ (.A(net2004),
    .B(_18364_),
    .Y(_20729_));
 AOI211x1_ASAP7_75t_R _29247_ (.A1(net1398),
    .A2(_20727_),
    .B(_20728_),
    .C(_20729_),
    .Y(_20730_));
 NAND3x1_ASAP7_75t_R _29248_ (.A(_20722_),
    .B(_20726_),
    .C(_20730_),
    .Y(_20731_));
 NOR2x1_ASAP7_75t_R _29249_ (.A(_20713_),
    .B(_20731_),
    .Y(_20732_));
 NAND2x2_ASAP7_75t_R _29250_ (.A(_20692_),
    .B(_20732_),
    .Y(_20733_));
 NOR2x2_ASAP7_75t_R _29251_ (.A(_20657_),
    .B(_20733_),
    .Y(_20734_));
 OAI21x1_ASAP7_75t_R _29252_ (.A1(_20625_),
    .A2(_20654_),
    .B(_20734_),
    .Y(_20735_));
 AOI22x1_ASAP7_75t_R _29253_ (.A1(_20640_),
    .A2(_17918_),
    .B1(_20623_),
    .B2(_17974_),
    .Y(_20736_));
 NOR2x1_ASAP7_75t_R _29254_ (.A(_20641_),
    .B(_20624_),
    .Y(_20737_));
 INVx1_ASAP7_75t_R _29255_ (.A(_20722_),
    .Y(_20738_));
 NAND2x1_ASAP7_75t_R _29256_ (.A(_20730_),
    .B(_20726_),
    .Y(_20739_));
 NOR2x1_ASAP7_75t_R _29257_ (.A(_20738_),
    .B(_20739_),
    .Y(_20740_));
 INVx1_ASAP7_75t_R _29258_ (.A(_20707_),
    .Y(_20741_));
 NAND2x1_ASAP7_75t_R _29259_ (.A(_20712_),
    .B(_20700_),
    .Y(_20742_));
 NOR2x1_ASAP7_75t_R _29260_ (.A(_20741_),
    .B(_20742_),
    .Y(_20743_));
 NAND2x1_ASAP7_75t_R _29261_ (.A(_20740_),
    .B(_20743_),
    .Y(_20744_));
 INVx1_ASAP7_75t_R _29262_ (.A(_20692_),
    .Y(_20745_));
 NOR2x2_ASAP7_75t_R _29263_ (.A(_20744_),
    .B(_20745_),
    .Y(_20746_));
 NAND2x2_ASAP7_75t_R _29264_ (.A(_18279_),
    .B(_20746_),
    .Y(_20747_));
 OAI21x1_ASAP7_75t_R _29265_ (.A1(_20736_),
    .A2(_20737_),
    .B(_20747_),
    .Y(_20748_));
 NAND2x1_ASAP7_75t_R _29266_ (.A(_20192_),
    .B(_18612_),
    .Y(_20749_));
 AO31x2_ASAP7_75t_R _29267_ (.A1(net2067),
    .A2(_18617_),
    .A3(_18651_),
    .B(net2414),
    .Y(_20750_));
 NAND3x1_ASAP7_75t_R _29268_ (.A(_18616_),
    .B(_20749_),
    .C(_20750_),
    .Y(_20751_));
 NOR2x1_ASAP7_75t_R _29269_ (.A(net2811),
    .B(net2578),
    .Y(_20752_));
 OA21x2_ASAP7_75t_R _29270_ (.A1(_19614_),
    .A2(_18650_),
    .B(_19046_),
    .Y(_20753_));
 NOR2x1_ASAP7_75t_R _29271_ (.A(_20752_),
    .B(_20753_),
    .Y(_20754_));
 AO21x1_ASAP7_75t_R _29272_ (.A1(net1388),
    .A2(_18547_),
    .B(net2579),
    .Y(_20755_));
 NAND3x1_ASAP7_75t_R _29273_ (.A(_20754_),
    .B(_20206_),
    .C(_20755_),
    .Y(_20756_));
 NOR2x1_ASAP7_75t_R _29274_ (.A(_20756_),
    .B(_20751_),
    .Y(_20757_));
 AO21x1_ASAP7_75t_R _29275_ (.A1(net2067),
    .A2(net2052),
    .B(_18625_),
    .Y(_20758_));
 NAND3x1_ASAP7_75t_R _29276_ (.A(_20758_),
    .B(_19632_),
    .C(_19635_),
    .Y(_20759_));
 OA21x2_ASAP7_75t_R _29277_ (.A1(_18537_),
    .A2(_18590_),
    .B(_18635_),
    .Y(_20760_));
 NOR2x1_ASAP7_75t_R _29278_ (.A(_18641_),
    .B(_18553_),
    .Y(_20761_));
 AOI21x1_ASAP7_75t_R _29279_ (.A1(_18687_),
    .A2(net2633),
    .B(_18641_),
    .Y(_20762_));
 OR3x1_ASAP7_75t_R _29280_ (.A(_20760_),
    .B(_20761_),
    .C(_20762_),
    .Y(_20763_));
 NOR2x1_ASAP7_75t_R _29281_ (.A(_20759_),
    .B(_20763_),
    .Y(_20764_));
 AND2x2_ASAP7_75t_R _29282_ (.A(_20764_),
    .B(_20757_),
    .Y(_20765_));
 INVx1_ASAP7_75t_R _29283_ (.A(_20765_),
    .Y(_20766_));
 AO21x1_ASAP7_75t_R _29284_ (.A1(net2052),
    .A2(net2633),
    .B(_18588_),
    .Y(_20767_));
 AO21x1_ASAP7_75t_R _29285_ (.A1(net2177),
    .A2(_18601_),
    .B(_18588_),
    .Y(_20768_));
 NAND2x1_ASAP7_75t_R _29286_ (.A(_18592_),
    .B(_19083_),
    .Y(_20769_));
 NAND3x1_ASAP7_75t_R _29287_ (.A(_20767_),
    .B(_20768_),
    .C(_20769_),
    .Y(_20770_));
 OAI21x1_ASAP7_75t_R _29288_ (.A1(_18569_),
    .A2(_19656_),
    .B(_18577_),
    .Y(_20771_));
 AO21x1_ASAP7_75t_R _29289_ (.A1(_19073_),
    .A2(_18992_),
    .B(_18569_),
    .Y(_20772_));
 OAI21x1_ASAP7_75t_R _29290_ (.A1(_18536_),
    .A2(_18569_),
    .B(_20772_),
    .Y(_20773_));
 NOR3x1_ASAP7_75t_R _29291_ (.A(_20770_),
    .B(_20771_),
    .C(_20773_),
    .Y(_20774_));
 AO21x1_ASAP7_75t_R _29292_ (.A1(_19060_),
    .A2(net2690),
    .B(_19107_),
    .Y(_20775_));
 OA211x2_ASAP7_75t_R _29293_ (.A1(net1472),
    .A2(net3380),
    .B(_18524_),
    .C(net2302),
    .Y(_20776_));
 AOI211x1_ASAP7_75t_R _29294_ (.A1(_19114_),
    .A2(net2690),
    .B(_20775_),
    .C(_20776_),
    .Y(_20777_));
 AO21x1_ASAP7_75t_R _29295_ (.A1(_18528_),
    .A2(net2386),
    .B(_18545_),
    .Y(_20778_));
 AO21x1_ASAP7_75t_R _29296_ (.A1(_18702_),
    .A2(net1965),
    .B(_18545_),
    .Y(_20779_));
 NAND2x1_ASAP7_75t_R _29297_ (.A(_18694_),
    .B(_19664_),
    .Y(_20780_));
 INVx1_ASAP7_75t_R _29298_ (.A(_19701_),
    .Y(_20781_));
 AND4x1_ASAP7_75t_R _29299_ (.A(_20778_),
    .B(_20779_),
    .C(_20780_),
    .D(_20781_),
    .Y(_20782_));
 AND2x2_ASAP7_75t_R _29300_ (.A(_20777_),
    .B(_20782_),
    .Y(_20783_));
 NAND2x1_ASAP7_75t_R _29301_ (.A(_20774_),
    .B(_20783_),
    .Y(_20784_));
 NOR2x1_ASAP7_75t_R _29302_ (.A(_20784_),
    .B(_20766_),
    .Y(_20785_));
 NAND2x1_ASAP7_75t_R _29303_ (.A(_18991_),
    .B(_20213_),
    .Y(_20786_));
 INVx1_ASAP7_75t_R _29304_ (.A(_19601_),
    .Y(_20787_));
 OA21x2_ASAP7_75t_R _29305_ (.A1(_18681_),
    .A2(_18590_),
    .B(_19598_),
    .Y(_20788_));
 OA21x2_ASAP7_75t_R _29306_ (.A1(_18636_),
    .A2(_19614_),
    .B(_19598_),
    .Y(_20789_));
 OR4x1_ASAP7_75t_R _29307_ (.A(_20786_),
    .B(_20787_),
    .C(_20788_),
    .D(_20789_),
    .Y(_20790_));
 AO21x1_ASAP7_75t_R _29308_ (.A1(net2089),
    .A2(net2504),
    .B(_18714_),
    .Y(_20791_));
 AO21x1_ASAP7_75t_R _29309_ (.A1(net3215),
    .A2(net2421),
    .B(_18714_),
    .Y(_20792_));
 AND3x1_ASAP7_75t_R _29310_ (.A(_20791_),
    .B(_20792_),
    .C(_20228_),
    .Y(_20793_));
 INVx1_ASAP7_75t_R _29311_ (.A(_20793_),
    .Y(_20794_));
 AO21x1_ASAP7_75t_R _29312_ (.A1(_18627_),
    .A2(net2421),
    .B(net3324),
    .Y(_20795_));
 OA21x2_ASAP7_75t_R _29313_ (.A1(net1965),
    .A2(net3324),
    .B(_20795_),
    .Y(_20796_));
 NAND2x1_ASAP7_75t_R _29314_ (.A(_18981_),
    .B(_20796_),
    .Y(_20797_));
 NOR3x1_ASAP7_75t_R _29315_ (.A(_20790_),
    .B(_20794_),
    .C(_20797_),
    .Y(_20798_));
 AO21x1_ASAP7_75t_R _29316_ (.A1(net2012),
    .A2(net1825),
    .B(_18655_),
    .Y(_20799_));
 NAND3x1_ASAP7_75t_R _29317_ (.A(_19742_),
    .B(_20250_),
    .C(_20799_),
    .Y(_20800_));
 NOR2x1_ASAP7_75t_R _29318_ (.A(_18666_),
    .B(net2012),
    .Y(_20801_));
 OA211x2_ASAP7_75t_R _29319_ (.A1(net1471),
    .A2(net1734),
    .B(_18671_),
    .C(_18558_),
    .Y(_20802_));
 NOR2x1_ASAP7_75t_R _29320_ (.A(_20801_),
    .B(_20802_),
    .Y(_20803_));
 AND4x1_ASAP7_75t_R _29321_ (.A(_20258_),
    .B(_18676_),
    .C(_19604_),
    .D(_19734_),
    .Y(_20804_));
 NAND2x1_ASAP7_75t_R _29322_ (.A(_20804_),
    .B(_20803_),
    .Y(_20805_));
 NOR2x1_ASAP7_75t_R _29323_ (.A(_20800_),
    .B(_20805_),
    .Y(_20806_));
 AO21x1_ASAP7_75t_R _29324_ (.A1(net3376),
    .A2(net3381),
    .B(net2545),
    .Y(_20807_));
 NAND2x1_ASAP7_75t_R _29325_ (.A(_18583_),
    .B(_18683_),
    .Y(_20808_));
 NAND3x1_ASAP7_75t_R _29326_ (.A(_20807_),
    .B(_20236_),
    .C(_20808_),
    .Y(_20809_));
 INVx1_ASAP7_75t_R _29327_ (.A(_20809_),
    .Y(_20810_));
 NAND2x1_ASAP7_75t_R _29328_ (.A(net1747),
    .B(_18696_),
    .Y(_20811_));
 AND3x1_ASAP7_75t_R _29329_ (.A(_19017_),
    .B(_20811_),
    .C(_18697_),
    .Y(_20812_));
 AO21x1_ASAP7_75t_R _29330_ (.A1(_18621_),
    .A2(net2028),
    .B(net2545),
    .Y(_20813_));
 AND3x1_ASAP7_75t_R _29331_ (.A(_20810_),
    .B(_20812_),
    .C(_20813_),
    .Y(_20814_));
 AND2x2_ASAP7_75t_R _29332_ (.A(_20806_),
    .B(_20814_),
    .Y(_20815_));
 NAND2x2_ASAP7_75t_R _29333_ (.A(_20815_),
    .B(_20798_),
    .Y(_20816_));
 INVx2_ASAP7_75t_R _29334_ (.A(_20816_),
    .Y(_20817_));
 NAND2x2_ASAP7_75t_R _29335_ (.A(_20785_),
    .B(_20817_),
    .Y(_20818_));
 XOR2x1_ASAP7_75t_R _29336_ (.A(_20818_),
    .Y(_20819_),
    .B(_20352_));
 NAND3x1_ASAP7_75t_R _29337_ (.A(_20735_),
    .B(_20748_),
    .C(_20819_),
    .Y(_20820_));
 AO21x1_ASAP7_75t_R _29338_ (.A1(_20735_),
    .A2(_20748_),
    .B(_20819_),
    .Y(_20821_));
 AOI21x1_ASAP7_75t_R _29339_ (.A1(_20820_),
    .A2(_20821_),
    .B(net390),
    .Y(_20822_));
 INVx1_ASAP7_75t_R _29340_ (.A(_20822_),
    .Y(_20823_));
 AOI21x1_ASAP7_75t_R _29341_ (.A1(_20462_),
    .A2(_20823_),
    .B(_00447_),
    .Y(_20824_));
 NOR3x1_ASAP7_75t_R _29342_ (.A(_20822_),
    .B(_14643_),
    .C(_20461_),
    .Y(_20825_));
 NOR2x1_ASAP7_75t_R _29343_ (.A(_20825_),
    .B(_20824_),
    .Y(_00126_));
 OAI21x1_ASAP7_75t_R _29344_ (.A1(net2879),
    .A2(_17605_),
    .B(_17861_),
    .Y(_20826_));
 AO21x1_ASAP7_75t_R _29345_ (.A1(_17834_),
    .A2(_19294_),
    .B(_17614_),
    .Y(_20827_));
 AO21x1_ASAP7_75t_R _29346_ (.A1(_17626_),
    .A2(_17695_),
    .B(_17614_),
    .Y(_20828_));
 NAND2x1_ASAP7_75t_R _29347_ (.A(_20827_),
    .B(_20828_),
    .Y(_20829_));
 AO21x1_ASAP7_75t_R _29348_ (.A1(net2630),
    .A2(_17538_),
    .B(_17589_),
    .Y(_20830_));
 AO21x1_ASAP7_75t_R _29349_ (.A1(_17639_),
    .A2(net1789),
    .B(_17589_),
    .Y(_20831_));
 NAND2x1_ASAP7_75t_R _29350_ (.A(_20830_),
    .B(_20831_),
    .Y(_20832_));
 NOR3x1_ASAP7_75t_R _29351_ (.A(_20826_),
    .B(_20829_),
    .C(_20832_),
    .Y(_20833_));
 AOI211x1_ASAP7_75t_R _29352_ (.A1(net2862),
    .A2(net1185),
    .B(_17566_),
    .C(net1103),
    .Y(_20834_));
 INVx1_ASAP7_75t_R _29353_ (.A(_20834_),
    .Y(_20835_));
 AO21x1_ASAP7_75t_R _29354_ (.A1(net2904),
    .A2(_17538_),
    .B(_17566_),
    .Y(_20836_));
 AO21x1_ASAP7_75t_R _29355_ (.A1(net936),
    .A2(net2202),
    .B(_17566_),
    .Y(_20837_));
 NAND3x1_ASAP7_75t_R _29356_ (.A(_20835_),
    .B(_20836_),
    .C(_20837_),
    .Y(_20838_));
 AND2x2_ASAP7_75t_R _29357_ (.A(_18766_),
    .B(_20519_),
    .Y(_20839_));
 AND2x2_ASAP7_75t_R _29358_ (.A(_19954_),
    .B(_17870_),
    .Y(_20840_));
 NAND2x1_ASAP7_75t_R _29359_ (.A(_20839_),
    .B(_20840_),
    .Y(_20841_));
 NOR2x1_ASAP7_75t_R _29360_ (.A(_20838_),
    .B(_20841_),
    .Y(_20842_));
 NAND2x1_ASAP7_75t_R _29361_ (.A(_20833_),
    .B(_20842_),
    .Y(_20843_));
 AO21x1_ASAP7_75t_R _29362_ (.A1(_17639_),
    .A2(net3193),
    .B(net2484),
    .Y(_20844_));
 AOI211x1_ASAP7_75t_R _29363_ (.A1(net1123),
    .A2(net1189),
    .B(net2484),
    .C(net1977),
    .Y(_20845_));
 INVx1_ASAP7_75t_R _29364_ (.A(_20845_),
    .Y(_20846_));
 NAND2x1_ASAP7_75t_R _29365_ (.A(_20844_),
    .B(_20846_),
    .Y(_20847_));
 AO21x1_ASAP7_75t_R _29366_ (.A1(net1082),
    .A2(_19294_),
    .B(_17629_),
    .Y(_20848_));
 INVx1_ASAP7_75t_R _29367_ (.A(_17636_),
    .Y(_20849_));
 NAND3x2_ASAP7_75t_R _29368_ (.B(_20848_),
    .C(_20849_),
    .Y(_20850_),
    .A(_20524_));
 NOR2x2_ASAP7_75t_R _29369_ (.A(_20850_),
    .B(_20847_),
    .Y(_20851_));
 AO21x1_ASAP7_75t_R _29370_ (.A1(net936),
    .A2(_17756_),
    .B(net2889),
    .Y(_20852_));
 AO21x1_ASAP7_75t_R _29371_ (.A1(_17626_),
    .A2(net2900),
    .B(net2889),
    .Y(_20853_));
 NAND2x1_ASAP7_75t_R _29372_ (.A(_20852_),
    .B(_20853_),
    .Y(_20854_));
 AO21x1_ASAP7_75t_R _29373_ (.A1(_17639_),
    .A2(net1789),
    .B(net2889),
    .Y(_20855_));
 OAI21x1_ASAP7_75t_R _29374_ (.A1(net3193),
    .A2(net2889),
    .B(_20855_),
    .Y(_20856_));
 NOR2x1_ASAP7_75t_R _29375_ (.A(_20854_),
    .B(_20856_),
    .Y(_20857_));
 AO21x1_ASAP7_75t_R _29376_ (.A1(_17845_),
    .A2(net941),
    .B(net2847),
    .Y(_20858_));
 AO21x1_ASAP7_75t_R _29377_ (.A1(net1789),
    .A2(_17834_),
    .B(net2847),
    .Y(_20859_));
 NAND2x1_ASAP7_75t_R _29378_ (.A(_17576_),
    .B(_17662_),
    .Y(_20860_));
 AND3x1_ASAP7_75t_R _29379_ (.A(_20858_),
    .B(_20859_),
    .C(_20860_),
    .Y(_20861_));
 AND2x2_ASAP7_75t_R _29380_ (.A(_20857_),
    .B(_20861_),
    .Y(_20862_));
 NAND2x2_ASAP7_75t_R _29381_ (.A(_20851_),
    .B(_20862_),
    .Y(_20863_));
 NOR2x2_ASAP7_75t_R _29382_ (.A(_20843_),
    .B(_20863_),
    .Y(_20864_));
 AO21x1_ASAP7_75t_R _29383_ (.A1(_17834_),
    .A2(_17575_),
    .B(_17744_),
    .Y(_20865_));
 INVx1_ASAP7_75t_R _29384_ (.A(_17747_),
    .Y(_20866_));
 NAND3x2_ASAP7_75t_R _29385_ (.B(_20865_),
    .C(_20866_),
    .Y(_20867_),
    .A(_19888_));
 AO21x1_ASAP7_75t_R _29386_ (.A1(net936),
    .A2(net2202),
    .B(_17759_),
    .Y(_20868_));
 AO21x1_ASAP7_75t_R _29387_ (.A1(_17639_),
    .A2(net2237),
    .B(_17759_),
    .Y(_20869_));
 NAND2x2_ASAP7_75t_R _29388_ (.A(_18825_),
    .B(_17678_),
    .Y(_20870_));
 NAND3x2_ASAP7_75t_R _29389_ (.B(_20869_),
    .C(_20870_),
    .Y(_20871_),
    .A(_20868_));
 NOR2x2_ASAP7_75t_R _29390_ (.A(_20867_),
    .B(_20871_),
    .Y(_20872_));
 AO21x1_ASAP7_75t_R _29391_ (.A1(_17758_),
    .A2(net2899),
    .B(_17777_),
    .Y(_20873_));
 NAND2x1_ASAP7_75t_R _29392_ (.A(_17787_),
    .B(_20873_),
    .Y(_20874_));
 AO21x1_ASAP7_75t_R _29393_ (.A1(_17576_),
    .A2(_17782_),
    .B(_17783_),
    .Y(_20875_));
 NOR2x2_ASAP7_75t_R _29394_ (.A(_20874_),
    .B(_20875_),
    .Y(_20876_));
 AO21x1_ASAP7_75t_R _29395_ (.A1(_17626_),
    .A2(net2451),
    .B(_17770_),
    .Y(_20877_));
 OAI21x1_ASAP7_75t_R _29396_ (.A1(net2909),
    .A2(net941),
    .B(_20877_),
    .Y(_20878_));
 OAI21x1_ASAP7_75t_R _29397_ (.A1(net2909),
    .A2(net1097),
    .B(_17836_),
    .Y(_20879_));
 NOR2x2_ASAP7_75t_R _29398_ (.A(_20878_),
    .B(_20879_),
    .Y(_20880_));
 NAND3x2_ASAP7_75t_R _29399_ (.B(_20876_),
    .C(_20880_),
    .Y(_20881_),
    .A(_20872_));
 AO21x1_ASAP7_75t_R _29400_ (.A1(net1081),
    .A2(_17551_),
    .B(_17691_),
    .Y(_20882_));
 OAI21x1_ASAP7_75t_R _29401_ (.A1(net2893),
    .A2(_17691_),
    .B(_20882_),
    .Y(_20883_));
 INVx1_ASAP7_75t_R _29402_ (.A(_17692_),
    .Y(_20884_));
 NAND2x1_ASAP7_75t_R _29403_ (.A(_20884_),
    .B(_20494_),
    .Y(_20885_));
 AOI211x1_ASAP7_75t_R _29404_ (.A1(_17801_),
    .A2(_17573_),
    .B(_20883_),
    .C(_20885_),
    .Y(_20886_));
 AO21x1_ASAP7_75t_R _29405_ (.A1(_17813_),
    .A2(net2630),
    .B(_17712_),
    .Y(_20887_));
 NAND2x2_ASAP7_75t_R _29406_ (.A(_17661_),
    .B(_17714_),
    .Y(_20888_));
 NAND3x2_ASAP7_75t_R _29407_ (.B(_17810_),
    .C(_20888_),
    .Y(_20889_),
    .A(_20887_));
 AO21x1_ASAP7_75t_R _29408_ (.A1(net936),
    .A2(net941),
    .B(_17725_),
    .Y(_20890_));
 AO21x1_ASAP7_75t_R _29409_ (.A1(_17647_),
    .A2(_17538_),
    .B(_17725_),
    .Y(_20891_));
 NAND3x2_ASAP7_75t_R _29410_ (.B(_20891_),
    .C(_19876_),
    .Y(_20892_),
    .A(_20890_));
 NOR2x2_ASAP7_75t_R _29411_ (.A(_20889_),
    .B(_20892_),
    .Y(_20893_));
 INVx1_ASAP7_75t_R _29412_ (.A(_19295_),
    .Y(_20894_));
 NOR2x2_ASAP7_75t_R _29413_ (.A(_20894_),
    .B(_17913_),
    .Y(_20895_));
 NAND3x2_ASAP7_75t_R _29414_ (.B(_20893_),
    .C(_20895_),
    .Y(_20896_),
    .A(_20886_));
 NOR2x2_ASAP7_75t_R _29415_ (.A(_20881_),
    .B(_20896_),
    .Y(_20897_));
 NAND2x2_ASAP7_75t_R _29416_ (.A(_20864_),
    .B(_20897_),
    .Y(_20898_));
 NOR2x2_ASAP7_75t_R _29417_ (.A(net2143),
    .B(_20898_),
    .Y(_20899_));
 AO21x1_ASAP7_75t_R _29418_ (.A1(net3184),
    .A2(net1348),
    .B(net3205),
    .Y(_20900_));
 AO21x1_ASAP7_75t_R _29419_ (.A1(_18147_),
    .A2(_18081_),
    .B(_17977_),
    .Y(_20901_));
 AO21x1_ASAP7_75t_R _29420_ (.A1(_18002_),
    .A2(net1367),
    .B(_17977_),
    .Y(_20902_));
 AND3x1_ASAP7_75t_R _29421_ (.A(_20900_),
    .B(_20901_),
    .C(_20902_),
    .Y(_20903_));
 AO21x1_ASAP7_75t_R _29422_ (.A1(_18931_),
    .A2(_18958_),
    .B(_17997_),
    .Y(_20904_));
 NAND2x1_ASAP7_75t_R _29423_ (.A(_19802_),
    .B(_18006_),
    .Y(_20905_));
 AND3x1_ASAP7_75t_R _29424_ (.A(_19861_),
    .B(_20904_),
    .C(_20905_),
    .Y(_20906_));
 AND2x2_ASAP7_75t_R _29425_ (.A(_20903_),
    .B(_20906_),
    .Y(_20907_));
 AO21x1_ASAP7_75t_R _29426_ (.A1(net1675),
    .A2(_18881_),
    .B(_18024_),
    .Y(_20908_));
 INVx1_ASAP7_75t_R _29427_ (.A(_18922_),
    .Y(_20909_));
 NAND3x1_ASAP7_75t_R _29428_ (.A(_20908_),
    .B(_19363_),
    .C(_20909_),
    .Y(_20910_));
 NAND2x1_ASAP7_75t_R _29429_ (.A(net1815),
    .B(net2718),
    .Y(_20911_));
 AO21x1_ASAP7_75t_R _29430_ (.A1(_18883_),
    .A2(_20911_),
    .B(_18012_),
    .Y(_20912_));
 NAND3x1_ASAP7_75t_R _29431_ (.A(_20912_),
    .B(_19359_),
    .C(_20550_),
    .Y(_20913_));
 OAI21x1_ASAP7_75t_R _29432_ (.A1(_19802_),
    .A2(_18900_),
    .B(_18020_),
    .Y(_20914_));
 OAI21x1_ASAP7_75t_R _29433_ (.A1(net3124),
    .A2(_18027_),
    .B(_20914_),
    .Y(_20915_));
 NOR3x1_ASAP7_75t_R _29434_ (.A(_20910_),
    .B(_20913_),
    .C(_20915_),
    .Y(_20916_));
 NAND2x1_ASAP7_75t_R _29435_ (.A(_20907_),
    .B(_20916_),
    .Y(_20917_));
 NOR2x1_ASAP7_75t_R _29436_ (.A(_19832_),
    .B(_19395_),
    .Y(_20918_));
 AOI211x1_ASAP7_75t_R _29437_ (.A1(net1061),
    .A2(net1117),
    .B(net1907),
    .C(net2057),
    .Y(_20919_));
 OA21x2_ASAP7_75t_R _29438_ (.A1(net2792),
    .A2(_18134_),
    .B(_18069_),
    .Y(_20920_));
 NOR2x1_ASAP7_75t_R _29439_ (.A(_20919_),
    .B(_20920_),
    .Y(_20921_));
 AO21x1_ASAP7_75t_R _29440_ (.A1(_18147_),
    .A2(_17987_),
    .B(net2181),
    .Y(_20922_));
 AND3x1_ASAP7_75t_R _29441_ (.A(_20918_),
    .B(_20921_),
    .C(_20922_),
    .Y(_20923_));
 OA21x2_ASAP7_75t_R _29442_ (.A1(net2877),
    .A2(net1857),
    .B(_18040_),
    .Y(_20924_));
 OA21x2_ASAP7_75t_R _29443_ (.A1(_18923_),
    .A2(_18869_),
    .B(_18040_),
    .Y(_20925_));
 NOR2x1_ASAP7_75t_R _29444_ (.A(_18039_),
    .B(_17980_),
    .Y(_20926_));
 OR3x1_ASAP7_75t_R _29445_ (.A(_20924_),
    .B(_20925_),
    .C(_20926_),
    .Y(_20927_));
 AOI22x1_ASAP7_75t_R _29446_ (.A1(_18061_),
    .A2(net1117),
    .B1(_18952_),
    .B2(net2792),
    .Y(_20928_));
 AO21x1_ASAP7_75t_R _29447_ (.A1(net3300),
    .A2(net2757),
    .B(_18054_),
    .Y(_20929_));
 AO21x1_ASAP7_75t_R _29448_ (.A1(net2821),
    .A2(net939),
    .B(_18054_),
    .Y(_20930_));
 NAND3x1_ASAP7_75t_R _29449_ (.A(_20928_),
    .B(_20929_),
    .C(_20930_),
    .Y(_20931_));
 NOR2x1_ASAP7_75t_R _29450_ (.A(_20927_),
    .B(_20931_),
    .Y(_20932_));
 NAND2x1_ASAP7_75t_R _29451_ (.A(_20923_),
    .B(_20932_),
    .Y(_20933_));
 NOR2x2_ASAP7_75t_R _29452_ (.A(_20917_),
    .B(_20933_),
    .Y(_20934_));
 AO21x1_ASAP7_75t_R _29453_ (.A1(_18883_),
    .A2(_17947_),
    .B(net2446),
    .Y(_20935_));
 NAND3x2_ASAP7_75t_R _29454_ (.B(_18149_),
    .C(_20935_),
    .Y(_20936_),
    .A(_19805_));
 AO21x1_ASAP7_75t_R _29455_ (.A1(net3188),
    .A2(net1839),
    .B(_18156_),
    .Y(_20937_));
 NAND2x2_ASAP7_75t_R _29456_ (.A(net2162),
    .B(net3202),
    .Y(_20938_));
 OAI21x1_ASAP7_75t_R _29457_ (.A1(_18134_),
    .A2(_18923_),
    .B(net2162),
    .Y(_20939_));
 NAND3x2_ASAP7_75t_R _29458_ (.B(_20938_),
    .C(_20939_),
    .Y(_20940_),
    .A(_20937_));
 NOR2x2_ASAP7_75t_R _29459_ (.A(_20936_),
    .B(_20940_),
    .Y(_20941_));
 AO21x1_ASAP7_75t_R _29460_ (.A1(_18147_),
    .A2(net2757),
    .B(_19423_),
    .Y(_20942_));
 NAND2x1_ASAP7_75t_R _29461_ (.A(net2244),
    .B(net3367),
    .Y(_20943_));
 AND4x2_ASAP7_75t_R _29462_ (.A(_20942_),
    .B(_20943_),
    .C(_18177_),
    .D(_18183_),
    .Y(_20944_));
 AO21x1_ASAP7_75t_R _29463_ (.A1(_18028_),
    .A2(_18010_),
    .B(_18169_),
    .Y(_20945_));
 OAI21x1_ASAP7_75t_R _29464_ (.A1(net974),
    .A2(_18169_),
    .B(_20945_),
    .Y(_20946_));
 OAI21x1_ASAP7_75t_R _29465_ (.A1(net3212),
    .A2(_18169_),
    .B(_18905_),
    .Y(_20947_));
 NOR2x2_ASAP7_75t_R _29466_ (.A(_20946_),
    .B(_20947_),
    .Y(_20948_));
 NAND3x2_ASAP7_75t_R _29467_ (.B(_20944_),
    .C(_20948_),
    .Y(_20949_),
    .A(_20941_));
 OA21x2_ASAP7_75t_R _29468_ (.A1(_18000_),
    .A2(_18130_),
    .B(_18123_),
    .Y(_20950_));
 OA21x2_ASAP7_75t_R _29469_ (.A1(_18900_),
    .A2(_18901_),
    .B(_18123_),
    .Y(_20951_));
 NOR2x1_ASAP7_75t_R _29470_ (.A(_18022_),
    .B(_18126_),
    .Y(_20952_));
 OR3x1_ASAP7_75t_R _29471_ (.A(_20950_),
    .B(_20951_),
    .C(_20952_),
    .Y(_20953_));
 AOI22x1_ASAP7_75t_R _29472_ (.A1(_18118_),
    .A2(net1057),
    .B1(net2680),
    .B2(_17925_),
    .Y(_20954_));
 AO21x1_ASAP7_75t_R _29473_ (.A1(net2944),
    .A2(_17958_),
    .B(_18864_),
    .Y(_20955_));
 NAND3x1_ASAP7_75t_R _29474_ (.A(_20954_),
    .B(_19767_),
    .C(_20955_),
    .Y(_20956_));
 NOR2x1_ASAP7_75t_R _29475_ (.A(_20953_),
    .B(_20956_),
    .Y(_20957_));
 AO21x1_ASAP7_75t_R _29476_ (.A1(_17984_),
    .A2(_17951_),
    .B(net2364),
    .Y(_20958_));
 AO21x1_ASAP7_75t_R _29477_ (.A1(net3307),
    .A2(_18958_),
    .B(net2364),
    .Y(_20959_));
 NAND2x1_ASAP7_75t_R _29478_ (.A(_20958_),
    .B(_20959_),
    .Y(_20960_));
 OA21x2_ASAP7_75t_R _29479_ (.A1(net3213),
    .A2(net1746),
    .B(_20403_),
    .Y(_20961_));
 NAND2x1_ASAP7_75t_R _29480_ (.A(_17965_),
    .B(_20961_),
    .Y(_20962_));
 NOR2x1_ASAP7_75t_R _29481_ (.A(_20960_),
    .B(_20962_),
    .Y(_20963_));
 NAND2x1_ASAP7_75t_R _29482_ (.A(_20957_),
    .B(_20963_),
    .Y(_20964_));
 NOR2x2_ASAP7_75t_R _29483_ (.A(_20949_),
    .B(_20964_),
    .Y(_20965_));
 NAND2x2_ASAP7_75t_R _29484_ (.A(_20934_),
    .B(_20965_),
    .Y(_20966_));
 NOR2x2_ASAP7_75t_R _29485_ (.A(_20642_),
    .B(_20966_),
    .Y(_20967_));
 NAND2x1_ASAP7_75t_R _29486_ (.A(_20899_),
    .B(_20967_),
    .Y(_20968_));
 OAI22x1_ASAP7_75t_R _29487_ (.A1(_20966_),
    .A2(_20642_),
    .B1(_20898_),
    .B2(net2143),
    .Y(_20969_));
 AO21x1_ASAP7_75t_R _29488_ (.A1(_19969_),
    .A2(net2499),
    .B(_18266_),
    .Y(_20970_));
 AO21x1_ASAP7_75t_R _29489_ (.A1(net2176),
    .A2(_18335_),
    .B(_18266_),
    .Y(_20971_));
 AND2x2_ASAP7_75t_R _29490_ (.A(_20970_),
    .B(_20971_),
    .Y(_20972_));
 NAND3x1_ASAP7_75t_R _29491_ (.A(_20972_),
    .B(_18274_),
    .C(_19484_),
    .Y(_20973_));
 AO21x1_ASAP7_75t_R _29492_ (.A1(net2963),
    .A2(net2437),
    .B(_18428_),
    .Y(_20974_));
 NAND2x1_ASAP7_75t_R _29493_ (.A(_18468_),
    .B(_18434_),
    .Y(_20975_));
 NOR2x1_ASAP7_75t_R _29494_ (.A(_18428_),
    .B(_19174_),
    .Y(_20976_));
 INVx1_ASAP7_75t_R _29495_ (.A(_20976_),
    .Y(_20977_));
 AND3x1_ASAP7_75t_R _29496_ (.A(_20974_),
    .B(_20975_),
    .C(_20977_),
    .Y(_20978_));
 AO21x2_ASAP7_75t_R _29497_ (.A1(net2701),
    .A2(net1482),
    .B(_18439_),
    .Y(_20979_));
 AO21x1_ASAP7_75t_R _29498_ (.A1(_18350_),
    .A2(_18460_),
    .B(net2989),
    .Y(_20980_));
 INVx1_ASAP7_75t_R _29499_ (.A(_19995_),
    .Y(_20981_));
 AND3x1_ASAP7_75t_R _29500_ (.A(_20979_),
    .B(_20980_),
    .C(_20981_),
    .Y(_20982_));
 NAND2x1_ASAP7_75t_R _29501_ (.A(_20978_),
    .B(_20982_),
    .Y(_20983_));
 NOR2x1_ASAP7_75t_R _29502_ (.A(_20973_),
    .B(_20983_),
    .Y(_20984_));
 AO21x1_ASAP7_75t_R _29503_ (.A1(net2699),
    .A2(net2251),
    .B(_18456_),
    .Y(_20985_));
 AO21x1_ASAP7_75t_R _29504_ (.A1(_18402_),
    .A2(net1606),
    .B(_18456_),
    .Y(_20986_));
 NAND2x1_ASAP7_75t_R _29505_ (.A(_19465_),
    .B(_19185_),
    .Y(_20987_));
 AND3x1_ASAP7_75t_R _29506_ (.A(_20985_),
    .B(_20986_),
    .C(_20987_),
    .Y(_20988_));
 NAND2x1_ASAP7_75t_R _29507_ (.A(_18474_),
    .B(_19964_),
    .Y(_20989_));
 OA211x2_ASAP7_75t_R _29508_ (.A1(_18280_),
    .A2(net1087),
    .B(_18469_),
    .C(net2980),
    .Y(_20990_));
 NOR2x1_ASAP7_75t_R _29509_ (.A(_20989_),
    .B(_20990_),
    .Y(_20991_));
 NAND2x1_ASAP7_75t_R _29510_ (.A(_20988_),
    .B(_20991_),
    .Y(_20992_));
 NOR2x1_ASAP7_75t_R _29511_ (.A(_18490_),
    .B(net2250),
    .Y(_20993_));
 AO21x1_ASAP7_75t_R _29512_ (.A1(_19170_),
    .A2(net2971),
    .B(_20993_),
    .Y(_20994_));
 NAND2x1_ASAP7_75t_R _29513_ (.A(_19156_),
    .B(_19472_),
    .Y(_20995_));
 AO21x1_ASAP7_75t_R _29514_ (.A1(_18381_),
    .A2(net2043),
    .B(net2595),
    .Y(_20996_));
 NAND2x1_ASAP7_75t_R _29515_ (.A(_20995_),
    .B(_20996_),
    .Y(_20997_));
 NOR2x2_ASAP7_75t_R _29516_ (.A(_20994_),
    .B(_20997_),
    .Y(_20998_));
 AO21x1_ASAP7_75t_R _29517_ (.A1(net2638),
    .A2(net3003),
    .B(net3282),
    .Y(_20999_));
 AND2x2_ASAP7_75t_R _29518_ (.A(_20999_),
    .B(_18486_),
    .Y(_21000_));
 AOI21x1_ASAP7_75t_R _29519_ (.A1(_18306_),
    .A2(_18483_),
    .B(_18499_),
    .Y(_21001_));
 NAND3x2_ASAP7_75t_R _29520_ (.B(_21000_),
    .C(_21001_),
    .Y(_21002_),
    .A(_20998_));
 NOR2x2_ASAP7_75t_R _29521_ (.A(_20992_),
    .B(_21002_),
    .Y(_21003_));
 NAND2x2_ASAP7_75t_R _29522_ (.A(_20984_),
    .B(_21003_),
    .Y(_21004_));
 AO21x1_ASAP7_75t_R _29523_ (.A1(net2452),
    .A2(net937),
    .B(_18364_),
    .Y(_21005_));
 AO21x1_ASAP7_75t_R _29524_ (.A1(net1606),
    .A2(net2095),
    .B(_18364_),
    .Y(_21006_));
 NAND2x1_ASAP7_75t_R _29525_ (.A(_18306_),
    .B(_18371_),
    .Y(_21007_));
 AND3x1_ASAP7_75t_R _29526_ (.A(_21005_),
    .B(_21006_),
    .C(_21007_),
    .Y(_21008_));
 AO21x1_ASAP7_75t_R _29527_ (.A1(_18381_),
    .A2(net3182),
    .B(_18354_),
    .Y(_21009_));
 AO21x1_ASAP7_75t_R _29528_ (.A1(net1335),
    .A2(net2967),
    .B(net3178),
    .Y(_21010_));
 NAND2x1_ASAP7_75t_R _29529_ (.A(_21009_),
    .B(_21010_),
    .Y(_21011_));
 AO21x1_ASAP7_75t_R _29530_ (.A1(_18402_),
    .A2(net2250),
    .B(_18354_),
    .Y(_21012_));
 OAI21x1_ASAP7_75t_R _29531_ (.A1(net2004),
    .A2(net3178),
    .B(_21012_),
    .Y(_21013_));
 NOR2x1_ASAP7_75t_R _29532_ (.A(_21011_),
    .B(_21013_),
    .Y(_21014_));
 NAND2x1_ASAP7_75t_R _29533_ (.A(_21008_),
    .B(_21014_),
    .Y(_21015_));
 AO21x1_ASAP7_75t_R _29534_ (.A1(net1954),
    .A2(net2788),
    .B(net2981),
    .Y(_21016_));
 AND3x1_ASAP7_75t_R _29535_ (.A(_20714_),
    .B(_18380_),
    .C(_21016_),
    .Y(_21017_));
 OA21x2_ASAP7_75t_R _29536_ (.A1(_19465_),
    .A2(_18257_),
    .B(_18398_),
    .Y(_21018_));
 OA211x2_ASAP7_75t_R _29537_ (.A1(net2999),
    .A2(_18237_),
    .B(_18398_),
    .C(_18272_),
    .Y(_21019_));
 NOR2x1_ASAP7_75t_R _29538_ (.A(_21018_),
    .B(_21019_),
    .Y(_21020_));
 NAND2x1_ASAP7_75t_R _29539_ (.A(_21017_),
    .B(_21020_),
    .Y(_21021_));
 NOR2x1_ASAP7_75t_R _29540_ (.A(_21015_),
    .B(_21021_),
    .Y(_21022_));
 AOI211x1_ASAP7_75t_R _29541_ (.A1(net2999),
    .A2(net2990),
    .B(net1579),
    .C(_18300_),
    .Y(_21023_));
 INVx1_ASAP7_75t_R _29542_ (.A(_21023_),
    .Y(_21024_));
 AO21x1_ASAP7_75t_R _29543_ (.A1(_18460_),
    .A2(net2010),
    .B(net2970),
    .Y(_21025_));
 AO21x1_ASAP7_75t_R _29544_ (.A1(net2634),
    .A2(net1335),
    .B(net2970),
    .Y(_21026_));
 AND3x1_ASAP7_75t_R _29545_ (.A(_21024_),
    .B(_21025_),
    .C(_21026_),
    .Y(_21027_));
 NAND2x1_ASAP7_75t_R _29546_ (.A(_20693_),
    .B(_19211_),
    .Y(_21028_));
 NAND2x2_ASAP7_75t_R _29547_ (.A(_18344_),
    .B(_18292_),
    .Y(_21029_));
 INVx1_ASAP7_75t_R _29548_ (.A(_21029_),
    .Y(_21030_));
 NOR3x1_ASAP7_75t_R _29549_ (.A(_21028_),
    .B(_20033_),
    .C(_21030_),
    .Y(_21031_));
 NAND2x1_ASAP7_75t_R _29550_ (.A(_21027_),
    .B(_21031_),
    .Y(_21032_));
 AO21x1_ASAP7_75t_R _29551_ (.A1(_18402_),
    .A2(net1606),
    .B(_18330_),
    .Y(_21033_));
 AO21x1_ASAP7_75t_R _29552_ (.A1(net2963),
    .A2(net2004),
    .B(_18330_),
    .Y(_21034_));
 AND3x1_ASAP7_75t_R _29553_ (.A(_21033_),
    .B(_21034_),
    .C(_19203_),
    .Y(_21035_));
 AO21x1_ASAP7_75t_R _29554_ (.A1(net1335),
    .A2(net2966),
    .B(_18330_),
    .Y(_21036_));
 AO21x1_ASAP7_75t_R _29555_ (.A1(_18381_),
    .A2(_18383_),
    .B(_18330_),
    .Y(_21037_));
 AND2x2_ASAP7_75t_R _29556_ (.A(_21036_),
    .B(_21037_),
    .Y(_21038_));
 AO21x1_ASAP7_75t_R _29557_ (.A1(_18381_),
    .A2(_18394_),
    .B(_18318_),
    .Y(_21039_));
 AO21x1_ASAP7_75t_R _29558_ (.A1(net2095),
    .A2(net2788),
    .B(_18318_),
    .Y(_21040_));
 AND2x2_ASAP7_75t_R _29559_ (.A(_21039_),
    .B(_21040_),
    .Y(_21041_));
 NAND3x1_ASAP7_75t_R _29560_ (.A(_21035_),
    .B(_21038_),
    .C(_21041_),
    .Y(_21042_));
 NOR2x1_ASAP7_75t_R _29561_ (.A(_21032_),
    .B(_21042_),
    .Y(_21043_));
 NAND2x1_ASAP7_75t_R _29562_ (.A(_21022_),
    .B(_21043_),
    .Y(_21044_));
 NOR2x2_ASAP7_75t_R _29563_ (.A(_21004_),
    .B(_21044_),
    .Y(_21045_));
 NAND2x2_ASAP7_75t_R _29564_ (.A(_18279_),
    .B(_21045_),
    .Y(_21046_));
 INVx1_ASAP7_75t_R _29565_ (.A(_21046_),
    .Y(_21047_));
 AO21x1_ASAP7_75t_R _29566_ (.A1(_20968_),
    .A2(_20969_),
    .B(_21047_),
    .Y(_21048_));
 XOR2x1_ASAP7_75t_R _29567_ (.A(_20967_),
    .Y(_21049_),
    .B(_20899_));
 NAND2x1_ASAP7_75t_R _29568_ (.A(_21047_),
    .B(_21049_),
    .Y(_21050_));
 AO21x1_ASAP7_75t_R _29569_ (.A1(_18547_),
    .A2(_18601_),
    .B(_18588_),
    .Y(_21051_));
 NAND2x2_ASAP7_75t_R _29570_ (.A(_18592_),
    .B(_18675_),
    .Y(_21052_));
 NAND2x1_ASAP7_75t_R _29571_ (.A(net2991),
    .B(_18592_),
    .Y(_21053_));
 AND3x1_ASAP7_75t_R _29572_ (.A(_21051_),
    .B(_21052_),
    .C(_21053_),
    .Y(_21054_));
 INVx1_ASAP7_75t_R _29573_ (.A(_19036_),
    .Y(_21055_));
 AOI211x1_ASAP7_75t_R _29574_ (.A1(_18564_),
    .A2(net3380),
    .B(_18569_),
    .C(net3007),
    .Y(_21056_));
 AOI211x1_ASAP7_75t_R _29575_ (.A1(_18570_),
    .A2(_21055_),
    .B(_21056_),
    .C(_19657_),
    .Y(_21057_));
 NAND2x1_ASAP7_75t_R _29576_ (.A(_21054_),
    .B(_21057_),
    .Y(_21058_));
 NAND2x1_ASAP7_75t_R _29577_ (.A(_19668_),
    .B(net2776),
    .Y(_21059_));
 NOR2x1_ASAP7_75t_R _29578_ (.A(_19107_),
    .B(_21059_),
    .Y(_21060_));
 AO221x1_ASAP7_75t_R _29579_ (.A1(net1472),
    .A2(net3380),
    .B1(net1565),
    .B2(_18536_),
    .C(_18525_),
    .Y(_21061_));
 NAND2x1_ASAP7_75t_R _29580_ (.A(_21060_),
    .B(_21061_),
    .Y(_21062_));
 AO21x1_ASAP7_75t_R _29581_ (.A1(_18674_),
    .A2(net1069),
    .B(net2631),
    .Y(_21063_));
 AO21x1_ASAP7_75t_R _29582_ (.A1(_21063_),
    .A2(net2405),
    .B(net2479),
    .Y(_21064_));
 AO21x1_ASAP7_75t_R _29583_ (.A1(_19073_),
    .A2(_18623_),
    .B(net2479),
    .Y(_21065_));
 AO21x1_ASAP7_75t_R _29584_ (.A1(net1307),
    .A2(net1388),
    .B(net2479),
    .Y(_21066_));
 NAND3x1_ASAP7_75t_R _29585_ (.A(_21064_),
    .B(_21065_),
    .C(_21066_),
    .Y(_21067_));
 NOR3x1_ASAP7_75t_R _29586_ (.A(_21058_),
    .B(_21062_),
    .C(_21067_),
    .Y(_21068_));
 OA21x2_ASAP7_75t_R _29587_ (.A1(_18590_),
    .A2(_19114_),
    .B(_18635_),
    .Y(_21069_));
 AOI211x1_ASAP7_75t_R _29588_ (.A1(net3090),
    .A2(net3380),
    .B(_18641_),
    .C(net2631),
    .Y(_21070_));
 AOI211x1_ASAP7_75t_R _29589_ (.A1(_18635_),
    .A2(_19614_),
    .B(_21069_),
    .C(_21070_),
    .Y(_21071_));
 AO21x1_ASAP7_75t_R _29590_ (.A1(net2633),
    .A2(net1965),
    .B(_18625_),
    .Y(_21072_));
 AND3x1_ASAP7_75t_R _29591_ (.A(_19067_),
    .B(_20180_),
    .C(_21072_),
    .Y(_21073_));
 NAND2x1_ASAP7_75t_R _29592_ (.A(_21071_),
    .B(_21073_),
    .Y(_21074_));
 AO21x1_ASAP7_75t_R _29593_ (.A1(net2028),
    .A2(_18992_),
    .B(net2414),
    .Y(_21075_));
 NAND2x1_ASAP7_75t_R _29594_ (.A(_19040_),
    .B(_21075_),
    .Y(_21076_));
 AO21x1_ASAP7_75t_R _29595_ (.A1(net2811),
    .A2(net1966),
    .B(net2415),
    .Y(_21077_));
 OAI21x1_ASAP7_75t_R _29596_ (.A1(_18627_),
    .A2(net2415),
    .B(_21077_),
    .Y(_21078_));
 NOR2x2_ASAP7_75t_R _29597_ (.A(_21076_),
    .B(_21078_),
    .Y(_21079_));
 AO21x1_ASAP7_75t_R _29598_ (.A1(net1307),
    .A2(_18548_),
    .B(net2579),
    .Y(_21080_));
 AND2x2_ASAP7_75t_R _29599_ (.A(_20206_),
    .B(_21080_),
    .Y(_21081_));
 AO21x1_ASAP7_75t_R _29600_ (.A1(_19647_),
    .A2(net1010),
    .B(_20752_),
    .Y(_21082_));
 INVx1_ASAP7_75t_R _29601_ (.A(_21082_),
    .Y(_21083_));
 NAND3x2_ASAP7_75t_R _29602_ (.B(_21081_),
    .C(_21083_),
    .Y(_21084_),
    .A(_21079_));
 NOR2x1_ASAP7_75t_R _29603_ (.A(_21074_),
    .B(_21084_),
    .Y(_21085_));
 NAND2x1_ASAP7_75t_R _29604_ (.A(_21068_),
    .B(_21085_),
    .Y(_21086_));
 AO21x1_ASAP7_75t_R _29605_ (.A1(_18651_),
    .A2(_18702_),
    .B(_18729_),
    .Y(_21087_));
 AND2x2_ASAP7_75t_R _29606_ (.A(_21087_),
    .B(_18733_),
    .Y(_21088_));
 AO21x1_ASAP7_75t_R _29607_ (.A1(_18600_),
    .A2(_18623_),
    .B(_18723_),
    .Y(_21089_));
 AO21x1_ASAP7_75t_R _29608_ (.A1(_18528_),
    .A2(_18548_),
    .B(_18723_),
    .Y(_21090_));
 AND2x2_ASAP7_75t_R _29609_ (.A(_21089_),
    .B(_21090_),
    .Y(_21091_));
 OA21x2_ASAP7_75t_R _29610_ (.A1(net2626),
    .A2(net2405),
    .B(_21091_),
    .Y(_21092_));
 NAND2x1_ASAP7_75t_R _29611_ (.A(_21088_),
    .B(_21092_),
    .Y(_21093_));
 AOI211x1_ASAP7_75t_R _29612_ (.A1(net1469),
    .A2(_18554_),
    .B(net2394),
    .C(net1563),
    .Y(_21094_));
 INVx1_ASAP7_75t_R _29613_ (.A(_21094_),
    .Y(_21095_));
 AO21x1_ASAP7_75t_R _29614_ (.A1(_18975_),
    .A2(net1965),
    .B(net2394),
    .Y(_21096_));
 AO21x1_ASAP7_75t_R _29615_ (.A1(net2386),
    .A2(_18547_),
    .B(net2394),
    .Y(_21097_));
 AND3x1_ASAP7_75t_R _29616_ (.A(_21095_),
    .B(_21096_),
    .C(_21097_),
    .Y(_21098_));
 NAND2x1_ASAP7_75t_R _29617_ (.A(_20257_),
    .B(_18718_),
    .Y(_21099_));
 AO21x1_ASAP7_75t_R _29618_ (.A1(net2504),
    .A2(_18992_),
    .B(_18712_),
    .Y(_21100_));
 NAND2x1_ASAP7_75t_R _29619_ (.A(_21099_),
    .B(_21100_),
    .Y(_21101_));
 AO21x1_ASAP7_75t_R _29620_ (.A1(_18651_),
    .A2(_18627_),
    .B(_18712_),
    .Y(_21102_));
 OAI21x1_ASAP7_75t_R _29621_ (.A1(net3376),
    .A2(_18712_),
    .B(_21102_),
    .Y(_21103_));
 AOI211x1_ASAP7_75t_R _29622_ (.A1(_18636_),
    .A2(_18718_),
    .B(_21101_),
    .C(_21103_),
    .Y(_21104_));
 NAND2x1_ASAP7_75t_R _29623_ (.A(_21098_),
    .B(_21104_),
    .Y(_21105_));
 NOR2x2_ASAP7_75t_R _29624_ (.A(_21093_),
    .B(_21105_),
    .Y(_21106_));
 AO21x1_ASAP7_75t_R _29625_ (.A1(_18992_),
    .A2(net2386),
    .B(_18682_),
    .Y(_21107_));
 AO21x1_ASAP7_75t_R _29626_ (.A1(_18553_),
    .A2(net1825),
    .B(_18682_),
    .Y(_21108_));
 NAND2x1_ASAP7_75t_R _29627_ (.A(_21107_),
    .B(_21108_),
    .Y(_21109_));
 OAI21x1_ASAP7_75t_R _29628_ (.A1(net2142),
    .A2(net2304),
    .B(_18698_),
    .Y(_21110_));
 AO21x1_ASAP7_75t_R _29629_ (.A1(_18702_),
    .A2(net1965),
    .B(net2182),
    .Y(_21111_));
 OAI21x1_ASAP7_75t_R _29630_ (.A1(_18627_),
    .A2(net2304),
    .B(_21111_),
    .Y(_21112_));
 NOR3x1_ASAP7_75t_R _29631_ (.A(_21109_),
    .B(_21110_),
    .C(_21112_),
    .Y(_21113_));
 AO21x1_ASAP7_75t_R _29632_ (.A1(net2012),
    .A2(net1726),
    .B(_18666_),
    .Y(_21114_));
 OA211x2_ASAP7_75t_R _29633_ (.A1(net2029),
    .A2(_18666_),
    .B(_21114_),
    .C(_18676_),
    .Y(_21115_));
 AO21x1_ASAP7_75t_R _29634_ (.A1(net2012),
    .A2(net2633),
    .B(_18655_),
    .Y(_21116_));
 NAND2x1_ASAP7_75t_R _29635_ (.A(net1732),
    .B(net2555),
    .Y(_21117_));
 AO21x1_ASAP7_75t_R _29636_ (.A1(_21117_),
    .A2(net2398),
    .B(_18655_),
    .Y(_21118_));
 AND4x1_ASAP7_75t_R _29637_ (.A(_21116_),
    .B(_19743_),
    .C(_21118_),
    .D(_20250_),
    .Y(_21119_));
 AND3x1_ASAP7_75t_R _29638_ (.A(_21113_),
    .B(_21115_),
    .C(_21119_),
    .Y(_21120_));
 NAND2x2_ASAP7_75t_R _29639_ (.A(_21106_),
    .B(_21120_),
    .Y(_21121_));
 NOR2x2_ASAP7_75t_R _29640_ (.A(_21086_),
    .B(_21121_),
    .Y(_21122_));
 NAND2x2_ASAP7_75t_R _29641_ (.A(_19120_),
    .B(_21122_),
    .Y(_21123_));
 XOR2x1_ASAP7_75t_R _29642_ (.A(_21123_),
    .Y(_21124_),
    .B(_20544_));
 INVx1_ASAP7_75t_R _29643_ (.A(_21124_),
    .Y(_21125_));
 AOI21x1_ASAP7_75t_R _29644_ (.A1(_21048_),
    .A2(_21050_),
    .B(_21125_),
    .Y(_21126_));
 INVx2_ASAP7_75t_R _29645_ (.A(_20899_),
    .Y(_21127_));
 NOR2x1_ASAP7_75t_R _29646_ (.A(_21046_),
    .B(_21127_),
    .Y(_21128_));
 NOR2x1_ASAP7_75t_R _29647_ (.A(_20899_),
    .B(_21047_),
    .Y(_21129_));
 OAI21x1_ASAP7_75t_R _29648_ (.A1(_21128_),
    .A2(_21129_),
    .B(_20967_),
    .Y(_21130_));
 NAND3x2_ASAP7_75t_R _29649_ (.B(_20965_),
    .C(_20934_),
    .Y(_21131_),
    .A(_17974_));
 XNOR2x2_ASAP7_75t_R _29650_ (.A(_20899_),
    .B(_21046_),
    .Y(_21132_));
 NAND2x1_ASAP7_75t_R _29651_ (.A(_21131_),
    .B(_21132_),
    .Y(_21133_));
 AOI21x1_ASAP7_75t_R _29652_ (.A1(_21130_),
    .A2(_21133_),
    .B(_21124_),
    .Y(_21134_));
 TAPCELL_ASAP7_75t_R TAP_820 ();
 OAI21x1_ASAP7_75t_R _29654_ (.A1(_21126_),
    .A2(_21134_),
    .B(net397),
    .Y(_21136_));
 TAPCELL_ASAP7_75t_R TAP_819 ();
 NOR2x1_ASAP7_75t_R _29656_ (.A(net397),
    .B(_00909_),
    .Y(_21138_));
 INVx2_ASAP7_75t_R _29657_ (.A(_21138_),
    .Y(_21139_));
 NAND3x2_ASAP7_75t_R _29658_ (.B(_14758_),
    .C(_21139_),
    .Y(_21140_),
    .A(_21136_));
 AO21x1_ASAP7_75t_R _29659_ (.A1(_21136_),
    .A2(_21139_),
    .B(_14758_),
    .Y(_21141_));
 NAND2x2_ASAP7_75t_R _29660_ (.A(_21140_),
    .B(_21141_),
    .Y(_00127_));
 AO21x1_ASAP7_75t_R _29661_ (.A1(_18553_),
    .A2(net2405),
    .B(net2394),
    .Y(_21142_));
 AO21x1_ASAP7_75t_R _29662_ (.A1(net1404),
    .A2(net2633),
    .B(net2394),
    .Y(_21143_));
 AO21x1_ASAP7_75t_R _29663_ (.A1(_18547_),
    .A2(net1570),
    .B(net2394),
    .Y(_21144_));
 NAND3x1_ASAP7_75t_R _29664_ (.A(_21142_),
    .B(_21143_),
    .C(_21144_),
    .Y(_21145_));
 AO21x1_ASAP7_75t_R _29665_ (.A1(_21063_),
    .A2(_18651_),
    .B(_18712_),
    .Y(_21146_));
 INVx1_ASAP7_75t_R _29666_ (.A(_19591_),
    .Y(_21147_));
 NAND3x1_ASAP7_75t_R _29667_ (.A(_21146_),
    .B(_21099_),
    .C(_21147_),
    .Y(_21148_));
 NOR2x1_ASAP7_75t_R _29668_ (.A(_21145_),
    .B(_21148_),
    .Y(_21149_));
 AO21x1_ASAP7_75t_R _29669_ (.A1(net2029),
    .A2(_18680_),
    .B(net2694),
    .Y(_21150_));
 INVx1_ASAP7_75t_R _29670_ (.A(_21150_),
    .Y(_21151_));
 NOR2x1_ASAP7_75t_R _29671_ (.A(net2694),
    .B(_18651_),
    .Y(_21152_));
 OR3x1_ASAP7_75t_R _29672_ (.A(_19759_),
    .B(_21151_),
    .C(_21152_),
    .Y(_21153_));
 AO21x1_ASAP7_75t_R _29673_ (.A1(net1404),
    .A2(net1823),
    .B(net2626),
    .Y(_21154_));
 AND2x2_ASAP7_75t_R _29674_ (.A(_18724_),
    .B(_21154_),
    .Y(_21155_));
 AO21x1_ASAP7_75t_R _29675_ (.A1(net2504),
    .A2(_19073_),
    .B(net2626),
    .Y(_21156_));
 AO21x1_ASAP7_75t_R _29676_ (.A1(_18528_),
    .A2(net2398),
    .B(net2626),
    .Y(_21157_));
 AND3x1_ASAP7_75t_R _29677_ (.A(_21156_),
    .B(_21157_),
    .C(_19595_),
    .Y(_21158_));
 NAND2x1_ASAP7_75t_R _29678_ (.A(_21155_),
    .B(_21158_),
    .Y(_21159_));
 NOR2x1_ASAP7_75t_R _29679_ (.A(_21153_),
    .B(_21159_),
    .Y(_21160_));
 NAND2x2_ASAP7_75t_R _29680_ (.A(_21149_),
    .B(_21160_),
    .Y(_21161_));
 AO21x1_ASAP7_75t_R _29681_ (.A1(_18627_),
    .A2(net1965),
    .B(net3006),
    .Y(_21162_));
 AO21x1_ASAP7_75t_R _29682_ (.A1(net2142),
    .A2(net2030),
    .B(net3006),
    .Y(_21163_));
 NOR2x1_ASAP7_75t_R _29683_ (.A(_18528_),
    .B(net3006),
    .Y(_21164_));
 INVx1_ASAP7_75t_R _29684_ (.A(_21164_),
    .Y(_21165_));
 AND3x2_ASAP7_75t_R _29685_ (.A(_21162_),
    .B(_21163_),
    .C(_21165_),
    .Y(_21166_));
 AO21x1_ASAP7_75t_R _29686_ (.A1(_18651_),
    .A2(net2405),
    .B(_18666_),
    .Y(_21167_));
 AO21x1_ASAP7_75t_R _29687_ (.A1(net1404),
    .A2(net1824),
    .B(_18666_),
    .Y(_21168_));
 AND2x2_ASAP7_75t_R _29688_ (.A(_21167_),
    .B(_21168_),
    .Y(_21169_));
 AO21x1_ASAP7_75t_R _29689_ (.A1(_19073_),
    .A2(net2142),
    .B(_18666_),
    .Y(_21170_));
 OA21x2_ASAP7_75t_R _29690_ (.A1(net1307),
    .A2(_18666_),
    .B(_21170_),
    .Y(_21171_));
 NAND3x2_ASAP7_75t_R _29691_ (.B(_21169_),
    .C(_21171_),
    .Y(_21172_),
    .A(_21166_));
 OA211x2_ASAP7_75t_R _29692_ (.A1(net3090),
    .A2(net3380),
    .B(_18696_),
    .C(net2101),
    .Y(_21173_));
 NAND2x1_ASAP7_75t_R _29693_ (.A(_18689_),
    .B(_19008_),
    .Y(_21174_));
 OA21x2_ASAP7_75t_R _29694_ (.A1(_18675_),
    .A2(_18681_),
    .B(_18683_),
    .Y(_21175_));
 OA21x2_ASAP7_75t_R _29695_ (.A1(_18572_),
    .A2(_19114_),
    .B(_18696_),
    .Y(_21176_));
 OR4x2_ASAP7_75t_R _29696_ (.A(_21173_),
    .B(_21174_),
    .C(_21175_),
    .D(_21176_),
    .Y(_21177_));
 NOR3x2_ASAP7_75t_R _29697_ (.B(_21172_),
    .C(_21177_),
    .Y(_21178_),
    .A(_21161_));
 OA21x2_ASAP7_75t_R _29698_ (.A1(net2615),
    .A2(net3379),
    .B(_19044_),
    .Y(_21179_));
 AO21x1_ASAP7_75t_R _29699_ (.A1(_18516_),
    .A2(net2633),
    .B(net2615),
    .Y(_21180_));
 AO21x1_ASAP7_75t_R _29700_ (.A1(_18553_),
    .A2(net2405),
    .B(net2615),
    .Y(_21181_));
 NAND2x1_ASAP7_75t_R _29701_ (.A(_21180_),
    .B(_21181_),
    .Y(_21182_));
 INVx1_ASAP7_75t_R _29702_ (.A(_21182_),
    .Y(_21183_));
 AO21x1_ASAP7_75t_R _29703_ (.A1(_19582_),
    .A2(net1965),
    .B(net2414),
    .Y(_21184_));
 NAND2x1_ASAP7_75t_R _29704_ (.A(_18613_),
    .B(_21184_),
    .Y(_21185_));
 INVx1_ASAP7_75t_R _29705_ (.A(_21185_),
    .Y(_21186_));
 AND3x1_ASAP7_75t_R _29706_ (.A(_21179_),
    .B(_21183_),
    .C(_21186_),
    .Y(_21187_));
 OA21x2_ASAP7_75t_R _29707_ (.A1(_18641_),
    .A2(_18584_),
    .B(_19052_),
    .Y(_21188_));
 NAND2x1_ASAP7_75t_R _29708_ (.A(_18614_),
    .B(_18635_),
    .Y(_21189_));
 AND3x1_ASAP7_75t_R _29709_ (.A(_20173_),
    .B(_20175_),
    .C(_21189_),
    .Y(_21190_));
 NAND2x1_ASAP7_75t_R _29710_ (.A(_21188_),
    .B(_21190_),
    .Y(_21191_));
 AO21x1_ASAP7_75t_R _29711_ (.A1(_19073_),
    .A2(net2142),
    .B(_18625_),
    .Y(_21192_));
 AO21x1_ASAP7_75t_R _29712_ (.A1(net1404),
    .A2(net2633),
    .B(_18625_),
    .Y(_21193_));
 OA211x2_ASAP7_75t_R _29713_ (.A1(net1307),
    .A2(_18625_),
    .B(_21192_),
    .C(_21193_),
    .Y(_21194_));
 INVx1_ASAP7_75t_R _29714_ (.A(_21194_),
    .Y(_21195_));
 NOR2x1_ASAP7_75t_R _29715_ (.A(_21191_),
    .B(_21195_),
    .Y(_21196_));
 NAND2x1_ASAP7_75t_R _29716_ (.A(_21187_),
    .B(_21196_),
    .Y(_21197_));
 OA21x2_ASAP7_75t_R _29717_ (.A1(_18572_),
    .A2(_20192_),
    .B(_18570_),
    .Y(_21198_));
 AO21x1_ASAP7_75t_R _29718_ (.A1(_18590_),
    .A2(_18570_),
    .B(_21198_),
    .Y(_21199_));
 NAND2x2_ASAP7_75t_R _29719_ (.A(_20188_),
    .B(_18576_),
    .Y(_21200_));
 AO21x1_ASAP7_75t_R _29720_ (.A1(_18528_),
    .A2(_18548_),
    .B(_18588_),
    .Y(_21201_));
 NAND2x2_ASAP7_75t_R _29721_ (.A(_18585_),
    .B(_18592_),
    .Y(_21202_));
 NAND3x2_ASAP7_75t_R _29722_ (.B(_21052_),
    .C(_21202_),
    .Y(_21203_),
    .A(_21201_));
 NOR3x2_ASAP7_75t_R _29723_ (.B(_21200_),
    .C(_21203_),
    .Y(_21204_),
    .A(_21199_));
 AND2x2_ASAP7_75t_R _29724_ (.A(_19110_),
    .B(_19698_),
    .Y(_21205_));
 AO21x1_ASAP7_75t_R _29725_ (.A1(net2177),
    .A2(_18601_),
    .B(net2479),
    .Y(_21206_));
 NOR2x1_ASAP7_75t_R _29726_ (.A(_18975_),
    .B(net2479),
    .Y(_21207_));
 INVx1_ASAP7_75t_R _29727_ (.A(_21207_),
    .Y(_21208_));
 AND4x2_ASAP7_75t_R _29728_ (.A(_18551_),
    .B(_19071_),
    .C(_21206_),
    .D(_21208_),
    .Y(_21209_));
 NAND3x2_ASAP7_75t_R _29729_ (.B(_21205_),
    .C(_21209_),
    .Y(_21210_),
    .A(_21204_));
 NOR2x2_ASAP7_75t_R _29730_ (.A(_21197_),
    .B(_21210_),
    .Y(_21211_));
 NAND3x2_ASAP7_75t_R _29731_ (.B(_19120_),
    .C(_21211_),
    .Y(_21212_),
    .A(_21178_));
 AO21x1_ASAP7_75t_R _29732_ (.A1(_18881_),
    .A2(_18883_),
    .B(_17997_),
    .Y(_21213_));
 AO21x1_ASAP7_75t_R _29733_ (.A1(_18014_),
    .A2(_18002_),
    .B(_17997_),
    .Y(_21214_));
 NAND3x1_ASAP7_75t_R _29734_ (.A(_21213_),
    .B(_21214_),
    .C(_20905_),
    .Y(_21215_));
 AO21x1_ASAP7_75t_R _29735_ (.A1(net3203),
    .A2(_18073_),
    .B(_17977_),
    .Y(_21216_));
 NAND2x1_ASAP7_75t_R _29736_ (.A(_18105_),
    .B(_19376_),
    .Y(_21217_));
 NAND3x1_ASAP7_75t_R _29737_ (.A(_17990_),
    .B(_21216_),
    .C(_21217_),
    .Y(_21218_));
 NOR2x1_ASAP7_75t_R _29738_ (.A(_21215_),
    .B(_21218_),
    .Y(_21219_));
 OAI21x1_ASAP7_75t_R _29739_ (.A1(_18134_),
    .A2(net2843),
    .B(net3196),
    .Y(_21220_));
 NAND2x1_ASAP7_75t_R _29740_ (.A(net3196),
    .B(_18110_),
    .Y(_21221_));
 NAND3x1_ASAP7_75t_R _29741_ (.A(_20914_),
    .B(_21220_),
    .C(_21221_),
    .Y(_21222_));
 AO21x1_ASAP7_75t_R _29742_ (.A1(_17980_),
    .A2(_17999_),
    .B(_18012_),
    .Y(_21223_));
 OAI21x1_ASAP7_75t_R _29743_ (.A1(net3216),
    .A2(_19855_),
    .B(_21223_),
    .Y(_21224_));
 AO21x1_ASAP7_75t_R _29744_ (.A1(net1348),
    .A2(net1622),
    .B(_18012_),
    .Y(_21225_));
 AO21x1_ASAP7_75t_R _29745_ (.A1(net1530),
    .A2(_18081_),
    .B(_18012_),
    .Y(_21226_));
 NAND2x1_ASAP7_75t_R _29746_ (.A(_21225_),
    .B(_21226_),
    .Y(_21227_));
 NOR3x1_ASAP7_75t_R _29747_ (.A(_21222_),
    .B(_21224_),
    .C(_21227_),
    .Y(_21228_));
 NAND2x1_ASAP7_75t_R _29748_ (.A(_21219_),
    .B(_21228_),
    .Y(_21229_));
 AOI22x1_ASAP7_75t_R _29749_ (.A1(_19403_),
    .A2(net1645),
    .B1(net2842),
    .B2(_18069_),
    .Y(_21230_));
 INVx1_ASAP7_75t_R _29750_ (.A(_19401_),
    .Y(_21231_));
 AOI211x1_ASAP7_75t_R _29751_ (.A1(net3366),
    .A2(_17953_),
    .B(net1910),
    .C(net1074),
    .Y(_21232_));
 NOR2x1_ASAP7_75t_R _29752_ (.A(_21231_),
    .B(_21232_),
    .Y(_21233_));
 NAND2x1_ASAP7_75t_R _29753_ (.A(_21230_),
    .B(_21233_),
    .Y(_21234_));
 NOR2x1_ASAP7_75t_R _29754_ (.A(_18076_),
    .B(_18942_),
    .Y(_21235_));
 AOI21x1_ASAP7_75t_R _29755_ (.A1(_18147_),
    .A2(_18010_),
    .B(_18074_),
    .Y(_21236_));
 AOI211x1_ASAP7_75t_R _29756_ (.A1(net1061),
    .A2(net1644),
    .B(net2057),
    .C(_18074_),
    .Y(_21237_));
 NOR2x1_ASAP7_75t_R _29757_ (.A(_21236_),
    .B(_21237_),
    .Y(_21238_));
 NAND2x1_ASAP7_75t_R _29758_ (.A(_21235_),
    .B(_21238_),
    .Y(_21239_));
 NOR2x1_ASAP7_75t_R _29759_ (.A(_21234_),
    .B(_21239_),
    .Y(_21240_));
 AO21x1_ASAP7_75t_R _29760_ (.A1(_18010_),
    .A2(net1348),
    .B(_18054_),
    .Y(_21241_));
 AO21x1_ASAP7_75t_R _29761_ (.A1(_18002_),
    .A2(net1145),
    .B(_18054_),
    .Y(_21242_));
 NAND2x1_ASAP7_75t_R _29762_ (.A(net3218),
    .B(_18952_),
    .Y(_21243_));
 NAND3x1_ASAP7_75t_R _29763_ (.A(_21241_),
    .B(_21242_),
    .C(_21243_),
    .Y(_21244_));
 AO31x2_ASAP7_75t_R _29764_ (.A1(_18958_),
    .A2(_18057_),
    .A3(_18883_),
    .B(_18039_),
    .Y(_21245_));
 NOR2x1_ASAP7_75t_R _29765_ (.A(_18039_),
    .B(_18028_),
    .Y(_21246_));
 NOR3x1_ASAP7_75t_R _29766_ (.A(_19382_),
    .B(_18962_),
    .C(_21246_),
    .Y(_21247_));
 NAND2x1_ASAP7_75t_R _29767_ (.A(_21245_),
    .B(_21247_),
    .Y(_21248_));
 NOR2x1_ASAP7_75t_R _29768_ (.A(_21244_),
    .B(_21248_),
    .Y(_21249_));
 NAND2x1_ASAP7_75t_R _29769_ (.A(_21240_),
    .B(_21249_),
    .Y(_21250_));
 NOR2x1_ASAP7_75t_R _29770_ (.A(_21250_),
    .B(_21229_),
    .Y(_21251_));
 AO21x1_ASAP7_75t_R _29771_ (.A1(net1622),
    .A2(net1070),
    .B(_19423_),
    .Y(_21252_));
 NAND2x1_ASAP7_75t_R _29772_ (.A(net2843),
    .B(_18175_),
    .Y(_21253_));
 NAND3x1_ASAP7_75t_R _29773_ (.A(_19788_),
    .B(_21252_),
    .C(_21253_),
    .Y(_21254_));
 NOR2x1_ASAP7_75t_R _29774_ (.A(_18169_),
    .B(_20430_),
    .Y(_21255_));
 AOI21x1_ASAP7_75t_R _29775_ (.A1(net1542),
    .A2(_18904_),
    .B(_21255_),
    .Y(_21256_));
 OA21x2_ASAP7_75t_R _29776_ (.A1(_18178_),
    .A2(_17952_),
    .B(_18165_),
    .Y(_21257_));
 NOR2x1_ASAP7_75t_R _29777_ (.A(_21257_),
    .B(_18902_),
    .Y(_21258_));
 NAND2x1_ASAP7_75t_R _29778_ (.A(_21256_),
    .B(_21258_),
    .Y(_21259_));
 NOR2x1_ASAP7_75t_R _29779_ (.A(_21254_),
    .B(_21259_),
    .Y(_21260_));
 OAI21x1_ASAP7_75t_R _29780_ (.A1(_18131_),
    .A2(_18000_),
    .B(_18155_),
    .Y(_21261_));
 OAI21x1_ASAP7_75t_R _29781_ (.A1(_18901_),
    .A2(_18178_),
    .B(_18155_),
    .Y(_21262_));
 NAND2x1_ASAP7_75t_R _29782_ (.A(_18155_),
    .B(_17925_),
    .Y(_21263_));
 NAND3x1_ASAP7_75t_R _29783_ (.A(_21261_),
    .B(_21262_),
    .C(_21263_),
    .Y(_21264_));
 AO21x1_ASAP7_75t_R _29784_ (.A1(_18881_),
    .A2(_17943_),
    .B(net2946),
    .Y(_21265_));
 OAI21x1_ASAP7_75t_R _29785_ (.A1(_17999_),
    .A2(net2446),
    .B(_21265_),
    .Y(_21266_));
 AO21x1_ASAP7_75t_R _29786_ (.A1(net2824),
    .A2(_18081_),
    .B(net2946),
    .Y(_21267_));
 AO21x1_ASAP7_75t_R _29787_ (.A1(_18052_),
    .A2(_17956_),
    .B(net2946),
    .Y(_21268_));
 NAND2x1_ASAP7_75t_R _29788_ (.A(_21267_),
    .B(_21268_),
    .Y(_21269_));
 NOR3x1_ASAP7_75t_R _29789_ (.A(_21264_),
    .B(_21266_),
    .C(_21269_),
    .Y(_21270_));
 NAND2x1_ASAP7_75t_R _29790_ (.A(_21270_),
    .B(_21260_),
    .Y(_21271_));
 AO21x1_ASAP7_75t_R _29791_ (.A1(net3186),
    .A2(_17958_),
    .B(_17931_),
    .Y(_21272_));
 AO21x1_ASAP7_75t_R _29792_ (.A1(_17980_),
    .A2(_18057_),
    .B(_17931_),
    .Y(_21273_));
 NAND2x1_ASAP7_75t_R _29793_ (.A(_18158_),
    .B(_17932_),
    .Y(_21274_));
 NAND3x1_ASAP7_75t_R _29794_ (.A(_21272_),
    .B(_21273_),
    .C(_21274_),
    .Y(_21275_));
 AO31x2_ASAP7_75t_R _29795_ (.A1(net1145),
    .A2(net1368),
    .A3(_18002_),
    .B(_17968_),
    .Y(_21276_));
 AOI211x1_ASAP7_75t_R _29796_ (.A1(net3366),
    .A2(_17953_),
    .B(net1074),
    .C(_17968_),
    .Y(_21277_));
 NOR2x1_ASAP7_75t_R _29797_ (.A(_21277_),
    .B(_20605_),
    .Y(_21278_));
 NAND2x1_ASAP7_75t_R _29798_ (.A(_21276_),
    .B(_21278_),
    .Y(_21279_));
 NOR2x1_ASAP7_75t_R _29799_ (.A(_21275_),
    .B(_21279_),
    .Y(_21280_));
 NOR2x1_ASAP7_75t_R _29800_ (.A(_20951_),
    .B(_18874_),
    .Y(_21281_));
 OA21x2_ASAP7_75t_R _29801_ (.A1(_18047_),
    .A2(_18923_),
    .B(_18123_),
    .Y(_21282_));
 OA21x2_ASAP7_75t_R _29802_ (.A1(_18158_),
    .A2(_18130_),
    .B(_18123_),
    .Y(_21283_));
 NOR2x1_ASAP7_75t_R _29803_ (.A(_21282_),
    .B(_21283_),
    .Y(_21284_));
 NAND2x1_ASAP7_75t_R _29804_ (.A(_21281_),
    .B(_21284_),
    .Y(_21285_));
 AND2x2_ASAP7_75t_R _29805_ (.A(_18116_),
    .B(_19769_),
    .Y(_21286_));
 AND2x2_ASAP7_75t_R _29806_ (.A(_20955_),
    .B(_18108_),
    .Y(_21287_));
 NAND2x1_ASAP7_75t_R _29807_ (.A(_21286_),
    .B(_21287_),
    .Y(_21288_));
 NOR2x1_ASAP7_75t_R _29808_ (.A(_21285_),
    .B(_21288_),
    .Y(_21289_));
 NAND2x1_ASAP7_75t_R _29809_ (.A(_21280_),
    .B(_21289_),
    .Y(_21290_));
 NOR2x1_ASAP7_75t_R _29810_ (.A(_21290_),
    .B(_21271_),
    .Y(_21291_));
 NAND2x2_ASAP7_75t_R _29811_ (.A(_21251_),
    .B(_21291_),
    .Y(_21292_));
 XNOR2x1_ASAP7_75t_R _29812_ (.B(_17905_),
    .Y(_21293_),
    .A(_21292_));
 XOR2x2_ASAP7_75t_R _29813_ (.A(_21212_),
    .B(_21293_),
    .Y(_21294_));
 AO21x1_ASAP7_75t_R _29814_ (.A1(net1482),
    .A2(net3247),
    .B(net2994),
    .Y(_21295_));
 OAI21x1_ASAP7_75t_R _29815_ (.A1(net2595),
    .A2(_19174_),
    .B(_21295_),
    .Y(_21296_));
 NAND2x1_ASAP7_75t_R _29816_ (.A(net2971),
    .B(_19170_),
    .Y(_21297_));
 NAND2x2_ASAP7_75t_R _29817_ (.A(_20115_),
    .B(_21297_),
    .Y(_21298_));
 AO21x1_ASAP7_75t_R _29818_ (.A1(net937),
    .A2(net2093),
    .B(_18479_),
    .Y(_21299_));
 AO21x1_ASAP7_75t_R _29819_ (.A1(net2473),
    .A2(_18335_),
    .B(_18479_),
    .Y(_21300_));
 NAND2x1_ASAP7_75t_R _29820_ (.A(_21299_),
    .B(_21300_),
    .Y(_21301_));
 NOR3x1_ASAP7_75t_R _29821_ (.A(_21296_),
    .B(_21298_),
    .C(_21301_),
    .Y(_21302_));
 AO21x1_ASAP7_75t_R _29822_ (.A1(net2964),
    .A2(net1482),
    .B(_18456_),
    .Y(_21303_));
 AO21x2_ASAP7_75t_R _29823_ (.A1(_18333_),
    .A2(net2437),
    .B(_18456_),
    .Y(_21304_));
 NAND2x2_ASAP7_75t_R _29824_ (.A(net2754),
    .B(_19185_),
    .Y(_21305_));
 NAND3x2_ASAP7_75t_R _29825_ (.B(_21304_),
    .C(_21305_),
    .Y(_21306_),
    .A(_21303_));
 AOI211x1_ASAP7_75t_R _29826_ (.A1(_18259_),
    .A2(_18469_),
    .B(_19464_),
    .C(_18466_),
    .Y(_21307_));
 OA21x2_ASAP7_75t_R _29827_ (.A1(_18444_),
    .A2(_18445_),
    .B(_18469_),
    .Y(_21308_));
 AO21x1_ASAP7_75t_R _29828_ (.A1(net2964),
    .A2(_18383_),
    .B(_18464_),
    .Y(_21309_));
 INVx1_ASAP7_75t_R _29829_ (.A(_21309_),
    .Y(_21310_));
 NOR2x1_ASAP7_75t_R _29830_ (.A(_21308_),
    .B(_21310_),
    .Y(_21311_));
 NAND2x1_ASAP7_75t_R _29831_ (.A(_21307_),
    .B(_21311_),
    .Y(_21312_));
 NOR2x1_ASAP7_75t_R _29832_ (.A(_21306_),
    .B(_21312_),
    .Y(_21313_));
 NAND2x1_ASAP7_75t_R _29833_ (.A(_21302_),
    .B(_21313_),
    .Y(_21314_));
 INVx1_ASAP7_75t_R _29834_ (.A(_18443_),
    .Y(_21315_));
 AO21x1_ASAP7_75t_R _29835_ (.A1(_18333_),
    .A2(_18419_),
    .B(_18439_),
    .Y(_21316_));
 NAND3x2_ASAP7_75t_R _29836_ (.B(_21315_),
    .C(_21316_),
    .Y(_21317_),
    .A(_20979_));
 NOR2x1_ASAP7_75t_R _29837_ (.A(_20976_),
    .B(_19157_),
    .Y(_21318_));
 NAND2x1_ASAP7_75t_R _29838_ (.A(_18254_),
    .B(_18434_),
    .Y(_21319_));
 AO21x1_ASAP7_75t_R _29839_ (.A1(net2963),
    .A2(net2407),
    .B(_18428_),
    .Y(_21320_));
 NAND2x1_ASAP7_75t_R _29840_ (.A(_21319_),
    .B(_21320_),
    .Y(_21321_));
 INVx1_ASAP7_75t_R _29841_ (.A(_21321_),
    .Y(_21322_));
 NAND2x1_ASAP7_75t_R _29842_ (.A(_21318_),
    .B(_21322_),
    .Y(_21323_));
 NOR2x1_ASAP7_75t_R _29843_ (.A(_21317_),
    .B(_21323_),
    .Y(_21324_));
 AO21x1_ASAP7_75t_R _29844_ (.A1(_18453_),
    .A2(net1482),
    .B(_18248_),
    .Y(_21325_));
 AO21x1_ASAP7_75t_R _29845_ (.A1(_18305_),
    .A2(_18333_),
    .B(_18248_),
    .Y(_21326_));
 NAND2x1_ASAP7_75t_R _29846_ (.A(_18247_),
    .B(_18401_),
    .Y(_21327_));
 NAND3x1_ASAP7_75t_R _29847_ (.A(_21325_),
    .B(_21326_),
    .C(_21327_),
    .Y(_21328_));
 NAND2x1_ASAP7_75t_R _29848_ (.A(net2533),
    .B(_18416_),
    .Y(_21329_));
 AO21x1_ASAP7_75t_R _29849_ (.A1(_18460_),
    .A2(net2437),
    .B(_18266_),
    .Y(_21330_));
 NAND2x1_ASAP7_75t_R _29850_ (.A(_21329_),
    .B(_21330_),
    .Y(_21331_));
 AO21x1_ASAP7_75t_R _29851_ (.A1(_18314_),
    .A2(_18442_),
    .B(_18266_),
    .Y(_21332_));
 NAND2x1_ASAP7_75t_R _29852_ (.A(_20658_),
    .B(_21332_),
    .Y(_21333_));
 NOR2x1_ASAP7_75t_R _29853_ (.A(_21331_),
    .B(_21333_),
    .Y(_21334_));
 INVx1_ASAP7_75t_R _29854_ (.A(_21334_),
    .Y(_21335_));
 NOR2x1_ASAP7_75t_R _29855_ (.A(_21328_),
    .B(_21335_),
    .Y(_21336_));
 NAND2x1_ASAP7_75t_R _29856_ (.A(_21324_),
    .B(_21336_),
    .Y(_21337_));
 NOR2x2_ASAP7_75t_R _29857_ (.A(_21314_),
    .B(_21337_),
    .Y(_21338_));
 AO31x2_ASAP7_75t_R _29858_ (.A1(net2095),
    .A2(net2050),
    .A3(_18335_),
    .B(_18364_),
    .Y(_21339_));
 NOR2x1_ASAP7_75t_R _29859_ (.A(_18364_),
    .B(_18381_),
    .Y(_21340_));
 NOR2x1_ASAP7_75t_R _29860_ (.A(_21340_),
    .B(_19544_),
    .Y(_21341_));
 NAND2x1_ASAP7_75t_R _29861_ (.A(_21339_),
    .B(_21341_),
    .Y(_21342_));
 AO21x1_ASAP7_75t_R _29862_ (.A1(_18314_),
    .A2(net1753),
    .B(_18354_),
    .Y(_21343_));
 NOR2x1_ASAP7_75t_R _29863_ (.A(_18327_),
    .B(_18354_),
    .Y(_21344_));
 AOI211x1_ASAP7_75t_R _29864_ (.A1(net3005),
    .A2(net1394),
    .B(_18354_),
    .C(net2975),
    .Y(_21345_));
 NOR2x1_ASAP7_75t_R _29865_ (.A(_21344_),
    .B(_21345_),
    .Y(_21346_));
 NAND2x1_ASAP7_75t_R _29866_ (.A(_21343_),
    .B(_21346_),
    .Y(_21347_));
 NOR2x2_ASAP7_75t_R _29867_ (.A(_21347_),
    .B(_21342_),
    .Y(_21348_));
 AOI21x1_ASAP7_75t_R _29868_ (.A1(net2849),
    .A2(_18398_),
    .B(_20719_),
    .Y(_21349_));
 INVx2_ASAP7_75t_R _29869_ (.A(_19539_),
    .Y(_21350_));
 AOI211x1_ASAP7_75t_R _29870_ (.A1(net3005),
    .A2(_18237_),
    .B(_18395_),
    .C(net1958),
    .Y(_21351_));
 NOR2x1_ASAP7_75t_R _29871_ (.A(_21351_),
    .B(_21350_),
    .Y(_21352_));
 NAND2x1_ASAP7_75t_R _29872_ (.A(_21349_),
    .B(_21352_),
    .Y(_21353_));
 AOI211x1_ASAP7_75t_R _29873_ (.A1(_18242_),
    .A2(net3246),
    .B(net2981),
    .C(_18282_),
    .Y(_21354_));
 INVx1_ASAP7_75t_R _29874_ (.A(_21354_),
    .Y(_21355_));
 AOI211x1_ASAP7_75t_R _29875_ (.A1(net3005),
    .A2(_18237_),
    .B(_18377_),
    .C(net2093),
    .Y(_21356_));
 AOI211x1_ASAP7_75t_R _29876_ (.A1(net1087),
    .A2(net1395),
    .B(_18377_),
    .C(net2499),
    .Y(_21357_));
 NOR2x1_ASAP7_75t_R _29877_ (.A(_21356_),
    .B(_21357_),
    .Y(_21358_));
 NAND2x1_ASAP7_75t_R _29878_ (.A(_21355_),
    .B(_21358_),
    .Y(_21359_));
 NOR2x1_ASAP7_75t_R _29879_ (.A(_21359_),
    .B(_21353_),
    .Y(_21360_));
 NAND2x2_ASAP7_75t_R _29880_ (.A(_21348_),
    .B(_21360_),
    .Y(_21361_));
 AO21x1_ASAP7_75t_R _29881_ (.A1(net2505),
    .A2(net2095),
    .B(net2982),
    .Y(_21362_));
 AO21x1_ASAP7_75t_R _29882_ (.A1(net2671),
    .A2(_18460_),
    .B(_18287_),
    .Y(_21363_));
 NAND3x2_ASAP7_75t_R _29883_ (.B(_21363_),
    .C(_21029_),
    .Y(_21364_),
    .A(_21362_));
 AO31x2_ASAP7_75t_R _29884_ (.A1(net2107),
    .A2(_18327_),
    .A3(net2506),
    .B(_18300_),
    .Y(_21365_));
 AO21x1_ASAP7_75t_R _29885_ (.A1(_18381_),
    .A2(net2964),
    .B(_18300_),
    .Y(_21366_));
 NAND3x1_ASAP7_75t_R _29886_ (.A(_21365_),
    .B(_21366_),
    .C(_18302_),
    .Y(_21367_));
 NOR2x1_ASAP7_75t_R _29887_ (.A(_21364_),
    .B(_21367_),
    .Y(_21368_));
 NAND2x1_ASAP7_75t_R _29888_ (.A(_18444_),
    .B(_18345_),
    .Y(_21369_));
 NAND3x1_ASAP7_75t_R _29889_ (.A(_21037_),
    .B(_19526_),
    .C(_21369_),
    .Y(_21370_));
 INVx1_ASAP7_75t_R _29890_ (.A(_21370_),
    .Y(_21371_));
 AO21x1_ASAP7_75t_R _29891_ (.A1(net2748),
    .A2(net2437),
    .B(_18318_),
    .Y(_21372_));
 NAND2x1_ASAP7_75t_R _29892_ (.A(_21372_),
    .B(_20028_),
    .Y(_21373_));
 AO21x1_ASAP7_75t_R _29893_ (.A1(net1335),
    .A2(net937),
    .B(_18318_),
    .Y(_21374_));
 AO21x1_ASAP7_75t_R _29894_ (.A1(net2945),
    .A2(net3182),
    .B(_18318_),
    .Y(_21375_));
 NAND2x1_ASAP7_75t_R _29895_ (.A(_21374_),
    .B(_21375_),
    .Y(_21376_));
 NOR2x1_ASAP7_75t_R _29896_ (.A(_21373_),
    .B(_21376_),
    .Y(_21377_));
 NAND2x1_ASAP7_75t_R _29897_ (.A(_21371_),
    .B(_21377_),
    .Y(_21378_));
 INVx1_ASAP7_75t_R _29898_ (.A(_21378_),
    .Y(_21379_));
 NAND2x1_ASAP7_75t_R _29899_ (.A(_21368_),
    .B(_21379_),
    .Y(_21380_));
 NOR2x1_ASAP7_75t_R _29900_ (.A(_21361_),
    .B(_21380_),
    .Y(_21381_));
 NAND2x2_ASAP7_75t_R _29901_ (.A(_21338_),
    .B(_21381_),
    .Y(_21382_));
 XOR2x1_ASAP7_75t_R _29902_ (.A(_20899_),
    .Y(_21383_),
    .B(_21382_));
 AO21x1_ASAP7_75t_R _29903_ (.A1(_21294_),
    .A2(_21383_),
    .B(net390),
    .Y(_21384_));
 NOR2x1_ASAP7_75t_R _29904_ (.A(_21383_),
    .B(_21294_),
    .Y(_21385_));
 NAND2x1_ASAP7_75t_R _29905_ (.A(_00908_),
    .B(net390),
    .Y(_21386_));
 OA21x2_ASAP7_75t_R _29906_ (.A1(_21384_),
    .A2(_21385_),
    .B(_21386_),
    .Y(_21387_));
 XOR2x2_ASAP7_75t_R _29907_ (.A(_21387_),
    .B(_14645_),
    .Y(_00128_));
 NOR2x2_ASAP7_75t_R _29908_ (.A(net2144),
    .B(_18205_),
    .Y(_21388_));
 NAND2x1_ASAP7_75t_R _29909_ (.A(_18192_),
    .B(_21388_),
    .Y(_21389_));
 NAND2x2_ASAP7_75t_R _29910_ (.A(_17918_),
    .B(_17796_),
    .Y(_21390_));
 NAND2x1_ASAP7_75t_R _29911_ (.A(_21390_),
    .B(_18193_),
    .Y(_21391_));
 INVx1_ASAP7_75t_R _29912_ (.A(_21301_),
    .Y(_21392_));
 NOR2x1_ASAP7_75t_R _29913_ (.A(_21298_),
    .B(_21296_),
    .Y(_21393_));
 NAND2x1_ASAP7_75t_R _29914_ (.A(_21392_),
    .B(_21393_),
    .Y(_21394_));
 INVx1_ASAP7_75t_R _29915_ (.A(_21306_),
    .Y(_21395_));
 AO21x1_ASAP7_75t_R _29916_ (.A1(net2753),
    .A2(net2251),
    .B(net3310),
    .Y(_21396_));
 NAND2x1_ASAP7_75t_R _29917_ (.A(_21309_),
    .B(_21396_),
    .Y(_21397_));
 AO21x1_ASAP7_75t_R _29918_ (.A1(net2457),
    .A2(net2347),
    .B(net3310),
    .Y(_21398_));
 OAI21x1_ASAP7_75t_R _29919_ (.A1(net2437),
    .A2(net3310),
    .B(_21398_),
    .Y(_21399_));
 NOR2x1_ASAP7_75t_R _29920_ (.A(_21397_),
    .B(_21399_),
    .Y(_21400_));
 NAND2x1_ASAP7_75t_R _29921_ (.A(_21395_),
    .B(_21400_),
    .Y(_21401_));
 NOR2x1_ASAP7_75t_R _29922_ (.A(_21394_),
    .B(_21401_),
    .Y(_21402_));
 AO21x1_ASAP7_75t_R _29923_ (.A1(net2699),
    .A2(net937),
    .B(_18428_),
    .Y(_21403_));
 NAND2x1_ASAP7_75t_R _29924_ (.A(_20977_),
    .B(_21403_),
    .Y(_21404_));
 NOR2x1_ASAP7_75t_R _29925_ (.A(_21404_),
    .B(_21321_),
    .Y(_21405_));
 INVx1_ASAP7_75t_R _29926_ (.A(_21317_),
    .Y(_21406_));
 NAND2x1_ASAP7_75t_R _29927_ (.A(_21405_),
    .B(_21406_),
    .Y(_21407_));
 INVx1_ASAP7_75t_R _29928_ (.A(_21328_),
    .Y(_21408_));
 NAND2x1_ASAP7_75t_R _29929_ (.A(_21408_),
    .B(_21334_),
    .Y(_21409_));
 NOR2x2_ASAP7_75t_R _29930_ (.A(_21409_),
    .B(_21407_),
    .Y(_21410_));
 NAND2x2_ASAP7_75t_R _29931_ (.A(_21402_),
    .B(_21410_),
    .Y(_21411_));
 NAND2x1_ASAP7_75t_R _29932_ (.A(_18302_),
    .B(_21366_),
    .Y(_21412_));
 INVx1_ASAP7_75t_R _29933_ (.A(_21365_),
    .Y(_21413_));
 NOR2x1_ASAP7_75t_R _29934_ (.A(_21412_),
    .B(_21413_),
    .Y(_21414_));
 INVx1_ASAP7_75t_R _29935_ (.A(_21364_),
    .Y(_21415_));
 NAND2x1_ASAP7_75t_R _29936_ (.A(_21414_),
    .B(_21415_),
    .Y(_21416_));
 NOR2x1_ASAP7_75t_R _29937_ (.A(_21378_),
    .B(_21416_),
    .Y(_21417_));
 INVx2_ASAP7_75t_R _29938_ (.A(_21361_),
    .Y(_21418_));
 NAND2x2_ASAP7_75t_R _29939_ (.A(_21417_),
    .B(_21418_),
    .Y(_21419_));
 NOR2x2_ASAP7_75t_R _29940_ (.A(_21411_),
    .B(_21419_),
    .Y(_21420_));
 AOI21x1_ASAP7_75t_R _29941_ (.A1(_21389_),
    .A2(_21391_),
    .B(_21420_),
    .Y(_21421_));
 NAND2x1_ASAP7_75t_R _29942_ (.A(_18192_),
    .B(_21390_),
    .Y(_21422_));
 NAND2x1_ASAP7_75t_R _29943_ (.A(_21388_),
    .B(_18193_),
    .Y(_21423_));
 AOI21x1_ASAP7_75t_R _29944_ (.A1(_21422_),
    .A2(_21423_),
    .B(_21382_),
    .Y(_21424_));
 OA21x2_ASAP7_75t_R _29945_ (.A1(_21421_),
    .A2(_21424_),
    .B(net2888),
    .Y(_21425_));
 NOR3x1_ASAP7_75t_R _29946_ (.A(_21421_),
    .B(_21424_),
    .C(net2888),
    .Y(_21426_));
 TAPCELL_ASAP7_75t_R TAP_818 ();
 OAI21x1_ASAP7_75t_R _29948_ (.A1(_21425_),
    .A2(_21426_),
    .B(net391),
    .Y(_21428_));
 NOR2x1_ASAP7_75t_R _29949_ (.A(net391),
    .B(_00907_),
    .Y(_21429_));
 INVx1_ASAP7_75t_R _29950_ (.A(_21429_),
    .Y(_21430_));
 NAND3x1_ASAP7_75t_R _29951_ (.A(_21428_),
    .B(_15432_),
    .C(_21430_),
    .Y(_21431_));
 AO21x1_ASAP7_75t_R _29952_ (.A1(_21428_),
    .A2(_21430_),
    .B(_15432_),
    .Y(_21432_));
 NAND2x1_ASAP7_75t_R _29953_ (.A(_21431_),
    .B(_21432_),
    .Y(_00089_));
 AND2x2_ASAP7_75t_R _29954_ (.A(net390),
    .B(_00906_),
    .Y(_21433_));
 AOI21x1_ASAP7_75t_R _29955_ (.A1(_18279_),
    .A2(_18506_),
    .B(_21382_),
    .Y(_21434_));
 NOR2x1_ASAP7_75t_R _29956_ (.A(_18451_),
    .B(_18503_),
    .Y(_21435_));
 INVx1_ASAP7_75t_R _29957_ (.A(_18393_),
    .Y(_21436_));
 NAND2x1_ASAP7_75t_R _29958_ (.A(_18400_),
    .B(_18407_),
    .Y(_21437_));
 NOR2x1_ASAP7_75t_R _29959_ (.A(_21436_),
    .B(_21437_),
    .Y(_21438_));
 NAND2x1_ASAP7_75t_R _29960_ (.A(_18375_),
    .B(_21438_),
    .Y(_21439_));
 INVx1_ASAP7_75t_R _29961_ (.A(_18312_),
    .Y(_21440_));
 INVx1_ASAP7_75t_R _29962_ (.A(_18348_),
    .Y(_21441_));
 NAND2x1_ASAP7_75t_R _29963_ (.A(_21440_),
    .B(_21441_),
    .Y(_21442_));
 NOR2x1_ASAP7_75t_R _29964_ (.A(_21439_),
    .B(_21442_),
    .Y(_21443_));
 NAND2x2_ASAP7_75t_R _29965_ (.A(_21435_),
    .B(_21443_),
    .Y(_21444_));
 NOR3x2_ASAP7_75t_R _29966_ (.B(net2342),
    .C(_20657_),
    .Y(_21445_),
    .A(_21444_));
 NOR2x2_ASAP7_75t_R _29967_ (.A(_21434_),
    .B(_21445_),
    .Y(_21446_));
 INVx3_ASAP7_75t_R _29968_ (.A(_21446_),
    .Y(_21447_));
 NOR2x2_ASAP7_75t_R _29969_ (.A(net3239),
    .B(_21447_),
    .Y(_21448_));
 NOR2x1_ASAP7_75t_R _29970_ (.A(_21446_),
    .B(net2820),
    .Y(_21449_));
 XOR2x2_ASAP7_75t_R _29971_ (.A(net2888),
    .B(_19679_),
    .Y(_21450_));
 OAI21x1_ASAP7_75t_R _29972_ (.A1(_21448_),
    .A2(_21449_),
    .B(_21450_),
    .Y(_21451_));
 NOR2x2_ASAP7_75t_R _29973_ (.A(net2820),
    .B(_21447_),
    .Y(_21452_));
 NOR2x1_ASAP7_75t_R _29974_ (.A(_21446_),
    .B(net3239),
    .Y(_21453_));
 XOR2x2_ASAP7_75t_R _29975_ (.A(net2888),
    .B(_19675_),
    .Y(_21454_));
 OAI21x1_ASAP7_75t_R _29976_ (.A1(_21452_),
    .A2(_21453_),
    .B(_21454_),
    .Y(_21455_));
 AOI21x1_ASAP7_75t_R _29977_ (.A1(_21451_),
    .A2(_21455_),
    .B(net390),
    .Y(_21456_));
 OAI21x1_ASAP7_75t_R _29978_ (.A1(_21433_),
    .A2(_21456_),
    .B(_15425_),
    .Y(_21457_));
 NOR2x1_ASAP7_75t_R _29979_ (.A(net391),
    .B(_00906_),
    .Y(_21458_));
 OAI21x1_ASAP7_75t_R _29980_ (.A1(_21453_),
    .A2(_21452_),
    .B(_21450_),
    .Y(_21459_));
 OAI21x1_ASAP7_75t_R _29981_ (.A1(_21448_),
    .A2(_21449_),
    .B(_21454_),
    .Y(_21460_));
 AOI21x1_ASAP7_75t_R _29982_ (.A1(_21459_),
    .A2(_21460_),
    .B(net390),
    .Y(_21461_));
 OAI21x1_ASAP7_75t_R _29983_ (.A1(_21458_),
    .A2(_21461_),
    .B(net3545),
    .Y(_21462_));
 NAND2x1_ASAP7_75t_R _29984_ (.A(_21462_),
    .B(_21457_),
    .Y(_00090_));
 TAPCELL_ASAP7_75t_R TAP_817 ();
 AND2x2_ASAP7_75t_R _29986_ (.A(net390),
    .B(_00905_),
    .Y(_21464_));
 INVx1_ASAP7_75t_R _29987_ (.A(_19575_),
    .Y(_21465_));
 NOR2x2_ASAP7_75t_R _29988_ (.A(_19576_),
    .B(_21465_),
    .Y(_21466_));
 XOR2x2_ASAP7_75t_R _29989_ (.A(_19675_),
    .B(_19252_),
    .Y(_21467_));
 XOR2x1_ASAP7_75t_R _29990_ (.A(_21467_),
    .Y(_21468_),
    .B(_19763_));
 NAND2x1_ASAP7_75t_R _29991_ (.A(_21466_),
    .B(_21468_),
    .Y(_21469_));
 NOR2x1_ASAP7_75t_R _29992_ (.A(_21466_),
    .B(_21468_),
    .Y(_21470_));
 INVx1_ASAP7_75t_R _29993_ (.A(_21470_),
    .Y(_21471_));
 AOI21x1_ASAP7_75t_R _29994_ (.A1(_21469_),
    .A2(_21471_),
    .B(net390),
    .Y(_21472_));
 OAI21x1_ASAP7_75t_R _29995_ (.A1(_21464_),
    .A2(_21472_),
    .B(_15427_),
    .Y(_21473_));
 INVx1_ASAP7_75t_R _29996_ (.A(_21466_),
    .Y(_21474_));
 INVx3_ASAP7_75t_R _29997_ (.A(_19763_),
    .Y(_21475_));
 XOR2x1_ASAP7_75t_R _29998_ (.A(net2528),
    .Y(_21476_),
    .B(_21475_));
 NOR2x1_ASAP7_75t_R _29999_ (.A(_21474_),
    .B(_21476_),
    .Y(_21477_));
 TAPCELL_ASAP7_75t_R TAP_816 ();
 OAI21x1_ASAP7_75t_R _30001_ (.A1(_21470_),
    .A2(_21477_),
    .B(net391),
    .Y(_21479_));
 INVx1_ASAP7_75t_R _30002_ (.A(_21464_),
    .Y(_21480_));
 NAND3x1_ASAP7_75t_R _30003_ (.A(_21479_),
    .B(_00442_),
    .C(_21480_),
    .Y(_21481_));
 NAND2x1_ASAP7_75t_R _30004_ (.A(_21481_),
    .B(_21473_),
    .Y(_00091_));
 TAPCELL_ASAP7_75t_R TAP_815 ();
 NOR2x1_ASAP7_75t_R _30006_ (.A(net391),
    .B(_00904_),
    .Y(_21483_));
 XOR2x2_ASAP7_75t_R _30007_ (.A(_19764_),
    .B(_20267_),
    .Y(_21484_));
 XOR2x2_ASAP7_75t_R _30008_ (.A(_19560_),
    .B(_21420_),
    .Y(_21485_));
 NOR2x2_ASAP7_75t_R _30009_ (.A(_19960_),
    .B(_19963_),
    .Y(_21486_));
 XNOR2x1_ASAP7_75t_R _30010_ (.B(_21486_),
    .Y(_21487_),
    .A(_21485_));
 NAND2x1_ASAP7_75t_R _30011_ (.A(_21484_),
    .B(_21487_),
    .Y(_21488_));
 XOR2x1_ASAP7_75t_R _30012_ (.A(_21486_),
    .Y(_21489_),
    .B(_21485_));
 INVx2_ASAP7_75t_R _30013_ (.A(_21484_),
    .Y(_21490_));
 NAND2x1_ASAP7_75t_R _30014_ (.A(_21489_),
    .B(_21490_),
    .Y(_21491_));
 AOI21x1_ASAP7_75t_R _30015_ (.A1(_21488_),
    .A2(_21491_),
    .B(net390),
    .Y(_21492_));
 OAI21x1_ASAP7_75t_R _30016_ (.A1(_21483_),
    .A2(_21492_),
    .B(_00441_),
    .Y(_21493_));
 TAPCELL_ASAP7_75t_R TAP_814 ();
 AND2x2_ASAP7_75t_R _30018_ (.A(net390),
    .B(_00904_),
    .Y(_21495_));
 NAND2x1_ASAP7_75t_R _30019_ (.A(_21484_),
    .B(_21489_),
    .Y(_21496_));
 NAND2x1_ASAP7_75t_R _30020_ (.A(_21490_),
    .B(_21487_),
    .Y(_21497_));
 AOI21x1_ASAP7_75t_R _30021_ (.A1(_21496_),
    .A2(_21497_),
    .B(net390),
    .Y(_21498_));
 OAI21x1_ASAP7_75t_R _30022_ (.A1(_21495_),
    .A2(_21498_),
    .B(_15433_),
    .Y(_21499_));
 NAND2x2_ASAP7_75t_R _30023_ (.A(_21493_),
    .B(_21499_),
    .Y(_00092_));
 NOR2x1_ASAP7_75t_R _30024_ (.A(net391),
    .B(_00903_),
    .Y(_21500_));
 INVx1_ASAP7_75t_R _30025_ (.A(_21500_),
    .Y(_21501_));
 XOR2x2_ASAP7_75t_R _30026_ (.A(_20049_),
    .B(_21420_),
    .Y(_21502_));
 INVx2_ASAP7_75t_R _30027_ (.A(_21502_),
    .Y(_21503_));
 NOR2x1_ASAP7_75t_R _30028_ (.A(_20437_),
    .B(_21503_),
    .Y(_21504_));
 NOR2x1_ASAP7_75t_R _30029_ (.A(net2276),
    .B(_20449_),
    .Y(_21505_));
 NOR2x1_ASAP7_75t_R _30030_ (.A(_19143_),
    .B(net2812),
    .Y(_21506_));
 NOR2x1_ASAP7_75t_R _30031_ (.A(_18742_),
    .B(_20275_),
    .Y(_21507_));
 OAI21x1_ASAP7_75t_R _30032_ (.A1(_21506_),
    .A2(_21507_),
    .B(_20818_),
    .Y(_21508_));
 INVx6_ASAP7_75t_R _30033_ (.A(_20818_),
    .Y(_21509_));
 OAI21x1_ASAP7_75t_R _30034_ (.A1(_20268_),
    .A2(_20276_),
    .B(_21509_),
    .Y(_21510_));
 NAND2x1_ASAP7_75t_R _30035_ (.A(_21508_),
    .B(_21510_),
    .Y(_21511_));
 OAI21x1_ASAP7_75t_R _30036_ (.A1(_21504_),
    .A2(_21505_),
    .B(_21511_),
    .Y(_21512_));
 NOR2x1_ASAP7_75t_R _30037_ (.A(_20449_),
    .B(_21503_),
    .Y(_21513_));
 NOR2x1_ASAP7_75t_R _30038_ (.A(net2276),
    .B(_20437_),
    .Y(_21514_));
 NAND2x1_ASAP7_75t_R _30039_ (.A(net2812),
    .B(_18742_),
    .Y(_21515_));
 NAND2x1_ASAP7_75t_R _30040_ (.A(net2885),
    .B(_20275_),
    .Y(_21516_));
 AOI21x1_ASAP7_75t_R _30041_ (.A1(_21515_),
    .A2(_21516_),
    .B(_20818_),
    .Y(_21517_));
 NAND2x1_ASAP7_75t_R _30042_ (.A(net2885),
    .B(net2812),
    .Y(_21518_));
 INVx1_ASAP7_75t_R _30043_ (.A(_21506_),
    .Y(_21519_));
 AOI21x1_ASAP7_75t_R _30044_ (.A1(_21518_),
    .A2(_21519_),
    .B(_21509_),
    .Y(_21520_));
 NOR2x1_ASAP7_75t_R _30045_ (.A(_21517_),
    .B(_21520_),
    .Y(_21521_));
 OAI21x1_ASAP7_75t_R _30046_ (.A1(_21513_),
    .A2(_21514_),
    .B(_21521_),
    .Y(_21522_));
 AOI21x1_ASAP7_75t_R _30047_ (.A1(_21512_),
    .A2(_21522_),
    .B(net390),
    .Y(_21523_));
 INVx1_ASAP7_75t_R _30048_ (.A(_21523_),
    .Y(_21524_));
 AOI21x1_ASAP7_75t_R _30049_ (.A1(_21501_),
    .A2(_21524_),
    .B(_00440_),
    .Y(_21525_));
 NOR3x1_ASAP7_75t_R _30050_ (.A(_21523_),
    .B(_15400_),
    .C(_21500_),
    .Y(_21526_));
 NOR2x1_ASAP7_75t_R _30051_ (.A(_21525_),
    .B(_21526_),
    .Y(_00093_));
 AND2x2_ASAP7_75t_R _30052_ (.A(net390),
    .B(_00902_),
    .Y(_21527_));
 XNOR2x2_ASAP7_75t_R _30053_ (.A(_20544_),
    .B(_20624_),
    .Y(_21528_));
 NAND2x2_ASAP7_75t_R _30054_ (.A(net2537),
    .B(_21528_),
    .Y(_21529_));
 NAND3x2_ASAP7_75t_R _30055_ (.B(_20147_),
    .C(_20159_),
    .Y(_21530_),
    .A(_20167_));
 INVx1_ASAP7_75t_R _30056_ (.A(_20122_),
    .Y(_21531_));
 NOR2x1_ASAP7_75t_R _30057_ (.A(_20130_),
    .B(_21531_),
    .Y(_21532_));
 NAND2x1_ASAP7_75t_R _30058_ (.A(_20107_),
    .B(_21532_),
    .Y(_21533_));
 NOR2x2_ASAP7_75t_R _30059_ (.A(_21530_),
    .B(_21533_),
    .Y(_21534_));
 XOR2x2_ASAP7_75t_R _30060_ (.A(_20624_),
    .B(_20544_),
    .Y(_21535_));
 NAND2x1_ASAP7_75t_R _30061_ (.A(_21534_),
    .B(_21535_),
    .Y(_21536_));
 XOR2x1_ASAP7_75t_R _30062_ (.A(net2168),
    .Y(_21537_),
    .B(net2800));
 AO21x1_ASAP7_75t_R _30063_ (.A1(_21529_),
    .A2(_21536_),
    .B(_21537_),
    .Y(_21538_));
 NAND3x1_ASAP7_75t_R _30064_ (.A(_21529_),
    .B(_21536_),
    .C(_21537_),
    .Y(_21539_));
 AOI21x1_ASAP7_75t_R _30065_ (.A1(_21538_),
    .A2(_21539_),
    .B(net390),
    .Y(_21540_));
 OAI21x1_ASAP7_75t_R _30066_ (.A1(_21527_),
    .A2(_21540_),
    .B(_15457_),
    .Y(_21541_));
 NOR2x1_ASAP7_75t_R _30067_ (.A(net391),
    .B(_00902_),
    .Y(_21542_));
 INVx2_ASAP7_75t_R _30068_ (.A(_21123_),
    .Y(_21543_));
 NAND2x2_ASAP7_75t_R _30069_ (.A(_21543_),
    .B(_21528_),
    .Y(_21544_));
 NAND2x1_ASAP7_75t_R _30070_ (.A(_21123_),
    .B(_21535_),
    .Y(_21545_));
 XOR2x1_ASAP7_75t_R _30071_ (.A(net2800),
    .Y(_21546_),
    .B(net2537));
 AO21x1_ASAP7_75t_R _30072_ (.A1(_21544_),
    .A2(_21545_),
    .B(_21546_),
    .Y(_21547_));
 NAND3x1_ASAP7_75t_R _30073_ (.A(_21544_),
    .B(_21545_),
    .C(_21546_),
    .Y(_21548_));
 AOI21x1_ASAP7_75t_R _30074_ (.A1(_21547_),
    .A2(_21548_),
    .B(net390),
    .Y(_21549_));
 OAI21x1_ASAP7_75t_R _30075_ (.A1(_21542_),
    .A2(_21549_),
    .B(_00439_),
    .Y(_21550_));
 NAND2x1_ASAP7_75t_R _30076_ (.A(_21550_),
    .B(_21541_),
    .Y(_00094_));
 TAPCELL_ASAP7_75t_R TAP_813 ();
 NOR2x2_ASAP7_75t_R _30078_ (.A(net391),
    .B(_00901_),
    .Y(_21552_));
 NAND2x2_ASAP7_75t_R _30079_ (.A(_21211_),
    .B(_21178_),
    .Y(_21553_));
 NOR2x2_ASAP7_75t_R _30080_ (.A(_19121_),
    .B(_21553_),
    .Y(_21554_));
 AOI21x1_ASAP7_75t_R _30081_ (.A1(_20969_),
    .A2(_20968_),
    .B(_21554_),
    .Y(_21555_));
 INVx1_ASAP7_75t_R _30082_ (.A(_21555_),
    .Y(_21556_));
 NAND2x1_ASAP7_75t_R _30083_ (.A(_20899_),
    .B(_21131_),
    .Y(_21557_));
 NAND2x1_ASAP7_75t_R _30084_ (.A(_20967_),
    .B(_21127_),
    .Y(_21558_));
 AOI21x1_ASAP7_75t_R _30085_ (.A1(_21557_),
    .A2(_21558_),
    .B(net2428),
    .Y(_21559_));
 INVx1_ASAP7_75t_R _30086_ (.A(_21559_),
    .Y(_21560_));
 XOR2x1_ASAP7_75t_R _30087_ (.A(net2168),
    .Y(_21561_),
    .B(_20734_));
 INVx1_ASAP7_75t_R _30088_ (.A(_21561_),
    .Y(_21562_));
 AOI21x1_ASAP7_75t_R _30089_ (.A1(_21556_),
    .A2(_21560_),
    .B(_21562_),
    .Y(_21563_));
 INVx1_ASAP7_75t_R _30090_ (.A(_21563_),
    .Y(_21564_));
 NAND3x1_ASAP7_75t_R _30091_ (.A(_21560_),
    .B(_21556_),
    .C(_21562_),
    .Y(_21565_));
 AOI21x1_ASAP7_75t_R _30092_ (.A1(_21564_),
    .A2(_21565_),
    .B(net390),
    .Y(_21566_));
 OAI21x1_ASAP7_75t_R _30093_ (.A1(_21552_),
    .A2(_21566_),
    .B(_00438_),
    .Y(_21567_));
 NOR3x1_ASAP7_75t_R _30094_ (.A(_21559_),
    .B(_21555_),
    .C(_21561_),
    .Y(_21568_));
 OAI21x1_ASAP7_75t_R _30095_ (.A1(_21563_),
    .A2(_21568_),
    .B(net391),
    .Y(_21569_));
 INVx1_ASAP7_75t_R _30096_ (.A(_21552_),
    .Y(_21570_));
 NAND3x1_ASAP7_75t_R _30097_ (.A(_21569_),
    .B(_15402_),
    .C(_21570_),
    .Y(_21571_));
 NAND2x1_ASAP7_75t_R _30098_ (.A(_21571_),
    .B(_21567_),
    .Y(_00095_));
 XOR2x1_ASAP7_75t_R _30099_ (.A(_21046_),
    .Y(_21572_),
    .B(_18742_));
 XOR2x1_ASAP7_75t_R _30100_ (.A(_21294_),
    .Y(_21573_),
    .B(_21572_));
 NOR2x1_ASAP7_75t_R _30101_ (.A(net391),
    .B(_00900_),
    .Y(_21574_));
 AO21x1_ASAP7_75t_R _30102_ (.A1(_21573_),
    .A2(net391),
    .B(_21574_),
    .Y(_21575_));
 XOR2x2_ASAP7_75t_R _30103_ (.A(_21575_),
    .B(_15411_),
    .Y(_00096_));
 TAPCELL_ASAP7_75t_R TAP_812 ();
 NOR2x2_ASAP7_75t_R _30105_ (.A(net391),
    .B(_00899_),
    .Y(_21577_));
 NAND2x2_ASAP7_75t_R _30106_ (.A(_19120_),
    .B(_19105_),
    .Y(_21578_));
 INVx5_ASAP7_75t_R _30107_ (.A(_21292_),
    .Y(_21579_));
 XOR2x1_ASAP7_75t_R _30108_ (.A(_21388_),
    .Y(_21580_),
    .B(_21579_));
 NAND2x2_ASAP7_75t_R _30109_ (.A(_21578_),
    .B(_21580_),
    .Y(_21581_));
 NOR2x2_ASAP7_75t_R _30110_ (.A(_19121_),
    .B(_19134_),
    .Y(_21582_));
 XOR2x1_ASAP7_75t_R _30111_ (.A(_21388_),
    .Y(_21583_),
    .B(net2363));
 NAND2x1_ASAP7_75t_R _30112_ (.A(_21582_),
    .B(_21583_),
    .Y(_21584_));
 AOI21x1_ASAP7_75t_R _30113_ (.A1(_21581_),
    .A2(_21584_),
    .B(_21446_),
    .Y(_21585_));
 INVx1_ASAP7_75t_R _30114_ (.A(_21585_),
    .Y(_21586_));
 NAND3x1_ASAP7_75t_R _30115_ (.A(_21581_),
    .B(_21584_),
    .C(_21446_),
    .Y(_21587_));
 AOI21x1_ASAP7_75t_R _30116_ (.A1(_21586_),
    .A2(_21587_),
    .B(net390),
    .Y(_21588_));
 OAI21x1_ASAP7_75t_R _30117_ (.A1(_21577_),
    .A2(_21588_),
    .B(net2208),
    .Y(_21589_));
 NAND2x1_ASAP7_75t_R _30118_ (.A(_21390_),
    .B(_21578_),
    .Y(_21590_));
 NAND2x1_ASAP7_75t_R _30119_ (.A(_21388_),
    .B(_21582_),
    .Y(_21591_));
 AO21x1_ASAP7_75t_R _30120_ (.A1(_21590_),
    .A2(_21591_),
    .B(_21579_),
    .Y(_21592_));
 NAND3x1_ASAP7_75t_R _30121_ (.A(_21590_),
    .B(_21591_),
    .C(_21579_),
    .Y(_21593_));
 AOI21x1_ASAP7_75t_R _30122_ (.A1(_21592_),
    .A2(_21593_),
    .B(_21447_),
    .Y(_21594_));
 OAI21x1_ASAP7_75t_R _30123_ (.A1(_21585_),
    .A2(_21594_),
    .B(net391),
    .Y(_21595_));
 INVx1_ASAP7_75t_R _30124_ (.A(_21577_),
    .Y(_21596_));
 NAND3x1_ASAP7_75t_R _30125_ (.A(_21595_),
    .B(_16287_),
    .C(_21596_),
    .Y(_21597_));
 NAND2x1_ASAP7_75t_R _30126_ (.A(_21589_),
    .B(_21597_),
    .Y(_00057_));
 NOR2x2_ASAP7_75t_R _30127_ (.A(net391),
    .B(_00898_),
    .Y(_21598_));
 AOI21x1_ASAP7_75t_R _30128_ (.A1(_18279_),
    .A2(_18506_),
    .B(net2342),
    .Y(_21599_));
 NOR3x1_ASAP7_75t_R _30129_ (.A(_21444_),
    .B(_21382_),
    .C(_20657_),
    .Y(_21600_));
 OAI21x1_ASAP7_75t_R _30130_ (.A1(_21599_),
    .A2(_21600_),
    .B(_19257_),
    .Y(_21601_));
 OAI21x1_ASAP7_75t_R _30131_ (.A1(_21434_),
    .A2(_21445_),
    .B(_19252_),
    .Y(_21602_));
 NAND2x2_ASAP7_75t_R _30132_ (.A(_21601_),
    .B(_21602_),
    .Y(_21603_));
 INVx1_ASAP7_75t_R _30133_ (.A(_21603_),
    .Y(_21604_));
 INVx1_ASAP7_75t_R _30134_ (.A(_18191_),
    .Y(_21605_));
 OAI21x1_ASAP7_75t_R _30135_ (.A1(_20642_),
    .A2(_21605_),
    .B(_21579_),
    .Y(_21606_));
 NAND3x2_ASAP7_75t_R _30136_ (.B(_21292_),
    .C(net2557),
    .Y(_21607_),
    .A(_18191_));
 NAND2x2_ASAP7_75t_R _30137_ (.A(_21606_),
    .B(_21607_),
    .Y(_21608_));
 XOR2x1_ASAP7_75t_R _30138_ (.A(_19676_),
    .Y(_21609_),
    .B(_21608_));
 NAND2x1_ASAP7_75t_R _30139_ (.A(_21609_),
    .B(_21604_),
    .Y(_21610_));
 INVx1_ASAP7_75t_R _30140_ (.A(_19676_),
    .Y(_21611_));
 NAND2x1_ASAP7_75t_R _30141_ (.A(_21608_),
    .B(_21611_),
    .Y(_21612_));
 INVx2_ASAP7_75t_R _30142_ (.A(_21608_),
    .Y(_21613_));
 NAND2x2_ASAP7_75t_R _30143_ (.A(_19676_),
    .B(_21613_),
    .Y(_21614_));
 NAND3x1_ASAP7_75t_R _30144_ (.A(net2822),
    .B(_21612_),
    .C(_21614_),
    .Y(_21615_));
 AOI21x1_ASAP7_75t_R _30145_ (.A1(_21610_),
    .A2(_21615_),
    .B(net390),
    .Y(_21616_));
 OAI21x1_ASAP7_75t_R _30146_ (.A1(_21598_),
    .A2(_21616_),
    .B(net1854),
    .Y(_21617_));
 AOI21x1_ASAP7_75t_R _30147_ (.A1(_21614_),
    .A2(_21612_),
    .B(net2822),
    .Y(_21618_));
 NOR2x1_ASAP7_75t_R _30148_ (.A(_21604_),
    .B(_21609_),
    .Y(_21619_));
 OAI21x1_ASAP7_75t_R _30149_ (.A1(_21618_),
    .A2(_21619_),
    .B(net391),
    .Y(_21620_));
 INVx1_ASAP7_75t_R _30150_ (.A(_21598_),
    .Y(_21621_));
 NAND3x2_ASAP7_75t_R _30151_ (.B(_16262_),
    .C(_21621_),
    .Y(_21622_),
    .A(_21620_));
 NAND2x2_ASAP7_75t_R _30152_ (.A(_21622_),
    .B(_21617_),
    .Y(_00058_));
 AND2x2_ASAP7_75t_R _30153_ (.A(net390),
    .B(_00897_),
    .Y(_21623_));
 NOR2x1_ASAP7_75t_R _30154_ (.A(net3317),
    .B(net1308),
    .Y(_21624_));
 INVx4_ASAP7_75t_R _30155_ (.A(net3317),
    .Y(_21625_));
 NAND2x1_ASAP7_75t_R _30156_ (.A(_18967_),
    .B(_18912_),
    .Y(_21626_));
 NOR2x2_ASAP7_75t_R _30157_ (.A(_20642_),
    .B(_21626_),
    .Y(_21627_));
 NOR2x1_ASAP7_75t_R _30158_ (.A(_21625_),
    .B(_21627_),
    .Y(_21628_));
 OAI21x1_ASAP7_75t_R _30159_ (.A1(_21624_),
    .A2(_21628_),
    .B(_19763_),
    .Y(_21629_));
 NAND2x1_ASAP7_75t_R _30160_ (.A(net3317),
    .B(_21627_),
    .Y(_21630_));
 NAND2x1_ASAP7_75t_R _30161_ (.A(_21625_),
    .B(net1308),
    .Y(_21631_));
 AO21x1_ASAP7_75t_R _30162_ (.A1(_21630_),
    .A2(_21631_),
    .B(_19763_),
    .Y(_21632_));
 XOR2x1_ASAP7_75t_R _30163_ (.A(_19252_),
    .Y(_21633_),
    .B(_19560_));
 AOI21x1_ASAP7_75t_R _30164_ (.A1(_21629_),
    .A2(_21632_),
    .B(_21633_),
    .Y(_21634_));
 AO21x1_ASAP7_75t_R _30165_ (.A1(_21630_),
    .A2(_21631_),
    .B(_21475_),
    .Y(_21635_));
 XOR2x1_ASAP7_75t_R _30166_ (.A(net1308),
    .Y(_21636_),
    .B(_21625_));
 NAND2x1_ASAP7_75t_R _30167_ (.A(_21475_),
    .B(_21636_),
    .Y(_21637_));
 INVx1_ASAP7_75t_R _30168_ (.A(_21633_),
    .Y(_21638_));
 AOI21x1_ASAP7_75t_R _30169_ (.A1(_21635_),
    .A2(_21637_),
    .B(_21638_),
    .Y(_21639_));
 OAI21x1_ASAP7_75t_R _30170_ (.A1(_21634_),
    .A2(_21639_),
    .B(net391),
    .Y(_21640_));
 INVx1_ASAP7_75t_R _30171_ (.A(_21640_),
    .Y(_21641_));
 OAI21x1_ASAP7_75t_R _30172_ (.A1(_21623_),
    .A2(_21641_),
    .B(_16286_),
    .Y(_21642_));
 INVx1_ASAP7_75t_R _30173_ (.A(_21623_),
    .Y(_21643_));
 NAND3x2_ASAP7_75t_R _30174_ (.B(net3485),
    .C(_21643_),
    .Y(_21644_),
    .A(_21640_));
 NAND2x2_ASAP7_75t_R _30175_ (.A(_21642_),
    .B(_21644_),
    .Y(_00059_));
 NOR2x1_ASAP7_75t_R _30176_ (.A(net391),
    .B(_00896_),
    .Y(_21645_));
 XOR2x2_ASAP7_75t_R _30177_ (.A(net2141),
    .B(_20049_),
    .Y(_21646_));
 INVx2_ASAP7_75t_R _30178_ (.A(_21646_),
    .Y(_21647_));
 NAND2x2_ASAP7_75t_R _30179_ (.A(_21485_),
    .B(_21647_),
    .Y(_21648_));
 INVx1_ASAP7_75t_R _30180_ (.A(_21485_),
    .Y(_21649_));
 NAND2x1_ASAP7_75t_R _30181_ (.A(_21646_),
    .B(_21649_),
    .Y(_21650_));
 NOR2x1_ASAP7_75t_R _30182_ (.A(_21292_),
    .B(_19574_),
    .Y(_21651_));
 NOR2x1_ASAP7_75t_R _30183_ (.A(_21579_),
    .B(_19457_),
    .Y(_21652_));
 OAI21x1_ASAP7_75t_R _30184_ (.A1(_21651_),
    .A2(_21652_),
    .B(_20275_),
    .Y(_21653_));
 NOR2x2_ASAP7_75t_R _30185_ (.A(_21579_),
    .B(_19574_),
    .Y(_21654_));
 NOR2x1_ASAP7_75t_R _30186_ (.A(_21292_),
    .B(_19457_),
    .Y(_21655_));
 OAI21x1_ASAP7_75t_R _30187_ (.A1(_21654_),
    .A2(_21655_),
    .B(_20267_),
    .Y(_21656_));
 NAND2x2_ASAP7_75t_R _30188_ (.A(_21653_),
    .B(_21656_),
    .Y(_21657_));
 AOI21x1_ASAP7_75t_R _30189_ (.A1(_21648_),
    .A2(_21650_),
    .B(_21657_),
    .Y(_21658_));
 INVx1_ASAP7_75t_R _30190_ (.A(_21658_),
    .Y(_21659_));
 NAND3x1_ASAP7_75t_R _30191_ (.A(_21657_),
    .B(_21648_),
    .C(_21650_),
    .Y(_21660_));
 AOI21x1_ASAP7_75t_R _30192_ (.A1(_21659_),
    .A2(_21660_),
    .B(net390),
    .Y(_21661_));
 OAI21x1_ASAP7_75t_R _30193_ (.A1(_21645_),
    .A2(_21661_),
    .B(net3490),
    .Y(_21662_));
 INVx1_ASAP7_75t_R _30194_ (.A(_21657_),
    .Y(_21663_));
 XOR2x1_ASAP7_75t_R _30195_ (.A(_21646_),
    .Y(_21664_),
    .B(_21485_));
 NOR2x1_ASAP7_75t_R _30196_ (.A(_21663_),
    .B(_21664_),
    .Y(_21665_));
 OAI21x1_ASAP7_75t_R _30197_ (.A1(_21658_),
    .A2(_21665_),
    .B(net391),
    .Y(_21666_));
 INVx1_ASAP7_75t_R _30198_ (.A(_21645_),
    .Y(_21667_));
 NAND3x1_ASAP7_75t_R _30199_ (.A(_21666_),
    .B(_16276_),
    .C(_21667_),
    .Y(_21668_));
 NAND2x1_ASAP7_75t_R _30200_ (.A(_21668_),
    .B(_21662_),
    .Y(_00060_));
 AND2x2_ASAP7_75t_R _30201_ (.A(net390),
    .B(_00895_),
    .Y(_21669_));
 XOR2x2_ASAP7_75t_R _30202_ (.A(_19962_),
    .B(_21292_),
    .Y(_21670_));
 XOR2x1_ASAP7_75t_R _30203_ (.A(_21670_),
    .Y(_21671_),
    .B(_21509_));
 XOR2x2_ASAP7_75t_R _30204_ (.A(_20352_),
    .B(_20170_),
    .Y(_21672_));
 XOR2x1_ASAP7_75t_R _30205_ (.A(_21672_),
    .Y(_21673_),
    .B(_21502_));
 NAND2x1_ASAP7_75t_R _30206_ (.A(_21671_),
    .B(_21673_),
    .Y(_21674_));
 XOR2x2_ASAP7_75t_R _30207_ (.A(_19962_),
    .B(_21579_),
    .Y(_21675_));
 XOR2x1_ASAP7_75t_R _30208_ (.A(_21675_),
    .Y(_21676_),
    .B(_21509_));
 XNOR2x1_ASAP7_75t_R _30209_ (.B(_21672_),
    .Y(_21677_),
    .A(_21502_));
 NAND2x1_ASAP7_75t_R _30210_ (.A(_21676_),
    .B(_21677_),
    .Y(_21678_));
 AOI21x1_ASAP7_75t_R _30211_ (.A1(_21674_),
    .A2(_21678_),
    .B(net390),
    .Y(_21679_));
 OAI21x1_ASAP7_75t_R _30212_ (.A1(_21669_),
    .A2(_21679_),
    .B(_16339_),
    .Y(_21680_));
 NOR2x1_ASAP7_75t_R _30213_ (.A(net391),
    .B(_00895_),
    .Y(_21681_));
 XOR2x1_ASAP7_75t_R _30214_ (.A(_21502_),
    .Y(_21682_),
    .B(_21509_));
 XOR2x1_ASAP7_75t_R _30215_ (.A(_21672_),
    .Y(_21683_),
    .B(_21675_));
 NAND2x1_ASAP7_75t_R _30216_ (.A(_21682_),
    .B(_21683_),
    .Y(_21684_));
 XOR2x1_ASAP7_75t_R _30217_ (.A(_21672_),
    .Y(_21685_),
    .B(_21670_));
 INVx1_ASAP7_75t_R _30218_ (.A(_21682_),
    .Y(_21686_));
 NAND2x1_ASAP7_75t_R _30219_ (.A(_21686_),
    .B(_21685_),
    .Y(_21687_));
 AOI21x1_ASAP7_75t_R _30220_ (.A1(_21684_),
    .A2(_21687_),
    .B(net390),
    .Y(_21688_));
 OAI21x1_ASAP7_75t_R _30221_ (.A1(_21681_),
    .A2(_21688_),
    .B(net3502),
    .Y(_21689_));
 NAND2x1_ASAP7_75t_R _30222_ (.A(_21689_),
    .B(_21680_),
    .Y(_00061_));
 TAPCELL_ASAP7_75t_R TAP_811 ();
 NAND2x1_ASAP7_75t_R _30224_ (.A(_00894_),
    .B(net390),
    .Y(_21691_));
 OAI22x1_ASAP7_75t_R _30225_ (.A1(_20733_),
    .A2(_20657_),
    .B1(_20543_),
    .B2(net2145),
    .Y(_21692_));
 NAND2x2_ASAP7_75t_R _30226_ (.A(_20544_),
    .B(_20734_),
    .Y(_21693_));
 AOI21x1_ASAP7_75t_R _30227_ (.A1(_21692_),
    .A2(_21693_),
    .B(net2167),
    .Y(_21694_));
 NAND3x2_ASAP7_75t_R _30228_ (.B(_21692_),
    .C(net2167),
    .Y(_21695_),
    .A(_21693_));
 INVx1_ASAP7_75t_R _30229_ (.A(_21695_),
    .Y(_21696_));
 NAND2x2_ASAP7_75t_R _30230_ (.A(_20448_),
    .B(_20170_),
    .Y(_21697_));
 NAND2x2_ASAP7_75t_R _30231_ (.A(net3238),
    .B(_21534_),
    .Y(_21698_));
 NAND2x2_ASAP7_75t_R _30232_ (.A(_21697_),
    .B(_21698_),
    .Y(_21699_));
 INVx1_ASAP7_75t_R _30233_ (.A(_21699_),
    .Y(_21700_));
 OAI21x1_ASAP7_75t_R _30234_ (.A1(_21694_),
    .A2(_21696_),
    .B(_21700_),
    .Y(_21701_));
 INVx1_ASAP7_75t_R _30235_ (.A(_21701_),
    .Y(_21702_));
 INVx1_ASAP7_75t_R _30236_ (.A(_21694_),
    .Y(_21703_));
 AND3x1_ASAP7_75t_R _30237_ (.A(_21695_),
    .B(_21703_),
    .C(_21699_),
    .Y(_21704_));
 TAPCELL_ASAP7_75t_R TAP_810 ();
 OAI21x1_ASAP7_75t_R _30239_ (.A1(_21702_),
    .A2(_21704_),
    .B(net391),
    .Y(_21706_));
 AOI21x1_ASAP7_75t_R _30240_ (.A1(_21691_),
    .A2(_21706_),
    .B(_16270_),
    .Y(_21707_));
 TAPCELL_ASAP7_75t_R TAP_809 ();
 OR2x2_ASAP7_75t_R _30242_ (.A(net391),
    .B(_00894_),
    .Y(_21709_));
 NAND3x1_ASAP7_75t_R _30243_ (.A(_21695_),
    .B(_21703_),
    .C(_21699_),
    .Y(_21710_));
 NAND3x1_ASAP7_75t_R _30244_ (.A(_21710_),
    .B(_21701_),
    .C(net391),
    .Y(_21711_));
 AOI21x1_ASAP7_75t_R _30245_ (.A1(_21709_),
    .A2(_21711_),
    .B(net3496),
    .Y(_21712_));
 NOR2x1_ASAP7_75t_R _30246_ (.A(_21712_),
    .B(_21707_),
    .Y(_00062_));
 XNOR2x2_ASAP7_75t_R _30247_ (.A(_20734_),
    .B(_20624_),
    .Y(_21713_));
 XOR2x1_ASAP7_75t_R _30248_ (.A(_21713_),
    .Y(_21714_),
    .B(_21554_));
 NAND2x1_ASAP7_75t_R _30249_ (.A(_21132_),
    .B(_21714_),
    .Y(_21715_));
 INVx1_ASAP7_75t_R _30250_ (.A(_21132_),
    .Y(_21716_));
 XOR2x1_ASAP7_75t_R _30251_ (.A(_21713_),
    .Y(_21717_),
    .B(net2428));
 TAPCELL_ASAP7_75t_R TAP_808 ();
 AOI21x1_ASAP7_75t_R _30253_ (.A1(_21716_),
    .A2(_21717_),
    .B(net390),
    .Y(_21719_));
 AND2x2_ASAP7_75t_R _30254_ (.A(net390),
    .B(_00893_),
    .Y(_21720_));
 AOI21x1_ASAP7_75t_R _30255_ (.A1(_21715_),
    .A2(_21719_),
    .B(_21720_),
    .Y(_21721_));
 XOR2x1_ASAP7_75t_R _30256_ (.A(_21721_),
    .Y(_00063_),
    .B(_16268_));
 NAND2x1_ASAP7_75t_R _30257_ (.A(_00892_),
    .B(net390),
    .Y(_21722_));
 XOR2x2_ASAP7_75t_R _30258_ (.A(_20967_),
    .B(_21046_),
    .Y(_21723_));
 NAND2x2_ASAP7_75t_R _30259_ (.A(_21382_),
    .B(_21723_),
    .Y(_21724_));
 INVx3_ASAP7_75t_R _30260_ (.A(_21723_),
    .Y(_21725_));
 NAND2x2_ASAP7_75t_R _30261_ (.A(_21420_),
    .B(_21725_),
    .Y(_21726_));
 XOR2x2_ASAP7_75t_R _30262_ (.A(net2885),
    .B(net2898),
    .Y(_21727_));
 AOI21x1_ASAP7_75t_R _30263_ (.A1(_21724_),
    .A2(_21726_),
    .B(_21727_),
    .Y(_21728_));
 NAND2x2_ASAP7_75t_R _30264_ (.A(_21420_),
    .B(_21723_),
    .Y(_21729_));
 NAND2x2_ASAP7_75t_R _30265_ (.A(_21382_),
    .B(_21725_),
    .Y(_21730_));
 INVx1_ASAP7_75t_R _30266_ (.A(_21727_),
    .Y(_21731_));
 AOI21x1_ASAP7_75t_R _30267_ (.A1(_21729_),
    .A2(_21730_),
    .B(_21731_),
    .Y(_21732_));
 OAI21x1_ASAP7_75t_R _30268_ (.A1(_21728_),
    .A2(_21732_),
    .B(net391),
    .Y(_21733_));
 AOI21x1_ASAP7_75t_R _30269_ (.A1(_21722_),
    .A2(_21733_),
    .B(_16291_),
    .Y(_21734_));
 OR2x2_ASAP7_75t_R _30270_ (.A(net391),
    .B(_00892_),
    .Y(_21735_));
 AOI21x1_ASAP7_75t_R _30271_ (.A1(_21724_),
    .A2(_21726_),
    .B(_21731_),
    .Y(_21736_));
 AOI21x1_ASAP7_75t_R _30272_ (.A1(_21729_),
    .A2(_21730_),
    .B(_21727_),
    .Y(_21737_));
 OAI21x1_ASAP7_75t_R _30273_ (.A1(_21736_),
    .A2(_21737_),
    .B(net391),
    .Y(_21738_));
 AOI21x1_ASAP7_75t_R _30274_ (.A1(_21735_),
    .A2(_21738_),
    .B(_00429_),
    .Y(_21739_));
 NOR2x1_ASAP7_75t_R _30275_ (.A(_21734_),
    .B(_21739_),
    .Y(_00064_));
 AND2x2_ASAP7_75t_R _30276_ (.A(net390),
    .B(_00891_),
    .Y(_21740_));
 NAND2x2_ASAP7_75t_R _30277_ (.A(_21578_),
    .B(_21613_),
    .Y(_21741_));
 XOR2x2_ASAP7_75t_R _30278_ (.A(_18507_),
    .B(_17905_),
    .Y(_21742_));
 AO21x1_ASAP7_75t_R _30279_ (.A1(_21607_),
    .A2(_21606_),
    .B(_21578_),
    .Y(_21743_));
 NAND3x1_ASAP7_75t_R _30280_ (.A(_21741_),
    .B(_21742_),
    .C(_21743_),
    .Y(_21744_));
 AO21x1_ASAP7_75t_R _30281_ (.A1(_21741_),
    .A2(_21743_),
    .B(_21742_),
    .Y(_21745_));
 TAPCELL_ASAP7_75t_R TAP_807 ();
 AOI21x1_ASAP7_75t_R _30283_ (.A1(_21744_),
    .A2(_21745_),
    .B(net390),
    .Y(_21747_));
 OAI21x1_ASAP7_75t_R _30284_ (.A1(_21740_),
    .A2(_21747_),
    .B(_05925_),
    .Y(_21748_));
 NOR2x1_ASAP7_75t_R _30285_ (.A(net397),
    .B(_00891_),
    .Y(_21749_));
 XOR2x1_ASAP7_75t_R _30286_ (.A(_18507_),
    .Y(_21750_),
    .B(net2898));
 NAND2x1_ASAP7_75t_R _30287_ (.A(_21582_),
    .B(_21750_),
    .Y(_21751_));
 NAND2x1_ASAP7_75t_R _30288_ (.A(_21578_),
    .B(_21742_),
    .Y(_21752_));
 AO21x1_ASAP7_75t_R _30289_ (.A1(_21751_),
    .A2(_21752_),
    .B(_21608_),
    .Y(_21753_));
 NAND3x1_ASAP7_75t_R _30290_ (.A(_21751_),
    .B(_21752_),
    .C(_21608_),
    .Y(_21754_));
 AOI21x1_ASAP7_75t_R _30291_ (.A1(_21753_),
    .A2(_21754_),
    .B(net390),
    .Y(_21755_));
 OAI21x1_ASAP7_75t_R _30292_ (.A1(_21749_),
    .A2(_21755_),
    .B(net2129),
    .Y(_21756_));
 NAND2x1_ASAP7_75t_R _30293_ (.A(_21756_),
    .B(_21748_),
    .Y(_00025_));
 NOR2x2_ASAP7_75t_R _30294_ (.A(net397),
    .B(_00890_),
    .Y(_21757_));
 OAI21x1_ASAP7_75t_R _30295_ (.A1(_17920_),
    .A2(_18231_),
    .B(_18968_),
    .Y(_21758_));
 NAND3x1_ASAP7_75t_R _30296_ (.A(_17919_),
    .B(_17921_),
    .C(_21627_),
    .Y(_21759_));
 NAND2x1_ASAP7_75t_R _30297_ (.A(_21758_),
    .B(_21759_),
    .Y(_21760_));
 XNOR2x1_ASAP7_75t_R _30298_ (.B(_21467_),
    .Y(_21761_),
    .A(_21608_));
 NAND2x1_ASAP7_75t_R _30299_ (.A(_21760_),
    .B(_21761_),
    .Y(_21762_));
 NOR2x1_ASAP7_75t_R _30300_ (.A(_21760_),
    .B(_21761_),
    .Y(_21763_));
 INVx1_ASAP7_75t_R _30301_ (.A(_21763_),
    .Y(_21764_));
 AOI21x1_ASAP7_75t_R _30302_ (.A1(_21762_),
    .A2(_21764_),
    .B(net390),
    .Y(_21765_));
 OAI21x1_ASAP7_75t_R _30303_ (.A1(_21757_),
    .A2(_21765_),
    .B(net1146),
    .Y(_21766_));
 XOR2x1_ASAP7_75t_R _30304_ (.A(_21467_),
    .Y(_21767_),
    .B(_21608_));
 INVx1_ASAP7_75t_R _30305_ (.A(_21758_),
    .Y(_21768_));
 NOR3x1_ASAP7_75t_R _30306_ (.A(_18231_),
    .B(_17920_),
    .C(_18968_),
    .Y(_21769_));
 NOR2x1_ASAP7_75t_R _30307_ (.A(_21768_),
    .B(_21769_),
    .Y(_21770_));
 NOR2x1_ASAP7_75t_R _30308_ (.A(_21767_),
    .B(_21770_),
    .Y(_21771_));
 OAI21x1_ASAP7_75t_R _30309_ (.A1(_21763_),
    .A2(_21771_),
    .B(net397),
    .Y(_21772_));
 INVx1_ASAP7_75t_R _30310_ (.A(_21757_),
    .Y(_21773_));
 NAND3x1_ASAP7_75t_R _30311_ (.A(_21772_),
    .B(_06397_),
    .C(_21773_),
    .Y(_21774_));
 NAND2x1_ASAP7_75t_R _30312_ (.A(_21766_),
    .B(_21774_),
    .Y(_00026_));
 TAPCELL_ASAP7_75t_R TAP_806 ();
 AND2x2_ASAP7_75t_R _30314_ (.A(net390),
    .B(_00889_),
    .Y(_21776_));
 NOR2x2_ASAP7_75t_R _30315_ (.A(_21475_),
    .B(_18971_),
    .Y(_21777_));
 NOR2x1_ASAP7_75t_R _30316_ (.A(_19763_),
    .B(_18969_),
    .Y(_21778_));
 XOR2x2_ASAP7_75t_R _30317_ (.A(_19560_),
    .B(_19574_),
    .Y(_21779_));
 INVx1_ASAP7_75t_R _30318_ (.A(_21779_),
    .Y(_21780_));
 OAI21x1_ASAP7_75t_R _30319_ (.A1(_21777_),
    .A2(_21778_),
    .B(_21780_),
    .Y(_21781_));
 NOR2x2_ASAP7_75t_R _30320_ (.A(_19763_),
    .B(_18971_),
    .Y(_21782_));
 NOR2x1_ASAP7_75t_R _30321_ (.A(_21475_),
    .B(_18969_),
    .Y(_21783_));
 OAI21x1_ASAP7_75t_R _30322_ (.A1(_21782_),
    .A2(_21783_),
    .B(_21779_),
    .Y(_21784_));
 AOI21x1_ASAP7_75t_R _30323_ (.A1(_21781_),
    .A2(_21784_),
    .B(net390),
    .Y(_21785_));
 OAI21x1_ASAP7_75t_R _30324_ (.A1(_21776_),
    .A2(_21785_),
    .B(_05848_),
    .Y(_21786_));
 NOR2x1_ASAP7_75t_R _30325_ (.A(net397),
    .B(_00889_),
    .Y(_21787_));
 OAI21x1_ASAP7_75t_R _30326_ (.A1(_21777_),
    .A2(_21778_),
    .B(_21779_),
    .Y(_21788_));
 OAI21x1_ASAP7_75t_R _30327_ (.A1(_21782_),
    .A2(_21783_),
    .B(_21780_),
    .Y(_21789_));
 AOI21x1_ASAP7_75t_R _30328_ (.A1(_21788_),
    .A2(_21789_),
    .B(net390),
    .Y(_21790_));
 OAI21x1_ASAP7_75t_R _30329_ (.A1(_21787_),
    .A2(_21790_),
    .B(net3396),
    .Y(_21791_));
 NAND2x1_ASAP7_75t_R _30330_ (.A(_21786_),
    .B(_21791_),
    .Y(_00027_));
 XOR2x1_ASAP7_75t_R _30331_ (.A(_19688_),
    .Y(_21792_),
    .B(_20267_));
 NOR2x1_ASAP7_75t_R _30332_ (.A(_21655_),
    .B(_21654_),
    .Y(_21793_));
 XOR2x1_ASAP7_75t_R _30333_ (.A(_19962_),
    .Y(_21794_),
    .B(net2986));
 XOR2x1_ASAP7_75t_R _30334_ (.A(_21793_),
    .Y(_21795_),
    .B(_21794_));
 TAPCELL_ASAP7_75t_R TAP_805 ();
 AOI21x1_ASAP7_75t_R _30336_ (.A1(_21792_),
    .A2(_21795_),
    .B(net390),
    .Y(_21797_));
 OR2x2_ASAP7_75t_R _30337_ (.A(_21795_),
    .B(_21792_),
    .Y(_21798_));
 AND2x2_ASAP7_75t_R _30338_ (.A(net390),
    .B(_00888_),
    .Y(_21799_));
 AOI21x1_ASAP7_75t_R _30339_ (.A1(_21797_),
    .A2(_21798_),
    .B(_21799_),
    .Y(_21800_));
 XOR2x1_ASAP7_75t_R _30340_ (.A(_21800_),
    .Y(_00028_),
    .B(_06189_));
 NOR2x1_ASAP7_75t_R _30341_ (.A(net397),
    .B(_00887_),
    .Y(_21801_));
 INVx1_ASAP7_75t_R _30342_ (.A(_21801_),
    .Y(_21802_));
 NOR2x1_ASAP7_75t_R _30343_ (.A(_20088_),
    .B(_21675_),
    .Y(_21803_));
 NOR2x1_ASAP7_75t_R _30344_ (.A(_20440_),
    .B(_21670_),
    .Y(_21804_));
 AOI22x1_ASAP7_75t_R _30345_ (.A1(_20169_),
    .A2(_20133_),
    .B1(_20435_),
    .B2(_20390_),
    .Y(_21805_));
 NOR2x1_ASAP7_75t_R _30346_ (.A(net3238),
    .B(_20170_),
    .Y(_21806_));
 OAI21x1_ASAP7_75t_R _30347_ (.A1(_21805_),
    .A2(_21806_),
    .B(_20818_),
    .Y(_21807_));
 NOR2x1_ASAP7_75t_R _30348_ (.A(_20448_),
    .B(_20170_),
    .Y(_21808_));
 NOR2x1_ASAP7_75t_R _30349_ (.A(_20436_),
    .B(_21534_),
    .Y(_21809_));
 OAI21x1_ASAP7_75t_R _30350_ (.A1(_21808_),
    .A2(_21809_),
    .B(_21509_),
    .Y(_21810_));
 NAND2x1_ASAP7_75t_R _30351_ (.A(_21807_),
    .B(_21810_),
    .Y(_21811_));
 OAI21x1_ASAP7_75t_R _30352_ (.A1(_21803_),
    .A2(_21804_),
    .B(_21811_),
    .Y(_21812_));
 NOR2x1_ASAP7_75t_R _30353_ (.A(_20440_),
    .B(_21675_),
    .Y(_21813_));
 NOR2x1_ASAP7_75t_R _30354_ (.A(_20088_),
    .B(_21670_),
    .Y(_21814_));
 AOI21x1_ASAP7_75t_R _30355_ (.A1(_21697_),
    .A2(_21698_),
    .B(net2800),
    .Y(_21815_));
 NAND2x1_ASAP7_75t_R _30356_ (.A(_20436_),
    .B(_20170_),
    .Y(_21816_));
 NAND2x1_ASAP7_75t_R _30357_ (.A(_20448_),
    .B(_21534_),
    .Y(_21817_));
 AOI21x1_ASAP7_75t_R _30358_ (.A1(_21816_),
    .A2(_21817_),
    .B(_21509_),
    .Y(_21818_));
 NOR2x1_ASAP7_75t_R _30359_ (.A(_21818_),
    .B(_21815_),
    .Y(_21819_));
 OAI21x1_ASAP7_75t_R _30360_ (.A1(_21813_),
    .A2(_21814_),
    .B(_21819_),
    .Y(_21820_));
 AOI21x1_ASAP7_75t_R _30361_ (.A1(_21812_),
    .A2(_21820_),
    .B(net390),
    .Y(_21821_));
 INVx1_ASAP7_75t_R _30362_ (.A(_21821_),
    .Y(_21822_));
 AOI21x1_ASAP7_75t_R _30363_ (.A1(_21802_),
    .A2(_21822_),
    .B(_00424_),
    .Y(_21823_));
 NOR3x1_ASAP7_75t_R _30364_ (.A(_21821_),
    .B(_05749_),
    .C(_21801_),
    .Y(_21824_));
 NOR2x1_ASAP7_75t_R _30365_ (.A(_21824_),
    .B(_21823_),
    .Y(_00029_));
 NOR2x2_ASAP7_75t_R _30366_ (.A(net397),
    .B(_00886_),
    .Y(_21825_));
 INVx1_ASAP7_75t_R _30367_ (.A(_21825_),
    .Y(_21826_));
 AOI22x1_ASAP7_75t_R _30368_ (.A1(_20746_),
    .A2(_18279_),
    .B1(_20623_),
    .B2(_17974_),
    .Y(_21827_));
 NOR2x1_ASAP7_75t_R _30369_ (.A(_20624_),
    .B(_20747_),
    .Y(_21828_));
 OAI21x1_ASAP7_75t_R _30370_ (.A1(_21827_),
    .A2(_21828_),
    .B(_21543_),
    .Y(_21829_));
 INVx1_ASAP7_75t_R _30371_ (.A(_21829_),
    .Y(_21830_));
 NOR2x1_ASAP7_75t_R _30372_ (.A(_20624_),
    .B(_20734_),
    .Y(_21831_));
 NOR2x1_ASAP7_75t_R _30373_ (.A(_20747_),
    .B(_20653_),
    .Y(_21832_));
 OAI21x1_ASAP7_75t_R _30374_ (.A1(_21831_),
    .A2(_21832_),
    .B(_21123_),
    .Y(_21833_));
 INVx1_ASAP7_75t_R _30375_ (.A(_21833_),
    .Y(_21834_));
 OAI21x1_ASAP7_75t_R _30376_ (.A1(_21830_),
    .A2(_21834_),
    .B(_20437_),
    .Y(_21835_));
 NAND3x1_ASAP7_75t_R _30377_ (.A(_21833_),
    .B(_21829_),
    .C(_20449_),
    .Y(_21836_));
 AOI21x1_ASAP7_75t_R _30378_ (.A1(_21835_),
    .A2(_21836_),
    .B(net390),
    .Y(_21837_));
 INVx1_ASAP7_75t_R _30379_ (.A(_21837_),
    .Y(_21838_));
 AOI21x1_ASAP7_75t_R _30380_ (.A1(_21826_),
    .A2(_21838_),
    .B(_00423_),
    .Y(_21839_));
 NOR3x1_ASAP7_75t_R _30381_ (.A(_21837_),
    .B(_06353_),
    .C(_21825_),
    .Y(_21840_));
 NOR2x1_ASAP7_75t_R _30382_ (.A(_21840_),
    .B(_21839_),
    .Y(_00030_));
 NAND2x1_ASAP7_75t_R _30383_ (.A(_00885_),
    .B(net390),
    .Y(_21841_));
 NAND2x2_ASAP7_75t_R _30384_ (.A(net2341),
    .B(_21528_),
    .Y(_21842_));
 NAND2x1_ASAP7_75t_R _30385_ (.A(_21535_),
    .B(_21725_),
    .Y(_21843_));
 AOI21x1_ASAP7_75t_R _30386_ (.A1(_21842_),
    .A2(_21843_),
    .B(_21554_),
    .Y(_21844_));
 NAND2x2_ASAP7_75t_R _30387_ (.A(_21535_),
    .B(net2341),
    .Y(_21845_));
 NAND2x1_ASAP7_75t_R _30388_ (.A(_21528_),
    .B(_21725_),
    .Y(_21846_));
 AOI21x1_ASAP7_75t_R _30389_ (.A1(_21845_),
    .A2(_21846_),
    .B(net2428),
    .Y(_21847_));
 OAI21x1_ASAP7_75t_R _30390_ (.A1(_21844_),
    .A2(_21847_),
    .B(net397),
    .Y(_21848_));
 AOI21x1_ASAP7_75t_R _30391_ (.A1(_21841_),
    .A2(_21848_),
    .B(_06342_),
    .Y(_21849_));
 OR2x2_ASAP7_75t_R _30392_ (.A(net397),
    .B(_00885_),
    .Y(_21850_));
 AOI21x1_ASAP7_75t_R _30393_ (.A1(_21845_),
    .A2(_21846_),
    .B(_21554_),
    .Y(_21851_));
 AOI21x1_ASAP7_75t_R _30394_ (.A1(_21842_),
    .A2(_21843_),
    .B(_21212_),
    .Y(_21852_));
 OAI21x1_ASAP7_75t_R _30395_ (.A1(_21851_),
    .A2(_21852_),
    .B(net397),
    .Y(_21853_));
 AOI21x1_ASAP7_75t_R _30396_ (.A1(_21850_),
    .A2(_21853_),
    .B(_00422_),
    .Y(_21854_));
 NOR2x1_ASAP7_75t_R _30397_ (.A(_21849_),
    .B(_21854_),
    .Y(_00031_));
 NOR2x1_ASAP7_75t_R _30398_ (.A(net397),
    .B(_00884_),
    .Y(_21855_));
 INVx1_ASAP7_75t_R _30399_ (.A(_21855_),
    .Y(_21856_));
 XOR2x1_ASAP7_75t_R _30400_ (.A(_19143_),
    .Y(_21857_),
    .B(net2363));
 XOR2x1_ASAP7_75t_R _30401_ (.A(_21857_),
    .Y(_21858_),
    .B(_21420_));
 XOR2x2_ASAP7_75t_R _30402_ (.A(_21858_),
    .B(_21049_),
    .Y(_21859_));
 NAND2x1_ASAP7_75t_R _30403_ (.A(_21859_),
    .B(net397),
    .Y(_21860_));
 AOI21x1_ASAP7_75t_R _30404_ (.A1(_21856_),
    .A2(_21860_),
    .B(net3386),
    .Y(_21861_));
 AOI211x1_ASAP7_75t_R _30405_ (.A1(_21859_),
    .A2(net397),
    .B(_21855_),
    .C(_06331_),
    .Y(_21862_));
 NOR2x1_ASAP7_75t_R _30406_ (.A(_21862_),
    .B(_21861_),
    .Y(_00032_));
 AND2x2_ASAP7_75t_R _30407_ (.A(_18753_),
    .B(_00883_),
    .Y(_21863_));
 INVx1_ASAP7_75t_R _30408_ (.A(_21863_),
    .Y(_21864_));
 INVx4_ASAP7_75t_R _30409_ (.A(net3278),
    .Y(_21865_));
 TAPCELL_ASAP7_75t_R TAP_804 ();
 INVx3_ASAP7_75t_R _30411_ (.A(_00546_),
    .Y(_21867_));
 OR3x2_ASAP7_75t_R _30412_ (.A(_21865_),
    .B(_21867_),
    .C(_00547_),
    .Y(_21868_));
 INVx1_ASAP7_75t_R _30413_ (.A(_21868_),
    .Y(_21869_));
 TAPCELL_ASAP7_75t_R TAP_803 ();
 TAPCELL_ASAP7_75t_R TAP_802 ();
 INVx4_ASAP7_75t_R _30416_ (.A(net2005),
    .Y(_21872_));
 NAND2x2_ASAP7_75t_R _30417_ (.A(_00550_),
    .B(_21872_),
    .Y(_21873_));
 TAPCELL_ASAP7_75t_R TAP_801 ();
 TAPCELL_ASAP7_75t_R TAP_800 ();
 CKINVDCx16_ASAP7_75t_R _30420_ (.A(net1169),
    .Y(_21876_));
 NAND2x2_ASAP7_75t_R _30421_ (.A(net1409),
    .B(_21876_),
    .Y(_21877_));
 NOR2x2_ASAP7_75t_R _30422_ (.A(_21873_),
    .B(_21877_),
    .Y(_21878_));
 NAND2x2_ASAP7_75t_R _30423_ (.A(net1407),
    .B(net1170),
    .Y(_21879_));
 TAPCELL_ASAP7_75t_R TAP_799 ();
 NOR2x2_ASAP7_75t_R _30425_ (.A(net995),
    .B(net1712),
    .Y(_21881_));
 TAPCELL_ASAP7_75t_R TAP_798 ();
 NAND2x2_ASAP7_75t_R _30427_ (.A(_00547_),
    .B(_00548_),
    .Y(_21883_));
 NAND2x2_ASAP7_75t_R _30428_ (.A(net3278),
    .B(_00546_),
    .Y(_21884_));
 NOR2x2_ASAP7_75t_R _30429_ (.A(_21883_),
    .B(net1904),
    .Y(_21885_));
 OA21x2_ASAP7_75t_R _30430_ (.A1(_21878_),
    .A2(_21881_),
    .B(_21885_),
    .Y(_21886_));
 CKINVDCx20_ASAP7_75t_R _30431_ (.A(net1406),
    .Y(_21887_));
 INVx3_ASAP7_75t_R _30432_ (.A(_00550_),
    .Y(_21888_));
 NOR2x2_ASAP7_75t_R _30433_ (.A(net2005),
    .B(_21888_),
    .Y(_21889_));
 NAND2x2_ASAP7_75t_R _30434_ (.A(_21887_),
    .B(net1648),
    .Y(_21890_));
 AND2x6_ASAP7_75t_R _30435_ (.A(_00547_),
    .B(_00548_),
    .Y(_21891_));
 INVx4_ASAP7_75t_R _30436_ (.A(_21884_),
    .Y(_21892_));
 NAND2x2_ASAP7_75t_R _30437_ (.A(_21891_),
    .B(_21892_),
    .Y(_21893_));
 NOR2x2_ASAP7_75t_R _30438_ (.A(_21890_),
    .B(_21893_),
    .Y(_21894_));
 NAND2x2_ASAP7_75t_R _30439_ (.A(_21872_),
    .B(_21888_),
    .Y(_21895_));
 TAPCELL_ASAP7_75t_R TAP_797 ();
 NOR2x2_ASAP7_75t_R _30441_ (.A(_21895_),
    .B(_21893_),
    .Y(_21897_));
 NOR3x2_ASAP7_75t_R _30442_ (.B(_21894_),
    .C(_21897_),
    .Y(_21898_),
    .A(_21886_));
 INVx2_ASAP7_75t_R _30443_ (.A(_00547_),
    .Y(_21899_));
 NOR2x2_ASAP7_75t_R _30444_ (.A(_00548_),
    .B(_21899_),
    .Y(_21900_));
 NAND2x2_ASAP7_75t_R _30445_ (.A(_21900_),
    .B(_21892_),
    .Y(_21901_));
 TAPCELL_ASAP7_75t_R TAP_796 ();
 TAPCELL_ASAP7_75t_R TAP_795 ();
 NAND2x2_ASAP7_75t_R _30448_ (.A(net2007),
    .B(_21888_),
    .Y(_21904_));
 TAPCELL_ASAP7_75t_R TAP_794 ();
 TAPCELL_ASAP7_75t_R TAP_793 ();
 NAND2x2_ASAP7_75t_R _30451_ (.A(net2005),
    .B(_00550_),
    .Y(_21907_));
 NOR2x2_ASAP7_75t_R _30452_ (.A(net1407),
    .B(net1039),
    .Y(_21908_));
 NOR2x2_ASAP7_75t_R _30453_ (.A(_21907_),
    .B(_21877_),
    .Y(_21909_));
 OAI21x1_ASAP7_75t_R _30454_ (.A1(_21908_),
    .A2(_21909_),
    .B(_21885_),
    .Y(_21910_));
 OA21x2_ASAP7_75t_R _30455_ (.A1(net1849),
    .A2(_21893_),
    .B(_21910_),
    .Y(_21911_));
 NAND3x2_ASAP7_75t_R _30456_ (.B(_21901_),
    .C(_21911_),
    .Y(_21912_),
    .A(_21898_));
 NOR2x2_ASAP7_75t_R _30457_ (.A(_21869_),
    .B(_21912_),
    .Y(_21913_));
 NAND3x2_ASAP7_75t_R _30458_ (.B(net3279),
    .C(_00546_),
    .Y(_21914_),
    .A(_21913_));
 NOR2x1_ASAP7_75t_R _30459_ (.A(net1710),
    .B(_21901_),
    .Y(_21915_));
 NOR2x2_ASAP7_75t_R _30460_ (.A(net1170),
    .B(_21887_),
    .Y(_21916_));
 NOR2x2_ASAP7_75t_R _30461_ (.A(net1407),
    .B(_21876_),
    .Y(_21917_));
 NOR2x2_ASAP7_75t_R _30462_ (.A(_21916_),
    .B(net2427),
    .Y(_21918_));
 NOR2x2_ASAP7_75t_R _30463_ (.A(_00550_),
    .B(_21872_),
    .Y(_21919_));
 NAND2x2_ASAP7_75t_R _30464_ (.A(_21919_),
    .B(_21916_),
    .Y(_21920_));
 TAPCELL_ASAP7_75t_R TAP_792 ();
 NAND2x2_ASAP7_75t_R _30466_ (.A(_21919_),
    .B(_21917_),
    .Y(_21922_));
 TAPCELL_ASAP7_75t_R TAP_791 ();
 AOI21x1_ASAP7_75t_R _30468_ (.A1(_21920_),
    .A2(net1048),
    .B(net1751),
    .Y(_21924_));
 NOR2x2_ASAP7_75t_R _30469_ (.A(net1411),
    .B(net1170),
    .Y(_21925_));
 INVx4_ASAP7_75t_R _30470_ (.A(net1040),
    .Y(_21926_));
 NAND2x2_ASAP7_75t_R _30471_ (.A(_21925_),
    .B(_21926_),
    .Y(_21927_));
 TAPCELL_ASAP7_75t_R TAP_790 ();
 NAND2x2_ASAP7_75t_R _30473_ (.A(_21926_),
    .B(net2426),
    .Y(_21929_));
 TAPCELL_ASAP7_75t_R TAP_789 ();
 AOI21x1_ASAP7_75t_R _30475_ (.A1(net3076),
    .A2(_21929_),
    .B(_21901_),
    .Y(_21931_));
 AOI211x1_ASAP7_75t_R _30476_ (.A1(_21915_),
    .A2(_21918_),
    .B(_21924_),
    .C(_21931_),
    .Y(_21932_));
 TAPCELL_ASAP7_75t_R TAP_788 ();
 NAND2x2_ASAP7_75t_R _30478_ (.A(_21889_),
    .B(_21916_),
    .Y(_21934_));
 TAPCELL_ASAP7_75t_R TAP_787 ();
 AO21x1_ASAP7_75t_R _30480_ (.A1(_21934_),
    .A2(_21890_),
    .B(net2497),
    .Y(_21936_));
 NOR2x2_ASAP7_75t_R _30481_ (.A(net2005),
    .B(_00550_),
    .Y(_21937_));
 NAND2x2_ASAP7_75t_R _30482_ (.A(net2608),
    .B(_21916_),
    .Y(_21938_));
 TAPCELL_ASAP7_75t_R TAP_786 ();
 NAND2x2_ASAP7_75t_R _30484_ (.A(net1255),
    .B(_21917_),
    .Y(_21940_));
 TAPCELL_ASAP7_75t_R TAP_785 ();
 AO21x1_ASAP7_75t_R _30486_ (.A1(net2258),
    .A2(_21940_),
    .B(net2497),
    .Y(_21942_));
 AND2x2_ASAP7_75t_R _30487_ (.A(_21936_),
    .B(_21942_),
    .Y(_21943_));
 INVx3_ASAP7_75t_R _30488_ (.A(_21908_),
    .Y(_21944_));
 NOR2x2_ASAP7_75t_R _30489_ (.A(_21944_),
    .B(_21893_),
    .Y(_21945_));
 TAPCELL_ASAP7_75t_R TAP_784 ();
 TAPCELL_ASAP7_75t_R TAP_783 ();
 TAPCELL_ASAP7_75t_R TAP_782 ();
 TAPCELL_ASAP7_75t_R TAP_781 ();
 AOI211x1_ASAP7_75t_R _30494_ (.A1(net1139),
    .A2(net1049),
    .B(net2497),
    .C(net1850),
    .Y(_21950_));
 NOR2x2_ASAP7_75t_R _30495_ (.A(_21945_),
    .B(_21950_),
    .Y(_21951_));
 NAND3x2_ASAP7_75t_R _30496_ (.B(_21943_),
    .C(_21951_),
    .Y(_21952_),
    .A(_21932_));
 NOR2x2_ASAP7_75t_R _30497_ (.A(_21887_),
    .B(net1039),
    .Y(_21953_));
 NAND2x2_ASAP7_75t_R _30498_ (.A(net1170),
    .B(_21887_),
    .Y(_21954_));
 NOR2x2_ASAP7_75t_R _30499_ (.A(net1040),
    .B(_21954_),
    .Y(_21955_));
 NAND2x1_ASAP7_75t_R _30500_ (.A(_00548_),
    .B(_21899_),
    .Y(_21956_));
 NOR2x2_ASAP7_75t_R _30501_ (.A(net1904),
    .B(_21956_),
    .Y(_21957_));
 OAI21x1_ASAP7_75t_R _30502_ (.A1(_21953_),
    .A2(_21955_),
    .B(_21957_),
    .Y(_21958_));
 TAPCELL_ASAP7_75t_R TAP_780 ();
 INVx1_ASAP7_75t_R _30504_ (.A(_00548_),
    .Y(_21960_));
 NOR2x2_ASAP7_75t_R _30505_ (.A(_00547_),
    .B(_21960_),
    .Y(_21961_));
 NAND2x2_ASAP7_75t_R _30506_ (.A(_21961_),
    .B(_21892_),
    .Y(_21962_));
 AO21x1_ASAP7_75t_R _30507_ (.A1(_21920_),
    .A2(net1633),
    .B(_21962_),
    .Y(_21963_));
 NAND2x1_ASAP7_75t_R _30508_ (.A(_21958_),
    .B(_21963_),
    .Y(_21964_));
 TAPCELL_ASAP7_75t_R TAP_779 ();
 INVx6_ASAP7_75t_R _30510_ (.A(_21879_),
    .Y(_21966_));
 NAND2x2_ASAP7_75t_R _30511_ (.A(net1256),
    .B(_21966_),
    .Y(_21967_));
 TAPCELL_ASAP7_75t_R TAP_778 ();
 NAND2x2_ASAP7_75t_R _30513_ (.A(_21887_),
    .B(_21937_),
    .Y(_21969_));
 TAPCELL_ASAP7_75t_R TAP_777 ();
 AO21x1_ASAP7_75t_R _30515_ (.A1(_21967_),
    .A2(_21969_),
    .B(_21962_),
    .Y(_21971_));
 AO21x1_ASAP7_75t_R _30516_ (.A1(_21934_),
    .A2(_21890_),
    .B(_21962_),
    .Y(_21972_));
 NAND2x1_ASAP7_75t_R _30517_ (.A(_21971_),
    .B(_21972_),
    .Y(_21973_));
 NOR2x1_ASAP7_75t_R _30518_ (.A(_21964_),
    .B(_21973_),
    .Y(_21974_));
 NOR2x2_ASAP7_75t_R _30519_ (.A(_00547_),
    .B(_00548_),
    .Y(_21975_));
 NAND2x2_ASAP7_75t_R _30520_ (.A(net3078),
    .B(_21892_),
    .Y(_21976_));
 TAPCELL_ASAP7_75t_R TAP_776 ();
 NOR2x2_ASAP7_75t_R _30522_ (.A(net1173),
    .B(net1041),
    .Y(_21978_));
 INVx2_ASAP7_75t_R _30523_ (.A(net3078),
    .Y(_21979_));
 NOR2x2_ASAP7_75t_R _30524_ (.A(net1905),
    .B(_21979_),
    .Y(_21980_));
 OAI21x1_ASAP7_75t_R _30525_ (.A1(_21978_),
    .A2(_21955_),
    .B(_21980_),
    .Y(_21981_));
 OAI21x1_ASAP7_75t_R _30526_ (.A1(net1048),
    .A2(_21976_),
    .B(_21981_),
    .Y(_21982_));
 NAND2x2_ASAP7_75t_R _30527_ (.A(net1652),
    .B(_21966_),
    .Y(_21983_));
 TAPCELL_ASAP7_75t_R TAP_775 ();
 NOR2x1_ASAP7_75t_R _30529_ (.A(_21976_),
    .B(_21983_),
    .Y(_21985_));
 TAPCELL_ASAP7_75t_R TAP_774 ();
 AOI211x1_ASAP7_75t_R _30531_ (.A1(_21887_),
    .A2(net1049),
    .B(_21976_),
    .C(_21895_),
    .Y(_21987_));
 NOR3x1_ASAP7_75t_R _30532_ (.A(_21982_),
    .B(_21985_),
    .C(_21987_),
    .Y(_21988_));
 NAND2x1_ASAP7_75t_R _30533_ (.A(_21974_),
    .B(_21988_),
    .Y(_21989_));
 NOR2x2_ASAP7_75t_R _30534_ (.A(_21952_),
    .B(_21989_),
    .Y(_21990_));
 NOR2x2_ASAP7_75t_R _30535_ (.A(_00546_),
    .B(_21865_),
    .Y(_21991_));
 NAND2x2_ASAP7_75t_R _30536_ (.A(_21991_),
    .B(_21900_),
    .Y(_21992_));
 TAPCELL_ASAP7_75t_R TAP_773 ();
 AOI211x1_ASAP7_75t_R _30538_ (.A1(_21969_),
    .A2(net1713),
    .B(_21992_),
    .C(net1049),
    .Y(_21994_));
 INVx5_ASAP7_75t_R _30539_ (.A(_21953_),
    .Y(_21995_));
 AO21x1_ASAP7_75t_R _30540_ (.A1(_21995_),
    .A2(_21927_),
    .B(_21992_),
    .Y(_21996_));
 NAND2x2_ASAP7_75t_R _30541_ (.A(_21925_),
    .B(_21919_),
    .Y(_21997_));
 TAPCELL_ASAP7_75t_R TAP_772 ();
 AO21x1_ASAP7_75t_R _30543_ (.A1(net1631),
    .A2(net1834),
    .B(_21992_),
    .Y(_21999_));
 NAND2x1_ASAP7_75t_R _30544_ (.A(_21996_),
    .B(_21999_),
    .Y(_22000_));
 NOR2x1_ASAP7_75t_R _30545_ (.A(_21994_),
    .B(_22000_),
    .Y(_22001_));
 NAND2x2_ASAP7_75t_R _30546_ (.A(net2763),
    .B(_21966_),
    .Y(_22002_));
 INVx4_ASAP7_75t_R _30547_ (.A(net2296),
    .Y(_22003_));
 NAND2x2_ASAP7_75t_R _30548_ (.A(_21991_),
    .B(_21891_),
    .Y(_22004_));
 INVx2_ASAP7_75t_R _30549_ (.A(_22004_),
    .Y(_22005_));
 OA21x2_ASAP7_75t_R _30550_ (.A1(_22003_),
    .A2(_21953_),
    .B(_22005_),
    .Y(_22006_));
 NAND2x2_ASAP7_75t_R _30551_ (.A(net1649),
    .B(_22005_),
    .Y(_22007_));
 NAND2x2_ASAP7_75t_R _30552_ (.A(net1412),
    .B(net1257),
    .Y(_22008_));
 TAPCELL_ASAP7_75t_R TAP_771 ();
 AO21x1_ASAP7_75t_R _30554_ (.A1(_21940_),
    .A2(_22008_),
    .B(_22004_),
    .Y(_22010_));
 OAI21x1_ASAP7_75t_R _30555_ (.A1(net1049),
    .A2(_22007_),
    .B(_22010_),
    .Y(_22011_));
 NOR2x1_ASAP7_75t_R _30556_ (.A(_22006_),
    .B(_22011_),
    .Y(_22012_));
 NAND2x1_ASAP7_75t_R _30557_ (.A(_22001_),
    .B(_22012_),
    .Y(_22013_));
 NOR2x2_ASAP7_75t_R _30558_ (.A(_21954_),
    .B(_21895_),
    .Y(_22014_));
 NAND2x2_ASAP7_75t_R _30559_ (.A(_21991_),
    .B(_21961_),
    .Y(_22015_));
 INVx2_ASAP7_75t_R _30560_ (.A(_22015_),
    .Y(_22016_));
 NAND2x1_ASAP7_75t_R _30561_ (.A(_22014_),
    .B(_22016_),
    .Y(_22017_));
 NAND2x2_ASAP7_75t_R _30562_ (.A(_21925_),
    .B(net1651),
    .Y(_22018_));
 NAND2x2_ASAP7_75t_R _30563_ (.A(net1410),
    .B(net1648),
    .Y(_22019_));
 TAPCELL_ASAP7_75t_R TAP_770 ();
 TAPCELL_ASAP7_75t_R TAP_769 ();
 AO21x1_ASAP7_75t_R _30566_ (.A1(_22018_),
    .A2(_22019_),
    .B(_22015_),
    .Y(_22022_));
 NAND2x1_ASAP7_75t_R _30567_ (.A(_22017_),
    .B(_22022_),
    .Y(_22023_));
 NAND2x2_ASAP7_75t_R _30568_ (.A(_21916_),
    .B(_21926_),
    .Y(_22024_));
 AO21x1_ASAP7_75t_R _30569_ (.A1(_22024_),
    .A2(net3280),
    .B(net2785),
    .Y(_22025_));
 OAI21x1_ASAP7_75t_R _30570_ (.A1(net1852),
    .A2(net2785),
    .B(_22025_),
    .Y(_22026_));
 NOR2x1_ASAP7_75t_R _30571_ (.A(_22023_),
    .B(_22026_),
    .Y(_22027_));
 NAND2x2_ASAP7_75t_R _30572_ (.A(_21975_),
    .B(_21991_),
    .Y(_22028_));
 TAPCELL_ASAP7_75t_R TAP_768 ();
 TAPCELL_ASAP7_75t_R TAP_767 ();
 AO21x1_ASAP7_75t_R _30575_ (.A1(net2258),
    .A2(_21940_),
    .B(net3156),
    .Y(_22031_));
 OAI21x1_ASAP7_75t_R _30576_ (.A1(net2556),
    .A2(net2337),
    .B(_22031_),
    .Y(_22032_));
 NOR2x1_ASAP7_75t_R _30577_ (.A(net1171),
    .B(net1851),
    .Y(_22033_));
 INVx4_ASAP7_75t_R _30578_ (.A(net3156),
    .Y(_22034_));
 NAND2x1_ASAP7_75t_R _30579_ (.A(_22033_),
    .B(_22034_),
    .Y(_22035_));
 TAPCELL_ASAP7_75t_R TAP_766 ();
 AOI211x1_ASAP7_75t_R _30581_ (.A1(_21887_),
    .A2(net1049),
    .B(net3156),
    .C(net1045),
    .Y(_22037_));
 INVx1_ASAP7_75t_R _30582_ (.A(_22037_),
    .Y(_22038_));
 NAND2x1_ASAP7_75t_R _30583_ (.A(_22035_),
    .B(_22038_),
    .Y(_22039_));
 NOR2x1_ASAP7_75t_R _30584_ (.A(_22032_),
    .B(_22039_),
    .Y(_22040_));
 NAND2x1_ASAP7_75t_R _30585_ (.A(_22027_),
    .B(_22040_),
    .Y(_22041_));
 NOR2x1_ASAP7_75t_R _30586_ (.A(_22013_),
    .B(_22041_),
    .Y(_22042_));
 NAND2x2_ASAP7_75t_R _30587_ (.A(_21990_),
    .B(_22042_),
    .Y(_22043_));
 NOR2x2_ASAP7_75t_R _30588_ (.A(_21876_),
    .B(net1043),
    .Y(_22044_));
 INVx3_ASAP7_75t_R _30589_ (.A(_21925_),
    .Y(_22045_));
 NOR2x2_ASAP7_75t_R _30590_ (.A(net1040),
    .B(_22045_),
    .Y(_22046_));
 TAPCELL_ASAP7_75t_R TAP_765 ();
 NAND2x2_ASAP7_75t_R _30592_ (.A(_00546_),
    .B(_21865_),
    .Y(_22048_));
 NOR2x2_ASAP7_75t_R _30593_ (.A(_22048_),
    .B(_21979_),
    .Y(_22049_));
 TAPCELL_ASAP7_75t_R TAP_764 ();
 OAI21x1_ASAP7_75t_R _30595_ (.A1(_22044_),
    .A2(net2038),
    .B(_22049_),
    .Y(_22051_));
 INVx1_ASAP7_75t_R _30596_ (.A(_22051_),
    .Y(_22052_));
 NOR2x2_ASAP7_75t_R _30597_ (.A(_21904_),
    .B(_22045_),
    .Y(_22053_));
 NOR2x2_ASAP7_75t_R _30598_ (.A(_21887_),
    .B(net1845),
    .Y(_22054_));
 OA21x2_ASAP7_75t_R _30599_ (.A1(_22053_),
    .A2(_22054_),
    .B(_22049_),
    .Y(_22055_));
 NOR2x1_ASAP7_75t_R _30600_ (.A(_22052_),
    .B(_22055_),
    .Y(_22056_));
 NAND2x2_ASAP7_75t_R _30601_ (.A(_21937_),
    .B(_21954_),
    .Y(_22057_));
 TAPCELL_ASAP7_75t_R TAP_763 ();
 NAND2x1_ASAP7_75t_R _30603_ (.A(_22057_),
    .B(net2365),
    .Y(_22059_));
 NOR2x2_ASAP7_75t_R _30604_ (.A(net3278),
    .B(_21867_),
    .Y(_22060_));
 NAND2x2_ASAP7_75t_R _30605_ (.A(_22060_),
    .B(_21961_),
    .Y(_22061_));
 INVx4_ASAP7_75t_R _30606_ (.A(_22061_),
    .Y(_22062_));
 OAI21x1_ASAP7_75t_R _30607_ (.A1(_22003_),
    .A2(_22059_),
    .B(_22062_),
    .Y(_22063_));
 NAND2x2_ASAP7_75t_R _30608_ (.A(net3079),
    .B(_22060_),
    .Y(_22064_));
 TAPCELL_ASAP7_75t_R TAP_762 ();
 TAPCELL_ASAP7_75t_R TAP_761 ();
 NOR2x1_ASAP7_75t_R _30611_ (.A(_22064_),
    .B(net2752),
    .Y(_22067_));
 INVx1_ASAP7_75t_R _30612_ (.A(_22067_),
    .Y(_22068_));
 NAND3x1_ASAP7_75t_R _30613_ (.A(_22056_),
    .B(_22063_),
    .C(_22068_),
    .Y(_22069_));
 NAND2x2_ASAP7_75t_R _30614_ (.A(_21900_),
    .B(_22060_),
    .Y(_22070_));
 TAPCELL_ASAP7_75t_R TAP_760 ();
 TAPCELL_ASAP7_75t_R TAP_759 ();
 AO21x1_ASAP7_75t_R _30617_ (.A1(_22024_),
    .A2(_21929_),
    .B(_22070_),
    .Y(_22073_));
 OA21x2_ASAP7_75t_R _30618_ (.A1(_21969_),
    .A2(_22070_),
    .B(_22073_),
    .Y(_22074_));
 NOR2x2_ASAP7_75t_R _30619_ (.A(_21879_),
    .B(net1040),
    .Y(_22075_));
 INVx3_ASAP7_75t_R _30620_ (.A(_22075_),
    .Y(_22076_));
 NAND2x2_ASAP7_75t_R _30621_ (.A(_22060_),
    .B(_21891_),
    .Y(_22077_));
 TAPCELL_ASAP7_75t_R TAP_758 ();
 AO21x1_ASAP7_75t_R _30623_ (.A1(_22076_),
    .A2(_21929_),
    .B(_22077_),
    .Y(_22079_));
 NAND2x2_ASAP7_75t_R _30624_ (.A(net1407),
    .B(net2762),
    .Y(_22080_));
 AO21x1_ASAP7_75t_R _30625_ (.A1(net1792),
    .A2(_22080_),
    .B(_22077_),
    .Y(_22081_));
 AND2x2_ASAP7_75t_R _30626_ (.A(_22079_),
    .B(_22081_),
    .Y(_22082_));
 NOR2x2_ASAP7_75t_R _30627_ (.A(net1712),
    .B(_22045_),
    .Y(_22083_));
 NOR2x2_ASAP7_75t_R _30628_ (.A(_21883_),
    .B(_22048_),
    .Y(_22084_));
 OA21x2_ASAP7_75t_R _30629_ (.A1(_22083_),
    .A2(_21878_),
    .B(_22084_),
    .Y(_22085_));
 AND3x1_ASAP7_75t_R _30630_ (.A(_22084_),
    .B(_21879_),
    .C(net1258),
    .Y(_22086_));
 NOR2x1_ASAP7_75t_R _30631_ (.A(_22085_),
    .B(_22086_),
    .Y(_22087_));
 NAND3x1_ASAP7_75t_R _30632_ (.A(_22074_),
    .B(_22082_),
    .C(_22087_),
    .Y(_22088_));
 NOR2x1_ASAP7_75t_R _30633_ (.A(_22069_),
    .B(_22088_),
    .Y(_22089_));
 NOR2x2_ASAP7_75t_R _30634_ (.A(net3278),
    .B(_00546_),
    .Y(_22090_));
 NAND2x2_ASAP7_75t_R _30635_ (.A(_22090_),
    .B(_21975_),
    .Y(_22091_));
 INVx4_ASAP7_75t_R _30636_ (.A(_22091_),
    .Y(_22092_));
 TAPCELL_ASAP7_75t_R TAP_757 ();
 AOI211x1_ASAP7_75t_R _30638_ (.A1(net1139),
    .A2(net1049),
    .B(_22091_),
    .C(net1040),
    .Y(_22094_));
 OA21x2_ASAP7_75t_R _30639_ (.A1(_22014_),
    .A2(_21889_),
    .B(_22092_),
    .Y(_22095_));
 AOI211x1_ASAP7_75t_R _30640_ (.A1(_22003_),
    .A2(_22092_),
    .B(_22094_),
    .C(_22095_),
    .Y(_22096_));
 TAPCELL_ASAP7_75t_R TAP_756 ();
 NAND2x1_ASAP7_75t_R _30642_ (.A(_21876_),
    .B(_21937_),
    .Y(_22098_));
 AO21x1_ASAP7_75t_R _30643_ (.A1(net1408),
    .A2(_21876_),
    .B(net1708),
    .Y(_22099_));
 NAND2x2_ASAP7_75t_R _30644_ (.A(_22090_),
    .B(_21961_),
    .Y(_22100_));
 TAPCELL_ASAP7_75t_R TAP_755 ();
 AOI21x1_ASAP7_75t_R _30646_ (.A1(_22098_),
    .A2(_22099_),
    .B(_22100_),
    .Y(_01067_));
 AO21x1_ASAP7_75t_R _30647_ (.A1(_22076_),
    .A2(_21927_),
    .B(net3080),
    .Y(_01068_));
 OAI21x1_ASAP7_75t_R _30648_ (.A1(net3080),
    .A2(_22080_),
    .B(_01068_),
    .Y(_01069_));
 NOR2x1_ASAP7_75t_R _30649_ (.A(_01067_),
    .B(_01069_),
    .Y(_01070_));
 NAND2x1_ASAP7_75t_R _30650_ (.A(_22096_),
    .B(_01070_),
    .Y(_01071_));
 NAND2x2_ASAP7_75t_R _30651_ (.A(_22090_),
    .B(_21891_),
    .Y(_01072_));
 INVx4_ASAP7_75t_R _30652_ (.A(_01072_),
    .Y(_01073_));
 TAPCELL_ASAP7_75t_R TAP_754 ();
 AOI211x1_ASAP7_75t_R _30654_ (.A1(_21887_),
    .A2(_21876_),
    .B(_01072_),
    .C(_21895_),
    .Y(_01075_));
 OA21x2_ASAP7_75t_R _30655_ (.A1(_22083_),
    .A2(_21878_),
    .B(_01073_),
    .Y(_01076_));
 AOI211x1_ASAP7_75t_R _30656_ (.A1(_21955_),
    .A2(_01073_),
    .B(_01075_),
    .C(_01076_),
    .Y(_01077_));
 NAND2x2_ASAP7_75t_R _30657_ (.A(_22090_),
    .B(_21900_),
    .Y(_01078_));
 CKINVDCx6p67_ASAP7_75t_R _30658_ (.A(_01078_),
    .Y(_01079_));
 TAPCELL_ASAP7_75t_R TAP_753 ();
 OAI21x1_ASAP7_75t_R _30660_ (.A1(_21881_),
    .A2(_21878_),
    .B(_01079_),
    .Y(_01081_));
 NOR2x2_ASAP7_75t_R _30661_ (.A(_21873_),
    .B(_21954_),
    .Y(_01082_));
 OAI21x1_ASAP7_75t_R _30662_ (.A1(_01082_),
    .A2(_22083_),
    .B(_01079_),
    .Y(_01083_));
 NAND2x1_ASAP7_75t_R _30663_ (.A(_01081_),
    .B(_01083_),
    .Y(_01084_));
 NOR2x2_ASAP7_75t_R _30664_ (.A(_21904_),
    .B(_21877_),
    .Y(_01085_));
 OA21x2_ASAP7_75t_R _30665_ (.A1(_01085_),
    .A2(_21955_),
    .B(_01079_),
    .Y(_01086_));
 INVx3_ASAP7_75t_R _30666_ (.A(net2258),
    .Y(_01087_));
 OA21x2_ASAP7_75t_R _30667_ (.A1(_01087_),
    .A2(_22014_),
    .B(_01079_),
    .Y(_01088_));
 NOR3x1_ASAP7_75t_R _30668_ (.A(_01084_),
    .B(_01086_),
    .C(_01088_),
    .Y(_01089_));
 NAND2x1_ASAP7_75t_R _30669_ (.A(_01077_),
    .B(_01089_),
    .Y(_01090_));
 NOR2x1_ASAP7_75t_R _30670_ (.A(_01071_),
    .B(_01090_),
    .Y(_01091_));
 NAND2x1_ASAP7_75t_R _30671_ (.A(_01091_),
    .B(_22089_),
    .Y(_01092_));
 NOR2x2_ASAP7_75t_R _30672_ (.A(_22043_),
    .B(_01092_),
    .Y(_01093_));
 NAND2x2_ASAP7_75t_R _30673_ (.A(net2789),
    .B(_01093_),
    .Y(_01094_));
 TAPCELL_ASAP7_75t_R TAP_752 ();
 CKINVDCx16_ASAP7_75t_R _30675_ (.A(net1686),
    .Y(_01096_));
 NOR2x2_ASAP7_75t_R _30676_ (.A(_00591_),
    .B(_01096_),
    .Y(_01097_));
 TAPCELL_ASAP7_75t_R TAP_751 ();
 NAND2x2_ASAP7_75t_R _30678_ (.A(_00587_),
    .B(_00588_),
    .Y(_01099_));
 TAPCELL_ASAP7_75t_R TAP_750 ();
 INVx4_ASAP7_75t_R _30680_ (.A(_00585_),
    .Y(_01101_));
 NAND2x2_ASAP7_75t_R _30681_ (.A(_00586_),
    .B(_01101_),
    .Y(_01102_));
 NOR2x2_ASAP7_75t_R _30682_ (.A(_01099_),
    .B(_01102_),
    .Y(_01103_));
 TAPCELL_ASAP7_75t_R TAP_749 ();
 TAPCELL_ASAP7_75t_R TAP_748 ();
 INVx4_ASAP7_75t_R _30685_ (.A(net2647),
    .Y(_01106_));
 NAND3x2_ASAP7_75t_R _30686_ (.B(net2326),
    .C(_01106_),
    .Y(_01107_),
    .A(_01103_));
 NAND2x2_ASAP7_75t_R _30687_ (.A(net2323),
    .B(net2650),
    .Y(_01108_));
 CKINVDCx12_ASAP7_75t_R _30688_ (.A(_01108_),
    .Y(_01109_));
 TAPCELL_ASAP7_75t_R TAP_747 ();
 NAND2x2_ASAP7_75t_R _30690_ (.A(net1594),
    .B(net1686),
    .Y(_01111_));
 CKINVDCx6p67_ASAP7_75t_R _30691_ (.A(_01111_),
    .Y(_01112_));
 NAND2x2_ASAP7_75t_R _30692_ (.A(_01109_),
    .B(_01112_),
    .Y(_01113_));
 TAPCELL_ASAP7_75t_R TAP_746 ();
 NAND2x2_ASAP7_75t_R _30694_ (.A(_01097_),
    .B(_01109_),
    .Y(_01115_));
 TAPCELL_ASAP7_75t_R TAP_745 ();
 INVx3_ASAP7_75t_R _30696_ (.A(_00586_),
    .Y(_01117_));
 NOR2x2_ASAP7_75t_R _30697_ (.A(_00585_),
    .B(_01117_),
    .Y(_01118_));
 AND2x6_ASAP7_75t_R _30698_ (.A(_00587_),
    .B(_00588_),
    .Y(_01119_));
 NAND2x2_ASAP7_75t_R _30699_ (.A(_01118_),
    .B(_01119_),
    .Y(_01120_));
 TAPCELL_ASAP7_75t_R TAP_744 ();
 AO21x1_ASAP7_75t_R _30701_ (.A1(_01113_),
    .A2(_01115_),
    .B(_01120_),
    .Y(_01122_));
 OAI21x1_ASAP7_75t_R _30702_ (.A1(_01097_),
    .A2(_01107_),
    .B(_01122_),
    .Y(_01123_));
 NOR2x2_ASAP7_75t_R _30703_ (.A(net2323),
    .B(_00590_),
    .Y(_01124_));
 NAND2x2_ASAP7_75t_R _30704_ (.A(_01124_),
    .B(_01097_),
    .Y(_01125_));
 TAPCELL_ASAP7_75t_R TAP_743 ();
 NOR2x2_ASAP7_75t_R _30706_ (.A(net1594),
    .B(net1686),
    .Y(_01127_));
 NAND2x2_ASAP7_75t_R _30707_ (.A(net1327),
    .B(net1196),
    .Y(_01128_));
 TAPCELL_ASAP7_75t_R TAP_742 ();
 TAPCELL_ASAP7_75t_R TAP_741 ();
 INVx2_ASAP7_75t_R _30710_ (.A(_00587_),
    .Y(_01131_));
 NOR2x2_ASAP7_75t_R _30711_ (.A(_00588_),
    .B(_01131_),
    .Y(_01132_));
 NAND2x2_ASAP7_75t_R _30712_ (.A(_01132_),
    .B(_01118_),
    .Y(_01133_));
 TAPCELL_ASAP7_75t_R TAP_740 ();
 AO21x1_ASAP7_75t_R _30714_ (.A1(net1572),
    .A2(net1122),
    .B(_01133_),
    .Y(_01135_));
 CKINVDCx20_ASAP7_75t_R _30715_ (.A(net1593),
    .Y(_01136_));
 NOR2x2_ASAP7_75t_R _30716_ (.A(net1682),
    .B(_01136_),
    .Y(_01137_));
 NAND2x2_ASAP7_75t_R _30717_ (.A(_01137_),
    .B(_01109_),
    .Y(_01138_));
 TAPCELL_ASAP7_75t_R TAP_739 ();
 AO21x1_ASAP7_75t_R _30719_ (.A1(_01115_),
    .A2(_01138_),
    .B(_01133_),
    .Y(_01140_));
 NAND2x1_ASAP7_75t_R _30720_ (.A(_01135_),
    .B(_01140_),
    .Y(_01141_));
 TAPCELL_ASAP7_75t_R TAP_738 ();
 NAND2x2_ASAP7_75t_R _30722_ (.A(net1134),
    .B(net1327),
    .Y(_01143_));
 OR2x2_ASAP7_75t_R _30723_ (.A(_01143_),
    .B(_01120_),
    .Y(_01144_));
 NOR2x2_ASAP7_75t_R _30724_ (.A(net2324),
    .B(_01106_),
    .Y(_01145_));
 NAND2x2_ASAP7_75t_R _30725_ (.A(_01137_),
    .B(_01145_),
    .Y(_01146_));
 TAPCELL_ASAP7_75t_R TAP_737 ();
 NAND2x2_ASAP7_75t_R _30727_ (.A(_01127_),
    .B(net1967),
    .Y(_01148_));
 TAPCELL_ASAP7_75t_R TAP_736 ();
 AO21x1_ASAP7_75t_R _30729_ (.A1(net3320),
    .A2(net940),
    .B(_01120_),
    .Y(_01150_));
 NAND2x1_ASAP7_75t_R _30730_ (.A(_01144_),
    .B(_01150_),
    .Y(_01151_));
 NOR3x1_ASAP7_75t_R _30731_ (.A(_01123_),
    .B(_01141_),
    .C(_01151_),
    .Y(_01152_));
 NAND2x2_ASAP7_75t_R _30732_ (.A(_00591_),
    .B(net1334),
    .Y(_01153_));
 INVx1_ASAP7_75t_R _30733_ (.A(_00588_),
    .Y(_01154_));
 NOR2x2_ASAP7_75t_R _30734_ (.A(_00587_),
    .B(_01154_),
    .Y(_01155_));
 NAND2x2_ASAP7_75t_R _30735_ (.A(_01155_),
    .B(_01118_),
    .Y(_01156_));
 TAPCELL_ASAP7_75t_R TAP_735 ();
 AO21x1_ASAP7_75t_R _30737_ (.A1(net1752),
    .A2(_01153_),
    .B(_01156_),
    .Y(_01158_));
 NAND2x2_ASAP7_75t_R _30738_ (.A(net2323),
    .B(_01106_),
    .Y(_01159_));
 NOR2x2_ASAP7_75t_R _30739_ (.A(net1134),
    .B(_01159_),
    .Y(_01160_));
 TAPCELL_ASAP7_75t_R TAP_734 ();
 NAND2x1_ASAP7_75t_R _30741_ (.A(_00588_),
    .B(_01131_),
    .Y(_01162_));
 NOR2x2_ASAP7_75t_R _30742_ (.A(_01162_),
    .B(_01102_),
    .Y(_01163_));
 TAPCELL_ASAP7_75t_R TAP_733 ();
 NAND2x1_ASAP7_75t_R _30744_ (.A(_01160_),
    .B(_01163_),
    .Y(_01165_));
 INVx4_ASAP7_75t_R _30745_ (.A(_01128_),
    .Y(_01166_));
 NAND2x1_ASAP7_75t_R _30746_ (.A(_01163_),
    .B(_01166_),
    .Y(_01167_));
 NAND3x1_ASAP7_75t_R _30747_ (.A(_01158_),
    .B(_01165_),
    .C(_01167_),
    .Y(_01168_));
 NOR2x2_ASAP7_75t_R _30748_ (.A(_00587_),
    .B(_00588_),
    .Y(_01169_));
 NAND2x2_ASAP7_75t_R _30749_ (.A(_01169_),
    .B(_01118_),
    .Y(_01170_));
 INVx5_ASAP7_75t_R _30750_ (.A(_01170_),
    .Y(_01171_));
 NAND2x2_ASAP7_75t_R _30751_ (.A(net1327),
    .B(_01112_),
    .Y(_01172_));
 INVx3_ASAP7_75t_R _30752_ (.A(_01172_),
    .Y(_01173_));
 NAND2x1_ASAP7_75t_R _30753_ (.A(_01171_),
    .B(_01173_),
    .Y(_01174_));
 TAPCELL_ASAP7_75t_R TAP_732 ();
 TAPCELL_ASAP7_75t_R TAP_731 ();
 AOI211x1_ASAP7_75t_R _30756_ (.A1(_00591_),
    .A2(_01096_),
    .B(_01170_),
    .C(net1433),
    .Y(_01177_));
 INVx3_ASAP7_75t_R _30757_ (.A(net1197),
    .Y(_01178_));
 NOR2x2_ASAP7_75t_R _30758_ (.A(net1914),
    .B(_01178_),
    .Y(_01179_));
 NOR2x2_ASAP7_75t_R _30759_ (.A(_01136_),
    .B(_01159_),
    .Y(_01180_));
 OA21x2_ASAP7_75t_R _30760_ (.A1(_01179_),
    .A2(_01180_),
    .B(_01171_),
    .Y(_01181_));
 NOR2x1_ASAP7_75t_R _30761_ (.A(_01177_),
    .B(_01181_),
    .Y(_01182_));
 NAND2x1_ASAP7_75t_R _30762_ (.A(_01174_),
    .B(_01182_),
    .Y(_01183_));
 NOR2x1_ASAP7_75t_R _30763_ (.A(_01168_),
    .B(_01183_),
    .Y(_01184_));
 NAND2x1_ASAP7_75t_R _30764_ (.A(_01152_),
    .B(_01184_),
    .Y(_01185_));
 INVx4_ASAP7_75t_R _30765_ (.A(net2323),
    .Y(_01186_));
 NOR2x2_ASAP7_75t_R _30766_ (.A(net2647),
    .B(_01186_),
    .Y(_01187_));
 NAND2x2_ASAP7_75t_R _30767_ (.A(_01137_),
    .B(_01187_),
    .Y(_01188_));
 TAPCELL_ASAP7_75t_R TAP_730 ();
 NOR2x2_ASAP7_75t_R _30769_ (.A(_00585_),
    .B(_00586_),
    .Y(_01190_));
 NAND2x2_ASAP7_75t_R _30770_ (.A(_01190_),
    .B(_01132_),
    .Y(_01191_));
 TAPCELL_ASAP7_75t_R TAP_729 ();
 AO21x1_ASAP7_75t_R _30772_ (.A1(net1275),
    .A2(net1266),
    .B(net3144),
    .Y(_01193_));
 NAND2x2_ASAP7_75t_R _30773_ (.A(net1327),
    .B(_01137_),
    .Y(_01194_));
 TAPCELL_ASAP7_75t_R TAP_728 ();
 AO21x1_ASAP7_75t_R _30775_ (.A1(net1572),
    .A2(net1076),
    .B(net3144),
    .Y(_01196_));
 INVx4_ASAP7_75t_R _30776_ (.A(_01191_),
    .Y(_01197_));
 NAND2x1_ASAP7_75t_R _30777_ (.A(net1972),
    .B(_01197_),
    .Y(_01198_));
 NAND3x1_ASAP7_75t_R _30778_ (.A(_01193_),
    .B(_01196_),
    .C(_01198_),
    .Y(_01199_));
 TAPCELL_ASAP7_75t_R TAP_727 ();
 TAPCELL_ASAP7_75t_R TAP_726 ();
 NAND2x2_ASAP7_75t_R _30781_ (.A(_01190_),
    .B(_01119_),
    .Y(_01202_));
 TAPCELL_ASAP7_75t_R TAP_725 ();
 CKINVDCx9p33_ASAP7_75t_R _30783_ (.A(net1332),
    .Y(_01204_));
 TAPCELL_ASAP7_75t_R TAP_724 ();
 AOI211x1_ASAP7_75t_R _30785_ (.A1(net2872),
    .A2(_01096_),
    .B(_01202_),
    .C(_01204_),
    .Y(_01206_));
 INVx1_ASAP7_75t_R _30786_ (.A(_01206_),
    .Y(_01207_));
 NAND2x2_ASAP7_75t_R _30787_ (.A(net1683),
    .B(_01136_),
    .Y(_01208_));
 NOR2x2_ASAP7_75t_R _30788_ (.A(net1427),
    .B(_01208_),
    .Y(_01209_));
 CKINVDCx5p33_ASAP7_75t_R _30789_ (.A(_01202_),
    .Y(_01210_));
 NAND2x1_ASAP7_75t_R _30790_ (.A(_01209_),
    .B(_01210_),
    .Y(_01211_));
 AO21x1_ASAP7_75t_R _30791_ (.A1(net3320),
    .A2(net940),
    .B(net3154),
    .Y(_01212_));
 NAND3x1_ASAP7_75t_R _30792_ (.A(_01207_),
    .B(_01211_),
    .C(_01212_),
    .Y(_01213_));
 NOR2x1_ASAP7_75t_R _30793_ (.A(_01199_),
    .B(_01213_),
    .Y(_01214_));
 NAND2x2_ASAP7_75t_R _30794_ (.A(_01190_),
    .B(_01169_),
    .Y(_01215_));
 NOR2x1_ASAP7_75t_R _30795_ (.A(net1426),
    .B(_01215_),
    .Y(_01216_));
 OAI21x1_ASAP7_75t_R _30796_ (.A1(net2872),
    .A2(net3289),
    .B(_01216_),
    .Y(_01217_));
 INVx8_ASAP7_75t_R _30797_ (.A(_01215_),
    .Y(_01218_));
 TAPCELL_ASAP7_75t_R TAP_723 ();
 NAND2x1_ASAP7_75t_R _30799_ (.A(_01160_),
    .B(_01218_),
    .Y(_01220_));
 NAND2x2_ASAP7_75t_R _30800_ (.A(net2648),
    .B(_01186_),
    .Y(_01221_));
 TAPCELL_ASAP7_75t_R TAP_722 ();
 TAPCELL_ASAP7_75t_R TAP_721 ();
 AO21x1_ASAP7_75t_R _30803_ (.A1(net1572),
    .A2(_01221_),
    .B(_01215_),
    .Y(_01224_));
 NAND3x1_ASAP7_75t_R _30804_ (.A(_01217_),
    .B(_01220_),
    .C(_01224_),
    .Y(_01225_));
 NAND2x2_ASAP7_75t_R _30805_ (.A(net1195),
    .B(_01109_),
    .Y(_01226_));
 TAPCELL_ASAP7_75t_R TAP_720 ();
 INVx3_ASAP7_75t_R _30807_ (.A(_01180_),
    .Y(_01228_));
 NAND2x2_ASAP7_75t_R _30808_ (.A(_01190_),
    .B(_01155_),
    .Y(_01229_));
 TAPCELL_ASAP7_75t_R TAP_719 ();
 AO31x2_ASAP7_75t_R _30810_ (.A1(_01226_),
    .A2(_01113_),
    .A3(_01228_),
    .B(_01229_),
    .Y(_01231_));
 AOI211x1_ASAP7_75t_R _30811_ (.A1(net1593),
    .A2(_01096_),
    .B(_01221_),
    .C(_01229_),
    .Y(_01232_));
 INVx6_ASAP7_75t_R _30812_ (.A(net2577),
    .Y(_01233_));
 INVx6_ASAP7_75t_R _30813_ (.A(_01229_),
    .Y(_01234_));
 OA21x2_ASAP7_75t_R _30814_ (.A1(_01233_),
    .A2(_01166_),
    .B(_01234_),
    .Y(_01235_));
 NOR2x1_ASAP7_75t_R _30815_ (.A(_01232_),
    .B(_01235_),
    .Y(_01236_));
 NAND2x1_ASAP7_75t_R _30816_ (.A(_01236_),
    .B(_01231_),
    .Y(_01237_));
 NOR2x1_ASAP7_75t_R _30817_ (.A(_01225_),
    .B(_01237_),
    .Y(_01238_));
 NAND2x2_ASAP7_75t_R _30818_ (.A(_01238_),
    .B(_01214_),
    .Y(_01239_));
 NOR2x2_ASAP7_75t_R _30819_ (.A(_01185_),
    .B(_01239_),
    .Y(_01240_));
 TAPCELL_ASAP7_75t_R TAP_718 ();
 AND2x6_ASAP7_75t_R _30821_ (.A(_00585_),
    .B(_00586_),
    .Y(_01242_));
 NAND2x2_ASAP7_75t_R _30822_ (.A(_01169_),
    .B(_01242_),
    .Y(_01243_));
 NOR2x2_ASAP7_75t_R _30823_ (.A(_01204_),
    .B(_01243_),
    .Y(_01244_));
 OAI21x1_ASAP7_75t_R _30824_ (.A1(net1341),
    .A2(net3289),
    .B(_01244_),
    .Y(_01245_));
 NAND2x2_ASAP7_75t_R _30825_ (.A(_01097_),
    .B(_01187_),
    .Y(_01246_));
 TAPCELL_ASAP7_75t_R TAP_717 ();
 NAND2x2_ASAP7_75t_R _30827_ (.A(net1134),
    .B(_01109_),
    .Y(_01248_));
 TAPCELL_ASAP7_75t_R TAP_716 ();
 AO21x1_ASAP7_75t_R _30829_ (.A1(net1158),
    .A2(_01248_),
    .B(_01243_),
    .Y(_01250_));
 INVx5_ASAP7_75t_R _30830_ (.A(_01243_),
    .Y(_01251_));
 NAND2x2_ASAP7_75t_R _30831_ (.A(net1967),
    .B(_01112_),
    .Y(_01252_));
 INVx1_ASAP7_75t_R _30832_ (.A(_01252_),
    .Y(_01253_));
 NAND2x1_ASAP7_75t_R _30833_ (.A(_01251_),
    .B(_01253_),
    .Y(_01254_));
 NAND3x1_ASAP7_75t_R _30834_ (.A(_01245_),
    .B(_01250_),
    .C(_01254_),
    .Y(_01255_));
 NAND2x2_ASAP7_75t_R _30835_ (.A(_01155_),
    .B(_01242_),
    .Y(_01256_));
 NOR2x2_ASAP7_75t_R _30836_ (.A(_01221_),
    .B(net3315),
    .Y(_01257_));
 TAPCELL_ASAP7_75t_R TAP_715 ();
 NAND2x2_ASAP7_75t_R _30838_ (.A(_01136_),
    .B(net1329),
    .Y(_01259_));
 TAPCELL_ASAP7_75t_R TAP_714 ();
 TAPCELL_ASAP7_75t_R TAP_713 ();
 AOI21x1_ASAP7_75t_R _30841_ (.A1(net2723),
    .A2(_01259_),
    .B(net3315),
    .Y(_01262_));
 AOI21x1_ASAP7_75t_R _30842_ (.A1(net1137),
    .A2(_01257_),
    .B(_01262_),
    .Y(_01263_));
 NOR2x1_ASAP7_75t_R _30843_ (.A(net1431),
    .B(net1196),
    .Y(_01264_));
 INVx3_ASAP7_75t_R _30844_ (.A(_01256_),
    .Y(_01265_));
 NAND2x2_ASAP7_75t_R _30845_ (.A(_01264_),
    .B(_01265_),
    .Y(_01266_));
 INVx1_ASAP7_75t_R _30846_ (.A(_01266_),
    .Y(_01267_));
 NOR2x2_ASAP7_75t_R _30847_ (.A(_01208_),
    .B(net1917),
    .Y(_01268_));
 NAND2x2_ASAP7_75t_R _30848_ (.A(net1593),
    .B(_01096_),
    .Y(_01269_));
 NOR2x2_ASAP7_75t_R _30849_ (.A(_01269_),
    .B(_01159_),
    .Y(_01270_));
 OA21x2_ASAP7_75t_R _30850_ (.A1(_01268_),
    .A2(_01270_),
    .B(_01265_),
    .Y(_01271_));
 NOR2x1_ASAP7_75t_R _30851_ (.A(_01267_),
    .B(_01271_),
    .Y(_01272_));
 NAND2x1_ASAP7_75t_R _30852_ (.A(_01263_),
    .B(_01272_),
    .Y(_01273_));
 NOR2x1_ASAP7_75t_R _30853_ (.A(_01255_),
    .B(_01273_),
    .Y(_01274_));
 TAPCELL_ASAP7_75t_R TAP_712 ();
 NAND2x2_ASAP7_75t_R _30855_ (.A(_01132_),
    .B(_01242_),
    .Y(_01276_));
 TAPCELL_ASAP7_75t_R TAP_711 ();
 NOR2x1_ASAP7_75t_R _30857_ (.A(net1915),
    .B(_01276_),
    .Y(_01278_));
 NOR2x2_ASAP7_75t_R _30858_ (.A(net1195),
    .B(_01112_),
    .Y(_01279_));
 TAPCELL_ASAP7_75t_R TAP_710 ();
 AOI21x1_ASAP7_75t_R _30860_ (.A1(_01226_),
    .A2(net1274),
    .B(_01276_),
    .Y(_01281_));
 TAPCELL_ASAP7_75t_R TAP_709 ();
 AOI21x1_ASAP7_75t_R _30862_ (.A1(net940),
    .A2(net1884),
    .B(_01276_),
    .Y(_01283_));
 AOI211x1_ASAP7_75t_R _30863_ (.A1(_01278_),
    .A2(_01279_),
    .B(_01281_),
    .C(_01283_),
    .Y(_01284_));
 INVx1_ASAP7_75t_R _30864_ (.A(_01284_),
    .Y(_01285_));
 NOR2x2_ASAP7_75t_R _30865_ (.A(net1196),
    .B(_01143_),
    .Y(_01286_));
 NAND2x2_ASAP7_75t_R _30866_ (.A(_01119_),
    .B(_01242_),
    .Y(_01287_));
 INVx4_ASAP7_75t_R _30867_ (.A(_01287_),
    .Y(_01288_));
 TAPCELL_ASAP7_75t_R TAP_708 ();
 TAPCELL_ASAP7_75t_R TAP_707 ();
 NOR2x1_ASAP7_75t_R _30870_ (.A(net1752),
    .B(_01287_),
    .Y(_01291_));
 NAND2x2_ASAP7_75t_R _30871_ (.A(_01136_),
    .B(_01145_),
    .Y(_01292_));
 NOR2x1_ASAP7_75t_R _30872_ (.A(_01292_),
    .B(_01287_),
    .Y(_01293_));
 AOI211x1_ASAP7_75t_R _30873_ (.A1(_01286_),
    .A2(_01288_),
    .B(_01291_),
    .C(_01293_),
    .Y(_01294_));
 TAPCELL_ASAP7_75t_R TAP_706 ();
 AOI211x1_ASAP7_75t_R _30875_ (.A1(net1341),
    .A2(net1277),
    .B(net1916),
    .C(net3145),
    .Y(_01296_));
 AO21x1_ASAP7_75t_R _30876_ (.A1(net1274),
    .A2(_01226_),
    .B(_01287_),
    .Y(_01297_));
 INVx1_ASAP7_75t_R _30877_ (.A(_01297_),
    .Y(_01298_));
 NOR2x1_ASAP7_75t_R _30878_ (.A(_01296_),
    .B(_01298_),
    .Y(_01299_));
 NAND2x1_ASAP7_75t_R _30879_ (.A(_01294_),
    .B(_01299_),
    .Y(_01300_));
 NOR2x1_ASAP7_75t_R _30880_ (.A(_01285_),
    .B(_01300_),
    .Y(_01301_));
 NAND2x1_ASAP7_75t_R _30881_ (.A(_01274_),
    .B(_01301_),
    .Y(_01302_));
 NAND2x2_ASAP7_75t_R _30882_ (.A(_01187_),
    .B(_01112_),
    .Y(_01303_));
 TAPCELL_ASAP7_75t_R TAP_705 ();
 NOR2x2_ASAP7_75t_R _30884_ (.A(_01136_),
    .B(net1426),
    .Y(_01305_));
 INVx5_ASAP7_75t_R _30885_ (.A(_01305_),
    .Y(_01306_));
 NOR2x2_ASAP7_75t_R _30886_ (.A(_00586_),
    .B(_01101_),
    .Y(_01307_));
 NAND2x2_ASAP7_75t_R _30887_ (.A(_01307_),
    .B(_01119_),
    .Y(_01308_));
 TAPCELL_ASAP7_75t_R TAP_704 ();
 AO21x1_ASAP7_75t_R _30889_ (.A1(_01303_),
    .A2(_01306_),
    .B(_01308_),
    .Y(_01310_));
 TAPCELL_ASAP7_75t_R TAP_703 ();
 TAPCELL_ASAP7_75t_R TAP_702 ();
 NAND2x2_ASAP7_75t_R _30892_ (.A(_01125_),
    .B(net1696),
    .Y(_01313_));
 NAND2x2_ASAP7_75t_R _30893_ (.A(net2316),
    .B(_01153_),
    .Y(_01314_));
 INVx4_ASAP7_75t_R _30894_ (.A(_01308_),
    .Y(_01315_));
 OAI21x1_ASAP7_75t_R _30895_ (.A1(_01313_),
    .A2(_01314_),
    .B(_01315_),
    .Y(_01316_));
 NAND2x1_ASAP7_75t_R _30896_ (.A(_01310_),
    .B(_01316_),
    .Y(_01317_));
 NAND2x2_ASAP7_75t_R _30897_ (.A(net1196),
    .B(_01187_),
    .Y(_01318_));
 TAPCELL_ASAP7_75t_R TAP_701 ();
 TAPCELL_ASAP7_75t_R TAP_700 ();
 NAND2x2_ASAP7_75t_R _30900_ (.A(_01208_),
    .B(_01109_),
    .Y(_01321_));
 NAND2x2_ASAP7_75t_R _30901_ (.A(_01132_),
    .B(_01307_),
    .Y(_01322_));
 TAPCELL_ASAP7_75t_R TAP_699 ();
 TAPCELL_ASAP7_75t_R TAP_698 ();
 AO31x2_ASAP7_75t_R _30904_ (.A1(net938),
    .A2(net1158),
    .A3(_01321_),
    .B(net2460),
    .Y(_01325_));
 NOR2x1_ASAP7_75t_R _30905_ (.A(net3341),
    .B(_01322_),
    .Y(_01326_));
 INVx6_ASAP7_75t_R _30906_ (.A(net1698),
    .Y(_01327_));
 NOR2x2_ASAP7_75t_R _30907_ (.A(_01269_),
    .B(_01221_),
    .Y(_01328_));
 INVx4_ASAP7_75t_R _30908_ (.A(_01322_),
    .Y(_01329_));
 OA21x2_ASAP7_75t_R _30909_ (.A1(_01327_),
    .A2(_01328_),
    .B(_01329_),
    .Y(_01330_));
 NOR2x1_ASAP7_75t_R _30910_ (.A(_01326_),
    .B(_01330_),
    .Y(_01331_));
 NAND2x1_ASAP7_75t_R _30911_ (.A(_01325_),
    .B(_01331_),
    .Y(_01332_));
 NOR2x1_ASAP7_75t_R _30912_ (.A(_01317_),
    .B(_01332_),
    .Y(_01333_));
 NAND2x2_ASAP7_75t_R _30913_ (.A(_01169_),
    .B(_01307_),
    .Y(_01334_));
 TAPCELL_ASAP7_75t_R TAP_697 ();
 AOI211x1_ASAP7_75t_R _30915_ (.A1(net2872),
    .A2(net1277),
    .B(_01334_),
    .C(net1432),
    .Y(_01336_));
 CKINVDCx6p67_ASAP7_75t_R _30916_ (.A(_01334_),
    .Y(_01337_));
 TAPCELL_ASAP7_75t_R TAP_696 ();
 OA21x2_ASAP7_75t_R _30918_ (.A1(_01179_),
    .A2(_01270_),
    .B(_01337_),
    .Y(_01339_));
 NOR2x1_ASAP7_75t_R _30919_ (.A(_01336_),
    .B(_01339_),
    .Y(_01340_));
 AO21x1_ASAP7_75t_R _30920_ (.A1(_01125_),
    .A2(net1293),
    .B(_01334_),
    .Y(_01341_));
 NAND2x1_ASAP7_75t_R _30921_ (.A(_01327_),
    .B(_01337_),
    .Y(_01342_));
 AND2x2_ASAP7_75t_R _30922_ (.A(_01341_),
    .B(_01342_),
    .Y(_01343_));
 NAND2x1_ASAP7_75t_R _30923_ (.A(_01340_),
    .B(_01343_),
    .Y(_01344_));
 NAND2x2_ASAP7_75t_R _30924_ (.A(_01155_),
    .B(_01307_),
    .Y(_01345_));
 NOR2x1_ASAP7_75t_R _30925_ (.A(_01125_),
    .B(_01345_),
    .Y(_01346_));
 INVx1_ASAP7_75t_R _30926_ (.A(_01346_),
    .Y(_01347_));
 NAND2x2_ASAP7_75t_R _30927_ (.A(net1593),
    .B(net1970),
    .Y(_01348_));
 AO21x1_ASAP7_75t_R _30928_ (.A1(_01348_),
    .A2(net1698),
    .B(_01345_),
    .Y(_01349_));
 NAND2x1_ASAP7_75t_R _30929_ (.A(_01347_),
    .B(_01349_),
    .Y(_01350_));
 INVx3_ASAP7_75t_R _30930_ (.A(_01345_),
    .Y(_01351_));
 NAND2x1_ASAP7_75t_R _30931_ (.A(_01187_),
    .B(_01351_),
    .Y(_01352_));
 AO21x1_ASAP7_75t_R _30932_ (.A1(_01138_),
    .A2(_01226_),
    .B(_01345_),
    .Y(_01353_));
 NAND2x1_ASAP7_75t_R _30933_ (.A(_01352_),
    .B(_01353_),
    .Y(_01354_));
 NOR2x1_ASAP7_75t_R _30934_ (.A(_01350_),
    .B(_01354_),
    .Y(_01355_));
 INVx1_ASAP7_75t_R _30935_ (.A(_01355_),
    .Y(_01356_));
 NOR2x1_ASAP7_75t_R _30936_ (.A(_01344_),
    .B(_01356_),
    .Y(_01357_));
 NAND2x2_ASAP7_75t_R _30937_ (.A(_01333_),
    .B(_01357_),
    .Y(_01358_));
 NOR2x2_ASAP7_75t_R _30938_ (.A(_01302_),
    .B(_01358_),
    .Y(_01359_));
 NAND2x2_ASAP7_75t_R _30939_ (.A(_01240_),
    .B(_01359_),
    .Y(_01360_));
 AO21x1_ASAP7_75t_R _30940_ (.A1(_01248_),
    .A2(net1915),
    .B(_01287_),
    .Y(_01361_));
 INVx1_ASAP7_75t_R _30941_ (.A(_01361_),
    .Y(_01362_));
 AO21x1_ASAP7_75t_R _30942_ (.A1(_01146_),
    .A2(_01252_),
    .B(_01287_),
    .Y(_01363_));
 NAND2x2_ASAP7_75t_R _30943_ (.A(net1328),
    .B(_01288_),
    .Y(_01364_));
 INVx1_ASAP7_75t_R _30944_ (.A(_01293_),
    .Y(_01365_));
 NAND3x2_ASAP7_75t_R _30945_ (.B(_01364_),
    .C(_01365_),
    .Y(_01366_),
    .A(_01363_));
 NOR2x2_ASAP7_75t_R _30946_ (.A(_01362_),
    .B(_01366_),
    .Y(_01367_));
 TAPCELL_ASAP7_75t_R TAP_695 ();
 OR3x2_ASAP7_75t_R _30948_ (.A(_01101_),
    .B(_01117_),
    .C(_00587_),
    .Y(_01369_));
 NAND3x2_ASAP7_75t_R _30949_ (.B(net3417),
    .C(_01369_),
    .Y(_01370_),
    .A(_01367_));
 NOR3x2_ASAP7_75t_R _30950_ (.B(_01101_),
    .C(_01117_),
    .Y(_01371_),
    .A(_01370_));
 OAI21x1_ASAP7_75t_R _30951_ (.A1(_01270_),
    .A2(_01160_),
    .B(_01337_),
    .Y(_01372_));
 NAND2x1_ASAP7_75t_R _30952_ (.A(_01179_),
    .B(_01337_),
    .Y(_01373_));
 NOR2x2_ASAP7_75t_R _30953_ (.A(net1688),
    .B(net1431),
    .Y(_01374_));
 NAND2x1_ASAP7_75t_R _30954_ (.A(_01374_),
    .B(_01337_),
    .Y(_01375_));
 NAND3x1_ASAP7_75t_R _30955_ (.A(_01372_),
    .B(_01373_),
    .C(_01375_),
    .Y(_01376_));
 TAPCELL_ASAP7_75t_R TAP_694 ();
 TAPCELL_ASAP7_75t_R TAP_693 ();
 AO21x1_ASAP7_75t_R _30958_ (.A1(net938),
    .A2(net1431),
    .B(net3240),
    .Y(_01379_));
 AO21x1_ASAP7_75t_R _30959_ (.A1(net2316),
    .A2(_01259_),
    .B(net3240),
    .Y(_01380_));
 NAND2x1_ASAP7_75t_R _30960_ (.A(_01379_),
    .B(_01380_),
    .Y(_01381_));
 NOR2x1_ASAP7_75t_R _30961_ (.A(_01143_),
    .B(_01334_),
    .Y(_01382_));
 INVx1_ASAP7_75t_R _30962_ (.A(_01382_),
    .Y(_01383_));
 NAND2x2_ASAP7_75t_R _30963_ (.A(_01097_),
    .B(_01145_),
    .Y(_01384_));
 TAPCELL_ASAP7_75t_R TAP_692 ();
 AO21x2_ASAP7_75t_R _30965_ (.A1(net1802),
    .A2(_01348_),
    .B(_01334_),
    .Y(_01386_));
 NAND2x1_ASAP7_75t_R _30966_ (.A(_01383_),
    .B(_01386_),
    .Y(_01387_));
 NOR3x1_ASAP7_75t_R _30967_ (.A(_01376_),
    .B(_01381_),
    .C(_01387_),
    .Y(_01388_));
 AO21x1_ASAP7_75t_R _30968_ (.A1(net1119),
    .A2(net940),
    .B(_01308_),
    .Y(_01389_));
 AO21x1_ASAP7_75t_R _30969_ (.A1(_01138_),
    .A2(net938),
    .B(_01308_),
    .Y(_01390_));
 TAPCELL_ASAP7_75t_R TAP_691 ();
 AO21x1_ASAP7_75t_R _30971_ (.A1(net1076),
    .A2(net1122),
    .B(_01308_),
    .Y(_01392_));
 NAND3x1_ASAP7_75t_R _30972_ (.A(_01389_),
    .B(_01390_),
    .C(_01392_),
    .Y(_01393_));
 NOR2x1_ASAP7_75t_R _30973_ (.A(net2124),
    .B(_01322_),
    .Y(_01394_));
 NOR2x2_ASAP7_75t_R _30974_ (.A(_01322_),
    .B(net2361),
    .Y(_01395_));
 AOI211x1_ASAP7_75t_R _30975_ (.A1(_01329_),
    .A2(_01374_),
    .B(_01394_),
    .C(_01395_),
    .Y(_01396_));
 NOR2x1_ASAP7_75t_R _30976_ (.A(_01322_),
    .B(net1802),
    .Y(_01397_));
 AOI211x1_ASAP7_75t_R _30977_ (.A1(_01328_),
    .A2(_01329_),
    .B(_01397_),
    .C(_01326_),
    .Y(_01398_));
 NAND2x1_ASAP7_75t_R _30978_ (.A(_01396_),
    .B(_01398_),
    .Y(_01399_));
 NOR2x1_ASAP7_75t_R _30979_ (.A(_01393_),
    .B(_01399_),
    .Y(_01400_));
 NAND2x1_ASAP7_75t_R _30980_ (.A(_01388_),
    .B(_01400_),
    .Y(_01401_));
 NOR2x2_ASAP7_75t_R _30981_ (.A(net1826),
    .B(_01243_),
    .Y(_01402_));
 AOI21x1_ASAP7_75t_R _30982_ (.A1(net1277),
    .A2(_01244_),
    .B(_01402_),
    .Y(_01403_));
 AOI21x1_ASAP7_75t_R _30983_ (.A1(_01318_),
    .A2(_01188_),
    .B(_01243_),
    .Y(_01404_));
 NOR2x2_ASAP7_75t_R _30984_ (.A(net1430),
    .B(_01269_),
    .Y(_01405_));
 NOR2x2_ASAP7_75t_R _30985_ (.A(net1431),
    .B(_01178_),
    .Y(_01406_));
 OA21x2_ASAP7_75t_R _30986_ (.A1(_01405_),
    .A2(_01406_),
    .B(_01251_),
    .Y(_01407_));
 NOR2x1_ASAP7_75t_R _30987_ (.A(_01404_),
    .B(_01407_),
    .Y(_01408_));
 NAND2x1_ASAP7_75t_R _30988_ (.A(_01403_),
    .B(_01408_),
    .Y(_01409_));
 NOR2x2_ASAP7_75t_R _30989_ (.A(net2393),
    .B(net3315),
    .Y(_01410_));
 AOI21x1_ASAP7_75t_R _30990_ (.A1(net1137),
    .A2(_01257_),
    .B(_01410_),
    .Y(_01411_));
 AO21x2_ASAP7_75t_R _30991_ (.A1(net2120),
    .A2(net1142),
    .B(net3315),
    .Y(_01412_));
 NAND3x1_ASAP7_75t_R _30992_ (.A(_01411_),
    .B(_01266_),
    .C(_01412_),
    .Y(_01413_));
 NOR2x1_ASAP7_75t_R _30993_ (.A(_01409_),
    .B(_01413_),
    .Y(_01414_));
 AO21x2_ASAP7_75t_R _30994_ (.A1(_01172_),
    .A2(_01194_),
    .B(_01276_),
    .Y(_01415_));
 CKINVDCx5p33_ASAP7_75t_R _30995_ (.A(_01276_),
    .Y(_01416_));
 NAND2x1_ASAP7_75t_R _30996_ (.A(net1969),
    .B(_01416_),
    .Y(_01417_));
 NAND2x2_ASAP7_75t_R _30997_ (.A(_01166_),
    .B(_01416_),
    .Y(_01418_));
 NAND3x1_ASAP7_75t_R _30998_ (.A(_01415_),
    .B(_01417_),
    .C(_01418_),
    .Y(_01419_));
 AO21x1_ASAP7_75t_R _30999_ (.A1(_01153_),
    .A2(net3138),
    .B(net3145),
    .Y(_01420_));
 AO21x1_ASAP7_75t_R _31000_ (.A1(_01303_),
    .A2(net938),
    .B(net3145),
    .Y(_01421_));
 NAND2x1_ASAP7_75t_R _31001_ (.A(_01420_),
    .B(_01421_),
    .Y(_01422_));
 AO21x2_ASAP7_75t_R _31002_ (.A1(_01303_),
    .A2(net1142),
    .B(_01276_),
    .Y(_01423_));
 AO21x1_ASAP7_75t_R _31003_ (.A1(net1274),
    .A2(_01306_),
    .B(net3417),
    .Y(_01424_));
 NAND2x1_ASAP7_75t_R _31004_ (.A(_01423_),
    .B(_01424_),
    .Y(_01425_));
 NOR3x1_ASAP7_75t_R _31005_ (.A(_01419_),
    .B(_01422_),
    .C(_01425_),
    .Y(_01426_));
 NAND2x1_ASAP7_75t_R _31006_ (.A(_01414_),
    .B(_01426_),
    .Y(_01427_));
 NOR2x2_ASAP7_75t_R _31007_ (.A(_01401_),
    .B(_01427_),
    .Y(_01428_));
 NOR2x2_ASAP7_75t_R _31008_ (.A(_01202_),
    .B(_01113_),
    .Y(_01429_));
 AOI211x1_ASAP7_75t_R _31009_ (.A1(net1341),
    .A2(net1277),
    .B(_01202_),
    .C(net1919),
    .Y(_01430_));
 NOR2x1_ASAP7_75t_R _31010_ (.A(_01429_),
    .B(_01430_),
    .Y(_01431_));
 AOI211x1_ASAP7_75t_R _31011_ (.A1(net1593),
    .A2(net1685),
    .B(_01202_),
    .C(_01204_),
    .Y(_01432_));
 AO21x2_ASAP7_75t_R _31012_ (.A1(net3321),
    .A2(_01252_),
    .B(_01202_),
    .Y(_01433_));
 INVx1_ASAP7_75t_R _31013_ (.A(_01433_),
    .Y(_01434_));
 NOR2x1_ASAP7_75t_R _31014_ (.A(_01432_),
    .B(_01434_),
    .Y(_01435_));
 NAND2x1_ASAP7_75t_R _31015_ (.A(_01431_),
    .B(_01435_),
    .Y(_01436_));
 TAPCELL_ASAP7_75t_R TAP_690 ();
 AO21x1_ASAP7_75t_R _31017_ (.A1(net2652),
    .A2(net2120),
    .B(net3144),
    .Y(_01438_));
 AOI21x1_ASAP7_75t_R _31018_ (.A1(net1294),
    .A2(_01172_),
    .B(_01191_),
    .Y(_01439_));
 NOR2x1_ASAP7_75t_R _31019_ (.A(_01128_),
    .B(_01191_),
    .Y(_01440_));
 AOI211x1_ASAP7_75t_R _31020_ (.A1(_01197_),
    .A2(_01327_),
    .B(_01439_),
    .C(_01440_),
    .Y(_01441_));
 NAND2x1_ASAP7_75t_R _31021_ (.A(_01438_),
    .B(_01441_),
    .Y(_01442_));
 NOR2x1_ASAP7_75t_R _31022_ (.A(_01436_),
    .B(_01442_),
    .Y(_01443_));
 AOI211x1_ASAP7_75t_R _31023_ (.A1(net1341),
    .A2(net1685),
    .B(net1919),
    .C(_01229_),
    .Y(_01444_));
 OA21x2_ASAP7_75t_R _31024_ (.A1(_01209_),
    .A2(_01305_),
    .B(_01234_),
    .Y(_01445_));
 NOR2x1_ASAP7_75t_R _31025_ (.A(_01444_),
    .B(_01445_),
    .Y(_01446_));
 NAND2x2_ASAP7_75t_R _31026_ (.A(net1329),
    .B(_01208_),
    .Y(_01447_));
 NOR2x1_ASAP7_75t_R _31027_ (.A(_01447_),
    .B(_01229_),
    .Y(_01448_));
 AOI21x1_ASAP7_75t_R _31028_ (.A1(_01269_),
    .A2(_01448_),
    .B(_01232_),
    .Y(_01449_));
 NAND2x1_ASAP7_75t_R _31029_ (.A(_01446_),
    .B(_01449_),
    .Y(_01450_));
 OA21x2_ASAP7_75t_R _31030_ (.A1(_01270_),
    .A2(_01160_),
    .B(_01218_),
    .Y(_01451_));
 OA21x2_ASAP7_75t_R _31031_ (.A1(_01209_),
    .A2(_01305_),
    .B(_01218_),
    .Y(_01452_));
 NAND2x2_ASAP7_75t_R _31032_ (.A(net1687),
    .B(net1330),
    .Y(_01453_));
 AOI21x1_ASAP7_75t_R _31033_ (.A1(_01453_),
    .A2(net1752),
    .B(_01215_),
    .Y(_01454_));
 OR3x1_ASAP7_75t_R _31034_ (.A(_01451_),
    .B(_01452_),
    .C(_01454_),
    .Y(_01455_));
 NOR2x1_ASAP7_75t_R _31035_ (.A(_01450_),
    .B(_01455_),
    .Y(_01456_));
 NAND2x1_ASAP7_75t_R _31036_ (.A(_01443_),
    .B(_01456_),
    .Y(_01457_));
 AO21x2_ASAP7_75t_R _31037_ (.A1(_01113_),
    .A2(_01226_),
    .B(_01120_),
    .Y(_01458_));
 AO21x1_ASAP7_75t_R _31038_ (.A1(net2522),
    .A2(net1884),
    .B(_01120_),
    .Y(_01459_));
 NAND2x2_ASAP7_75t_R _31039_ (.A(_01103_),
    .B(_01270_),
    .Y(_01460_));
 NAND3x1_ASAP7_75t_R _31040_ (.A(_01458_),
    .B(_01459_),
    .C(_01460_),
    .Y(_01461_));
 AO21x1_ASAP7_75t_R _31041_ (.A1(net2120),
    .A2(_01318_),
    .B(_01133_),
    .Y(_01462_));
 AO21x1_ASAP7_75t_R _31042_ (.A1(_01138_),
    .A2(_01226_),
    .B(_01133_),
    .Y(_01463_));
 AND2x2_ASAP7_75t_R _31043_ (.A(_01462_),
    .B(_01463_),
    .Y(_01464_));
 AO21x1_ASAP7_75t_R _31044_ (.A1(net3321),
    .A2(net1802),
    .B(_01133_),
    .Y(_01465_));
 AO21x1_ASAP7_75t_R _31045_ (.A1(_01172_),
    .A2(_01128_),
    .B(_01133_),
    .Y(_01466_));
 AND2x2_ASAP7_75t_R _31046_ (.A(_01465_),
    .B(_01466_),
    .Y(_01467_));
 NAND2x1_ASAP7_75t_R _31047_ (.A(_01464_),
    .B(_01467_),
    .Y(_01468_));
 NOR2x1_ASAP7_75t_R _31048_ (.A(_01461_),
    .B(_01468_),
    .Y(_01469_));
 INVx1_ASAP7_75t_R _31049_ (.A(_01181_),
    .Y(_01470_));
 NAND2x1_ASAP7_75t_R _31050_ (.A(_01305_),
    .B(_01171_),
    .Y(_01471_));
 AO21x1_ASAP7_75t_R _31051_ (.A1(net3138),
    .A2(_01292_),
    .B(_01170_),
    .Y(_01472_));
 NAND3x1_ASAP7_75t_R _31052_ (.A(_01470_),
    .B(_01471_),
    .C(_01472_),
    .Y(_01473_));
 NOR2x2_ASAP7_75t_R _31053_ (.A(net1431),
    .B(net1135),
    .Y(_01474_));
 AOI221x1_ASAP7_75t_R _31054_ (.A1(net2872),
    .A2(net3289),
    .B1(_01204_),
    .B2(_01221_),
    .C(_01156_),
    .Y(_01475_));
 AO21x1_ASAP7_75t_R _31055_ (.A1(_01474_),
    .A2(_01163_),
    .B(_01475_),
    .Y(_01476_));
 NOR2x1_ASAP7_75t_R _31056_ (.A(_01473_),
    .B(_01476_),
    .Y(_01477_));
 NAND2x1_ASAP7_75t_R _31057_ (.A(_01469_),
    .B(_01477_),
    .Y(_01478_));
 NOR2x2_ASAP7_75t_R _31058_ (.A(_01457_),
    .B(_01478_),
    .Y(_01479_));
 NAND2x2_ASAP7_75t_R _31059_ (.A(_01428_),
    .B(_01479_),
    .Y(_01480_));
 OA21x2_ASAP7_75t_R _31060_ (.A1(_01360_),
    .A2(_01371_),
    .B(_01480_),
    .Y(_01481_));
 NOR3x2_ASAP7_75t_R _31061_ (.B(net2689),
    .C(_01371_),
    .Y(_01482_),
    .A(_01480_));
 NOR2x2_ASAP7_75t_R _31062_ (.A(_01481_),
    .B(_01482_),
    .Y(_01483_));
 NAND2x1_ASAP7_75t_R _31063_ (.A(net2362),
    .B(_01483_),
    .Y(_01484_));
 INVx1_ASAP7_75t_R _31064_ (.A(_01482_),
    .Y(_01485_));
 INVx1_ASAP7_75t_R _31065_ (.A(_01481_),
    .Y(_01486_));
 AO21x1_ASAP7_75t_R _31066_ (.A1(_01485_),
    .A2(_01486_),
    .B(net2362),
    .Y(_01487_));
 TAPCELL_ASAP7_75t_R TAP_689 ();
 TAPCELL_ASAP7_75t_R TAP_688 ();
 TAPCELL_ASAP7_75t_R TAP_687 ();
 NOR2x2_ASAP7_75t_R _31070_ (.A(net2623),
    .B(_00638_),
    .Y(_01491_));
 TAPCELL_ASAP7_75t_R TAP_686 ();
 TAPCELL_ASAP7_75t_R TAP_685 ();
 CKINVDCx14_ASAP7_75t_R _31073_ (.A(net1896),
    .Y(_01494_));
 NOR2x2_ASAP7_75t_R _31074_ (.A(net1635),
    .B(_01494_),
    .Y(_01495_));
 NAND2x2_ASAP7_75t_R _31075_ (.A(_01491_),
    .B(_01495_),
    .Y(_01496_));
 TAPCELL_ASAP7_75t_R TAP_684 ();
 CKINVDCx20_ASAP7_75t_R _31077_ (.A(net1635),
    .Y(_01498_));
 NAND2x2_ASAP7_75t_R _31078_ (.A(net1896),
    .B(_01498_),
    .Y(_01499_));
 NAND2x2_ASAP7_75t_R _31079_ (.A(net1575),
    .B(_01499_),
    .Y(_01500_));
 NAND2x2_ASAP7_75t_R _31080_ (.A(_00635_),
    .B(_00636_),
    .Y(_01501_));
 TAPCELL_ASAP7_75t_R TAP_683 ();
 NAND2x2_ASAP7_75t_R _31082_ (.A(net2777),
    .B(_00634_),
    .Y(_01503_));
 NOR2x2_ASAP7_75t_R _31083_ (.A(_01501_),
    .B(_01503_),
    .Y(_01504_));
 CKINVDCx6p67_ASAP7_75t_R _31084_ (.A(_01504_),
    .Y(_01505_));
 AO21x1_ASAP7_75t_R _31085_ (.A1(net3415),
    .A2(_01500_),
    .B(_01505_),
    .Y(_01506_));
 INVx1_ASAP7_75t_R _31086_ (.A(_01506_),
    .Y(_01507_));
 TAPCELL_ASAP7_75t_R TAP_682 ();
 INVx4_ASAP7_75t_R _31088_ (.A(net2623),
    .Y(_01509_));
 NAND2x2_ASAP7_75t_R _31089_ (.A(net3129),
    .B(_01509_),
    .Y(_01510_));
 NOR2x2_ASAP7_75t_R _31090_ (.A(_01510_),
    .B(net1641),
    .Y(_01511_));
 NAND2x1_ASAP7_75t_R _31091_ (.A(_01504_),
    .B(_01511_),
    .Y(_01512_));
 NAND2x2_ASAP7_75t_R _31092_ (.A(net1637),
    .B(net1900),
    .Y(_01513_));
 NOR2x2_ASAP7_75t_R _31093_ (.A(net1025),
    .B(net2073),
    .Y(_01514_));
 NAND2x2_ASAP7_75t_R _31094_ (.A(net1635),
    .B(_01494_),
    .Y(_01515_));
 NOR2x2_ASAP7_75t_R _31095_ (.A(_01515_),
    .B(_01510_),
    .Y(_01516_));
 OAI21x1_ASAP7_75t_R _31096_ (.A1(_01514_),
    .A2(_01516_),
    .B(_01504_),
    .Y(_01517_));
 NAND2x1_ASAP7_75t_R _31097_ (.A(_01512_),
    .B(_01517_),
    .Y(_01518_));
 NOR2x2_ASAP7_75t_R _31098_ (.A(_01507_),
    .B(_01518_),
    .Y(_01519_));
 INVx3_ASAP7_75t_R _31099_ (.A(_00638_),
    .Y(_01520_));
 NAND2x2_ASAP7_75t_R _31100_ (.A(net2624),
    .B(_01520_),
    .Y(_01521_));
 TAPCELL_ASAP7_75t_R TAP_681 ();
 TAPCELL_ASAP7_75t_R TAP_680 ();
 NAND2x2_ASAP7_75t_R _31103_ (.A(net2623),
    .B(_00638_),
    .Y(_01524_));
 NOR2x2_ASAP7_75t_R _31104_ (.A(net1635),
    .B(_01524_),
    .Y(_01525_));
 NOR2x2_ASAP7_75t_R _31105_ (.A(_01515_),
    .B(_01524_),
    .Y(_01526_));
 OAI21x1_ASAP7_75t_R _31106_ (.A1(_01525_),
    .A2(_01526_),
    .B(_01504_),
    .Y(_01527_));
 OA21x2_ASAP7_75t_R _31107_ (.A1(net2379),
    .A2(_01505_),
    .B(_01527_),
    .Y(_01528_));
 INVx2_ASAP7_75t_R _31108_ (.A(_00635_),
    .Y(_01529_));
 NOR2x2_ASAP7_75t_R _31109_ (.A(_00636_),
    .B(_01529_),
    .Y(_01530_));
 INVx3_ASAP7_75t_R _31110_ (.A(_01503_),
    .Y(_01531_));
 NAND2x2_ASAP7_75t_R _31111_ (.A(_01530_),
    .B(_01531_),
    .Y(_01532_));
 TAPCELL_ASAP7_75t_R TAP_679 ();
 NAND3x2_ASAP7_75t_R _31113_ (.B(_01528_),
    .C(net2334),
    .Y(_01534_),
    .A(_01519_));
 INVx2_ASAP7_75t_R _31114_ (.A(net2777),
    .Y(_01535_));
 NOR2x2_ASAP7_75t_R _31115_ (.A(_00634_),
    .B(_01535_),
    .Y(_01536_));
 AND3x2_ASAP7_75t_R _31116_ (.A(_01529_),
    .B(net2777),
    .C(_00634_),
    .Y(_01537_));
 NOR3x2_ASAP7_75t_R _31117_ (.B(_01536_),
    .C(_01537_),
    .Y(_01538_),
    .A(_01534_));
 NAND2x2_ASAP7_75t_R _31118_ (.A(net2779),
    .B(_01538_),
    .Y(_01539_));
 NAND2x2_ASAP7_75t_R _31119_ (.A(_01498_),
    .B(net1573),
    .Y(_01540_));
 TAPCELL_ASAP7_75t_R TAP_678 ();
 TAPCELL_ASAP7_75t_R TAP_677 ();
 NAND2x2_ASAP7_75t_R _31122_ (.A(_01536_),
    .B(_01530_),
    .Y(_01543_));
 TAPCELL_ASAP7_75t_R TAP_676 ();
 TAPCELL_ASAP7_75t_R TAP_675 ();
 TAPCELL_ASAP7_75t_R TAP_674 ();
 AOI211x1_ASAP7_75t_R _31126_ (.A1(_01540_),
    .A2(net2080),
    .B(_01543_),
    .C(net1263),
    .Y(_01547_));
 TAPCELL_ASAP7_75t_R TAP_673 ();
 NOR2x2_ASAP7_75t_R _31128_ (.A(net1240),
    .B(net3153),
    .Y(_01549_));
 INVx4_ASAP7_75t_R _31129_ (.A(_01543_),
    .Y(_01550_));
 NAND2x1_ASAP7_75t_R _31130_ (.A(_01549_),
    .B(_01550_),
    .Y(_01551_));
 NOR2x2_ASAP7_75t_R _31131_ (.A(net3129),
    .B(_01509_),
    .Y(_01552_));
 NAND2x2_ASAP7_75t_R _31132_ (.A(net3416),
    .B(_01552_),
    .Y(_01553_));
 TAPCELL_ASAP7_75t_R TAP_672 ();
 NOR2x2_ASAP7_75t_R _31134_ (.A(net1635),
    .B(net1896),
    .Y(_01555_));
 NAND2x2_ASAP7_75t_R _31135_ (.A(_01555_),
    .B(_01552_),
    .Y(_01556_));
 TAPCELL_ASAP7_75t_R TAP_671 ();
 AO21x1_ASAP7_75t_R _31137_ (.A1(net2062),
    .A2(net2254),
    .B(_01543_),
    .Y(_01558_));
 NAND2x1_ASAP7_75t_R _31138_ (.A(_01551_),
    .B(_01558_),
    .Y(_01559_));
 NOR2x1_ASAP7_75t_R _31139_ (.A(_01547_),
    .B(_01559_),
    .Y(_01560_));
 NAND2x2_ASAP7_75t_R _31140_ (.A(_01498_),
    .B(_01494_),
    .Y(_01561_));
 NOR2x2_ASAP7_75t_R _31141_ (.A(net2073),
    .B(_01561_),
    .Y(_01562_));
 INVx2_ASAP7_75t_R _31142_ (.A(_00634_),
    .Y(_01563_));
 NAND2x1_ASAP7_75t_R _31143_ (.A(net2778),
    .B(_01563_),
    .Y(_01564_));
 NOR2x2_ASAP7_75t_R _31144_ (.A(_01501_),
    .B(_01564_),
    .Y(_01565_));
 TAPCELL_ASAP7_75t_R TAP_670 ();
 OAI21x1_ASAP7_75t_R _31146_ (.A1(_01516_),
    .A2(_01562_),
    .B(_01565_),
    .Y(_01567_));
 TAPCELL_ASAP7_75t_R TAP_669 ();
 NAND2x2_ASAP7_75t_R _31148_ (.A(net1636),
    .B(net1575),
    .Y(_01569_));
 INVx3_ASAP7_75t_R _31149_ (.A(_01501_),
    .Y(_01570_));
 NAND2x2_ASAP7_75t_R _31150_ (.A(_01536_),
    .B(_01570_),
    .Y(_01571_));
 TAPCELL_ASAP7_75t_R TAP_668 ();
 AO21x1_ASAP7_75t_R _31152_ (.A1(net1104),
    .A2(_01569_),
    .B(_01571_),
    .Y(_01573_));
 NAND2x2_ASAP7_75t_R _31153_ (.A(_01567_),
    .B(_01573_),
    .Y(_01574_));
 NOR2x2_ASAP7_75t_R _31154_ (.A(_01498_),
    .B(net1241),
    .Y(_01575_));
 INVx4_ASAP7_75t_R _31155_ (.A(_01513_),
    .Y(_01576_));
 NAND2x2_ASAP7_75t_R _31156_ (.A(_01552_),
    .B(_01576_),
    .Y(_01577_));
 NOR2x1_ASAP7_75t_R _31157_ (.A(_01571_),
    .B(net2572),
    .Y(_01578_));
 AO21x1_ASAP7_75t_R _31158_ (.A1(_01565_),
    .A2(_01575_),
    .B(_01578_),
    .Y(_01579_));
 NOR2x1_ASAP7_75t_R _31159_ (.A(_01574_),
    .B(_01579_),
    .Y(_01580_));
 NAND2x1_ASAP7_75t_R _31160_ (.A(_01560_),
    .B(_01580_),
    .Y(_01581_));
 NOR2x2_ASAP7_75t_R _31161_ (.A(net1899),
    .B(net1241),
    .Y(_01582_));
 INVx1_ASAP7_75t_R _31162_ (.A(_01582_),
    .Y(_01583_));
 INVx1_ASAP7_75t_R _31163_ (.A(_00636_),
    .Y(_01584_));
 NOR2x2_ASAP7_75t_R _31164_ (.A(_00635_),
    .B(_01584_),
    .Y(_01585_));
 NAND2x2_ASAP7_75t_R _31165_ (.A(_01536_),
    .B(_01585_),
    .Y(_01586_));
 TAPCELL_ASAP7_75t_R TAP_667 ();
 AO21x1_ASAP7_75t_R _31167_ (.A1(_01583_),
    .A2(net2381),
    .B(net2348),
    .Y(_01588_));
 NOR2x2_ASAP7_75t_R _31168_ (.A(net2623),
    .B(_01520_),
    .Y(_01589_));
 NAND2x2_ASAP7_75t_R _31169_ (.A(_01555_),
    .B(net1887),
    .Y(_01590_));
 TAPCELL_ASAP7_75t_R TAP_666 ();
 NAND2x2_ASAP7_75t_R _31171_ (.A(net1638),
    .B(_01589_),
    .Y(_01592_));
 TAPCELL_ASAP7_75t_R TAP_665 ();
 AO21x1_ASAP7_75t_R _31173_ (.A1(net1597),
    .A2(net3255),
    .B(net2348),
    .Y(_01594_));
 NOR2x1_ASAP7_75t_R _31174_ (.A(net2795),
    .B(_01586_),
    .Y(_01595_));
 INVx1_ASAP7_75t_R _31175_ (.A(_01595_),
    .Y(_01596_));
 AND3x1_ASAP7_75t_R _31176_ (.A(_01588_),
    .B(_01594_),
    .C(_01596_),
    .Y(_01597_));
 INVx3_ASAP7_75t_R _31177_ (.A(_01575_),
    .Y(_01598_));
 CKINVDCx6p67_ASAP7_75t_R _31178_ (.A(_01524_),
    .Y(_01599_));
 NAND2x2_ASAP7_75t_R _31179_ (.A(_01555_),
    .B(_01599_),
    .Y(_01600_));
 TAPCELL_ASAP7_75t_R TAP_664 ();
 NOR2x2_ASAP7_75t_R _31181_ (.A(_00635_),
    .B(_00636_),
    .Y(_01602_));
 NAND2x2_ASAP7_75t_R _31182_ (.A(_01602_),
    .B(_01536_),
    .Y(_01603_));
 TAPCELL_ASAP7_75t_R TAP_663 ();
 AO21x1_ASAP7_75t_R _31184_ (.A1(_01598_),
    .A2(_01600_),
    .B(net2275),
    .Y(_01605_));
 NOR2x2_ASAP7_75t_R _31185_ (.A(net1896),
    .B(_01498_),
    .Y(_01606_));
 NAND2x2_ASAP7_75t_R _31186_ (.A(_01606_),
    .B(_01552_),
    .Y(_01607_));
 AO21x1_ASAP7_75t_R _31187_ (.A1(net2366),
    .A2(net2256),
    .B(_01603_),
    .Y(_01608_));
 NAND2x1_ASAP7_75t_R _31188_ (.A(_01605_),
    .B(_01608_),
    .Y(_01609_));
 TAPCELL_ASAP7_75t_R TAP_662 ();
 TAPCELL_ASAP7_75t_R TAP_661 ();
 NAND2x2_ASAP7_75t_R _31191_ (.A(_01491_),
    .B(_01606_),
    .Y(_01612_));
 TAPCELL_ASAP7_75t_R TAP_660 ();
 AO21x1_ASAP7_75t_R _31193_ (.A1(net2795),
    .A2(_01612_),
    .B(_01603_),
    .Y(_01614_));
 OAI21x1_ASAP7_75t_R _31194_ (.A1(net1597),
    .A2(net2275),
    .B(_01614_),
    .Y(_01615_));
 NOR2x1_ASAP7_75t_R _31195_ (.A(_01609_),
    .B(_01615_),
    .Y(_01616_));
 NAND2x1_ASAP7_75t_R _31196_ (.A(_01597_),
    .B(_01616_),
    .Y(_01617_));
 NOR2x1_ASAP7_75t_R _31197_ (.A(_01581_),
    .B(_01617_),
    .Y(_01618_));
 NOR2x2_ASAP7_75t_R _31198_ (.A(net1240),
    .B(net1400),
    .Y(_01619_));
 NAND2x1_ASAP7_75t_R _31199_ (.A(_00636_),
    .B(_01529_),
    .Y(_01620_));
 NOR2x2_ASAP7_75t_R _31200_ (.A(_01503_),
    .B(_01620_),
    .Y(_01621_));
 NAND2x2_ASAP7_75t_R _31201_ (.A(_01619_),
    .B(_01621_),
    .Y(_01622_));
 TAPCELL_ASAP7_75t_R TAP_659 ();
 NAND2x2_ASAP7_75t_R _31203_ (.A(_01585_),
    .B(_01531_),
    .Y(_01624_));
 TAPCELL_ASAP7_75t_R TAP_658 ();
 AO21x1_ASAP7_75t_R _31205_ (.A1(net2366),
    .A2(net1613),
    .B(_01624_),
    .Y(_01626_));
 NAND2x1_ASAP7_75t_R _31206_ (.A(_01622_),
    .B(_01626_),
    .Y(_01627_));
 NOR2x1_ASAP7_75t_R _31207_ (.A(net2077),
    .B(_01576_),
    .Y(_01628_));
 INVx1_ASAP7_75t_R _31208_ (.A(_01628_),
    .Y(_01629_));
 NAND2x2_ASAP7_75t_R _31209_ (.A(_01491_),
    .B(_01576_),
    .Y(_01630_));
 TAPCELL_ASAP7_75t_R TAP_657 ();
 AO21x1_ASAP7_75t_R _31211_ (.A1(_01630_),
    .A2(_01540_),
    .B(_01624_),
    .Y(_01632_));
 OAI21x1_ASAP7_75t_R _31212_ (.A1(_01624_),
    .A2(_01629_),
    .B(_01632_),
    .Y(_01633_));
 NOR2x1_ASAP7_75t_R _31213_ (.A(_01627_),
    .B(_01633_),
    .Y(_01634_));
 NOR2x2_ASAP7_75t_R _31214_ (.A(_01499_),
    .B(net2376),
    .Y(_01635_));
 NAND2x2_ASAP7_75t_R _31215_ (.A(_01602_),
    .B(_01531_),
    .Y(_01636_));
 INVx4_ASAP7_75t_R _31216_ (.A(_01636_),
    .Y(_01637_));
 NAND2x1_ASAP7_75t_R _31217_ (.A(_01635_),
    .B(_01637_),
    .Y(_01638_));
 OAI21x1_ASAP7_75t_R _31218_ (.A1(_01525_),
    .A2(_01526_),
    .B(_01637_),
    .Y(_01639_));
 NAND2x1_ASAP7_75t_R _31219_ (.A(_01638_),
    .B(_01639_),
    .Y(_01640_));
 NAND2x2_ASAP7_75t_R _31220_ (.A(net1887),
    .B(_01576_),
    .Y(_01641_));
 NOR2x1_ASAP7_75t_R _31221_ (.A(_01636_),
    .B(_01641_),
    .Y(_01642_));
 TAPCELL_ASAP7_75t_R TAP_656 ();
 INVx11_ASAP7_75t_R _31223_ (.A(net1574),
    .Y(_01644_));
 TAPCELL_ASAP7_75t_R TAP_655 ();
 TAPCELL_ASAP7_75t_R TAP_654 ();
 AOI211x1_ASAP7_75t_R _31226_ (.A1(_01498_),
    .A2(net1263),
    .B(_01644_),
    .C(net2746),
    .Y(_01647_));
 NOR3x1_ASAP7_75t_R _31227_ (.A(_01640_),
    .B(_01642_),
    .C(_01647_),
    .Y(_01648_));
 NAND2x1_ASAP7_75t_R _31228_ (.A(_01634_),
    .B(_01648_),
    .Y(_01649_));
 TAPCELL_ASAP7_75t_R TAP_653 ();
 TAPCELL_ASAP7_75t_R TAP_652 ();
 AO21x1_ASAP7_75t_R _31231_ (.A1(net1104),
    .A2(net1457),
    .B(_01505_),
    .Y(_01652_));
 OA21x2_ASAP7_75t_R _31232_ (.A1(_01505_),
    .A2(_01629_),
    .B(_01652_),
    .Y(_01653_));
 TAPCELL_ASAP7_75t_R TAP_651 ();
 AOI211x1_ASAP7_75t_R _31234_ (.A1(net1120),
    .A2(net1263),
    .B(_01505_),
    .C(net2379),
    .Y(_01655_));
 AOI21x1_ASAP7_75t_R _31235_ (.A1(_01504_),
    .A2(_01525_),
    .B(_01655_),
    .Y(_01656_));
 INVx5_ASAP7_75t_R _31236_ (.A(_01532_),
    .Y(_01657_));
 TAPCELL_ASAP7_75t_R TAP_650 ();
 TAPCELL_ASAP7_75t_R TAP_649 ();
 AOI21x1_ASAP7_75t_R _31239_ (.A1(net2366),
    .A2(net1613),
    .B(_01532_),
    .Y(_01660_));
 AOI21x1_ASAP7_75t_R _31240_ (.A1(_01590_),
    .A2(_01641_),
    .B(_01532_),
    .Y(_01661_));
 AOI211x1_ASAP7_75t_R _31241_ (.A1(_01525_),
    .A2(_01657_),
    .B(_01660_),
    .C(_01661_),
    .Y(_01662_));
 NAND3x2_ASAP7_75t_R _31242_ (.B(_01656_),
    .C(_01662_),
    .Y(_01663_),
    .A(_01653_));
 NOR2x2_ASAP7_75t_R _31243_ (.A(_01649_),
    .B(_01663_),
    .Y(_01664_));
 NAND2x2_ASAP7_75t_R _31244_ (.A(_01618_),
    .B(_01664_),
    .Y(_01665_));
 TAPCELL_ASAP7_75t_R TAP_648 ();
 NOR2x2_ASAP7_75t_R _31246_ (.A(net2777),
    .B(_01563_),
    .Y(_01667_));
 NAND2x2_ASAP7_75t_R _31247_ (.A(_01585_),
    .B(_01667_),
    .Y(_01668_));
 TAPCELL_ASAP7_75t_R TAP_647 ();
 NAND2x2_ASAP7_75t_R _31249_ (.A(_01606_),
    .B(net2585),
    .Y(_01670_));
 TAPCELL_ASAP7_75t_R TAP_646 ();
 AO21x2_ASAP7_75t_R _31251_ (.A1(net3135),
    .A2(_01500_),
    .B(_01668_),
    .Y(_01672_));
 OA21x2_ASAP7_75t_R _31252_ (.A1(net2572),
    .A2(_01668_),
    .B(_01672_),
    .Y(_01673_));
 NAND2x2_ASAP7_75t_R _31253_ (.A(net1639),
    .B(_01552_),
    .Y(_01674_));
 NAND2x2_ASAP7_75t_R _31254_ (.A(_01602_),
    .B(_01667_),
    .Y(_01675_));
 TAPCELL_ASAP7_75t_R TAP_645 ();
 AO21x1_ASAP7_75t_R _31256_ (.A1(net2254),
    .A2(_01674_),
    .B(_01675_),
    .Y(_01677_));
 NAND2x2_ASAP7_75t_R _31257_ (.A(_01515_),
    .B(_01599_),
    .Y(_01678_));
 OR2x2_ASAP7_75t_R _31258_ (.A(_01675_),
    .B(_01678_),
    .Y(_01679_));
 NOR2x2_ASAP7_75t_R _31259_ (.A(net1025),
    .B(_01644_),
    .Y(_01680_));
 INVx3_ASAP7_75t_R _31260_ (.A(_01675_),
    .Y(_01681_));
 NAND2x1_ASAP7_75t_R _31261_ (.A(_01680_),
    .B(_01681_),
    .Y(_01682_));
 AND3x1_ASAP7_75t_R _31262_ (.A(_01677_),
    .B(_01679_),
    .C(_01682_),
    .Y(_01683_));
 NAND2x1_ASAP7_75t_R _31263_ (.A(_01673_),
    .B(_01683_),
    .Y(_01684_));
 NAND2x2_ASAP7_75t_R _31264_ (.A(_01570_),
    .B(_01667_),
    .Y(_01685_));
 TAPCELL_ASAP7_75t_R TAP_644 ();
 NAND2x2_ASAP7_75t_R _31266_ (.A(_01499_),
    .B(net3146),
    .Y(_01687_));
 NOR2x2_ASAP7_75t_R _31267_ (.A(_01513_),
    .B(_01524_),
    .Y(_01688_));
 CKINVDCx6p67_ASAP7_75t_R _31268_ (.A(_01688_),
    .Y(_01689_));
 TAPCELL_ASAP7_75t_R TAP_643 ();
 NAND2x2_ASAP7_75t_R _31270_ (.A(net3416),
    .B(_01599_),
    .Y(_01691_));
 TAPCELL_ASAP7_75t_R TAP_642 ();
 AO21x1_ASAP7_75t_R _31272_ (.A1(_01689_),
    .A2(_01691_),
    .B(_01685_),
    .Y(_01693_));
 OA21x2_ASAP7_75t_R _31273_ (.A1(_01685_),
    .A2(_01687_),
    .B(_01693_),
    .Y(_01694_));
 AOI211x1_ASAP7_75t_R _31274_ (.A1(net1640),
    .A2(net1898),
    .B(_01685_),
    .C(_01644_),
    .Y(_01695_));
 INVx4_ASAP7_75t_R _31275_ (.A(_01685_),
    .Y(_01696_));
 OA21x2_ASAP7_75t_R _31276_ (.A1(_01562_),
    .A2(_01516_),
    .B(_01696_),
    .Y(_01697_));
 NOR2x1_ASAP7_75t_R _31277_ (.A(_01695_),
    .B(_01697_),
    .Y(_01698_));
 NAND2x2_ASAP7_75t_R _31278_ (.A(_01606_),
    .B(_01599_),
    .Y(_01699_));
 TAPCELL_ASAP7_75t_R TAP_641 ();
 NAND2x2_ASAP7_75t_R _31280_ (.A(_01530_),
    .B(_01667_),
    .Y(_01701_));
 TAPCELL_ASAP7_75t_R TAP_640 ();
 AO31x2_ASAP7_75t_R _31282_ (.A1(_01540_),
    .A2(_01691_),
    .A3(_01699_),
    .B(_01701_),
    .Y(_01703_));
 NAND3x1_ASAP7_75t_R _31283_ (.A(_01694_),
    .B(_01698_),
    .C(_01703_),
    .Y(_01704_));
 NOR2x1_ASAP7_75t_R _31284_ (.A(_01684_),
    .B(_01704_),
    .Y(_01705_));
 NOR2x2_ASAP7_75t_R _31285_ (.A(net2777),
    .B(_00634_),
    .Y(_01706_));
 NAND2x2_ASAP7_75t_R _31286_ (.A(_01706_),
    .B(_01530_),
    .Y(_01707_));
 TAPCELL_ASAP7_75t_R TAP_639 ();
 AO21x1_ASAP7_75t_R _31288_ (.A1(net2366),
    .A2(_01691_),
    .B(net3256),
    .Y(_01709_));
 AO21x1_ASAP7_75t_R _31289_ (.A1(net1104),
    .A2(net1457),
    .B(_01707_),
    .Y(_01710_));
 INVx5_ASAP7_75t_R _31290_ (.A(_01707_),
    .Y(_01711_));
 NAND2x1_ASAP7_75t_R _31291_ (.A(_01589_),
    .B(_01711_),
    .Y(_01712_));
 AND3x1_ASAP7_75t_R _31292_ (.A(_01709_),
    .B(_01710_),
    .C(_01712_),
    .Y(_01713_));
 TAPCELL_ASAP7_75t_R TAP_638 ();
 NAND2x2_ASAP7_75t_R _31294_ (.A(_01706_),
    .B(_01570_),
    .Y(_01715_));
 TAPCELL_ASAP7_75t_R TAP_637 ();
 AOI211x1_ASAP7_75t_R _31296_ (.A1(_01498_),
    .A2(_01494_),
    .B(_01715_),
    .C(_01644_),
    .Y(_01717_));
 INVx1_ASAP7_75t_R _31297_ (.A(_01717_),
    .Y(_01718_));
 NOR2x2_ASAP7_75t_R _31298_ (.A(net1241),
    .B(_01499_),
    .Y(_01719_));
 INVx2_ASAP7_75t_R _31299_ (.A(_01715_),
    .Y(_01720_));
 NAND2x1_ASAP7_75t_R _31300_ (.A(_01719_),
    .B(_01720_),
    .Y(_01721_));
 TAPCELL_ASAP7_75t_R TAP_636 ();
 AO21x1_ASAP7_75t_R _31302_ (.A1(net2524),
    .A2(net1597),
    .B(_01715_),
    .Y(_01723_));
 AND3x1_ASAP7_75t_R _31303_ (.A(_01718_),
    .B(_01721_),
    .C(_01723_),
    .Y(_01724_));
 NAND2x1_ASAP7_75t_R _31304_ (.A(_01713_),
    .B(_01724_),
    .Y(_01725_));
 TAPCELL_ASAP7_75t_R TAP_635 ();
 AO21x2_ASAP7_75t_R _31306_ (.A1(_01561_),
    .A2(net1025),
    .B(net1241),
    .Y(_01727_));
 NAND2x2_ASAP7_75t_R _31307_ (.A(_01706_),
    .B(_01585_),
    .Y(_01728_));
 TAPCELL_ASAP7_75t_R TAP_634 ();
 AOI21x1_ASAP7_75t_R _31309_ (.A1(_01674_),
    .A2(_01727_),
    .B(net3175),
    .Y(_01730_));
 AOI211x1_ASAP7_75t_R _31310_ (.A1(net1640),
    .A2(_01494_),
    .B(_01728_),
    .C(net2071),
    .Y(_01731_));
 NAND2x2_ASAP7_75t_R _31311_ (.A(_01494_),
    .B(net1576),
    .Y(_01732_));
 NOR2x1_ASAP7_75t_R _31312_ (.A(_01732_),
    .B(net3175),
    .Y(_01733_));
 NOR3x1_ASAP7_75t_R _31313_ (.A(_01730_),
    .B(_01731_),
    .C(_01733_),
    .Y(_01734_));
 NAND2x2_ASAP7_75t_R _31314_ (.A(_01602_),
    .B(_01706_),
    .Y(_01735_));
 AO21x1_ASAP7_75t_R _31315_ (.A1(_01691_),
    .A2(_01600_),
    .B(_01735_),
    .Y(_01736_));
 INVx4_ASAP7_75t_R _31316_ (.A(_01735_),
    .Y(_01737_));
 NAND2x2_ASAP7_75t_R _31317_ (.A(_01526_),
    .B(_01737_),
    .Y(_01738_));
 NOR2x1_ASAP7_75t_R _31318_ (.A(_01735_),
    .B(net2572),
    .Y(_01739_));
 INVx1_ASAP7_75t_R _31319_ (.A(_01739_),
    .Y(_01740_));
 NAND3x1_ASAP7_75t_R _31320_ (.A(_01736_),
    .B(_01738_),
    .C(_01740_),
    .Y(_01741_));
 TAPCELL_ASAP7_75t_R TAP_633 ();
 TAPCELL_ASAP7_75t_R TAP_632 ();
 AO21x1_ASAP7_75t_R _31323_ (.A1(net2524),
    .A2(net3261),
    .B(_01735_),
    .Y(_01744_));
 NOR2x1_ASAP7_75t_R _31324_ (.A(_01735_),
    .B(net2728),
    .Y(_01745_));
 INVx1_ASAP7_75t_R _31325_ (.A(_01745_),
    .Y(_01746_));
 NAND2x2_ASAP7_75t_R _31326_ (.A(_01511_),
    .B(_01737_),
    .Y(_01747_));
 NAND3x1_ASAP7_75t_R _31327_ (.A(_01744_),
    .B(_01746_),
    .C(_01747_),
    .Y(_01748_));
 NOR2x1_ASAP7_75t_R _31328_ (.A(_01741_),
    .B(_01748_),
    .Y(_01749_));
 NAND2x1_ASAP7_75t_R _31329_ (.A(_01734_),
    .B(_01749_),
    .Y(_01750_));
 NOR2x1_ASAP7_75t_R _31330_ (.A(_01725_),
    .B(_01750_),
    .Y(_01751_));
 NAND2x1_ASAP7_75t_R _31331_ (.A(_01705_),
    .B(_01751_),
    .Y(_01752_));
 NOR2x2_ASAP7_75t_R _31332_ (.A(_01665_),
    .B(_01752_),
    .Y(_01753_));
 NAND2x2_ASAP7_75t_R _31333_ (.A(_01539_),
    .B(_01753_),
    .Y(_01754_));
 TAPCELL_ASAP7_75t_R TAP_631 ();
 INVx2_ASAP7_75t_R _31335_ (.A(_00596_),
    .Y(_01756_));
 NOR2x2_ASAP7_75t_R _31336_ (.A(net3273),
    .B(_01756_),
    .Y(_01757_));
 TAPCELL_ASAP7_75t_R TAP_630 ();
 INVx4_ASAP7_75t_R _31338_ (.A(_00594_),
    .Y(_01759_));
 NOR2x2_ASAP7_75t_R _31339_ (.A(net3262),
    .B(_01759_),
    .Y(_01760_));
 NAND2x2_ASAP7_75t_R _31340_ (.A(_01757_),
    .B(_01760_),
    .Y(_01761_));
 INVx6_ASAP7_75t_R _31341_ (.A(_01761_),
    .Y(_01762_));
 TAPCELL_ASAP7_75t_R TAP_629 ();
 TAPCELL_ASAP7_75t_R TAP_628 ();
 NAND2x2_ASAP7_75t_R _31344_ (.A(net1363),
    .B(net1454),
    .Y(_01765_));
 TAPCELL_ASAP7_75t_R TAP_627 ();
 TAPCELL_ASAP7_75t_R TAP_626 ();
 NAND2x2_ASAP7_75t_R _31347_ (.A(net2486),
    .B(_00598_),
    .Y(_01768_));
 NOR2x2_ASAP7_75t_R _31348_ (.A(_01765_),
    .B(net1299),
    .Y(_01769_));
 CKINVDCx20_ASAP7_75t_R _31349_ (.A(net1358),
    .Y(_01770_));
 TAPCELL_ASAP7_75t_R TAP_625 ();
 INVx2_ASAP7_75t_R _31351_ (.A(_00598_),
    .Y(_01772_));
 NOR2x2_ASAP7_75t_R _31352_ (.A(net2487),
    .B(_01772_),
    .Y(_01773_));
 NAND2x2_ASAP7_75t_R _31353_ (.A(_01770_),
    .B(net1459),
    .Y(_01774_));
 NOR2x2_ASAP7_75t_R _31354_ (.A(net2486),
    .B(_00598_),
    .Y(_01775_));
 CKINVDCx16_ASAP7_75t_R _31355_ (.A(net1447),
    .Y(_01776_));
 NOR2x2_ASAP7_75t_R _31356_ (.A(net1358),
    .B(_01776_),
    .Y(_01777_));
 NAND2x2_ASAP7_75t_R _31357_ (.A(net1126),
    .B(_01777_),
    .Y(_01778_));
 TAPCELL_ASAP7_75t_R TAP_624 ();
 NOR2x2_ASAP7_75t_R _31359_ (.A(_00595_),
    .B(_00596_),
    .Y(_01780_));
 NAND2x2_ASAP7_75t_R _31360_ (.A(_01780_),
    .B(_01760_),
    .Y(_01781_));
 AO21x1_ASAP7_75t_R _31361_ (.A1(_01774_),
    .A2(net3275),
    .B(_01781_),
    .Y(_01782_));
 TAPCELL_ASAP7_75t_R TAP_623 ();
 NOR2x2_ASAP7_75t_R _31363_ (.A(_01770_),
    .B(net1299),
    .Y(_01784_));
 INVx3_ASAP7_75t_R _31364_ (.A(_01784_),
    .Y(_01785_));
 NAND2x2_ASAP7_75t_R _31365_ (.A(net1448),
    .B(_01770_),
    .Y(_01786_));
 INVx4_ASAP7_75t_R _31366_ (.A(net2486),
    .Y(_01787_));
 NOR2x2_ASAP7_75t_R _31367_ (.A(net3133),
    .B(_01787_),
    .Y(_01788_));
 TAPCELL_ASAP7_75t_R TAP_622 ();
 NAND2x2_ASAP7_75t_R _31369_ (.A(net3258),
    .B(net1557),
    .Y(_01790_));
 AO21x1_ASAP7_75t_R _31370_ (.A1(_01785_),
    .A2(_01790_),
    .B(_01781_),
    .Y(_01791_));
 NAND2x1_ASAP7_75t_R _31371_ (.A(_01782_),
    .B(_01791_),
    .Y(_01792_));
 TAPCELL_ASAP7_75t_R TAP_621 ();
 TAPCELL_ASAP7_75t_R TAP_620 ();
 NAND2x2_ASAP7_75t_R _31374_ (.A(net1359),
    .B(net1133),
    .Y(_01795_));
 AO21x1_ASAP7_75t_R _31375_ (.A1(net3275),
    .A2(_01795_),
    .B(_01761_),
    .Y(_01796_));
 NAND2x2_ASAP7_75t_R _31376_ (.A(_01773_),
    .B(_01777_),
    .Y(_01797_));
 TAPCELL_ASAP7_75t_R TAP_619 ();
 NAND2x2_ASAP7_75t_R _31378_ (.A(net1364),
    .B(net1463),
    .Y(_01799_));
 TAPCELL_ASAP7_75t_R TAP_618 ();
 AO21x1_ASAP7_75t_R _31380_ (.A1(net2239),
    .A2(_01799_),
    .B(_01761_),
    .Y(_01801_));
 NAND2x1_ASAP7_75t_R _31381_ (.A(_01796_),
    .B(_01801_),
    .Y(_01802_));
 AOI211x1_ASAP7_75t_R _31382_ (.A1(_01762_),
    .A2(net3272),
    .B(_01792_),
    .C(_01802_),
    .Y(_01803_));
 NOR2x2_ASAP7_75t_R _31383_ (.A(net1363),
    .B(net1447),
    .Y(_01804_));
 INVx3_ASAP7_75t_R _31384_ (.A(_01804_),
    .Y(_01805_));
 NOR2x2_ASAP7_75t_R _31385_ (.A(net1299),
    .B(_01805_),
    .Y(_01806_));
 NAND2x2_ASAP7_75t_R _31386_ (.A(_00595_),
    .B(_00596_),
    .Y(_01807_));
 INVx3_ASAP7_75t_R _31387_ (.A(_01807_),
    .Y(_01808_));
 NAND2x2_ASAP7_75t_R _31388_ (.A(_01760_),
    .B(_01808_),
    .Y(_01809_));
 CKINVDCx5p33_ASAP7_75t_R _31389_ (.A(_01809_),
    .Y(_01810_));
 TAPCELL_ASAP7_75t_R TAP_617 ();
 OA21x2_ASAP7_75t_R _31391_ (.A1(_01806_),
    .A2(net3271),
    .B(_01810_),
    .Y(_01812_));
 INVx1_ASAP7_75t_R _31392_ (.A(_01812_),
    .Y(_01813_));
 NOR2x2_ASAP7_75t_R _31393_ (.A(net1454),
    .B(_01770_),
    .Y(_01814_));
 NAND2x2_ASAP7_75t_R _31394_ (.A(_01814_),
    .B(net1556),
    .Y(_01815_));
 INVx4_ASAP7_75t_R _31395_ (.A(net3132),
    .Y(_01816_));
 NAND2x1_ASAP7_75t_R _31396_ (.A(_01810_),
    .B(_01816_),
    .Y(_01817_));
 INVx3_ASAP7_75t_R _31397_ (.A(_01765_),
    .Y(_01818_));
 NAND2x2_ASAP7_75t_R _31398_ (.A(net2299),
    .B(_01818_),
    .Y(_01819_));
 TAPCELL_ASAP7_75t_R TAP_616 ();
 NAND2x2_ASAP7_75t_R _31400_ (.A(_01814_),
    .B(net2299),
    .Y(_01821_));
 AO21x1_ASAP7_75t_R _31401_ (.A1(_01819_),
    .A2(_01821_),
    .B(_01809_),
    .Y(_01822_));
 NAND3x1_ASAP7_75t_R _31402_ (.A(_01813_),
    .B(_01817_),
    .C(_01822_),
    .Y(_01823_));
 NAND2x2_ASAP7_75t_R _31403_ (.A(_01777_),
    .B(net1553),
    .Y(_01824_));
 NAND2x2_ASAP7_75t_R _31404_ (.A(_01804_),
    .B(net1556),
    .Y(_01825_));
 INVx2_ASAP7_75t_R _31405_ (.A(_00595_),
    .Y(_01826_));
 NOR2x2_ASAP7_75t_R _31406_ (.A(_00596_),
    .B(_01826_),
    .Y(_01827_));
 NAND2x2_ASAP7_75t_R _31407_ (.A(_01760_),
    .B(_01827_),
    .Y(_01828_));
 AO21x1_ASAP7_75t_R _31408_ (.A1(_01824_),
    .A2(net1244),
    .B(_01828_),
    .Y(_01829_));
 CKINVDCx9p33_ASAP7_75t_R _31409_ (.A(_01768_),
    .Y(_01830_));
 NAND2x2_ASAP7_75t_R _31410_ (.A(_01814_),
    .B(_01830_),
    .Y(_01831_));
 NAND2x2_ASAP7_75t_R _31411_ (.A(_01804_),
    .B(_01830_),
    .Y(_01832_));
 AO21x1_ASAP7_75t_R _31412_ (.A1(_01831_),
    .A2(_01832_),
    .B(_01828_),
    .Y(_01833_));
 AND2x2_ASAP7_75t_R _31413_ (.A(_01829_),
    .B(_01833_),
    .Y(_01834_));
 AO21x2_ASAP7_75t_R _31414_ (.A1(net2707),
    .A2(_01821_),
    .B(_01828_),
    .Y(_01835_));
 NAND2x2_ASAP7_75t_R _31415_ (.A(net1130),
    .B(_01818_),
    .Y(_01836_));
 NAND2x2_ASAP7_75t_R _31416_ (.A(_01804_),
    .B(net1127),
    .Y(_01837_));
 AO21x1_ASAP7_75t_R _31417_ (.A1(_01836_),
    .A2(_01837_),
    .B(_01828_),
    .Y(_01838_));
 AND2x2_ASAP7_75t_R _31418_ (.A(_01835_),
    .B(_01838_),
    .Y(_01839_));
 NAND2x1_ASAP7_75t_R _31419_ (.A(_01834_),
    .B(_01839_),
    .Y(_01840_));
 NOR2x1_ASAP7_75t_R _31420_ (.A(_01823_),
    .B(_01840_),
    .Y(_01841_));
 NAND2x1_ASAP7_75t_R _31421_ (.A(_01803_),
    .B(_01841_),
    .Y(_01842_));
 NOR2x2_ASAP7_75t_R _31422_ (.A(net1299),
    .B(_01786_),
    .Y(_01843_));
 NAND2x2_ASAP7_75t_R _31423_ (.A(_00596_),
    .B(_01826_),
    .Y(_01844_));
 NOR2x2_ASAP7_75t_R _31424_ (.A(net3262),
    .B(_00594_),
    .Y(_01845_));
 INVx3_ASAP7_75t_R _31425_ (.A(_01845_),
    .Y(_01846_));
 NOR2x2_ASAP7_75t_R _31426_ (.A(_01844_),
    .B(_01846_),
    .Y(_01847_));
 OA21x2_ASAP7_75t_R _31427_ (.A1(_01843_),
    .A2(_01784_),
    .B(_01847_),
    .Y(_01848_));
 TAPCELL_ASAP7_75t_R TAP_615 ();
 NAND2x2_ASAP7_75t_R _31429_ (.A(net2486),
    .B(_01772_),
    .Y(_01850_));
 NAND2x2_ASAP7_75t_R _31430_ (.A(_01845_),
    .B(_01757_),
    .Y(_01851_));
 AOI211x1_ASAP7_75t_R _31431_ (.A1(net1361),
    .A2(net1451),
    .B(_01850_),
    .C(_01851_),
    .Y(_01852_));
 NOR2x1_ASAP7_75t_R _31432_ (.A(_01848_),
    .B(_01852_),
    .Y(_01853_));
 AOI21x1_ASAP7_75t_R _31433_ (.A1(_01774_),
    .A2(_01819_),
    .B(_01851_),
    .Y(_01854_));
 INVx3_ASAP7_75t_R _31434_ (.A(_01837_),
    .Y(_01855_));
 TAPCELL_ASAP7_75t_R TAP_614 ();
 CKINVDCx14_ASAP7_75t_R _31436_ (.A(net1127),
    .Y(_01857_));
 NOR2x2_ASAP7_75t_R _31437_ (.A(net950),
    .B(_01857_),
    .Y(_01858_));
 OA21x2_ASAP7_75t_R _31438_ (.A1(_01855_),
    .A2(_01858_),
    .B(_01847_),
    .Y(_01859_));
 NOR2x1_ASAP7_75t_R _31439_ (.A(_01854_),
    .B(_01859_),
    .Y(_01860_));
 NAND2x1_ASAP7_75t_R _31440_ (.A(_01853_),
    .B(_01860_),
    .Y(_01861_));
 NOR2x2_ASAP7_75t_R _31441_ (.A(_01770_),
    .B(_01850_),
    .Y(_01862_));
 NAND2x2_ASAP7_75t_R _31442_ (.A(_01845_),
    .B(_01780_),
    .Y(_01863_));
 INVx3_ASAP7_75t_R _31443_ (.A(_01863_),
    .Y(_01864_));
 TAPCELL_ASAP7_75t_R TAP_613 ();
 AOI211x1_ASAP7_75t_R _31445_ (.A1(_01770_),
    .A2(_01776_),
    .B(_01863_),
    .C(net1300),
    .Y(_01866_));
 AOI21x1_ASAP7_75t_R _31446_ (.A1(_01862_),
    .A2(_01864_),
    .B(_01866_),
    .Y(_01867_));
 AO21x1_ASAP7_75t_R _31447_ (.A1(_01836_),
    .A2(net3275),
    .B(_01863_),
    .Y(_01868_));
 NAND2x2_ASAP7_75t_R _31448_ (.A(net1359),
    .B(_01776_),
    .Y(_01869_));
 NAND2x2_ASAP7_75t_R _31449_ (.A(net3133),
    .B(_01787_),
    .Y(_01870_));
 NOR2x2_ASAP7_75t_R _31450_ (.A(_01869_),
    .B(_01870_),
    .Y(_01871_));
 NAND2x1_ASAP7_75t_R _31451_ (.A(_01871_),
    .B(_01864_),
    .Y(_01872_));
 AND2x2_ASAP7_75t_R _31452_ (.A(_01868_),
    .B(_01872_),
    .Y(_01873_));
 NAND2x1_ASAP7_75t_R _31453_ (.A(_01867_),
    .B(_01873_),
    .Y(_01874_));
 NOR2x1_ASAP7_75t_R _31454_ (.A(_01861_),
    .B(_01874_),
    .Y(_01875_));
 NOR2x2_ASAP7_75t_R _31455_ (.A(net2685),
    .B(_01846_),
    .Y(_01876_));
 NAND2x2_ASAP7_75t_R _31456_ (.A(_01776_),
    .B(net1556),
    .Y(_01877_));
 NAND2x2_ASAP7_75t_R _31457_ (.A(_01845_),
    .B(_01808_),
    .Y(_01878_));
 AOI21x1_ASAP7_75t_R _31458_ (.A1(_01877_),
    .A2(_01824_),
    .B(_01878_),
    .Y(_01879_));
 AOI21x1_ASAP7_75t_R _31459_ (.A1(_01769_),
    .A2(_01876_),
    .B(_01879_),
    .Y(_01880_));
 TAPCELL_ASAP7_75t_R TAP_612 ();
 NOR2x2_ASAP7_75t_R _31461_ (.A(_01770_),
    .B(_01870_),
    .Y(_01882_));
 AOI211x1_ASAP7_75t_R _31462_ (.A1(net1362),
    .A2(net1451),
    .B(_01878_),
    .C(_01857_),
    .Y(_01883_));
 AOI21x1_ASAP7_75t_R _31463_ (.A1(_01882_),
    .A2(_01876_),
    .B(_01883_),
    .Y(_01884_));
 NAND2x1_ASAP7_75t_R _31464_ (.A(_01880_),
    .B(_01884_),
    .Y(_01885_));
 INVx3_ASAP7_75t_R _31465_ (.A(_01795_),
    .Y(_01886_));
 NAND2x2_ASAP7_75t_R _31466_ (.A(net3273),
    .B(_01756_),
    .Y(_01887_));
 NOR2x2_ASAP7_75t_R _31467_ (.A(_01887_),
    .B(_01846_),
    .Y(_01888_));
 OA21x2_ASAP7_75t_R _31468_ (.A1(_01855_),
    .A2(_01886_),
    .B(_01888_),
    .Y(_01889_));
 NOR2x2_ASAP7_75t_R _31469_ (.A(_01786_),
    .B(_01850_),
    .Y(_01890_));
 OA21x2_ASAP7_75t_R _31470_ (.A1(_01890_),
    .A2(_01843_),
    .B(_01888_),
    .Y(_01891_));
 NAND2x2_ASAP7_75t_R _31471_ (.A(_01804_),
    .B(net2299),
    .Y(_01892_));
 TAPCELL_ASAP7_75t_R TAP_611 ();
 NAND2x2_ASAP7_75t_R _31473_ (.A(_01845_),
    .B(_01827_),
    .Y(_01894_));
 TAPCELL_ASAP7_75t_R TAP_610 ();
 NOR2x1_ASAP7_75t_R _31475_ (.A(net3168),
    .B(_01894_),
    .Y(_01896_));
 OR3x1_ASAP7_75t_R _31476_ (.A(_01889_),
    .B(_01891_),
    .C(_01896_),
    .Y(_01897_));
 NOR2x1_ASAP7_75t_R _31477_ (.A(_01885_),
    .B(_01897_),
    .Y(_01898_));
 NAND2x1_ASAP7_75t_R _31478_ (.A(_01875_),
    .B(_01898_),
    .Y(_01899_));
 NOR2x1_ASAP7_75t_R _31479_ (.A(_01842_),
    .B(_01899_),
    .Y(_01900_));
 TAPCELL_ASAP7_75t_R TAP_609 ();
 TAPCELL_ASAP7_75t_R TAP_608 ();
 NAND2x2_ASAP7_75t_R _31482_ (.A(net3262),
    .B(_01759_),
    .Y(_01903_));
 NOR2x2_ASAP7_75t_R _31483_ (.A(_01807_),
    .B(_01903_),
    .Y(_01904_));
 CKINVDCx5p33_ASAP7_75t_R _31484_ (.A(_01904_),
    .Y(_01905_));
 TAPCELL_ASAP7_75t_R TAP_607 ();
 AO21x1_ASAP7_75t_R _31486_ (.A1(_01831_),
    .A2(net1458),
    .B(_01905_),
    .Y(_01907_));
 NAND2x2_ASAP7_75t_R _31487_ (.A(net1132),
    .B(_01814_),
    .Y(_01908_));
 AO21x1_ASAP7_75t_R _31488_ (.A1(_01908_),
    .A2(_01837_),
    .B(_01905_),
    .Y(_01909_));
 TAPCELL_ASAP7_75t_R TAP_606 ();
 INVx2_ASAP7_75t_R _31490_ (.A(_01774_),
    .Y(_01911_));
 NAND2x1_ASAP7_75t_R _31491_ (.A(_01904_),
    .B(_01911_),
    .Y(_01912_));
 NAND3x1_ASAP7_75t_R _31492_ (.A(_01907_),
    .B(_01909_),
    .C(_01912_),
    .Y(_01913_));
 INVx3_ASAP7_75t_R _31493_ (.A(net3262),
    .Y(_01914_));
 NOR2x2_ASAP7_75t_R _31494_ (.A(_00594_),
    .B(_01914_),
    .Y(_01915_));
 NAND2x2_ASAP7_75t_R _31495_ (.A(_01915_),
    .B(_01827_),
    .Y(_01916_));
 TAPCELL_ASAP7_75t_R TAP_605 ();
 NOR2x1_ASAP7_75t_R _31497_ (.A(_01837_),
    .B(_01916_),
    .Y(_01918_));
 AOI21x1_ASAP7_75t_R _31498_ (.A1(net2709),
    .A2(_01821_),
    .B(_01916_),
    .Y(_01919_));
 NOR2x1_ASAP7_75t_R _31499_ (.A(_01918_),
    .B(_01919_),
    .Y(_01920_));
 AO21x1_ASAP7_75t_R _31500_ (.A1(_01831_),
    .A2(_01832_),
    .B(_01916_),
    .Y(_01921_));
 TAPCELL_ASAP7_75t_R TAP_604 ();
 AO21x1_ASAP7_75t_R _31502_ (.A1(net3332),
    .A2(_01824_),
    .B(_01916_),
    .Y(_01923_));
 NAND3x1_ASAP7_75t_R _31503_ (.A(_01920_),
    .B(_01921_),
    .C(_01923_),
    .Y(_01924_));
 NOR2x1_ASAP7_75t_R _31504_ (.A(_01913_),
    .B(_01924_),
    .Y(_01925_));
 NAND2x2_ASAP7_75t_R _31505_ (.A(_01757_),
    .B(_01915_),
    .Y(_01926_));
 AO21x1_ASAP7_75t_R _31506_ (.A1(net3275),
    .A2(net2371),
    .B(net2215),
    .Y(_01927_));
 TAPCELL_ASAP7_75t_R TAP_603 ();
 AO21x1_ASAP7_75t_R _31508_ (.A1(net1458),
    .A2(net1299),
    .B(net2215),
    .Y(_01929_));
 NOR2x2_ASAP7_75t_R _31509_ (.A(_01844_),
    .B(_01903_),
    .Y(_01930_));
 NAND2x1_ASAP7_75t_R _31510_ (.A(_01871_),
    .B(_01930_),
    .Y(_01931_));
 NAND3x1_ASAP7_75t_R _31511_ (.A(_01927_),
    .B(_01929_),
    .C(_01931_),
    .Y(_01932_));
 TAPCELL_ASAP7_75t_R TAP_602 ();
 NAND2x2_ASAP7_75t_R _31513_ (.A(net1361),
    .B(net1558),
    .Y(_01934_));
 NAND2x2_ASAP7_75t_R _31514_ (.A(_01776_),
    .B(_01830_),
    .Y(_01935_));
 NAND2x2_ASAP7_75t_R _31515_ (.A(_01780_),
    .B(_01915_),
    .Y(_01936_));
 AO31x2_ASAP7_75t_R _31516_ (.A1(net1245),
    .A2(_01934_),
    .A3(_01935_),
    .B(_01936_),
    .Y(_01937_));
 NAND2x2_ASAP7_75t_R _31517_ (.A(net954),
    .B(net1127),
    .Y(_01938_));
 AO21x1_ASAP7_75t_R _31518_ (.A1(net2707),
    .A2(_01938_),
    .B(_01936_),
    .Y(_01939_));
 INVx3_ASAP7_75t_R _31519_ (.A(_01936_),
    .Y(_01940_));
 NAND2x1_ASAP7_75t_R _31520_ (.A(_01882_),
    .B(_01940_),
    .Y(_01941_));
 AND2x2_ASAP7_75t_R _31521_ (.A(_01939_),
    .B(_01941_),
    .Y(_01942_));
 NAND2x1_ASAP7_75t_R _31522_ (.A(_01937_),
    .B(_01942_),
    .Y(_01943_));
 NOR2x1_ASAP7_75t_R _31523_ (.A(_01932_),
    .B(_01943_),
    .Y(_01944_));
 NAND2x2_ASAP7_75t_R _31524_ (.A(_01925_),
    .B(_01944_),
    .Y(_01945_));
 NAND2x2_ASAP7_75t_R _31525_ (.A(_01777_),
    .B(_01830_),
    .Y(_01946_));
 NAND2x2_ASAP7_75t_R _31526_ (.A(net3262),
    .B(_00594_),
    .Y(_01947_));
 INVx4_ASAP7_75t_R _31527_ (.A(_01947_),
    .Y(_01948_));
 NAND2x2_ASAP7_75t_R _31528_ (.A(_01757_),
    .B(_01948_),
    .Y(_01949_));
 AO21x2_ASAP7_75t_R _31529_ (.A1(_01946_),
    .A2(_01785_),
    .B(_01949_),
    .Y(_01950_));
 AO21x1_ASAP7_75t_R _31530_ (.A1(_01824_),
    .A2(net1458),
    .B(_01949_),
    .Y(_01951_));
 NAND2x2_ASAP7_75t_R _31531_ (.A(_01765_),
    .B(net1462),
    .Y(_01952_));
 AO21x1_ASAP7_75t_R _31532_ (.A1(_01908_),
    .A2(_01952_),
    .B(net3125),
    .Y(_01953_));
 NAND3x1_ASAP7_75t_R _31533_ (.A(_01950_),
    .B(_01951_),
    .C(_01953_),
    .Y(_01954_));
 NAND2x2_ASAP7_75t_R _31534_ (.A(_01780_),
    .B(_01948_),
    .Y(_01955_));
 TAPCELL_ASAP7_75t_R TAP_601 ();
 NOR2x1_ASAP7_75t_R _31536_ (.A(_01955_),
    .B(_01935_),
    .Y(_01957_));
 AOI21x1_ASAP7_75t_R _31537_ (.A1(_01825_),
    .A2(net3131),
    .B(_01955_),
    .Y(_01958_));
 NOR2x1_ASAP7_75t_R _31538_ (.A(_01957_),
    .B(_01958_),
    .Y(_01959_));
 AO21x1_ASAP7_75t_R _31539_ (.A1(net2239),
    .A2(net3168),
    .B(_01955_),
    .Y(_01960_));
 TAPCELL_ASAP7_75t_R TAP_600 ();
 AO21x1_ASAP7_75t_R _31541_ (.A1(net2307),
    .A2(net3275),
    .B(_01955_),
    .Y(_01962_));
 NAND3x1_ASAP7_75t_R _31542_ (.A(_01959_),
    .B(_01960_),
    .C(_01962_),
    .Y(_01963_));
 NOR2x1_ASAP7_75t_R _31543_ (.A(_01954_),
    .B(_01963_),
    .Y(_01964_));
 NAND2x2_ASAP7_75t_R _31544_ (.A(net1556),
    .B(_01818_),
    .Y(_01965_));
 TAPCELL_ASAP7_75t_R TAP_599 ();
 NAND2x2_ASAP7_75t_R _31546_ (.A(_01808_),
    .B(_01948_),
    .Y(_01967_));
 TAPCELL_ASAP7_75t_R TAP_598 ();
 AO21x1_ASAP7_75t_R _31548_ (.A1(_01965_),
    .A2(net1458),
    .B(_01967_),
    .Y(_01969_));
 NOR2x2_ASAP7_75t_R _31549_ (.A(net2684),
    .B(_01947_),
    .Y(_01970_));
 OA211x2_ASAP7_75t_R _31550_ (.A1(net1359),
    .A2(net1449),
    .B(_01970_),
    .C(net1128),
    .Y(_01971_));
 INVx1_ASAP7_75t_R _31551_ (.A(_01971_),
    .Y(_01972_));
 NAND2x1_ASAP7_75t_R _31552_ (.A(_01969_),
    .B(_01972_),
    .Y(_01973_));
 NOR2x2_ASAP7_75t_R _31553_ (.A(_01947_),
    .B(_01887_),
    .Y(_01974_));
 TAPCELL_ASAP7_75t_R TAP_597 ();
 NAND2x2_ASAP7_75t_R _31555_ (.A(_01825_),
    .B(net3253),
    .Y(_01976_));
 NAND2x2_ASAP7_75t_R _31556_ (.A(_01827_),
    .B(_01948_),
    .Y(_01977_));
 AOI211x1_ASAP7_75t_R _31557_ (.A1(_01770_),
    .A2(_01776_),
    .B(_01977_),
    .C(net1301),
    .Y(_01978_));
 AOI21x1_ASAP7_75t_R _31558_ (.A1(_01974_),
    .A2(_01976_),
    .B(_01978_),
    .Y(_01979_));
 TAPCELL_ASAP7_75t_R TAP_596 ();
 AO21x1_ASAP7_75t_R _31560_ (.A1(_01795_),
    .A2(net2369),
    .B(_01977_),
    .Y(_01981_));
 OA21x2_ASAP7_75t_R _31561_ (.A1(_01870_),
    .A2(_01977_),
    .B(_01981_),
    .Y(_01982_));
 NAND2x1_ASAP7_75t_R _31562_ (.A(_01979_),
    .B(_01982_),
    .Y(_01983_));
 NOR2x1_ASAP7_75t_R _31563_ (.A(_01973_),
    .B(_01983_),
    .Y(_01984_));
 NAND2x1_ASAP7_75t_R _31564_ (.A(_01964_),
    .B(_01984_),
    .Y(_01985_));
 NOR2x2_ASAP7_75t_R _31565_ (.A(_01945_),
    .B(_01985_),
    .Y(_01986_));
 NAND2x2_ASAP7_75t_R _31566_ (.A(_01900_),
    .B(_01986_),
    .Y(_01987_));
 TAPCELL_ASAP7_75t_R TAP_595 ();
 XOR2x1_ASAP7_75t_R _31568_ (.A(_01754_),
    .Y(_01989_),
    .B(net2710));
 AOI21x1_ASAP7_75t_R _31569_ (.A1(_01484_),
    .A2(_01487_),
    .B(_01989_),
    .Y(_01990_));
 INVx2_ASAP7_75t_R _31570_ (.A(_01094_),
    .Y(_01991_));
 NAND2x1_ASAP7_75t_R _31571_ (.A(_01991_),
    .B(_01483_),
    .Y(_01992_));
 AO21x1_ASAP7_75t_R _31572_ (.A1(_01485_),
    .A2(_01486_),
    .B(_01991_),
    .Y(_01993_));
 INVx1_ASAP7_75t_R _31573_ (.A(_01989_),
    .Y(_01994_));
 AOI21x1_ASAP7_75t_R _31574_ (.A1(_01992_),
    .A2(_01993_),
    .B(_01994_),
    .Y(_01995_));
 OAI21x1_ASAP7_75t_R _31575_ (.A1(_01990_),
    .A2(_01995_),
    .B(net395),
    .Y(_01996_));
 NAND2x2_ASAP7_75t_R _31576_ (.A(_01996_),
    .B(_21864_),
    .Y(_01997_));
 XOR2x1_ASAP7_75t_R _31577_ (.A(_01997_),
    .Y(_00113_),
    .B(_00484_));
 AND2x2_ASAP7_75t_R _31578_ (.A(_18753_),
    .B(_00882_),
    .Y(_01998_));
 AO31x2_ASAP7_75t_R _31579_ (.A1(net1122),
    .A2(net1119),
    .A3(net2723),
    .B(net3144),
    .Y(_01999_));
 AOI211x1_ASAP7_75t_R _31580_ (.A1(net1341),
    .A2(net1277),
    .B(net1919),
    .C(net3144),
    .Y(_02000_));
 INVx1_ASAP7_75t_R _31581_ (.A(_02000_),
    .Y(_02001_));
 NAND2x1_ASAP7_75t_R _31582_ (.A(_01374_),
    .B(_01197_),
    .Y(_02002_));
 NAND3x1_ASAP7_75t_R _31583_ (.A(_01999_),
    .B(_02001_),
    .C(_02002_),
    .Y(_02003_));
 AO21x1_ASAP7_75t_R _31584_ (.A1(_01113_),
    .A2(_01226_),
    .B(net3154),
    .Y(_02004_));
 AO21x1_ASAP7_75t_R _31585_ (.A1(net1266),
    .A2(net2731),
    .B(net3154),
    .Y(_02005_));
 AND2x2_ASAP7_75t_R _31586_ (.A(_02004_),
    .B(_02005_),
    .Y(_02006_));
 AOI211x1_ASAP7_75t_R _31587_ (.A1(net1341),
    .A2(_01096_),
    .B(net3154),
    .C(_01204_),
    .Y(_02007_));
 AOI21x1_ASAP7_75t_R _31588_ (.A1(_01210_),
    .A2(_01327_),
    .B(_02007_),
    .Y(_02008_));
 NAND2x1_ASAP7_75t_R _31589_ (.A(_02006_),
    .B(_02008_),
    .Y(_02009_));
 NOR2x1_ASAP7_75t_R _31590_ (.A(_02003_),
    .B(_02009_),
    .Y(_02010_));
 TAPCELL_ASAP7_75t_R TAP_594 ();
 AO21x1_ASAP7_75t_R _31592_ (.A1(net1119),
    .A2(_01348_),
    .B(_01229_),
    .Y(_02012_));
 AO21x2_ASAP7_75t_R _31593_ (.A1(net2723),
    .A2(net3341),
    .B(_01229_),
    .Y(_02013_));
 TAPCELL_ASAP7_75t_R TAP_593 ();
 NAND2x1_ASAP7_75t_R _31595_ (.A(_01268_),
    .B(_01234_),
    .Y(_02015_));
 NAND3x1_ASAP7_75t_R _31596_ (.A(_02012_),
    .B(_02013_),
    .C(_02015_),
    .Y(_02016_));
 AOI211x1_ASAP7_75t_R _31597_ (.A1(net2872),
    .A2(net3289),
    .B(net1920),
    .C(_01215_),
    .Y(_02017_));
 NAND2x1_ASAP7_75t_R _31598_ (.A(_01218_),
    .B(_01327_),
    .Y(_02018_));
 AO21x1_ASAP7_75t_R _31599_ (.A1(net3138),
    .A2(net1122),
    .B(_01215_),
    .Y(_02019_));
 NAND2x1_ASAP7_75t_R _31600_ (.A(_02018_),
    .B(_02019_),
    .Y(_02020_));
 NOR3x1_ASAP7_75t_R _31601_ (.A(_02016_),
    .B(_02017_),
    .C(_02020_),
    .Y(_02021_));
 NAND2x1_ASAP7_75t_R _31602_ (.A(_02010_),
    .B(_02021_),
    .Y(_02022_));
 NOR2x2_ASAP7_75t_R _31603_ (.A(_01208_),
    .B(_01221_),
    .Y(_02023_));
 OA21x2_ASAP7_75t_R _31604_ (.A1(_01328_),
    .A2(_02023_),
    .B(_01103_),
    .Y(_02024_));
 AO21x1_ASAP7_75t_R _31605_ (.A1(_01166_),
    .A2(_01103_),
    .B(_02024_),
    .Y(_02025_));
 NAND2x1_ASAP7_75t_R _31606_ (.A(_01209_),
    .B(_01103_),
    .Y(_02026_));
 OAI21x1_ASAP7_75t_R _31607_ (.A1(_01097_),
    .A2(_01107_),
    .B(_02026_),
    .Y(_02027_));
 AO21x1_ASAP7_75t_R _31608_ (.A1(_01348_),
    .A2(_01204_),
    .B(_01133_),
    .Y(_02028_));
 AO21x1_ASAP7_75t_R _31609_ (.A1(_01228_),
    .A2(_01115_),
    .B(_01133_),
    .Y(_02029_));
 NAND2x1_ASAP7_75t_R _31610_ (.A(_02028_),
    .B(_02029_),
    .Y(_02030_));
 NOR3x1_ASAP7_75t_R _31611_ (.A(_02025_),
    .B(_02027_),
    .C(_02030_),
    .Y(_02031_));
 NAND2x2_ASAP7_75t_R _31612_ (.A(net3142),
    .B(_01109_),
    .Y(_02032_));
 AO21x1_ASAP7_75t_R _31613_ (.A1(_01138_),
    .A2(_02032_),
    .B(_01156_),
    .Y(_02033_));
 AO21x1_ASAP7_75t_R _31614_ (.A1(_01348_),
    .A2(net1696),
    .B(_01156_),
    .Y(_02034_));
 NAND2x1_ASAP7_75t_R _31615_ (.A(_01270_),
    .B(_01163_),
    .Y(_02035_));
 NAND3x1_ASAP7_75t_R _31616_ (.A(_02033_),
    .B(_02034_),
    .C(_02035_),
    .Y(_02036_));
 AO21x1_ASAP7_75t_R _31617_ (.A1(net2522),
    .A2(net940),
    .B(_01170_),
    .Y(_02037_));
 AO21x1_ASAP7_75t_R _31618_ (.A1(net3138),
    .A2(net1076),
    .B(_01170_),
    .Y(_02038_));
 AND2x2_ASAP7_75t_R _31619_ (.A(_02037_),
    .B(_02038_),
    .Y(_02039_));
 AO21x1_ASAP7_75t_R _31620_ (.A1(_01113_),
    .A2(_01115_),
    .B(_01170_),
    .Y(_02040_));
 OA21x2_ASAP7_75t_R _31621_ (.A1(net1158),
    .A2(_01170_),
    .B(_02040_),
    .Y(_02041_));
 NAND2x1_ASAP7_75t_R _31622_ (.A(_02039_),
    .B(_02041_),
    .Y(_02042_));
 NOR2x1_ASAP7_75t_R _31623_ (.A(_02036_),
    .B(_02042_),
    .Y(_02043_));
 NAND2x1_ASAP7_75t_R _31624_ (.A(_02031_),
    .B(_02043_),
    .Y(_02044_));
 NOR2x1_ASAP7_75t_R _31625_ (.A(_02022_),
    .B(_02044_),
    .Y(_02045_));
 AO21x1_ASAP7_75t_R _31626_ (.A1(net1158),
    .A2(_01303_),
    .B(net3417),
    .Y(_02046_));
 AO21x1_ASAP7_75t_R _31627_ (.A1(_01292_),
    .A2(net3138),
    .B(net3417),
    .Y(_02047_));
 NAND2x1_ASAP7_75t_R _31628_ (.A(_01305_),
    .B(_01416_),
    .Y(_02048_));
 AND3x1_ASAP7_75t_R _31629_ (.A(_02046_),
    .B(_02047_),
    .C(_02048_),
    .Y(_02049_));
 AO21x1_ASAP7_75t_R _31630_ (.A1(_01292_),
    .A2(_01204_),
    .B(net3145),
    .Y(_02050_));
 NOR2x2_ASAP7_75t_R _31631_ (.A(net1196),
    .B(net1914),
    .Y(_02051_));
 NAND2x1_ASAP7_75t_R _31632_ (.A(_02051_),
    .B(_01288_),
    .Y(_02052_));
 AND3x1_ASAP7_75t_R _31633_ (.A(_01297_),
    .B(_02050_),
    .C(_02052_),
    .Y(_02053_));
 AND2x2_ASAP7_75t_R _31634_ (.A(_02049_),
    .B(_02053_),
    .Y(_02054_));
 AO21x1_ASAP7_75t_R _31635_ (.A1(_01113_),
    .A2(_02032_),
    .B(net3315),
    .Y(_02055_));
 NAND2x1_ASAP7_75t_R _31636_ (.A(_02051_),
    .B(_01265_),
    .Y(_02056_));
 AND2x2_ASAP7_75t_R _31637_ (.A(_02055_),
    .B(_02056_),
    .Y(_02057_));
 INVx1_ASAP7_75t_R _31638_ (.A(_01248_),
    .Y(_02058_));
 AOI21x1_ASAP7_75t_R _31639_ (.A1(_01251_),
    .A2(_02058_),
    .B(_01404_),
    .Y(_02059_));
 AOI211x1_ASAP7_75t_R _31640_ (.A1(net2872),
    .A2(net3289),
    .B(_01243_),
    .C(_01204_),
    .Y(_02060_));
 NOR2x2_ASAP7_75t_R _31641_ (.A(net3142),
    .B(_01221_),
    .Y(_02061_));
 OA21x2_ASAP7_75t_R _31642_ (.A1(_01327_),
    .A2(_02061_),
    .B(_01251_),
    .Y(_02062_));
 NOR2x1_ASAP7_75t_R _31643_ (.A(_02060_),
    .B(_02062_),
    .Y(_02063_));
 AND3x1_ASAP7_75t_R _31644_ (.A(_02057_),
    .B(_02059_),
    .C(_02063_),
    .Y(_02064_));
 NAND2x1_ASAP7_75t_R _31645_ (.A(_02054_),
    .B(_02064_),
    .Y(_02065_));
 AOI211x1_ASAP7_75t_R _31646_ (.A1(net1595),
    .A2(net1686),
    .B(_01345_),
    .C(net1431),
    .Y(_02066_));
 OA21x2_ASAP7_75t_R _31647_ (.A1(_01268_),
    .A2(_01160_),
    .B(_01351_),
    .Y(_02067_));
 NOR2x1_ASAP7_75t_R _31648_ (.A(_02066_),
    .B(_02067_),
    .Y(_02068_));
 AO21x1_ASAP7_75t_R _31649_ (.A1(net1119),
    .A2(net940),
    .B(net3240),
    .Y(_02069_));
 AND2x2_ASAP7_75t_R _31650_ (.A(_02069_),
    .B(_01347_),
    .Y(_02070_));
 NAND2x1_ASAP7_75t_R _31651_ (.A(_02068_),
    .B(_02070_),
    .Y(_02071_));
 OA21x2_ASAP7_75t_R _31652_ (.A1(_01160_),
    .A2(_01374_),
    .B(_01337_),
    .Y(_02072_));
 OA21x2_ASAP7_75t_R _31653_ (.A1(_01328_),
    .A2(_02023_),
    .B(_01337_),
    .Y(_02073_));
 OR3x1_ASAP7_75t_R _31654_ (.A(_02072_),
    .B(_02073_),
    .C(_01382_),
    .Y(_02074_));
 NOR2x1_ASAP7_75t_R _31655_ (.A(_02071_),
    .B(_02074_),
    .Y(_02075_));
 AO21x1_ASAP7_75t_R _31656_ (.A1(_01113_),
    .A2(net938),
    .B(net2460),
    .Y(_02076_));
 AO21x1_ASAP7_75t_R _31657_ (.A1(net1119),
    .A2(_01348_),
    .B(net2460),
    .Y(_02077_));
 AO21x1_ASAP7_75t_R _31658_ (.A1(net2544),
    .A2(net1122),
    .B(net2460),
    .Y(_02078_));
 NAND3x2_ASAP7_75t_R _31659_ (.B(_02077_),
    .C(_02078_),
    .Y(_02079_),
    .A(_02076_));
 NAND2x2_ASAP7_75t_R _31660_ (.A(_02051_),
    .B(_01315_),
    .Y(_02080_));
 AO21x1_ASAP7_75t_R _31661_ (.A1(_01138_),
    .A2(_01226_),
    .B(_01308_),
    .Y(_02081_));
 NAND2x2_ASAP7_75t_R _31662_ (.A(_02080_),
    .B(_02081_),
    .Y(_02082_));
 NOR2x1_ASAP7_75t_R _31663_ (.A(_01221_),
    .B(_01308_),
    .Y(_02083_));
 INVx1_ASAP7_75t_R _31664_ (.A(_02083_),
    .Y(_02084_));
 AO21x1_ASAP7_75t_R _31665_ (.A1(net3138),
    .A2(net1076),
    .B(_01308_),
    .Y(_02085_));
 NAND2x2_ASAP7_75t_R _31666_ (.A(_02084_),
    .B(_02085_),
    .Y(_02086_));
 NOR3x2_ASAP7_75t_R _31667_ (.B(_02082_),
    .C(_02086_),
    .Y(_02087_),
    .A(_02079_));
 NAND2x2_ASAP7_75t_R _31668_ (.A(_02075_),
    .B(_02087_),
    .Y(_02088_));
 NOR2x2_ASAP7_75t_R _31669_ (.A(_02065_),
    .B(_02088_),
    .Y(_02089_));
 NAND2x2_ASAP7_75t_R _31670_ (.A(_02045_),
    .B(_02089_),
    .Y(_02090_));
 NOR2x2_ASAP7_75t_R _31671_ (.A(_01371_),
    .B(_02090_),
    .Y(_02091_));
 INVx3_ASAP7_75t_R _31672_ (.A(_02091_),
    .Y(_02092_));
 XOR2x1_ASAP7_75t_R _31673_ (.A(_01483_),
    .Y(_02093_),
    .B(_02092_));
 AO21x1_ASAP7_75t_R _31674_ (.A1(net2239),
    .A2(net3168),
    .B(_01967_),
    .Y(_02094_));
 TAPCELL_ASAP7_75t_R TAP_592 ();
 AO21x1_ASAP7_75t_R _31676_ (.A1(_01819_),
    .A2(_01821_),
    .B(_01967_),
    .Y(_02096_));
 NAND2x2_ASAP7_75t_R _31677_ (.A(_02094_),
    .B(_02096_),
    .Y(_02097_));
 NAND2x1_ASAP7_75t_R _31678_ (.A(net1554),
    .B(_01970_),
    .Y(_02098_));
 NOR2x2_ASAP7_75t_R _31679_ (.A(net1360),
    .B(net1298),
    .Y(_02099_));
 INVx3_ASAP7_75t_R _31680_ (.A(_02099_),
    .Y(_02100_));
 AO21x2_ASAP7_75t_R _31681_ (.A1(_02100_),
    .A2(_01935_),
    .B(_01967_),
    .Y(_02101_));
 NAND2x2_ASAP7_75t_R _31682_ (.A(_02098_),
    .B(_02101_),
    .Y(_02102_));
 NOR2x2_ASAP7_75t_R _31683_ (.A(_01857_),
    .B(_01967_),
    .Y(_02103_));
 NOR3x2_ASAP7_75t_R _31684_ (.B(_02102_),
    .C(_02103_),
    .Y(_02104_),
    .A(_02097_));
 OR3x2_ASAP7_75t_R _31685_ (.A(_01914_),
    .B(_01759_),
    .C(_00595_),
    .Y(_02105_));
 NAND3x2_ASAP7_75t_R _31686_ (.B(_01977_),
    .C(_02105_),
    .Y(_02106_),
    .A(_02104_));
 NOR3x2_ASAP7_75t_R _31687_ (.B(_01914_),
    .C(_01759_),
    .Y(_02107_),
    .A(_02106_));
 TAPCELL_ASAP7_75t_R TAP_591 ();
 NAND2x2_ASAP7_75t_R _31689_ (.A(_01862_),
    .B(_01847_),
    .Y(_02109_));
 CKINVDCx9p33_ASAP7_75t_R _31690_ (.A(_01769_),
    .Y(_02110_));
 TAPCELL_ASAP7_75t_R TAP_590 ();
 AO21x1_ASAP7_75t_R _31692_ (.A1(_02110_),
    .A2(_01832_),
    .B(_01851_),
    .Y(_02112_));
 NAND2x2_ASAP7_75t_R _31693_ (.A(_02109_),
    .B(_02112_),
    .Y(_02113_));
 NOR2x2_ASAP7_75t_R _31694_ (.A(_01869_),
    .B(_01857_),
    .Y(_02114_));
 OA21x2_ASAP7_75t_R _31695_ (.A1(_01855_),
    .A2(_02114_),
    .B(_01847_),
    .Y(_02115_));
 NOR3x2_ASAP7_75t_R _31696_ (.B(_01854_),
    .C(_02115_),
    .Y(_02116_),
    .A(_02113_));
 NOR2x2_ASAP7_75t_R _31697_ (.A(net955),
    .B(_01850_),
    .Y(_02117_));
 NAND2x1_ASAP7_75t_R _31698_ (.A(_02117_),
    .B(_01864_),
    .Y(_02118_));
 TAPCELL_ASAP7_75t_R TAP_589 ();
 AO21x1_ASAP7_75t_R _31700_ (.A1(net2175),
    .A2(_02100_),
    .B(net2494),
    .Y(_02120_));
 NAND2x1_ASAP7_75t_R _31701_ (.A(_02118_),
    .B(_02120_),
    .Y(_02121_));
 AO21x1_ASAP7_75t_R _31702_ (.A1(net2563),
    .A2(net2218),
    .B(net2494),
    .Y(_02122_));
 AO21x1_ASAP7_75t_R _31703_ (.A1(net2239),
    .A2(net3169),
    .B(_01863_),
    .Y(_02123_));
 NOR2x2_ASAP7_75t_R _31704_ (.A(_01786_),
    .B(_01857_),
    .Y(_02124_));
 NAND2x1_ASAP7_75t_R _31705_ (.A(_02124_),
    .B(_01864_),
    .Y(_02125_));
 NAND3x1_ASAP7_75t_R _31706_ (.A(_02122_),
    .B(_02123_),
    .C(_02125_),
    .Y(_02126_));
 NOR2x1_ASAP7_75t_R _31707_ (.A(_02121_),
    .B(_02126_),
    .Y(_02127_));
 NAND2x2_ASAP7_75t_R _31708_ (.A(_02116_),
    .B(_02127_),
    .Y(_02128_));
 NAND2x2_ASAP7_75t_R _31709_ (.A(_01869_),
    .B(_01830_),
    .Y(_02129_));
 AO21x1_ASAP7_75t_R _31710_ (.A1(_02129_),
    .A2(_01790_),
    .B(_01781_),
    .Y(_02130_));
 INVx4_ASAP7_75t_R _31711_ (.A(_01781_),
    .Y(_02131_));
 NAND2x1_ASAP7_75t_R _31712_ (.A(_01858_),
    .B(_02131_),
    .Y(_02132_));
 AND2x2_ASAP7_75t_R _31713_ (.A(_02130_),
    .B(_02132_),
    .Y(_02133_));
 NAND2x2_ASAP7_75t_R _31714_ (.A(net1131),
    .B(net3258),
    .Y(_02134_));
 AND2x2_ASAP7_75t_R _31715_ (.A(net2218),
    .B(_02134_),
    .Y(_02135_));
 INVx1_ASAP7_75t_R _31716_ (.A(_02135_),
    .Y(_02136_));
 OAI21x1_ASAP7_75t_R _31717_ (.A1(net3274),
    .A2(_02136_),
    .B(_01762_),
    .Y(_02137_));
 AND2x2_ASAP7_75t_R _31718_ (.A(_02133_),
    .B(_02137_),
    .Y(_02138_));
 TAPCELL_ASAP7_75t_R TAP_588 ();
 NAND2x1_ASAP7_75t_R _31720_ (.A(_00594_),
    .B(_01914_),
    .Y(_02140_));
 NOR2x2_ASAP7_75t_R _31721_ (.A(_02140_),
    .B(_01887_),
    .Y(_02141_));
 NAND2x1_ASAP7_75t_R _31722_ (.A(net1129),
    .B(_02141_),
    .Y(_02142_));
 TAPCELL_ASAP7_75t_R TAP_587 ();
 TAPCELL_ASAP7_75t_R TAP_586 ();
 TAPCELL_ASAP7_75t_R TAP_585 ();
 AO21x1_ASAP7_75t_R _31726_ (.A1(net2175),
    .A2(_01946_),
    .B(_01828_),
    .Y(_02146_));
 OAI21x1_ASAP7_75t_R _31727_ (.A1(net1116),
    .A2(_02142_),
    .B(_02146_),
    .Y(_02147_));
 AO21x1_ASAP7_75t_R _31728_ (.A1(_02110_),
    .A2(_01946_),
    .B(_01809_),
    .Y(_02148_));
 NAND2x1_ASAP7_75t_R _31729_ (.A(_01776_),
    .B(net1465),
    .Y(_02149_));
 AO21x1_ASAP7_75t_R _31730_ (.A1(_02149_),
    .A2(_01938_),
    .B(_01809_),
    .Y(_02150_));
 INVx1_ASAP7_75t_R _31731_ (.A(_01790_),
    .Y(_02151_));
 NAND2x1_ASAP7_75t_R _31732_ (.A(_02151_),
    .B(_01810_),
    .Y(_02152_));
 NAND3x1_ASAP7_75t_R _31733_ (.A(_02148_),
    .B(_02150_),
    .C(_02152_),
    .Y(_02153_));
 NOR2x1_ASAP7_75t_R _31734_ (.A(_02147_),
    .B(_02153_),
    .Y(_02154_));
 NAND2x2_ASAP7_75t_R _31735_ (.A(_02138_),
    .B(_02154_),
    .Y(_02155_));
 TAPCELL_ASAP7_75t_R TAP_584 ();
 AO21x1_ASAP7_75t_R _31737_ (.A1(net1413),
    .A2(_01946_),
    .B(net3128),
    .Y(_02157_));
 TAPCELL_ASAP7_75t_R TAP_583 ();
 TAPCELL_ASAP7_75t_R TAP_582 ();
 AO21x1_ASAP7_75t_R _31740_ (.A1(net2619),
    .A2(_01908_),
    .B(net3128),
    .Y(_02160_));
 TAPCELL_ASAP7_75t_R TAP_581 ();
 NAND2x1_ASAP7_75t_R _31742_ (.A(net1460),
    .B(_01888_),
    .Y(_02162_));
 AND3x1_ASAP7_75t_R _31743_ (.A(_02157_),
    .B(_02160_),
    .C(_02162_),
    .Y(_02163_));
 TAPCELL_ASAP7_75t_R TAP_580 ();
 TAPCELL_ASAP7_75t_R TAP_579 ();
 TAPCELL_ASAP7_75t_R TAP_578 ();
 TAPCELL_ASAP7_75t_R TAP_577 ();
 AOI211x1_ASAP7_75t_R _31748_ (.A1(_01770_),
    .A2(_01776_),
    .B(_01878_),
    .C(_01857_),
    .Y(_02168_));
 INVx1_ASAP7_75t_R _31749_ (.A(_02168_),
    .Y(_02169_));
 NAND2x1_ASAP7_75t_R _31750_ (.A(_01843_),
    .B(_01876_),
    .Y(_02170_));
 TAPCELL_ASAP7_75t_R TAP_576 ();
 AO21x1_ASAP7_75t_R _31752_ (.A1(_01821_),
    .A2(net1138),
    .B(_01878_),
    .Y(_02172_));
 AND3x1_ASAP7_75t_R _31753_ (.A(_02169_),
    .B(_02170_),
    .C(_02172_),
    .Y(_02173_));
 NAND2x2_ASAP7_75t_R _31754_ (.A(_02163_),
    .B(_02173_),
    .Y(_02174_));
 NOR3x2_ASAP7_75t_R _31755_ (.B(_02155_),
    .C(_02174_),
    .Y(_02175_),
    .A(_02128_));
 NOR2x1_ASAP7_75t_R _31756_ (.A(_01804_),
    .B(_01938_),
    .Y(_02176_));
 INVx3_ASAP7_75t_R _31757_ (.A(_01892_),
    .Y(_02177_));
 OA21x2_ASAP7_75t_R _31758_ (.A1(_02176_),
    .A2(_02177_),
    .B(_01940_),
    .Y(_02178_));
 TAPCELL_ASAP7_75t_R TAP_575 ();
 AO21x1_ASAP7_75t_R _31760_ (.A1(_02110_),
    .A2(_01935_),
    .B(net2194),
    .Y(_02180_));
 OAI21x1_ASAP7_75t_R _31761_ (.A1(_01877_),
    .A2(net2194),
    .B(_02180_),
    .Y(_02181_));
 NOR2x1_ASAP7_75t_R _31762_ (.A(_02178_),
    .B(_02181_),
    .Y(_02182_));
 NOR2x1_ASAP7_75t_R _31763_ (.A(_01870_),
    .B(net2549),
    .Y(_02183_));
 NAND2x1_ASAP7_75t_R _31764_ (.A(net3259),
    .B(_02183_),
    .Y(_02184_));
 NOR2x1_ASAP7_75t_R _31765_ (.A(net3275),
    .B(net3170),
    .Y(_02185_));
 INVx2_ASAP7_75t_R _31766_ (.A(_02185_),
    .Y(_02186_));
 AO21x1_ASAP7_75t_R _31767_ (.A1(_01935_),
    .A2(_01850_),
    .B(net2215),
    .Y(_02187_));
 AND3x1_ASAP7_75t_R _31768_ (.A(_02184_),
    .B(_02186_),
    .C(_02187_),
    .Y(_02188_));
 NAND2x1_ASAP7_75t_R _31769_ (.A(_02182_),
    .B(_02188_),
    .Y(_02189_));
 NOR2x2_ASAP7_75t_R _31770_ (.A(net1299),
    .B(_01777_),
    .Y(_02190_));
 INVx1_ASAP7_75t_R _31771_ (.A(_02190_),
    .Y(_02191_));
 NAND2x1_ASAP7_75t_R _31772_ (.A(_01770_),
    .B(net1556),
    .Y(_02192_));
 TAPCELL_ASAP7_75t_R TAP_574 ();
 AO21x1_ASAP7_75t_R _31774_ (.A1(_02191_),
    .A2(_02192_),
    .B(net2140),
    .Y(_02194_));
 INVx1_ASAP7_75t_R _31775_ (.A(_01918_),
    .Y(_02195_));
 AO21x1_ASAP7_75t_R _31776_ (.A1(_01821_),
    .A2(net1138),
    .B(net2140),
    .Y(_02196_));
 AND3x1_ASAP7_75t_R _31777_ (.A(_02194_),
    .B(_02195_),
    .C(_02196_),
    .Y(_02197_));
 NAND2x1_ASAP7_75t_R _31778_ (.A(_02117_),
    .B(_01904_),
    .Y(_02198_));
 AO21x1_ASAP7_75t_R _31779_ (.A1(_02110_),
    .A2(net2175),
    .B(_01905_),
    .Y(_02199_));
 NAND2x1_ASAP7_75t_R _31780_ (.A(_02198_),
    .B(_02199_),
    .Y(_02200_));
 AO21x1_ASAP7_75t_R _31781_ (.A1(net1138),
    .A2(_01908_),
    .B(_01905_),
    .Y(_02201_));
 AOI22x1_ASAP7_75t_R _31782_ (.A1(_01814_),
    .A2(net2299),
    .B1(net1454),
    .B2(net1127),
    .Y(_02202_));
 NOR2x1_ASAP7_75t_R _31783_ (.A(_01905_),
    .B(_02202_),
    .Y(_02203_));
 INVx1_ASAP7_75t_R _31784_ (.A(_02203_),
    .Y(_02204_));
 NAND2x1_ASAP7_75t_R _31785_ (.A(_02201_),
    .B(_02204_),
    .Y(_02205_));
 NOR2x1_ASAP7_75t_R _31786_ (.A(_02200_),
    .B(_02205_),
    .Y(_02206_));
 NAND2x1_ASAP7_75t_R _31787_ (.A(_02197_),
    .B(_02206_),
    .Y(_02207_));
 NOR2x2_ASAP7_75t_R _31788_ (.A(_02189_),
    .B(_02207_),
    .Y(_02208_));
 AO21x1_ASAP7_75t_R _31789_ (.A1(net2619),
    .A2(_01908_),
    .B(_01967_),
    .Y(_02209_));
 OA21x2_ASAP7_75t_R _31790_ (.A1(_01967_),
    .A2(_01952_),
    .B(_02209_),
    .Y(_02210_));
 NAND2x2_ASAP7_75t_R _31791_ (.A(_01765_),
    .B(_01805_),
    .Y(_02211_));
 AND3x1_ASAP7_75t_R _31792_ (.A(_02211_),
    .B(_01974_),
    .C(net1459),
    .Y(_02212_));
 NAND2x1_ASAP7_75t_R _31793_ (.A(net1555),
    .B(_01974_),
    .Y(_02213_));
 NAND2x1_ASAP7_75t_R _31794_ (.A(_02099_),
    .B(_01974_),
    .Y(_02214_));
 OAI21x1_ASAP7_75t_R _31795_ (.A1(_02211_),
    .A2(_02213_),
    .B(_02214_),
    .Y(_02215_));
 NOR2x1_ASAP7_75t_R _31796_ (.A(_02212_),
    .B(_02215_),
    .Y(_02216_));
 OA21x2_ASAP7_75t_R _31797_ (.A1(_01806_),
    .A2(_01843_),
    .B(_01970_),
    .Y(_02217_));
 AOI211x1_ASAP7_75t_R _31798_ (.A1(net1116),
    .A2(net1450),
    .B(_01967_),
    .C(_01850_),
    .Y(_02218_));
 NOR2x1_ASAP7_75t_R _31799_ (.A(_02217_),
    .B(_02218_),
    .Y(_02219_));
 NAND3x1_ASAP7_75t_R _31800_ (.A(_02210_),
    .B(_02216_),
    .C(_02219_),
    .Y(_02220_));
 NOR2x1_ASAP7_75t_R _31801_ (.A(_01955_),
    .B(_01819_),
    .Y(_02221_));
 TAPCELL_ASAP7_75t_R TAP_573 ();
 AOI21x1_ASAP7_75t_R _31803_ (.A1(net2370),
    .A2(_01795_),
    .B(net2352),
    .Y(_02223_));
 NOR2x1_ASAP7_75t_R _31804_ (.A(_02221_),
    .B(_02223_),
    .Y(_02224_));
 AO21x1_ASAP7_75t_R _31805_ (.A1(net1116),
    .A2(net1449),
    .B(net1299),
    .Y(_02225_));
 TAPCELL_ASAP7_75t_R TAP_572 ();
 AO21x1_ASAP7_75t_R _31807_ (.A1(_02225_),
    .A2(net1527),
    .B(net2352),
    .Y(_02227_));
 AND2x2_ASAP7_75t_R _31808_ (.A(_02224_),
    .B(_02227_),
    .Y(_02228_));
 NOR2x1_ASAP7_75t_R _31809_ (.A(_01870_),
    .B(net2262),
    .Y(_02229_));
 TAPCELL_ASAP7_75t_R TAP_571 ();
 AOI211x1_ASAP7_75t_R _31811_ (.A1(net1116),
    .A2(_01776_),
    .B(net3125),
    .C(_01857_),
    .Y(_02231_));
 AOI21x1_ASAP7_75t_R _31812_ (.A1(_01765_),
    .A2(_02229_),
    .B(_02231_),
    .Y(_02232_));
 AO21x1_ASAP7_75t_R _31813_ (.A1(net1413),
    .A2(net1527),
    .B(net3125),
    .Y(_02233_));
 AND2x2_ASAP7_75t_R _31814_ (.A(_02233_),
    .B(_01950_),
    .Y(_02234_));
 NAND3x1_ASAP7_75t_R _31815_ (.A(_02228_),
    .B(_02232_),
    .C(_02234_),
    .Y(_02235_));
 NOR2x1_ASAP7_75t_R _31816_ (.A(_02220_),
    .B(_02235_),
    .Y(_02236_));
 NAND2x2_ASAP7_75t_R _31817_ (.A(_02208_),
    .B(_02236_),
    .Y(_02237_));
 INVx1_ASAP7_75t_R _31818_ (.A(_02237_),
    .Y(_02238_));
 NAND2x2_ASAP7_75t_R _31819_ (.A(_02175_),
    .B(_02238_),
    .Y(_02239_));
 INVx2_ASAP7_75t_R _31820_ (.A(_01987_),
    .Y(_02240_));
 OAI21x1_ASAP7_75t_R _31821_ (.A1(_02107_),
    .A2(_02239_),
    .B(_02240_),
    .Y(_02241_));
 INVx1_ASAP7_75t_R _31822_ (.A(_02155_),
    .Y(_02242_));
 NOR2x1_ASAP7_75t_R _31823_ (.A(_02174_),
    .B(_02128_),
    .Y(_02243_));
 NAND2x1_ASAP7_75t_R _31824_ (.A(_02242_),
    .B(_02243_),
    .Y(_02244_));
 NOR2x2_ASAP7_75t_R _31825_ (.A(_02237_),
    .B(_02244_),
    .Y(_02245_));
 NOR2x1_ASAP7_75t_R _31826_ (.A(_01915_),
    .B(_02106_),
    .Y(_02246_));
 NAND2x2_ASAP7_75t_R _31827_ (.A(net3263),
    .B(_02246_),
    .Y(_02247_));
 NAND3x2_ASAP7_75t_R _31828_ (.B(_01987_),
    .C(_02247_),
    .Y(_02248_),
    .A(_02245_));
 NAND2x2_ASAP7_75t_R _31829_ (.A(_02241_),
    .B(_02248_),
    .Y(_02249_));
 NAND2x1_ASAP7_75t_R _31830_ (.A(_22083_),
    .B(_01073_),
    .Y(_02250_));
 AO21x1_ASAP7_75t_R _31831_ (.A1(_21967_),
    .A2(_21969_),
    .B(_01072_),
    .Y(_02251_));
 NAND2x1_ASAP7_75t_R _31832_ (.A(_02250_),
    .B(_02251_),
    .Y(_02252_));
 OAI21x1_ASAP7_75t_R _31833_ (.A1(net3083),
    .A2(net2038),
    .B(_01073_),
    .Y(_02253_));
 AO21x1_ASAP7_75t_R _31834_ (.A1(_21920_),
    .A2(net1792),
    .B(_01072_),
    .Y(_02254_));
 NAND2x1_ASAP7_75t_R _31835_ (.A(_02254_),
    .B(_02253_),
    .Y(_02255_));
 NOR2x1_ASAP7_75t_R _31836_ (.A(_02252_),
    .B(_02255_),
    .Y(_02256_));
 OA21x2_ASAP7_75t_R _31837_ (.A1(net2038),
    .A2(_21909_),
    .B(_01079_),
    .Y(_02257_));
 AOI211x1_ASAP7_75t_R _31838_ (.A1(net1139),
    .A2(net1049),
    .B(net2425),
    .C(net1847),
    .Y(_02258_));
 NAND2x2_ASAP7_75t_R _31839_ (.A(net1651),
    .B(_21917_),
    .Y(_02259_));
 TAPCELL_ASAP7_75t_R TAP_570 ();
 OAI21x1_ASAP7_75t_R _31841_ (.A1(_21925_),
    .A2(_21966_),
    .B(net1256),
    .Y(_02261_));
 AOI21x1_ASAP7_75t_R _31842_ (.A1(net1038),
    .A2(_02261_),
    .B(net3152),
    .Y(_02262_));
 NOR3x1_ASAP7_75t_R _31843_ (.A(_02257_),
    .B(_02258_),
    .C(_02262_),
    .Y(_02263_));
 NAND2x1_ASAP7_75t_R _31844_ (.A(_02263_),
    .B(_02256_),
    .Y(_02264_));
 AO21x1_ASAP7_75t_R _31845_ (.A1(net1038),
    .A2(_22019_),
    .B(net3081),
    .Y(_02265_));
 INVx3_ASAP7_75t_R _31846_ (.A(_22100_),
    .Y(_02266_));
 INVx1_ASAP7_75t_R _31847_ (.A(_02261_),
    .Y(_02267_));
 NAND2x1_ASAP7_75t_R _31848_ (.A(_02266_),
    .B(_02267_),
    .Y(_02268_));
 NOR2x2_ASAP7_75t_R _31849_ (.A(_21904_),
    .B(_21954_),
    .Y(_02269_));
 NAND2x1_ASAP7_75t_R _31850_ (.A(_02269_),
    .B(_02266_),
    .Y(_02270_));
 AND3x1_ASAP7_75t_R _31851_ (.A(_02265_),
    .B(_02268_),
    .C(_02270_),
    .Y(_02271_));
 AO21x1_ASAP7_75t_R _31852_ (.A1(net1048),
    .A2(_22080_),
    .B(_22091_),
    .Y(_02272_));
 NAND2x2_ASAP7_75t_R _31853_ (.A(_21925_),
    .B(net1255),
    .Y(_02273_));
 TAPCELL_ASAP7_75t_R TAP_569 ();
 AO21x1_ASAP7_75t_R _31855_ (.A1(_21940_),
    .A2(_02273_),
    .B(_22091_),
    .Y(_02275_));
 NAND2x2_ASAP7_75t_R _31856_ (.A(net3167),
    .B(_22092_),
    .Y(_02276_));
 AND3x1_ASAP7_75t_R _31857_ (.A(_02272_),
    .B(_02275_),
    .C(_02276_),
    .Y(_02277_));
 NAND2x1_ASAP7_75t_R _31858_ (.A(_02271_),
    .B(_02277_),
    .Y(_02278_));
 NOR2x1_ASAP7_75t_R _31859_ (.A(_02264_),
    .B(_02278_),
    .Y(_02279_));
 AO21x1_ASAP7_75t_R _31860_ (.A1(net3155),
    .A2(net2510),
    .B(_22064_),
    .Y(_02280_));
 AO21x1_ASAP7_75t_R _31861_ (.A1(net991),
    .A2(_21940_),
    .B(_22064_),
    .Y(_02281_));
 OAI21x1_ASAP7_75t_R _31862_ (.A1(_22044_),
    .A2(_02269_),
    .B(_22049_),
    .Y(_02282_));
 AND3x1_ASAP7_75t_R _31863_ (.A(_02280_),
    .B(_02281_),
    .C(_02282_),
    .Y(_02283_));
 TAPCELL_ASAP7_75t_R TAP_568 ();
 AOI211x1_ASAP7_75t_R _31865_ (.A1(net1139),
    .A2(net1049),
    .B(_22061_),
    .C(net1040),
    .Y(_02285_));
 NOR2x2_ASAP7_75t_R _31866_ (.A(_21887_),
    .B(net1714),
    .Y(_02286_));
 OA21x2_ASAP7_75t_R _31867_ (.A1(_22083_),
    .A2(_02286_),
    .B(_22062_),
    .Y(_02287_));
 AOI211x1_ASAP7_75t_R _31868_ (.A1(_01085_),
    .A2(_22062_),
    .B(_02285_),
    .C(_02287_),
    .Y(_02288_));
 NAND2x1_ASAP7_75t_R _31869_ (.A(_02283_),
    .B(_02288_),
    .Y(_02289_));
 AO21x1_ASAP7_75t_R _31870_ (.A1(net2293),
    .A2(_21920_),
    .B(_22070_),
    .Y(_02290_));
 AO21x1_ASAP7_75t_R _31871_ (.A1(_22019_),
    .A2(_21895_),
    .B(_22070_),
    .Y(_02291_));
 INVx2_ASAP7_75t_R _31872_ (.A(_22070_),
    .Y(_02292_));
 NAND2x1_ASAP7_75t_R _31873_ (.A(_21955_),
    .B(_02292_),
    .Y(_02293_));
 AND3x1_ASAP7_75t_R _31874_ (.A(_02290_),
    .B(_02291_),
    .C(_02293_),
    .Y(_02294_));
 NAND2x1_ASAP7_75t_R _31875_ (.A(net1926),
    .B(_22084_),
    .Y(_02295_));
 NAND2x1_ASAP7_75t_R _31876_ (.A(_22084_),
    .B(_21955_),
    .Y(_02296_));
 OAI21x1_ASAP7_75t_R _31877_ (.A1(_21917_),
    .A2(_02295_),
    .B(_02296_),
    .Y(_02297_));
 OA21x2_ASAP7_75t_R _31878_ (.A1(_01082_),
    .A2(_21878_),
    .B(_22084_),
    .Y(_02298_));
 NOR2x1_ASAP7_75t_R _31879_ (.A(_02273_),
    .B(_22077_),
    .Y(_02299_));
 NOR3x1_ASAP7_75t_R _31880_ (.A(_02297_),
    .B(_02298_),
    .C(_02299_),
    .Y(_02300_));
 NAND2x1_ASAP7_75t_R _31881_ (.A(_02294_),
    .B(_02300_),
    .Y(_02301_));
 NOR2x1_ASAP7_75t_R _31882_ (.A(_02289_),
    .B(_02301_),
    .Y(_02302_));
 NAND2x2_ASAP7_75t_R _31883_ (.A(_02279_),
    .B(_02302_),
    .Y(_02303_));
 NOR2x2_ASAP7_75t_R _31884_ (.A(net2637),
    .B(net1851),
    .Y(_02304_));
 INVx3_ASAP7_75t_R _31885_ (.A(_02304_),
    .Y(_02305_));
 NOR2x1_ASAP7_75t_R _31886_ (.A(_21962_),
    .B(_02305_),
    .Y(_02306_));
 AOI211x1_ASAP7_75t_R _31887_ (.A1(net1139),
    .A2(_21876_),
    .B(_21962_),
    .C(net1042),
    .Y(_02307_));
 NOR2x1_ASAP7_75t_R _31888_ (.A(_02306_),
    .B(_02307_),
    .Y(_02308_));
 OA21x2_ASAP7_75t_R _31889_ (.A1(_22083_),
    .A2(_02286_),
    .B(_21980_),
    .Y(_02309_));
 AOI211x1_ASAP7_75t_R _31890_ (.A1(_21887_),
    .A2(_21876_),
    .B(_21976_),
    .C(_21895_),
    .Y(_02310_));
 NOR2x1_ASAP7_75t_R _31891_ (.A(_02309_),
    .B(_02310_),
    .Y(_02311_));
 INVx1_ASAP7_75t_R _31892_ (.A(_22033_),
    .Y(_02312_));
 OA21x2_ASAP7_75t_R _31893_ (.A1(_02312_),
    .A2(_21976_),
    .B(_21981_),
    .Y(_02313_));
 NAND3x1_ASAP7_75t_R _31894_ (.A(_02308_),
    .B(_02311_),
    .C(_02313_),
    .Y(_02314_));
 AOI211x1_ASAP7_75t_R _31895_ (.A1(_21887_),
    .A2(_21876_),
    .B(_21893_),
    .C(net1849),
    .Y(_02315_));
 NOR2x2_ASAP7_75t_R _31896_ (.A(_00551_),
    .B(net1708),
    .Y(_02316_));
 OAI21x1_ASAP7_75t_R _31897_ (.A1(_21937_),
    .A2(_02316_),
    .B(_21885_),
    .Y(_02317_));
 INVx1_ASAP7_75t_R _31898_ (.A(_02317_),
    .Y(_02318_));
 NOR3x1_ASAP7_75t_R _31899_ (.A(_02315_),
    .B(_21945_),
    .C(_02318_),
    .Y(_02319_));
 AO21x1_ASAP7_75t_R _31900_ (.A1(net1829),
    .A2(net1633),
    .B(net1751),
    .Y(_02320_));
 AO21x1_ASAP7_75t_R _31901_ (.A1(_21890_),
    .A2(_21940_),
    .B(net1751),
    .Y(_02321_));
 INVx1_ASAP7_75t_R _31902_ (.A(_21900_),
    .Y(_02322_));
 NOR2x2_ASAP7_75t_R _31903_ (.A(net1906),
    .B(_02322_),
    .Y(_02323_));
 NAND2x1_ASAP7_75t_R _31904_ (.A(_21953_),
    .B(_02323_),
    .Y(_02324_));
 AND3x1_ASAP7_75t_R _31905_ (.A(_02320_),
    .B(_02321_),
    .C(_02324_),
    .Y(_02325_));
 NAND2x1_ASAP7_75t_R _31906_ (.A(_02319_),
    .B(_02325_),
    .Y(_02326_));
 NOR2x1_ASAP7_75t_R _31907_ (.A(_02314_),
    .B(_02326_),
    .Y(_02327_));
 AO21x1_ASAP7_75t_R _31908_ (.A1(net991),
    .A2(_21940_),
    .B(_22004_),
    .Y(_02328_));
 NAND2x1_ASAP7_75t_R _31909_ (.A(_22007_),
    .B(_02328_),
    .Y(_02329_));
 AO21x1_ASAP7_75t_R _31910_ (.A1(_22024_),
    .A2(_21927_),
    .B(_22004_),
    .Y(_02330_));
 OAI21x1_ASAP7_75t_R _31911_ (.A1(_22004_),
    .A2(_02305_),
    .B(_02330_),
    .Y(_02331_));
 NOR2x1_ASAP7_75t_R _31912_ (.A(_02329_),
    .B(_02331_),
    .Y(_02332_));
 AO21x1_ASAP7_75t_R _31913_ (.A1(_22076_),
    .A2(net1792),
    .B(net3151),
    .Y(_02333_));
 AO21x1_ASAP7_75t_R _31914_ (.A1(net1038),
    .A2(_22019_),
    .B(net3151),
    .Y(_02334_));
 AO21x1_ASAP7_75t_R _31915_ (.A1(_21967_),
    .A2(_02273_),
    .B(net3151),
    .Y(_02335_));
 AND3x1_ASAP7_75t_R _31916_ (.A(_02333_),
    .B(_02334_),
    .C(_02335_),
    .Y(_02336_));
 NAND2x1_ASAP7_75t_R _31917_ (.A(_02332_),
    .B(_02336_),
    .Y(_02337_));
 AO21x1_ASAP7_75t_R _31918_ (.A1(net1038),
    .A2(_22018_),
    .B(net3075),
    .Y(_02338_));
 NAND2x1_ASAP7_75t_R _31919_ (.A(_22017_),
    .B(_02338_),
    .Y(_02339_));
 NOR2x2_ASAP7_75t_R _31920_ (.A(net1044),
    .B(_22015_),
    .Y(_02340_));
 INVx1_ASAP7_75t_R _31921_ (.A(_02340_),
    .Y(_02341_));
 AO21x1_ASAP7_75t_R _31922_ (.A1(net1829),
    .A2(net1048),
    .B(net3075),
    .Y(_02342_));
 OAI21x1_ASAP7_75t_R _31923_ (.A1(_21966_),
    .A2(_02341_),
    .B(_02342_),
    .Y(_02343_));
 NOR2x1_ASAP7_75t_R _31924_ (.A(_02339_),
    .B(_02343_),
    .Y(_02344_));
 TAPCELL_ASAP7_75t_R TAP_567 ();
 AO21x1_ASAP7_75t_R _31926_ (.A1(_22024_),
    .A2(_21927_),
    .B(net2556),
    .Y(_02346_));
 OAI21x1_ASAP7_75t_R _31927_ (.A1(net1829),
    .A2(net2556),
    .B(_02346_),
    .Y(_02347_));
 NOR2x2_ASAP7_75t_R _31928_ (.A(_21895_),
    .B(_22028_),
    .Y(_02348_));
 INVx1_ASAP7_75t_R _31929_ (.A(_02348_),
    .Y(_02349_));
 AO21x1_ASAP7_75t_R _31930_ (.A1(net1038),
    .A2(net3155),
    .B(net2556),
    .Y(_02350_));
 OAI21x1_ASAP7_75t_R _31931_ (.A1(_21966_),
    .A2(_02349_),
    .B(_02350_),
    .Y(_02351_));
 NOR2x1_ASAP7_75t_R _31932_ (.A(_02347_),
    .B(_02351_),
    .Y(_02352_));
 NAND2x1_ASAP7_75t_R _31933_ (.A(_02344_),
    .B(_02352_),
    .Y(_02353_));
 NOR2x1_ASAP7_75t_R _31934_ (.A(_02337_),
    .B(_02353_),
    .Y(_02354_));
 NAND2x1_ASAP7_75t_R _31935_ (.A(_02327_),
    .B(_02354_),
    .Y(_02355_));
 NOR2x2_ASAP7_75t_R _31936_ (.A(_02355_),
    .B(_02303_),
    .Y(_02356_));
 NAND2x2_ASAP7_75t_R _31937_ (.A(_21914_),
    .B(_02356_),
    .Y(_02357_));
 AO21x1_ASAP7_75t_R _31938_ (.A1(_01691_),
    .A2(_01674_),
    .B(_01701_),
    .Y(_02358_));
 AO21x1_ASAP7_75t_R _31939_ (.A1(_01592_),
    .A2(_01644_),
    .B(_01701_),
    .Y(_02359_));
 AND2x2_ASAP7_75t_R _31940_ (.A(_02358_),
    .B(_02359_),
    .Y(_02360_));
 NAND2x2_ASAP7_75t_R _31941_ (.A(net1887),
    .B(net3416),
    .Y(_02361_));
 TAPCELL_ASAP7_75t_R TAP_566 ();
 NAND2x2_ASAP7_75t_R _31943_ (.A(_01555_),
    .B(_01491_),
    .Y(_02363_));
 TAPCELL_ASAP7_75t_R TAP_565 ();
 AO31x2_ASAP7_75t_R _31945_ (.A1(net2524),
    .A2(net1605),
    .A3(_02363_),
    .B(_01685_),
    .Y(_02365_));
 AO21x1_ASAP7_75t_R _31946_ (.A1(_01691_),
    .A2(_01687_),
    .B(_01685_),
    .Y(_02366_));
 NAND3x1_ASAP7_75t_R _31947_ (.A(_02360_),
    .B(_02365_),
    .C(_02366_),
    .Y(_02367_));
 AND2x6_ASAP7_75t_R _31948_ (.A(_01585_),
    .B(_01667_),
    .Y(_02368_));
 NAND2x2_ASAP7_75t_R _31949_ (.A(_01562_),
    .B(_02368_),
    .Y(_02369_));
 AO21x1_ASAP7_75t_R _31950_ (.A1(net3135),
    .A2(_01641_),
    .B(_01668_),
    .Y(_02370_));
 NAND2x1_ASAP7_75t_R _31951_ (.A(_02369_),
    .B(_02370_),
    .Y(_02371_));
 INVx2_ASAP7_75t_R _31952_ (.A(_01525_),
    .Y(_02372_));
 AO21x1_ASAP7_75t_R _31953_ (.A1(_01699_),
    .A2(_02372_),
    .B(_01668_),
    .Y(_02373_));
 OAI21x1_ASAP7_75t_R _31954_ (.A1(net2366),
    .A2(_01668_),
    .B(_02373_),
    .Y(_02374_));
 NOR2x1_ASAP7_75t_R _31955_ (.A(_02371_),
    .B(_02374_),
    .Y(_02375_));
 TAPCELL_ASAP7_75t_R TAP_564 ();
 AO21x1_ASAP7_75t_R _31957_ (.A1(net2729),
    .A2(net3149),
    .B(net2733),
    .Y(_02377_));
 AO21x1_ASAP7_75t_R _31958_ (.A1(net3137),
    .A2(_01590_),
    .B(net2733),
    .Y(_02378_));
 NAND2x1_ASAP7_75t_R _31959_ (.A(_02377_),
    .B(_02378_),
    .Y(_02379_));
 AO21x1_ASAP7_75t_R _31960_ (.A1(_01689_),
    .A2(_01691_),
    .B(net2733),
    .Y(_02380_));
 OAI21x1_ASAP7_75t_R _31961_ (.A1(net2064),
    .A2(net2733),
    .B(_02380_),
    .Y(_02381_));
 NOR2x1_ASAP7_75t_R _31962_ (.A(_02379_),
    .B(_02381_),
    .Y(_02382_));
 NAND2x1_ASAP7_75t_R _31963_ (.A(_02375_),
    .B(_02382_),
    .Y(_02383_));
 NOR2x1_ASAP7_75t_R _31964_ (.A(_02367_),
    .B(_02383_),
    .Y(_02384_));
 AOI21x1_ASAP7_75t_R _31965_ (.A1(_02363_),
    .A2(net1104),
    .B(_01735_),
    .Y(_02385_));
 AOI21x1_ASAP7_75t_R _31966_ (.A1(_01674_),
    .A2(net2066),
    .B(_01735_),
    .Y(_02386_));
 AOI211x1_ASAP7_75t_R _31967_ (.A1(_01562_),
    .A2(_01737_),
    .B(_02385_),
    .C(_02386_),
    .Y(_02387_));
 INVx2_ASAP7_75t_R _31968_ (.A(_01728_),
    .Y(_02388_));
 AOI21x1_ASAP7_75t_R _31969_ (.A1(net3255),
    .A2(net3266),
    .B(net3175),
    .Y(_02389_));
 OAI21x1_ASAP7_75t_R _31970_ (.A1(_01555_),
    .A2(_01576_),
    .B(_01491_),
    .Y(_02390_));
 NOR2x2_ASAP7_75t_R _31971_ (.A(_01728_),
    .B(_02390_),
    .Y(_02391_));
 AOI211x1_ASAP7_75t_R _31972_ (.A1(net3257),
    .A2(_02388_),
    .B(_02389_),
    .C(_02391_),
    .Y(_02392_));
 NAND2x1_ASAP7_75t_R _31973_ (.A(_02387_),
    .B(_02392_),
    .Y(_02393_));
 NOR2x1_ASAP7_75t_R _31974_ (.A(_01590_),
    .B(_01715_),
    .Y(_02394_));
 TAPCELL_ASAP7_75t_R TAP_563 ();
 AOI211x1_ASAP7_75t_R _31976_ (.A1(net1120),
    .A2(_01494_),
    .B(_01715_),
    .C(_01644_),
    .Y(_02396_));
 NOR2x1_ASAP7_75t_R _31977_ (.A(_02394_),
    .B(_02396_),
    .Y(_02397_));
 AO21x1_ASAP7_75t_R _31978_ (.A1(_01689_),
    .A2(_01600_),
    .B(_01715_),
    .Y(_02398_));
 AO21x2_ASAP7_75t_R _31979_ (.A1(_01607_),
    .A2(net2254),
    .B(_01715_),
    .Y(_02399_));
 AND2x2_ASAP7_75t_R _31980_ (.A(_02398_),
    .B(_02399_),
    .Y(_02400_));
 NAND2x1_ASAP7_75t_R _31981_ (.A(_02397_),
    .B(_02400_),
    .Y(_02401_));
 AOI211x1_ASAP7_75t_R _31982_ (.A1(net1120),
    .A2(net1263),
    .B(net3256),
    .C(net2376),
    .Y(_02402_));
 INVx1_ASAP7_75t_R _31983_ (.A(_02402_),
    .Y(_02403_));
 AO21x1_ASAP7_75t_R _31984_ (.A1(_02390_),
    .A2(net1605),
    .B(net3256),
    .Y(_02404_));
 NAND2x1_ASAP7_75t_R _31985_ (.A(_01582_),
    .B(_01711_),
    .Y(_02405_));
 NAND3x1_ASAP7_75t_R _31986_ (.A(_02403_),
    .B(_02404_),
    .C(_02405_),
    .Y(_02406_));
 NOR3x1_ASAP7_75t_R _31987_ (.A(_02393_),
    .B(_02401_),
    .C(_02406_),
    .Y(_02407_));
 NAND2x1_ASAP7_75t_R _31988_ (.A(_02384_),
    .B(_02407_),
    .Y(_02408_));
 AO21x1_ASAP7_75t_R _31989_ (.A1(net3267),
    .A2(net2254),
    .B(_01636_),
    .Y(_02409_));
 AND2x2_ASAP7_75t_R _31990_ (.A(_02409_),
    .B(_01639_),
    .Y(_02410_));
 AOI211x1_ASAP7_75t_R _31991_ (.A1(_01498_),
    .A2(net1897),
    .B(net2746),
    .C(net2078),
    .Y(_02411_));
 AOI211x1_ASAP7_75t_R _31992_ (.A1(_01498_),
    .A2(_01494_),
    .B(_01644_),
    .C(net2746),
    .Y(_02412_));
 NOR2x1_ASAP7_75t_R _31993_ (.A(_02411_),
    .B(_02412_),
    .Y(_02413_));
 NOR2x2_ASAP7_75t_R _31994_ (.A(net1399),
    .B(net2379),
    .Y(_02414_));
 OA21x2_ASAP7_75t_R _31995_ (.A1(_01688_),
    .A2(_01525_),
    .B(_01621_),
    .Y(_02415_));
 AOI21x1_ASAP7_75t_R _31996_ (.A1(_01621_),
    .A2(_02414_),
    .B(_02415_),
    .Y(_02416_));
 NAND3x1_ASAP7_75t_R _31997_ (.A(_02410_),
    .B(_02413_),
    .C(_02416_),
    .Y(_02417_));
 AO21x1_ASAP7_75t_R _31998_ (.A1(net2572),
    .A2(net2062),
    .B(net2334),
    .Y(_02418_));
 NAND2x2_ASAP7_75t_R _31999_ (.A(_01498_),
    .B(_01589_),
    .Y(_02419_));
 AO21x1_ASAP7_75t_R _32000_ (.A1(_02419_),
    .A2(_01496_),
    .B(net2334),
    .Y(_02420_));
 OAI21x1_ASAP7_75t_R _32001_ (.A1(_01688_),
    .A2(_01526_),
    .B(_01657_),
    .Y(_02421_));
 AND3x1_ASAP7_75t_R _32002_ (.A(_02418_),
    .B(_02420_),
    .C(_02421_),
    .Y(_02422_));
 NAND2x1_ASAP7_75t_R _32003_ (.A(_01512_),
    .B(_01506_),
    .Y(_02423_));
 NOR2x1_ASAP7_75t_R _32004_ (.A(net1025),
    .B(net2379),
    .Y(_02424_));
 NOR2x2_ASAP7_75t_R _32005_ (.A(_01515_),
    .B(net2376),
    .Y(_02425_));
 OAI21x1_ASAP7_75t_R _32006_ (.A1(_02424_),
    .A2(_02425_),
    .B(_01504_),
    .Y(_02426_));
 NAND2x2_ASAP7_75t_R _32007_ (.A(_01504_),
    .B(_01635_),
    .Y(_02427_));
 NAND2x1_ASAP7_75t_R _32008_ (.A(_01525_),
    .B(_01504_),
    .Y(_02428_));
 NAND3x1_ASAP7_75t_R _32009_ (.A(_02426_),
    .B(_02427_),
    .C(_02428_),
    .Y(_02429_));
 NOR2x1_ASAP7_75t_R _32010_ (.A(_02423_),
    .B(_02429_),
    .Y(_02430_));
 NAND2x1_ASAP7_75t_R _32011_ (.A(_02422_),
    .B(_02430_),
    .Y(_02431_));
 NOR2x1_ASAP7_75t_R _32012_ (.A(_02417_),
    .B(_02431_),
    .Y(_02432_));
 AO21x1_ASAP7_75t_R _32013_ (.A1(net3265),
    .A2(_01590_),
    .B(net2794),
    .Y(_02433_));
 NAND2x1_ASAP7_75t_R _32014_ (.A(_01596_),
    .B(_02433_),
    .Y(_02434_));
 AO21x1_ASAP7_75t_R _32015_ (.A1(net2572),
    .A2(net2062),
    .B(net2794),
    .Y(_02435_));
 TAPCELL_ASAP7_75t_R TAP_562 ();
 NOR2x2_ASAP7_75t_R _32017_ (.A(net1242),
    .B(_01586_),
    .Y(_02437_));
 NAND2x2_ASAP7_75t_R _32018_ (.A(net1026),
    .B(_02437_),
    .Y(_02438_));
 NAND2x1_ASAP7_75t_R _32019_ (.A(_02435_),
    .B(_02438_),
    .Y(_02439_));
 NOR2x1_ASAP7_75t_R _32020_ (.A(_02434_),
    .B(_02439_),
    .Y(_02440_));
 NOR2x2_ASAP7_75t_R _32021_ (.A(_01644_),
    .B(_01603_),
    .Y(_02441_));
 NAND2x1_ASAP7_75t_R _32022_ (.A(net1026),
    .B(_02441_),
    .Y(_02442_));
 AO21x1_ASAP7_75t_R _32023_ (.A1(net2572),
    .A2(_01583_),
    .B(_01603_),
    .Y(_02443_));
 AO21x1_ASAP7_75t_R _32024_ (.A1(net2524),
    .A2(net3265),
    .B(_01603_),
    .Y(_02444_));
 AND3x1_ASAP7_75t_R _32025_ (.A(_02442_),
    .B(_02443_),
    .C(_02444_),
    .Y(_02445_));
 NAND2x1_ASAP7_75t_R _32026_ (.A(_02440_),
    .B(_02445_),
    .Y(_02446_));
 NOR2x2_ASAP7_75t_R _32027_ (.A(net2376),
    .B(_01561_),
    .Y(_02447_));
 OA21x2_ASAP7_75t_R _32028_ (.A1(_02447_),
    .A2(_01688_),
    .B(_01550_),
    .Y(_02448_));
 INVx1_ASAP7_75t_R _32029_ (.A(_02363_),
    .Y(_02449_));
 OA21x2_ASAP7_75t_R _32030_ (.A1(_02449_),
    .A2(_01680_),
    .B(_01550_),
    .Y(_02450_));
 AOI211x1_ASAP7_75t_R _32031_ (.A1(_01498_),
    .A2(_01494_),
    .B(_01543_),
    .C(net2076),
    .Y(_02451_));
 NOR3x1_ASAP7_75t_R _32032_ (.A(_02448_),
    .B(_02450_),
    .C(_02451_),
    .Y(_02452_));
 NOR2x2_ASAP7_75t_R _32033_ (.A(net2072),
    .B(_01499_),
    .Y(_02453_));
 OAI21x1_ASAP7_75t_R _32034_ (.A1(_01514_),
    .A2(_02453_),
    .B(_01565_),
    .Y(_02454_));
 NAND2x2_ASAP7_75t_R _32035_ (.A(_02454_),
    .B(_01567_),
    .Y(_02455_));
 NAND2x1_ASAP7_75t_R _32036_ (.A(_01565_),
    .B(_02414_),
    .Y(_02456_));
 NOR2x2_ASAP7_75t_R _32037_ (.A(net1241),
    .B(_01561_),
    .Y(_02457_));
 OAI21x1_ASAP7_75t_R _32038_ (.A1(_01526_),
    .A2(_02457_),
    .B(_01565_),
    .Y(_02458_));
 NAND2x1_ASAP7_75t_R _32039_ (.A(_02456_),
    .B(_02458_),
    .Y(_02459_));
 INVx1_ASAP7_75t_R _32040_ (.A(_01496_),
    .Y(_02460_));
 INVx3_ASAP7_75t_R _32041_ (.A(_01612_),
    .Y(_02461_));
 OA21x2_ASAP7_75t_R _32042_ (.A1(_02460_),
    .A2(_02461_),
    .B(_01565_),
    .Y(_02462_));
 NOR3x1_ASAP7_75t_R _32043_ (.A(_02455_),
    .B(_02459_),
    .C(_02462_),
    .Y(_02463_));
 NAND2x1_ASAP7_75t_R _32044_ (.A(_02452_),
    .B(_02463_),
    .Y(_02464_));
 NOR2x1_ASAP7_75t_R _32045_ (.A(_02446_),
    .B(_02464_),
    .Y(_02465_));
 NAND2x1_ASAP7_75t_R _32046_ (.A(_02432_),
    .B(_02465_),
    .Y(_02466_));
 AOI211x1_ASAP7_75t_R _32047_ (.A1(_01538_),
    .A2(net2780),
    .B(_02408_),
    .C(_02466_),
    .Y(_02467_));
 XNOR2x2_ASAP7_75t_R _32048_ (.A(_02357_),
    .B(_02467_),
    .Y(_02468_));
 XOR2x1_ASAP7_75t_R _32049_ (.A(_02249_),
    .Y(_02469_),
    .B(_02468_));
 NAND2x1_ASAP7_75t_R _32050_ (.A(_02469_),
    .B(_02093_),
    .Y(_02470_));
 XOR2x1_ASAP7_75t_R _32051_ (.A(_01483_),
    .Y(_02471_),
    .B(net2041));
 XOR2x2_ASAP7_75t_R _32052_ (.A(_02467_),
    .B(_02357_),
    .Y(_02472_));
 XOR2x1_ASAP7_75t_R _32053_ (.A(_02249_),
    .Y(_02473_),
    .B(_02472_));
 NAND2x1_ASAP7_75t_R _32054_ (.A(_02471_),
    .B(_02473_),
    .Y(_02474_));
 AOI21x1_ASAP7_75t_R _32055_ (.A1(_02470_),
    .A2(_02474_),
    .B(_18753_),
    .Y(_02475_));
 OAI21x1_ASAP7_75t_R _32056_ (.A1(_01998_),
    .A2(_02475_),
    .B(_10171_),
    .Y(_02476_));
 NOR2x1_ASAP7_75t_R _32057_ (.A(net395),
    .B(_00882_),
    .Y(_02477_));
 NAND2x1_ASAP7_75t_R _32058_ (.A(_02471_),
    .B(_02469_),
    .Y(_02478_));
 NAND2x1_ASAP7_75t_R _32059_ (.A(_02093_),
    .B(_02473_),
    .Y(_02479_));
 AOI21x1_ASAP7_75t_R _32060_ (.A1(_02478_),
    .A2(_02479_),
    .B(_18753_),
    .Y(_02480_));
 OAI21x1_ASAP7_75t_R _32061_ (.A1(_02477_),
    .A2(_02480_),
    .B(_00483_),
    .Y(_02481_));
 NAND2x2_ASAP7_75t_R _32062_ (.A(_02481_),
    .B(_02476_),
    .Y(_00114_));
 NOR2x1_ASAP7_75t_R _32063_ (.A(net395),
    .B(_00881_),
    .Y(_02482_));
 NOR2x2_ASAP7_75t_R _32064_ (.A(net3275),
    .B(_01977_),
    .Y(_02483_));
 AOI21x1_ASAP7_75t_R _32065_ (.A1(net2286),
    .A2(net2239),
    .B(_01977_),
    .Y(_02484_));
 NOR2x1_ASAP7_75t_R _32066_ (.A(_02483_),
    .B(_02484_),
    .Y(_02485_));
 TAPCELL_ASAP7_75t_R TAP_561 ();
 AO21x1_ASAP7_75t_R _32068_ (.A1(_02110_),
    .A2(net2175),
    .B(_01977_),
    .Y(_02487_));
 AO21x1_ASAP7_75t_R _32069_ (.A1(net2560),
    .A2(net1527),
    .B(_01977_),
    .Y(_02488_));
 NAND3x1_ASAP7_75t_R _32070_ (.A(_02485_),
    .B(_02487_),
    .C(_02488_),
    .Y(_02489_));
 TAPCELL_ASAP7_75t_R TAP_560 ();
 OA21x2_ASAP7_75t_R _32072_ (.A1(_01890_),
    .A2(_01862_),
    .B(_01970_),
    .Y(_02491_));
 NOR2x1_ASAP7_75t_R _32073_ (.A(_02491_),
    .B(_02217_),
    .Y(_02492_));
 INVx1_ASAP7_75t_R _32074_ (.A(_02103_),
    .Y(_02493_));
 AND2x2_ASAP7_75t_R _32075_ (.A(_02094_),
    .B(_02493_),
    .Y(_02494_));
 NAND2x1_ASAP7_75t_R _32076_ (.A(_02492_),
    .B(_02494_),
    .Y(_02495_));
 NOR2x1_ASAP7_75t_R _32077_ (.A(_02489_),
    .B(_02495_),
    .Y(_02496_));
 AO21x1_ASAP7_75t_R _32078_ (.A1(_01946_),
    .A2(_01832_),
    .B(net3125),
    .Y(_02497_));
 INVx2_ASAP7_75t_R _32079_ (.A(_01949_),
    .Y(_02498_));
 NAND2x1_ASAP7_75t_R _32080_ (.A(_01769_),
    .B(_02498_),
    .Y(_02499_));
 NAND2x2_ASAP7_75t_R _32081_ (.A(net1556),
    .B(_01805_),
    .Y(_02500_));
 INVx1_ASAP7_75t_R _32082_ (.A(_02500_),
    .Y(_02501_));
 NAND2x1_ASAP7_75t_R _32083_ (.A(_02498_),
    .B(_02501_),
    .Y(_02502_));
 NAND3x1_ASAP7_75t_R _32084_ (.A(_02497_),
    .B(_02499_),
    .C(_02502_),
    .Y(_02503_));
 TAPCELL_ASAP7_75t_R TAP_559 ();
 INVx1_ASAP7_75t_R _32086_ (.A(_01958_),
    .Y(_02505_));
 OAI21x1_ASAP7_75t_R _32087_ (.A1(net2352),
    .A2(_02225_),
    .B(_02505_),
    .Y(_02506_));
 AO21x1_ASAP7_75t_R _32088_ (.A1(net2619),
    .A2(_01795_),
    .B(net2352),
    .Y(_02507_));
 AO21x1_ASAP7_75t_R _32089_ (.A1(_01799_),
    .A2(net1138),
    .B(net2352),
    .Y(_02508_));
 NAND2x1_ASAP7_75t_R _32090_ (.A(_02507_),
    .B(_02508_),
    .Y(_02509_));
 NOR3x1_ASAP7_75t_R _32091_ (.A(_02503_),
    .B(_02506_),
    .C(_02509_),
    .Y(_02510_));
 NAND2x1_ASAP7_75t_R _32092_ (.A(_02496_),
    .B(_02510_),
    .Y(_02511_));
 AOI211x1_ASAP7_75t_R _32093_ (.A1(_01770_),
    .A2(_01776_),
    .B(net2140),
    .C(_01870_),
    .Y(_02512_));
 INVx1_ASAP7_75t_R _32094_ (.A(_02512_),
    .Y(_02513_));
 AO21x1_ASAP7_75t_R _32095_ (.A1(_02110_),
    .A2(net1157),
    .B(net2140),
    .Y(_02514_));
 AO21x1_ASAP7_75t_R _32096_ (.A1(net2307),
    .A2(_01837_),
    .B(net2140),
    .Y(_02515_));
 NAND3x1_ASAP7_75t_R _32097_ (.A(_02513_),
    .B(_02514_),
    .C(_02515_),
    .Y(_02516_));
 NAND2x1_ASAP7_75t_R _32098_ (.A(_01904_),
    .B(_02114_),
    .Y(_02517_));
 NAND2x1_ASAP7_75t_R _32099_ (.A(_01904_),
    .B(_02124_),
    .Y(_02518_));
 NAND2x1_ASAP7_75t_R _32100_ (.A(net1465),
    .B(_01904_),
    .Y(_02519_));
 AND3x1_ASAP7_75t_R _32101_ (.A(_02517_),
    .B(_02518_),
    .C(_02519_),
    .Y(_02520_));
 NOR2x1_ASAP7_75t_R _32102_ (.A(_02500_),
    .B(_01905_),
    .Y(_02521_));
 NAND2x1_ASAP7_75t_R _32103_ (.A(_01904_),
    .B(_01806_),
    .Y(_02522_));
 OAI21x1_ASAP7_75t_R _32104_ (.A1(net2175),
    .A2(_01905_),
    .B(_02522_),
    .Y(_02523_));
 NOR2x1_ASAP7_75t_R _32105_ (.A(_02521_),
    .B(_02523_),
    .Y(_02524_));
 NAND2x1_ASAP7_75t_R _32106_ (.A(_02520_),
    .B(_02524_),
    .Y(_02525_));
 NOR2x1_ASAP7_75t_R _32107_ (.A(_02516_),
    .B(_02525_),
    .Y(_02526_));
 AOI211x1_ASAP7_75t_R _32108_ (.A1(net1116),
    .A2(net1456),
    .B(net2194),
    .C(_01857_),
    .Y(_02527_));
 INVx1_ASAP7_75t_R _32109_ (.A(_02527_),
    .Y(_02528_));
 AO21x1_ASAP7_75t_R _32110_ (.A1(net2560),
    .A2(_01935_),
    .B(net2194),
    .Y(_02529_));
 TAPCELL_ASAP7_75t_R TAP_558 ();
 AO21x1_ASAP7_75t_R _32112_ (.A1(net1253),
    .A2(_01821_),
    .B(net2194),
    .Y(_02531_));
 NAND3x1_ASAP7_75t_R _32113_ (.A(_02528_),
    .B(_02529_),
    .C(_02531_),
    .Y(_02532_));
 AO21x1_ASAP7_75t_R _32114_ (.A1(net1253),
    .A2(net2286),
    .B(net2549),
    .Y(_02533_));
 AND2x2_ASAP7_75t_R _32115_ (.A(_02533_),
    .B(_02186_),
    .Y(_02534_));
 NOR2x2_ASAP7_75t_R _32116_ (.A(net1299),
    .B(net2215),
    .Y(_02535_));
 NOR2x1_ASAP7_75t_R _32117_ (.A(net2384),
    .B(_01824_),
    .Y(_02536_));
 NOR2x1_ASAP7_75t_R _32118_ (.A(net2384),
    .B(net3254),
    .Y(_02537_));
 AOI211x1_ASAP7_75t_R _32119_ (.A1(_02535_),
    .A2(net950),
    .B(_02536_),
    .C(_02537_),
    .Y(_02538_));
 NAND2x1_ASAP7_75t_R _32120_ (.A(_02534_),
    .B(_02538_),
    .Y(_02539_));
 NOR2x1_ASAP7_75t_R _32121_ (.A(_02532_),
    .B(_02539_),
    .Y(_02540_));
 NAND2x1_ASAP7_75t_R _32122_ (.A(_02526_),
    .B(_02540_),
    .Y(_02541_));
 NOR2x1_ASAP7_75t_R _32123_ (.A(_02511_),
    .B(_02541_),
    .Y(_02542_));
 AO21x1_ASAP7_75t_R _32124_ (.A1(net2306),
    .A2(net2372),
    .B(net2458),
    .Y(_02543_));
 NOR2x2_ASAP7_75t_R _32125_ (.A(_01870_),
    .B(_01786_),
    .Y(_02544_));
 NAND2x1_ASAP7_75t_R _32126_ (.A(_02544_),
    .B(_01888_),
    .Y(_02545_));
 AND2x2_ASAP7_75t_R _32127_ (.A(_02543_),
    .B(_02545_),
    .Y(_02546_));
 NOR2x1_ASAP7_75t_R _32128_ (.A(_01850_),
    .B(net3128),
    .Y(_02547_));
 NOR2x1_ASAP7_75t_R _32129_ (.A(_01894_),
    .B(_01832_),
    .Y(_02548_));
 NOR2x1_ASAP7_75t_R _32130_ (.A(_01894_),
    .B(_01831_),
    .Y(_02549_));
 AOI211x1_ASAP7_75t_R _32131_ (.A1(_02547_),
    .A2(net952),
    .B(_02548_),
    .C(_02549_),
    .Y(_02550_));
 NAND2x1_ASAP7_75t_R _32132_ (.A(_02546_),
    .B(_02550_),
    .Y(_02551_));
 AO31x2_ASAP7_75t_R _32133_ (.A1(_02110_),
    .A2(_01877_),
    .A3(_01832_),
    .B(_01878_),
    .Y(_02552_));
 AOI211x1_ASAP7_75t_R _32134_ (.A1(net1116),
    .A2(_01776_),
    .B(_01878_),
    .C(_01857_),
    .Y(_02553_));
 INVx1_ASAP7_75t_R _32135_ (.A(_02553_),
    .Y(_02554_));
 NAND2x1_ASAP7_75t_R _32136_ (.A(_01876_),
    .B(_02177_),
    .Y(_02555_));
 NAND3x1_ASAP7_75t_R _32137_ (.A(_02552_),
    .B(_02554_),
    .C(_02555_),
    .Y(_02556_));
 NOR2x1_ASAP7_75t_R _32138_ (.A(_02551_),
    .B(_02556_),
    .Y(_02557_));
 AO21x1_ASAP7_75t_R _32139_ (.A1(net1527),
    .A2(_01934_),
    .B(_01863_),
    .Y(_02558_));
 NAND2x2_ASAP7_75t_R _32140_ (.A(_01770_),
    .B(net1127),
    .Y(_02559_));
 AO21x1_ASAP7_75t_R _32141_ (.A1(net1138),
    .A2(_02559_),
    .B(_01863_),
    .Y(_02560_));
 AND2x2_ASAP7_75t_R _32142_ (.A(_02558_),
    .B(_02560_),
    .Y(_02561_));
 NAND2x1_ASAP7_75t_R _32143_ (.A(net2330),
    .B(_01847_),
    .Y(_02562_));
 OA21x2_ASAP7_75t_R _32144_ (.A1(_02544_),
    .A2(_01882_),
    .B(_01847_),
    .Y(_02563_));
 NOR2x1_ASAP7_75t_R _32145_ (.A(_02563_),
    .B(_01859_),
    .Y(_02564_));
 AND3x1_ASAP7_75t_R _32146_ (.A(_02561_),
    .B(_02562_),
    .C(_02564_),
    .Y(_02565_));
 NAND2x1_ASAP7_75t_R _32147_ (.A(_02557_),
    .B(_02565_),
    .Y(_02566_));
 AO21x1_ASAP7_75t_R _32148_ (.A1(_01799_),
    .A2(_01857_),
    .B(_01828_),
    .Y(_02567_));
 AO21x1_ASAP7_75t_R _32149_ (.A1(_01946_),
    .A2(_01934_),
    .B(_01828_),
    .Y(_02568_));
 NAND2x1_ASAP7_75t_R _32150_ (.A(_02567_),
    .B(_02568_),
    .Y(_02569_));
 AO21x1_ASAP7_75t_R _32151_ (.A1(net1253),
    .A2(net2219),
    .B(_01809_),
    .Y(_02570_));
 AO21x1_ASAP7_75t_R _32152_ (.A1(_01946_),
    .A2(_01790_),
    .B(_01809_),
    .Y(_02571_));
 NAND2x1_ASAP7_75t_R _32153_ (.A(_01855_),
    .B(_01810_),
    .Y(_02572_));
 NAND3x1_ASAP7_75t_R _32154_ (.A(_02570_),
    .B(_02571_),
    .C(_02572_),
    .Y(_02573_));
 NOR2x1_ASAP7_75t_R _32155_ (.A(_02569_),
    .B(_02573_),
    .Y(_02574_));
 AO21x1_ASAP7_75t_R _32156_ (.A1(net2175),
    .A2(_02100_),
    .B(_01761_),
    .Y(_02575_));
 AO21x1_ASAP7_75t_R _32157_ (.A1(net1138),
    .A2(_01799_),
    .B(_01761_),
    .Y(_02576_));
 NAND2x1_ASAP7_75t_R _32158_ (.A(_01816_),
    .B(_01762_),
    .Y(_02577_));
 AND3x1_ASAP7_75t_R _32159_ (.A(_02575_),
    .B(_02576_),
    .C(_02577_),
    .Y(_02578_));
 NAND2x1_ASAP7_75t_R _32160_ (.A(net1451),
    .B(_01830_),
    .Y(_02579_));
 TAPCELL_ASAP7_75t_R TAP_557 ();
 AO21x1_ASAP7_75t_R _32162_ (.A1(net1527),
    .A2(_02579_),
    .B(_01781_),
    .Y(_02581_));
 AO21x1_ASAP7_75t_R _32163_ (.A1(_01821_),
    .A2(net1138),
    .B(_01781_),
    .Y(_02582_));
 AO21x1_ASAP7_75t_R _32164_ (.A1(net2619),
    .A2(_01908_),
    .B(_01781_),
    .Y(_02583_));
 AND3x1_ASAP7_75t_R _32165_ (.A(_02581_),
    .B(_02582_),
    .C(_02583_),
    .Y(_02584_));
 NAND3x1_ASAP7_75t_R _32166_ (.A(_02574_),
    .B(_02578_),
    .C(_02584_),
    .Y(_02585_));
 NOR2x1_ASAP7_75t_R _32167_ (.A(_02566_),
    .B(_02585_),
    .Y(_02586_));
 NAND2x1_ASAP7_75t_R _32168_ (.A(_02542_),
    .B(_02586_),
    .Y(_02587_));
 NOR2x2_ASAP7_75t_R _32169_ (.A(_02107_),
    .B(_02587_),
    .Y(_02588_));
 INVx2_ASAP7_75t_R _32170_ (.A(_02588_),
    .Y(_02589_));
 AO21x1_ASAP7_75t_R _32171_ (.A1(net2651),
    .A2(_01226_),
    .B(_01133_),
    .Y(_02590_));
 AO21x1_ASAP7_75t_R _32172_ (.A1(_01348_),
    .A2(net1697),
    .B(_01133_),
    .Y(_02591_));
 INVx1_ASAP7_75t_R _32173_ (.A(_01153_),
    .Y(_02592_));
 INVx2_ASAP7_75t_R _32174_ (.A(_01133_),
    .Y(_02593_));
 NAND2x1_ASAP7_75t_R _32175_ (.A(_02592_),
    .B(_02593_),
    .Y(_02594_));
 AND3x1_ASAP7_75t_R _32176_ (.A(_02590_),
    .B(_02591_),
    .C(_02594_),
    .Y(_02595_));
 AO21x1_ASAP7_75t_R _32177_ (.A1(_01306_),
    .A2(_01226_),
    .B(_01120_),
    .Y(_02596_));
 AO21x1_ASAP7_75t_R _32178_ (.A1(_01153_),
    .A2(_01221_),
    .B(_01120_),
    .Y(_02597_));
 AND3x1_ASAP7_75t_R _32179_ (.A(_02596_),
    .B(_02597_),
    .C(_01107_),
    .Y(_02598_));
 AND2x2_ASAP7_75t_R _32180_ (.A(_02595_),
    .B(_02598_),
    .Y(_02599_));
 INVx2_ASAP7_75t_R _32181_ (.A(_01125_),
    .Y(_02600_));
 OA21x2_ASAP7_75t_R _32182_ (.A1(_02600_),
    .A2(_01233_),
    .B(_01163_),
    .Y(_02601_));
 AND3x1_ASAP7_75t_R _32183_ (.A(_01163_),
    .B(_01187_),
    .C(net1136),
    .Y(_02602_));
 TAPCELL_ASAP7_75t_R TAP_556 ();
 NOR2x1_ASAP7_75t_R _32185_ (.A(net1802),
    .B(_01156_),
    .Y(_02604_));
 OR3x1_ASAP7_75t_R _32186_ (.A(_02601_),
    .B(_02602_),
    .C(_02604_),
    .Y(_02605_));
 OA21x2_ASAP7_75t_R _32187_ (.A1(_01268_),
    .A2(_01180_),
    .B(_01171_),
    .Y(_02606_));
 NOR2x1_ASAP7_75t_R _32188_ (.A(_01177_),
    .B(_02606_),
    .Y(_02607_));
 TAPCELL_ASAP7_75t_R TAP_555 ();
 AO21x1_ASAP7_75t_R _32190_ (.A1(net1752),
    .A2(_01252_),
    .B(_01170_),
    .Y(_02609_));
 AO21x1_ASAP7_75t_R _32191_ (.A1(net2723),
    .A2(net1572),
    .B(_01170_),
    .Y(_02610_));
 NAND2x1_ASAP7_75t_R _32192_ (.A(_02023_),
    .B(_01171_),
    .Y(_02611_));
 AND3x1_ASAP7_75t_R _32193_ (.A(_02609_),
    .B(_02610_),
    .C(_02611_),
    .Y(_02612_));
 NAND2x1_ASAP7_75t_R _32194_ (.A(_02607_),
    .B(_02612_),
    .Y(_02613_));
 NOR2x1_ASAP7_75t_R _32195_ (.A(_02605_),
    .B(_02613_),
    .Y(_02614_));
 NAND2x1_ASAP7_75t_R _32196_ (.A(_02599_),
    .B(_02614_),
    .Y(_02615_));
 OA21x2_ASAP7_75t_R _32197_ (.A1(_01179_),
    .A2(_01268_),
    .B(_01234_),
    .Y(_02616_));
 OA21x2_ASAP7_75t_R _32198_ (.A1(_01328_),
    .A2(_02023_),
    .B(_01234_),
    .Y(_02617_));
 OR3x1_ASAP7_75t_R _32199_ (.A(_02616_),
    .B(_02617_),
    .C(_01448_),
    .Y(_02618_));
 INVx2_ASAP7_75t_R _32200_ (.A(net1827),
    .Y(_02619_));
 NAND2x1_ASAP7_75t_R _32201_ (.A(_01218_),
    .B(_02619_),
    .Y(_02620_));
 AO21x1_ASAP7_75t_R _32202_ (.A1(net1294),
    .A2(_01128_),
    .B(_01215_),
    .Y(_02621_));
 NAND2x1_ASAP7_75t_R _32203_ (.A(_02620_),
    .B(_02621_),
    .Y(_02622_));
 INVx2_ASAP7_75t_R _32204_ (.A(_01279_),
    .Y(_02623_));
 AND2x2_ASAP7_75t_R _32205_ (.A(_01216_),
    .B(_02623_),
    .Y(_02624_));
 OR3x1_ASAP7_75t_R _32206_ (.A(_02622_),
    .B(_01451_),
    .C(_02624_),
    .Y(_02625_));
 NOR2x1_ASAP7_75t_R _32207_ (.A(_02618_),
    .B(_02625_),
    .Y(_02626_));
 AO21x1_ASAP7_75t_R _32208_ (.A1(net2522),
    .A2(_01384_),
    .B(net3144),
    .Y(_02627_));
 AO21x1_ASAP7_75t_R _32209_ (.A1(net2723),
    .A2(_01259_),
    .B(net3144),
    .Y(_02628_));
 AND2x2_ASAP7_75t_R _32210_ (.A(_02627_),
    .B(_02628_),
    .Y(_02629_));
 AO21x1_ASAP7_75t_R _32211_ (.A1(net2121),
    .A2(net2731),
    .B(_01191_),
    .Y(_02630_));
 AO21x1_ASAP7_75t_R _32212_ (.A1(net1275),
    .A2(_01226_),
    .B(_01191_),
    .Y(_02631_));
 NAND2x1_ASAP7_75t_R _32213_ (.A(_01405_),
    .B(_01197_),
    .Y(_02632_));
 AND3x1_ASAP7_75t_R _32214_ (.A(_02630_),
    .B(_02631_),
    .C(_02632_),
    .Y(_02633_));
 NAND2x1_ASAP7_75t_R _32215_ (.A(_02629_),
    .B(_02633_),
    .Y(_02634_));
 NAND2x2_ASAP7_75t_R _32216_ (.A(_01233_),
    .B(_01210_),
    .Y(_02635_));
 AO21x1_ASAP7_75t_R _32217_ (.A1(net3322),
    .A2(net1827),
    .B(_01202_),
    .Y(_02636_));
 NAND2x1_ASAP7_75t_R _32218_ (.A(_02636_),
    .B(_02635_),
    .Y(_02637_));
 TAPCELL_ASAP7_75t_R TAP_554 ();
 AO21x1_ASAP7_75t_R _32220_ (.A1(net1275),
    .A2(_01226_),
    .B(_01202_),
    .Y(_02639_));
 INVx1_ASAP7_75t_R _32221_ (.A(_02639_),
    .Y(_02640_));
 NOR2x1_ASAP7_75t_R _32222_ (.A(net1918),
    .B(net3154),
    .Y(_02641_));
 OR3x1_ASAP7_75t_R _32223_ (.A(_02637_),
    .B(_02640_),
    .C(_02641_),
    .Y(_02642_));
 NOR2x2_ASAP7_75t_R _32224_ (.A(_02634_),
    .B(_02642_),
    .Y(_02643_));
 NAND2x2_ASAP7_75t_R _32225_ (.A(_02643_),
    .B(_02626_),
    .Y(_02644_));
 NOR2x2_ASAP7_75t_R _32226_ (.A(_02615_),
    .B(_02644_),
    .Y(_02645_));
 OAI21x1_ASAP7_75t_R _32227_ (.A1(net3315),
    .A2(_01228_),
    .B(_01412_),
    .Y(_02646_));
 AO21x1_ASAP7_75t_R _32228_ (.A1(net1803),
    .A2(_01348_),
    .B(net3316),
    .Y(_02647_));
 OAI21x1_ASAP7_75t_R _32229_ (.A1(net1122),
    .A2(net3316),
    .B(_02647_),
    .Y(_02648_));
 NOR2x2_ASAP7_75t_R _32230_ (.A(_01321_),
    .B(net3316),
    .Y(_02649_));
 NOR3x2_ASAP7_75t_R _32231_ (.B(_02648_),
    .C(_02649_),
    .Y(_02650_),
    .A(_02646_));
 TAPCELL_ASAP7_75t_R TAP_553 ();
 AO21x1_ASAP7_75t_R _32233_ (.A1(_01113_),
    .A2(_01138_),
    .B(_01243_),
    .Y(_02652_));
 TAPCELL_ASAP7_75t_R TAP_552 ();
 TAPCELL_ASAP7_75t_R PHY_551 ();
 AO21x1_ASAP7_75t_R _32236_ (.A1(net2122),
    .A2(_01188_),
    .B(_01243_),
    .Y(_02655_));
 AO21x1_ASAP7_75t_R _32237_ (.A1(_01194_),
    .A2(net3341),
    .B(_01243_),
    .Y(_02656_));
 AND4x2_ASAP7_75t_R _32238_ (.A(_02652_),
    .B(_02655_),
    .C(_02656_),
    .D(_01254_),
    .Y(_02657_));
 AO21x1_ASAP7_75t_R _32239_ (.A1(net2120),
    .A2(_01226_),
    .B(net3417),
    .Y(_02658_));
 AO21x1_ASAP7_75t_R _32240_ (.A1(_01348_),
    .A2(net1698),
    .B(net3417),
    .Y(_02659_));
 NAND3x2_ASAP7_75t_R _32241_ (.B(_01415_),
    .C(_02659_),
    .Y(_02660_),
    .A(_02658_));
 TAPCELL_ASAP7_75t_R PHY_550 ();
 TAPCELL_ASAP7_75t_R PHY_549 ();
 AO21x1_ASAP7_75t_R _32244_ (.A1(net2120),
    .A2(net1142),
    .B(net3145),
    .Y(_02663_));
 AO21x1_ASAP7_75t_R _32245_ (.A1(net1274),
    .A2(_01138_),
    .B(net3145),
    .Y(_02664_));
 AO21x2_ASAP7_75t_R _32246_ (.A1(net1803),
    .A2(_01447_),
    .B(_01287_),
    .Y(_02665_));
 NAND3x2_ASAP7_75t_R _32247_ (.B(_02664_),
    .C(_02665_),
    .Y(_02666_),
    .A(_02663_));
 NOR2x2_ASAP7_75t_R _32248_ (.A(_02660_),
    .B(_02666_),
    .Y(_02667_));
 NAND3x2_ASAP7_75t_R _32249_ (.B(_02657_),
    .C(_02667_),
    .Y(_02668_),
    .A(_02650_));
 TAPCELL_ASAP7_75t_R PHY_548 ();
 AO21x1_ASAP7_75t_R _32251_ (.A1(net2361),
    .A2(net1142),
    .B(_01345_),
    .Y(_02670_));
 OA21x2_ASAP7_75t_R _32252_ (.A1(_01345_),
    .A2(_01138_),
    .B(_02670_),
    .Y(_02671_));
 AO21x1_ASAP7_75t_R _32253_ (.A1(net1866),
    .A2(net940),
    .B(net3240),
    .Y(_02672_));
 AO21x1_ASAP7_75t_R _32254_ (.A1(net1572),
    .A2(net1076),
    .B(net3240),
    .Y(_02673_));
 AND3x2_ASAP7_75t_R _32255_ (.A(_02671_),
    .B(_02672_),
    .C(_02673_),
    .Y(_02674_));
 AO21x1_ASAP7_75t_R _32256_ (.A1(net1802),
    .A2(_01259_),
    .B(_01308_),
    .Y(_02675_));
 NOR2x1_ASAP7_75t_R _32257_ (.A(net2651),
    .B(_01308_),
    .Y(_02676_));
 INVx1_ASAP7_75t_R _32258_ (.A(_02676_),
    .Y(_02677_));
 NOR2x1_ASAP7_75t_R _32259_ (.A(net2361),
    .B(_01308_),
    .Y(_02678_));
 INVx1_ASAP7_75t_R _32260_ (.A(_02678_),
    .Y(_02679_));
 AND3x1_ASAP7_75t_R _32261_ (.A(_02675_),
    .B(_02677_),
    .C(_02679_),
    .Y(_02680_));
 AO21x1_ASAP7_75t_R _32262_ (.A1(net2361),
    .A2(_01226_),
    .B(_01322_),
    .Y(_02681_));
 AO21x1_ASAP7_75t_R _32263_ (.A1(net1293),
    .A2(net3341),
    .B(_01322_),
    .Y(_02682_));
 INVx1_ASAP7_75t_R _32264_ (.A(_01397_),
    .Y(_02683_));
 AND3x1_ASAP7_75t_R _32265_ (.A(_02681_),
    .B(_02682_),
    .C(_02683_),
    .Y(_02684_));
 AND2x2_ASAP7_75t_R _32266_ (.A(_02680_),
    .B(_02684_),
    .Y(_02685_));
 AO21x1_ASAP7_75t_R _32267_ (.A1(net1266),
    .A2(net938),
    .B(_01334_),
    .Y(_02686_));
 AO21x1_ASAP7_75t_R _32268_ (.A1(_01348_),
    .A2(net1076),
    .B(_01334_),
    .Y(_02687_));
 NAND2x1_ASAP7_75t_R _32269_ (.A(_01406_),
    .B(_01337_),
    .Y(_02688_));
 AND3x2_ASAP7_75t_R _32270_ (.A(_02686_),
    .B(_02687_),
    .C(_02688_),
    .Y(_02689_));
 NAND3x2_ASAP7_75t_R _32271_ (.B(_02685_),
    .C(_02689_),
    .Y(_02690_),
    .A(_02674_));
 NOR2x2_ASAP7_75t_R _32272_ (.A(_02668_),
    .B(_02690_),
    .Y(_02691_));
 NAND2x2_ASAP7_75t_R _32273_ (.A(_02645_),
    .B(_02691_),
    .Y(_02692_));
 NAND2x1_ASAP7_75t_R _32274_ (.A(_02316_),
    .B(_22092_),
    .Y(_02693_));
 AO21x1_ASAP7_75t_R _32275_ (.A1(net991),
    .A2(_02273_),
    .B(_22091_),
    .Y(_02694_));
 NAND2x1_ASAP7_75t_R _32276_ (.A(_02693_),
    .B(_02694_),
    .Y(_02695_));
 NAND2x1_ASAP7_75t_R _32277_ (.A(_22054_),
    .B(_22092_),
    .Y(_02696_));
 AO21x1_ASAP7_75t_R _32278_ (.A1(_22076_),
    .A2(net3280),
    .B(_22091_),
    .Y(_02697_));
 NAND2x1_ASAP7_75t_R _32279_ (.A(_02696_),
    .B(_02697_),
    .Y(_02698_));
 NOR2x1_ASAP7_75t_R _32280_ (.A(_02695_),
    .B(_02698_),
    .Y(_02699_));
 TAPCELL_ASAP7_75t_R PHY_547 ();
 AO21x1_ASAP7_75t_R _32282_ (.A1(net1038),
    .A2(net2365),
    .B(net3081),
    .Y(_02701_));
 TAPCELL_ASAP7_75t_R PHY_546 ();
 AO21x1_ASAP7_75t_R _32284_ (.A1(net1048),
    .A2(net1792),
    .B(net3081),
    .Y(_02703_));
 OR2x2_ASAP7_75t_R _32285_ (.A(_22057_),
    .B(net3081),
    .Y(_02704_));
 AND3x1_ASAP7_75t_R _32286_ (.A(_02701_),
    .B(_02703_),
    .C(_02704_),
    .Y(_02705_));
 NAND2x1_ASAP7_75t_R _32287_ (.A(_02699_),
    .B(_02705_),
    .Y(_02706_));
 TAPCELL_ASAP7_75t_R PHY_545 ();
 AO21x1_ASAP7_75t_R _32289_ (.A1(net1048),
    .A2(net1792),
    .B(net3143),
    .Y(_02708_));
 AO21x1_ASAP7_75t_R _32290_ (.A1(_22024_),
    .A2(_21944_),
    .B(net3143),
    .Y(_02709_));
 NAND2x1_ASAP7_75t_R _32291_ (.A(_02708_),
    .B(_02709_),
    .Y(_02710_));
 AO21x1_ASAP7_75t_R _32292_ (.A1(_21967_),
    .A2(_21969_),
    .B(net3152),
    .Y(_02711_));
 AO21x1_ASAP7_75t_R _32293_ (.A1(net2265),
    .A2(net2365),
    .B(net3143),
    .Y(_02712_));
 NAND2x1_ASAP7_75t_R _32294_ (.A(_02711_),
    .B(_02712_),
    .Y(_02713_));
 NOR2x1_ASAP7_75t_R _32295_ (.A(net2005),
    .B(_21877_),
    .Y(_02714_));
 OAI21x1_ASAP7_75t_R _32296_ (.A1(_02316_),
    .A2(_02714_),
    .B(_01073_),
    .Y(_02715_));
 AO21x1_ASAP7_75t_R _32297_ (.A1(_21944_),
    .A2(net1848),
    .B(_01072_),
    .Y(_02716_));
 NAND2x1_ASAP7_75t_R _32298_ (.A(_02715_),
    .B(_02716_),
    .Y(_02717_));
 OR3x1_ASAP7_75t_R _32299_ (.A(_02710_),
    .B(_02713_),
    .C(_02717_),
    .Y(_02718_));
 NOR2x2_ASAP7_75t_R _32300_ (.A(_02706_),
    .B(_02718_),
    .Y(_02719_));
 AO21x1_ASAP7_75t_R _32301_ (.A1(_21890_),
    .A2(_22008_),
    .B(_22077_),
    .Y(_02720_));
 NAND2x1_ASAP7_75t_R _32302_ (.A(_22084_),
    .B(_02286_),
    .Y(_02721_));
 NOR2x2_ASAP7_75t_R _32303_ (.A(net1046),
    .B(net2427),
    .Y(_02722_));
 NAND2x1_ASAP7_75t_R _32304_ (.A(_22084_),
    .B(_02722_),
    .Y(_02723_));
 AND4x1_ASAP7_75t_R _32305_ (.A(_02720_),
    .B(_02721_),
    .C(_02295_),
    .D(_02723_),
    .Y(_02724_));
 TAPCELL_ASAP7_75t_R PHY_544 ();
 AO21x1_ASAP7_75t_R _32307_ (.A1(net2752),
    .A2(net991),
    .B(_22070_),
    .Y(_02726_));
 AO21x1_ASAP7_75t_R _32308_ (.A1(net2510),
    .A2(_22019_),
    .B(_22070_),
    .Y(_02727_));
 NAND2x1_ASAP7_75t_R _32309_ (.A(_21908_),
    .B(_02292_),
    .Y(_02728_));
 AND3x1_ASAP7_75t_R _32310_ (.A(_02726_),
    .B(_02727_),
    .C(_02728_),
    .Y(_02729_));
 AND2x2_ASAP7_75t_R _32311_ (.A(_02724_),
    .B(_02729_),
    .Y(_02730_));
 TAPCELL_ASAP7_75t_R PHY_543 ();
 AO21x1_ASAP7_75t_R _32313_ (.A1(net991),
    .A2(net2420),
    .B(_22061_),
    .Y(_02732_));
 OA21x2_ASAP7_75t_R _32314_ (.A1(net1038),
    .A2(_22061_),
    .B(_02732_),
    .Y(_02733_));
 OA211x2_ASAP7_75t_R _32315_ (.A1(_21887_),
    .A2(_21876_),
    .B(_22062_),
    .C(net1926),
    .Y(_02734_));
 INVx1_ASAP7_75t_R _32316_ (.A(_02734_),
    .Y(_02735_));
 NAND2x1_ASAP7_75t_R _32317_ (.A(_02733_),
    .B(_02735_),
    .Y(_02736_));
 AO21x1_ASAP7_75t_R _32318_ (.A1(net1048),
    .A2(_22080_),
    .B(_22064_),
    .Y(_02737_));
 AND2x2_ASAP7_75t_R _32319_ (.A(_02737_),
    .B(_22051_),
    .Y(_02738_));
 AO21x1_ASAP7_75t_R _32320_ (.A1(net2365),
    .A2(_21983_),
    .B(_22064_),
    .Y(_02739_));
 AO21x1_ASAP7_75t_R _32321_ (.A1(_21967_),
    .A2(net2420),
    .B(_22064_),
    .Y(_02740_));
 NAND2x1_ASAP7_75t_R _32322_ (.A(_01082_),
    .B(_22049_),
    .Y(_02741_));
 AND3x1_ASAP7_75t_R _32323_ (.A(_02739_),
    .B(_02740_),
    .C(_02741_),
    .Y(_02742_));
 NAND2x1_ASAP7_75t_R _32324_ (.A(_02738_),
    .B(_02742_),
    .Y(_02743_));
 NOR2x2_ASAP7_75t_R _32325_ (.A(_02736_),
    .B(_02743_),
    .Y(_02744_));
 NAND3x2_ASAP7_75t_R _32326_ (.B(_02730_),
    .C(_02744_),
    .Y(_02745_),
    .A(_02719_));
 AO21x1_ASAP7_75t_R _32327_ (.A1(net991),
    .A2(_22019_),
    .B(net2556),
    .Y(_02746_));
 NAND2x2_ASAP7_75t_R _32328_ (.A(net2802),
    .B(_22034_),
    .Y(_02747_));
 AND3x2_ASAP7_75t_R _32329_ (.A(_02746_),
    .B(_22035_),
    .C(_02747_),
    .Y(_02748_));
 AO21x1_ASAP7_75t_R _32330_ (.A1(_02312_),
    .A2(_22024_),
    .B(net2512),
    .Y(_02749_));
 AO21x1_ASAP7_75t_R _32331_ (.A1(_21983_),
    .A2(net2337),
    .B(net2512),
    .Y(_02750_));
 AO21x1_ASAP7_75t_R _32332_ (.A1(net991),
    .A2(net2420),
    .B(net2512),
    .Y(_02751_));
 AND2x2_ASAP7_75t_R _32333_ (.A(_02750_),
    .B(_02751_),
    .Y(_02752_));
 NAND3x2_ASAP7_75t_R _32334_ (.B(_02749_),
    .C(_02752_),
    .Y(_02753_),
    .A(_02748_));
 AO21x1_ASAP7_75t_R _32335_ (.A1(net3172),
    .A2(_21929_),
    .B(net3148),
    .Y(_02754_));
 AO21x1_ASAP7_75t_R _32336_ (.A1(net2267),
    .A2(_21969_),
    .B(net3148),
    .Y(_02755_));
 AND2x2_ASAP7_75t_R _32337_ (.A(_02754_),
    .B(_02755_),
    .Y(_02756_));
 AO21x1_ASAP7_75t_R _32338_ (.A1(net3172),
    .A2(net3280),
    .B(net3151),
    .Y(_02757_));
 INVx3_ASAP7_75t_R _32339_ (.A(_21992_),
    .Y(_02758_));
 NOR2x1_ASAP7_75t_R _32340_ (.A(net2267),
    .B(_21992_),
    .Y(_02759_));
 NOR2x1_ASAP7_75t_R _32341_ (.A(_02273_),
    .B(_21992_),
    .Y(_02760_));
 AOI211x1_ASAP7_75t_R _32342_ (.A1(_01087_),
    .A2(_02758_),
    .B(_02759_),
    .C(_02760_),
    .Y(_02761_));
 AND3x1_ASAP7_75t_R _32343_ (.A(_02756_),
    .B(_02757_),
    .C(_02761_),
    .Y(_02762_));
 INVx1_ASAP7_75t_R _32344_ (.A(_02762_),
    .Y(_02763_));
 NOR2x2_ASAP7_75t_R _32345_ (.A(_02753_),
    .B(_02763_),
    .Y(_02764_));
 INVx1_ASAP7_75t_R _32346_ (.A(_02273_),
    .Y(_02765_));
 OA211x2_ASAP7_75t_R _32347_ (.A1(net1139),
    .A2(net1049),
    .B(_21957_),
    .C(_21889_),
    .Y(_02766_));
 OA21x2_ASAP7_75t_R _32348_ (.A1(_02722_),
    .A2(net2589),
    .B(_21957_),
    .Y(_02767_));
 AOI211x1_ASAP7_75t_R _32349_ (.A1(_02765_),
    .A2(_21957_),
    .B(_02766_),
    .C(_02767_),
    .Y(_02768_));
 AO21x1_ASAP7_75t_R _32350_ (.A1(net1630),
    .A2(_21927_),
    .B(_21901_),
    .Y(_02769_));
 AO21x1_ASAP7_75t_R _32351_ (.A1(_21967_),
    .A2(net2258),
    .B(_21901_),
    .Y(_02770_));
 AO21x1_ASAP7_75t_R _32352_ (.A1(_22018_),
    .A2(_22019_),
    .B(_21901_),
    .Y(_02771_));
 NAND3x2_ASAP7_75t_R _32353_ (.B(_02770_),
    .C(_02771_),
    .Y(_02772_),
    .A(_02769_));
 AO21x1_ASAP7_75t_R _32354_ (.A1(_22024_),
    .A2(_21929_),
    .B(net2495),
    .Y(_02773_));
 AO21x2_ASAP7_75t_R _32355_ (.A1(_02259_),
    .A2(_22057_),
    .B(_21893_),
    .Y(_02774_));
 AO21x1_ASAP7_75t_R _32356_ (.A1(net1048),
    .A2(net1792),
    .B(_21893_),
    .Y(_02775_));
 NAND3x2_ASAP7_75t_R _32357_ (.B(_02774_),
    .C(_02775_),
    .Y(_02776_),
    .A(_02773_));
 NOR2x2_ASAP7_75t_R _32358_ (.A(_02772_),
    .B(_02776_),
    .Y(_02777_));
 AO21x1_ASAP7_75t_R _32359_ (.A1(_21877_),
    .A2(_21954_),
    .B(_21904_),
    .Y(_02778_));
 AO21x1_ASAP7_75t_R _32360_ (.A1(_02778_),
    .A2(_21995_),
    .B(_21976_),
    .Y(_02779_));
 INVx1_ASAP7_75t_R _32361_ (.A(_21985_),
    .Y(_02780_));
 AO21x1_ASAP7_75t_R _32362_ (.A1(net991),
    .A2(_02273_),
    .B(_21976_),
    .Y(_02781_));
 AND3x2_ASAP7_75t_R _32363_ (.A(_02779_),
    .B(_02780_),
    .C(_02781_),
    .Y(_02782_));
 NAND3x2_ASAP7_75t_R _32364_ (.B(_02777_),
    .C(_02782_),
    .Y(_02783_),
    .A(_02768_));
 INVx1_ASAP7_75t_R _32365_ (.A(_02783_),
    .Y(_02784_));
 NAND2x2_ASAP7_75t_R _32366_ (.A(_02764_),
    .B(_02784_),
    .Y(_02785_));
 NOR2x2_ASAP7_75t_R _32367_ (.A(_02745_),
    .B(_02785_),
    .Y(_02786_));
 XOR2x2_ASAP7_75t_R _32368_ (.A(_02692_),
    .B(_02786_),
    .Y(_02787_));
 INVx2_ASAP7_75t_R _32369_ (.A(_02787_),
    .Y(_02788_));
 NAND2x1_ASAP7_75t_R _32370_ (.A(_02589_),
    .B(_02788_),
    .Y(_02789_));
 NAND2x1_ASAP7_75t_R _32371_ (.A(_02588_),
    .B(_02787_),
    .Y(_02790_));
 AO21x1_ASAP7_75t_R _32372_ (.A1(net1613),
    .A2(net1612),
    .B(_01505_),
    .Y(_02791_));
 AO21x1_ASAP7_75t_R _32373_ (.A1(_01691_),
    .A2(_01699_),
    .B(_01505_),
    .Y(_02792_));
 TAPCELL_ASAP7_75t_R PHY_542 ();
 AO21x2_ASAP7_75t_R _32375_ (.A1(net1605),
    .A2(_01500_),
    .B(_01505_),
    .Y(_02794_));
 NAND3x2_ASAP7_75t_R _32376_ (.B(_02792_),
    .C(_02794_),
    .Y(_02795_),
    .A(_02791_));
 AOI211x1_ASAP7_75t_R _32377_ (.A1(_01498_),
    .A2(net1263),
    .B(net2334),
    .C(net2079),
    .Y(_02796_));
 INVx1_ASAP7_75t_R _32378_ (.A(_02796_),
    .Y(_02797_));
 INVx2_ASAP7_75t_R _32379_ (.A(_01569_),
    .Y(_02798_));
 NAND2x2_ASAP7_75t_R _32380_ (.A(_02798_),
    .B(_01657_),
    .Y(_02799_));
 AO21x1_ASAP7_75t_R _32381_ (.A1(net1613),
    .A2(_01600_),
    .B(net2334),
    .Y(_02800_));
 NAND3x2_ASAP7_75t_R _32382_ (.B(_02799_),
    .C(_02800_),
    .Y(_02801_),
    .A(_02797_));
 NOR2x2_ASAP7_75t_R _32383_ (.A(_02795_),
    .B(_02801_),
    .Y(_02802_));
 AO21x1_ASAP7_75t_R _32384_ (.A1(net1605),
    .A2(net3255),
    .B(_01624_),
    .Y(_02803_));
 NAND2x2_ASAP7_75t_R _32385_ (.A(_01499_),
    .B(_01599_),
    .Y(_02804_));
 AO21x1_ASAP7_75t_R _32386_ (.A1(_02804_),
    .A2(net2380),
    .B(_01624_),
    .Y(_02805_));
 OA211x2_ASAP7_75t_R _32387_ (.A1(_01624_),
    .A2(net2538),
    .B(_02803_),
    .C(_02805_),
    .Y(_02806_));
 AO21x1_ASAP7_75t_R _32388_ (.A1(net2366),
    .A2(net2063),
    .B(net2746),
    .Y(_02807_));
 AO21x1_ASAP7_75t_R _32389_ (.A1(net1457),
    .A2(_02363_),
    .B(_01636_),
    .Y(_02808_));
 INVx1_ASAP7_75t_R _32390_ (.A(_01642_),
    .Y(_02809_));
 NAND2x1_ASAP7_75t_R _32391_ (.A(_01575_),
    .B(_01637_),
    .Y(_02810_));
 AND4x2_ASAP7_75t_R _32392_ (.A(_02807_),
    .B(_02808_),
    .C(_02809_),
    .D(_02810_),
    .Y(_02811_));
 NAND3x2_ASAP7_75t_R _32393_ (.B(_02806_),
    .C(_02811_),
    .Y(_02812_),
    .A(_02802_));
 AO21x1_ASAP7_75t_R _32394_ (.A1(net3149),
    .A2(net2538),
    .B(_01543_),
    .Y(_02813_));
 NOR2x1_ASAP7_75t_R _32395_ (.A(net2818),
    .B(_01543_),
    .Y(_02814_));
 INVx1_ASAP7_75t_R _32396_ (.A(_02814_),
    .Y(_02815_));
 NAND2x1_ASAP7_75t_R _32397_ (.A(_02457_),
    .B(_01550_),
    .Y(_02816_));
 NAND2x1_ASAP7_75t_R _32398_ (.A(_02425_),
    .B(_01550_),
    .Y(_02817_));
 AND4x1_ASAP7_75t_R _32399_ (.A(_02813_),
    .B(_02815_),
    .C(_02816_),
    .D(_02817_),
    .Y(_02818_));
 AO21x1_ASAP7_75t_R _32400_ (.A1(net2819),
    .A2(_01540_),
    .B(_01571_),
    .Y(_02819_));
 NAND2x1_ASAP7_75t_R _32401_ (.A(_01565_),
    .B(_02425_),
    .Y(_02820_));
 NAND2x1_ASAP7_75t_R _32402_ (.A(_01565_),
    .B(_01719_),
    .Y(_02821_));
 AND3x1_ASAP7_75t_R _32403_ (.A(_02819_),
    .B(_02820_),
    .C(_02821_),
    .Y(_02822_));
 AND2x2_ASAP7_75t_R _32404_ (.A(_02818_),
    .B(_02822_),
    .Y(_02823_));
 AO21x1_ASAP7_75t_R _32405_ (.A1(net3149),
    .A2(net3255),
    .B(_01603_),
    .Y(_02824_));
 INVx1_ASAP7_75t_R _32406_ (.A(_01603_),
    .Y(_02825_));
 NAND2x1_ASAP7_75t_R _32407_ (.A(_02457_),
    .B(_02825_),
    .Y(_02826_));
 AND3x1_ASAP7_75t_R _32408_ (.A(_01608_),
    .B(_02824_),
    .C(_02826_),
    .Y(_02827_));
 AO21x1_ASAP7_75t_R _32409_ (.A1(net2366),
    .A2(net2256),
    .B(net2348),
    .Y(_02828_));
 INVx2_ASAP7_75t_R _32410_ (.A(_01586_),
    .Y(_02829_));
 NAND2x1_ASAP7_75t_R _32411_ (.A(_01526_),
    .B(_02829_),
    .Y(_02830_));
 AND2x2_ASAP7_75t_R _32412_ (.A(_02828_),
    .B(_02830_),
    .Y(_02831_));
 AO21x1_ASAP7_75t_R _32413_ (.A1(_01641_),
    .A2(_01590_),
    .B(net2794),
    .Y(_02832_));
 AO21x1_ASAP7_75t_R _32414_ (.A1(net1104),
    .A2(net3149),
    .B(net2794),
    .Y(_02833_));
 AND2x2_ASAP7_75t_R _32415_ (.A(_02832_),
    .B(_02833_),
    .Y(_02834_));
 AND3x1_ASAP7_75t_R _32416_ (.A(_02827_),
    .B(_02831_),
    .C(_02834_),
    .Y(_02835_));
 NAND2x1_ASAP7_75t_R _32417_ (.A(_02823_),
    .B(_02835_),
    .Y(_02836_));
 NOR2x2_ASAP7_75t_R _32418_ (.A(_02812_),
    .B(_02836_),
    .Y(_02837_));
 AO21x1_ASAP7_75t_R _32419_ (.A1(net1597),
    .A2(net3255),
    .B(_01701_),
    .Y(_02838_));
 INVx1_ASAP7_75t_R _32420_ (.A(_01701_),
    .Y(_02839_));
 NAND2x1_ASAP7_75t_R _32421_ (.A(_02798_),
    .B(_02839_),
    .Y(_02840_));
 NAND2x1_ASAP7_75t_R _32422_ (.A(_01525_),
    .B(_02839_),
    .Y(_02841_));
 NAND3x1_ASAP7_75t_R _32423_ (.A(_02838_),
    .B(_02840_),
    .C(_02841_),
    .Y(_02842_));
 OA21x2_ASAP7_75t_R _32424_ (.A1(_01635_),
    .A2(_01589_),
    .B(_01696_),
    .Y(_02843_));
 NOR2x1_ASAP7_75t_R _32425_ (.A(_02804_),
    .B(_01685_),
    .Y(_02844_));
 AOI21x1_ASAP7_75t_R _32426_ (.A1(_01569_),
    .A2(_01687_),
    .B(_01685_),
    .Y(_02845_));
 OR3x1_ASAP7_75t_R _32427_ (.A(_02843_),
    .B(_02844_),
    .C(_02845_),
    .Y(_02846_));
 NOR2x1_ASAP7_75t_R _32428_ (.A(_02842_),
    .B(_02846_),
    .Y(_02847_));
 AO21x1_ASAP7_75t_R _32429_ (.A1(net2062),
    .A2(_01674_),
    .B(_01675_),
    .Y(_02848_));
 AND2x2_ASAP7_75t_R _32430_ (.A(_02848_),
    .B(_01679_),
    .Y(_02849_));
 AO21x1_ASAP7_75t_R _32431_ (.A1(net3135),
    .A2(_01641_),
    .B(_01675_),
    .Y(_02850_));
 AO21x1_ASAP7_75t_R _32432_ (.A1(_01630_),
    .A2(net2728),
    .B(_01675_),
    .Y(_02851_));
 NAND2x1_ASAP7_75t_R _32433_ (.A(_02453_),
    .B(_01681_),
    .Y(_02852_));
 AND3x1_ASAP7_75t_R _32434_ (.A(_02850_),
    .B(_02851_),
    .C(_02852_),
    .Y(_02853_));
 NAND2x1_ASAP7_75t_R _32435_ (.A(_02849_),
    .B(_02853_),
    .Y(_02854_));
 NAND2x2_ASAP7_75t_R _32436_ (.A(_02453_),
    .B(_02368_),
    .Y(_02855_));
 AO21x1_ASAP7_75t_R _32437_ (.A1(net2728),
    .A2(_01612_),
    .B(_01668_),
    .Y(_02856_));
 NAND2x1_ASAP7_75t_R _32438_ (.A(_02855_),
    .B(_02856_),
    .Y(_02857_));
 OA211x2_ASAP7_75t_R _32439_ (.A1(_01498_),
    .A2(_01494_),
    .B(_02368_),
    .C(net3146),
    .Y(_02858_));
 OR2x2_ASAP7_75t_R _32440_ (.A(_02857_),
    .B(_02858_),
    .Y(_02859_));
 NOR2x1_ASAP7_75t_R _32441_ (.A(_02854_),
    .B(_02859_),
    .Y(_02860_));
 NAND2x1_ASAP7_75t_R _32442_ (.A(_02847_),
    .B(_02860_),
    .Y(_02861_));
 AO21x1_ASAP7_75t_R _32443_ (.A1(net3135),
    .A2(net2818),
    .B(_01728_),
    .Y(_02862_));
 AO21x1_ASAP7_75t_R _32444_ (.A1(net2062),
    .A2(net2254),
    .B(_01728_),
    .Y(_02863_));
 OR2x2_ASAP7_75t_R _32445_ (.A(_01500_),
    .B(_01728_),
    .Y(_02864_));
 NAND3x2_ASAP7_75t_R _32446_ (.B(_02863_),
    .C(_02864_),
    .Y(_02865_),
    .A(_02862_));
 AO21x1_ASAP7_75t_R _32447_ (.A1(net1457),
    .A2(_02363_),
    .B(_01735_),
    .Y(_02866_));
 NAND2x2_ASAP7_75t_R _32448_ (.A(_01747_),
    .B(_02866_),
    .Y(_02867_));
 NOR2x1_ASAP7_75t_R _32449_ (.A(_01735_),
    .B(_01674_),
    .Y(_02868_));
 INVx1_ASAP7_75t_R _32450_ (.A(_02868_),
    .Y(_02869_));
 AO21x1_ASAP7_75t_R _32451_ (.A1(_01689_),
    .A2(_01600_),
    .B(_01735_),
    .Y(_02870_));
 NAND2x2_ASAP7_75t_R _32452_ (.A(_02869_),
    .B(_02870_),
    .Y(_02871_));
 NOR3x2_ASAP7_75t_R _32453_ (.B(_02867_),
    .C(_02871_),
    .Y(_02872_),
    .A(_02865_));
 AO21x1_ASAP7_75t_R _32454_ (.A1(_02419_),
    .A2(net3149),
    .B(_01715_),
    .Y(_02873_));
 OAI21x1_ASAP7_75t_R _32455_ (.A1(net2524),
    .A2(_01715_),
    .B(_02873_),
    .Y(_02874_));
 OR3x2_ASAP7_75t_R _32456_ (.A(_01715_),
    .B(_01494_),
    .C(net2376),
    .Y(_02875_));
 AO21x1_ASAP7_75t_R _32457_ (.A1(_01691_),
    .A2(_01600_),
    .B(_01715_),
    .Y(_02876_));
 NAND3x2_ASAP7_75t_R _32458_ (.B(_02399_),
    .C(_02876_),
    .Y(_02877_),
    .A(_02875_));
 NOR2x2_ASAP7_75t_R _32459_ (.A(_02874_),
    .B(_02877_),
    .Y(_02878_));
 AOI211x1_ASAP7_75t_R _32460_ (.A1(net1120),
    .A2(net1263),
    .B(_01707_),
    .C(net1238),
    .Y(_02879_));
 INVx1_ASAP7_75t_R _32461_ (.A(_02879_),
    .Y(_02880_));
 TAPCELL_ASAP7_75t_R PHY_541 ();
 AO21x1_ASAP7_75t_R _32463_ (.A1(net2062),
    .A2(net2255),
    .B(_01707_),
    .Y(_02882_));
 AO21x1_ASAP7_75t_R _32464_ (.A1(net2524),
    .A2(net3266),
    .B(_01707_),
    .Y(_02883_));
 AO21x1_ASAP7_75t_R _32465_ (.A1(_01630_),
    .A2(_01540_),
    .B(_01707_),
    .Y(_02884_));
 AND4x2_ASAP7_75t_R _32466_ (.A(_02880_),
    .B(_02882_),
    .C(_02883_),
    .D(_02884_),
    .Y(_02885_));
 NAND3x2_ASAP7_75t_R _32467_ (.B(_02878_),
    .C(_02885_),
    .Y(_02886_),
    .A(_02872_));
 NOR2x2_ASAP7_75t_R _32468_ (.A(_02861_),
    .B(_02886_),
    .Y(_02887_));
 NAND2x2_ASAP7_75t_R _32469_ (.A(_02837_),
    .B(_02887_),
    .Y(_02888_));
 XOR2x1_ASAP7_75t_R _32470_ (.A(net2041),
    .Y(_02889_),
    .B(net3268));
 NAND3x1_ASAP7_75t_R _32471_ (.A(_02789_),
    .B(_02790_),
    .C(_02889_),
    .Y(_02890_));
 AO21x1_ASAP7_75t_R _32472_ (.A1(_02789_),
    .A2(_02790_),
    .B(_02889_),
    .Y(_02891_));
 AOI21x1_ASAP7_75t_R _32473_ (.A1(_02890_),
    .A2(_02891_),
    .B(_18753_),
    .Y(_02892_));
 OAI21x1_ASAP7_75t_R _32474_ (.A1(_02482_),
    .A2(_02892_),
    .B(_00482_),
    .Y(_02893_));
 AND2x2_ASAP7_75t_R _32475_ (.A(_18753_),
    .B(_00881_),
    .Y(_02894_));
 NAND2x1_ASAP7_75t_R _32476_ (.A(net3268),
    .B(_02788_),
    .Y(_02895_));
 INVx1_ASAP7_75t_R _32477_ (.A(_02888_),
    .Y(_02896_));
 NAND2x1_ASAP7_75t_R _32478_ (.A(_02896_),
    .B(_02787_),
    .Y(_02897_));
 XOR2x1_ASAP7_75t_R _32479_ (.A(net2041),
    .Y(_02898_),
    .B(_02588_));
 NAND3x1_ASAP7_75t_R _32480_ (.A(_02895_),
    .B(_02897_),
    .C(_02898_),
    .Y(_02899_));
 AO21x1_ASAP7_75t_R _32481_ (.A1(_02895_),
    .A2(_02897_),
    .B(_02898_),
    .Y(_02900_));
 AOI21x1_ASAP7_75t_R _32482_ (.A1(_02899_),
    .A2(_02900_),
    .B(_18753_),
    .Y(_02901_));
 INVx2_ASAP7_75t_R _32483_ (.A(_00482_),
    .Y(_02902_));
 OAI21x1_ASAP7_75t_R _32484_ (.A1(_02894_),
    .A2(_02901_),
    .B(_02902_),
    .Y(_02903_));
 NAND2x2_ASAP7_75t_R _32485_ (.A(_02903_),
    .B(_02893_),
    .Y(_00115_));
 NOR2x1_ASAP7_75t_R _32486_ (.A(net396),
    .B(_00880_),
    .Y(_02904_));
 AOI21x1_ASAP7_75t_R _32487_ (.A1(net3274),
    .A2(_01876_),
    .B(_01879_),
    .Y(_02905_));
 AO21x1_ASAP7_75t_R _32488_ (.A1(_01952_),
    .A2(_01908_),
    .B(_01878_),
    .Y(_02906_));
 AO21x1_ASAP7_75t_R _32489_ (.A1(_01946_),
    .A2(_01832_),
    .B(_01878_),
    .Y(_02907_));
 NAND3x1_ASAP7_75t_R _32490_ (.A(_02905_),
    .B(_02906_),
    .C(_02907_),
    .Y(_02908_));
 AO21x1_ASAP7_75t_R _32491_ (.A1(net2306),
    .A2(_02559_),
    .B(net2458),
    .Y(_02909_));
 NAND2x1_ASAP7_75t_R _32492_ (.A(_01871_),
    .B(_01888_),
    .Y(_02910_));
 AND3x1_ASAP7_75t_R _32493_ (.A(_02909_),
    .B(_02910_),
    .C(_02545_),
    .Y(_02911_));
 AO21x1_ASAP7_75t_R _32494_ (.A1(net3277),
    .A2(net1245),
    .B(net2458),
    .Y(_02912_));
 AO21x1_ASAP7_75t_R _32495_ (.A1(_01946_),
    .A2(_01832_),
    .B(net2458),
    .Y(_02913_));
 INVx1_ASAP7_75t_R _32496_ (.A(_02549_),
    .Y(_02914_));
 AND3x1_ASAP7_75t_R _32497_ (.A(_02912_),
    .B(_02913_),
    .C(_02914_),
    .Y(_02915_));
 NAND2x1_ASAP7_75t_R _32498_ (.A(_02911_),
    .B(_02915_),
    .Y(_02916_));
 NOR2x1_ASAP7_75t_R _32499_ (.A(_02908_),
    .B(_02916_),
    .Y(_02917_));
 INVx3_ASAP7_75t_R _32500_ (.A(net1245),
    .Y(_02918_));
 OA21x2_ASAP7_75t_R _32501_ (.A1(_02918_),
    .A2(_01890_),
    .B(_01847_),
    .Y(_02919_));
 NOR2x1_ASAP7_75t_R _32502_ (.A(_02134_),
    .B(_01851_),
    .Y(_02920_));
 OA21x2_ASAP7_75t_R _32503_ (.A1(_02544_),
    .A2(_01871_),
    .B(_01847_),
    .Y(_02921_));
 OR3x1_ASAP7_75t_R _32504_ (.A(_02919_),
    .B(_02920_),
    .C(_02921_),
    .Y(_02922_));
 NOR2x1_ASAP7_75t_R _32505_ (.A(_01857_),
    .B(_01863_),
    .Y(_02923_));
 INVx1_ASAP7_75t_R _32506_ (.A(_02923_),
    .Y(_02924_));
 OA21x2_ASAP7_75t_R _32507_ (.A1(net1453),
    .A2(_02924_),
    .B(_02123_),
    .Y(_02925_));
 NAND2x1_ASAP7_75t_R _32508_ (.A(_01862_),
    .B(_01864_),
    .Y(_02926_));
 AO21x1_ASAP7_75t_R _32509_ (.A1(_02110_),
    .A2(_01832_),
    .B(_01863_),
    .Y(_02927_));
 NAND3x1_ASAP7_75t_R _32510_ (.A(_02925_),
    .B(_02926_),
    .C(_02927_),
    .Y(_02928_));
 NOR2x1_ASAP7_75t_R _32511_ (.A(_02922_),
    .B(_02928_),
    .Y(_02929_));
 NAND2x2_ASAP7_75t_R _32512_ (.A(_02917_),
    .B(_02929_),
    .Y(_02930_));
 AO21x1_ASAP7_75t_R _32513_ (.A1(_01799_),
    .A2(net2286),
    .B(_01828_),
    .Y(_02931_));
 OA21x2_ASAP7_75t_R _32514_ (.A1(_01828_),
    .A2(_01795_),
    .B(_02931_),
    .Y(_02932_));
 NOR2x1_ASAP7_75t_R _32515_ (.A(_02190_),
    .B(_01886_),
    .Y(_02933_));
 NOR2x1_ASAP7_75t_R _32516_ (.A(net1459),
    .B(net1554),
    .Y(_02934_));
 AO21x1_ASAP7_75t_R _32517_ (.A1(_02933_),
    .A2(_02934_),
    .B(_01809_),
    .Y(_02935_));
 NAND2x1_ASAP7_75t_R _32518_ (.A(_02099_),
    .B(_02141_),
    .Y(_02936_));
 NAND3x1_ASAP7_75t_R _32519_ (.A(_02932_),
    .B(_02935_),
    .C(_02936_),
    .Y(_02937_));
 INVx1_ASAP7_75t_R _32520_ (.A(_02937_),
    .Y(_02938_));
 AO21x1_ASAP7_75t_R _32521_ (.A1(net3275),
    .A2(_01908_),
    .B(_01761_),
    .Y(_02939_));
 OA21x2_ASAP7_75t_R _32522_ (.A1(net2239),
    .A2(_01761_),
    .B(_02939_),
    .Y(_02940_));
 OA211x2_ASAP7_75t_R _32523_ (.A1(_01770_),
    .A2(_01776_),
    .B(_01762_),
    .C(net1554),
    .Y(_02941_));
 INVx1_ASAP7_75t_R _32524_ (.A(_02941_),
    .Y(_02942_));
 NAND2x1_ASAP7_75t_R _32525_ (.A(_02940_),
    .B(_02942_),
    .Y(_02943_));
 OA21x2_ASAP7_75t_R _32526_ (.A1(_01862_),
    .A2(_01890_),
    .B(_02131_),
    .Y(_02944_));
 OA21x2_ASAP7_75t_R _32527_ (.A1(_02124_),
    .A2(_01858_),
    .B(_02131_),
    .Y(_02945_));
 AOI211x1_ASAP7_75t_R _32528_ (.A1(_01770_),
    .A2(_01776_),
    .B(_01781_),
    .C(_01870_),
    .Y(_02946_));
 NOR2x1_ASAP7_75t_R _32529_ (.A(_01781_),
    .B(_02129_),
    .Y(_02947_));
 OR4x1_ASAP7_75t_R _32530_ (.A(_02944_),
    .B(_02945_),
    .C(_02946_),
    .D(_02947_),
    .Y(_02948_));
 NOR2x1_ASAP7_75t_R _32531_ (.A(_02943_),
    .B(_02948_),
    .Y(_02949_));
 NAND2x2_ASAP7_75t_R _32532_ (.A(_02938_),
    .B(_02949_),
    .Y(_02950_));
 NOR2x2_ASAP7_75t_R _32533_ (.A(_02930_),
    .B(_02950_),
    .Y(_02951_));
 AO21x1_ASAP7_75t_R _32534_ (.A1(net1316),
    .A2(_01832_),
    .B(net2653),
    .Y(_02952_));
 AO21x1_ASAP7_75t_R _32535_ (.A1(_01908_),
    .A2(net2371),
    .B(net2653),
    .Y(_02953_));
 NOR2x1_ASAP7_75t_R _32536_ (.A(net2708),
    .B(net2653),
    .Y(_02954_));
 INVx1_ASAP7_75t_R _32537_ (.A(_02954_),
    .Y(_02955_));
 NAND3x1_ASAP7_75t_R _32538_ (.A(_02952_),
    .B(_02953_),
    .C(_02955_),
    .Y(_02956_));
 OA21x2_ASAP7_75t_R _32539_ (.A1(_01816_),
    .A2(_01843_),
    .B(_01904_),
    .Y(_02957_));
 NOR2x1_ASAP7_75t_R _32540_ (.A(net2708),
    .B(_01905_),
    .Y(_02958_));
 OA21x2_ASAP7_75t_R _32541_ (.A1(_01855_),
    .A2(_02124_),
    .B(_01904_),
    .Y(_02959_));
 OR3x1_ASAP7_75t_R _32542_ (.A(_02957_),
    .B(_02958_),
    .C(_02959_),
    .Y(_02960_));
 NOR2x1_ASAP7_75t_R _32543_ (.A(_02956_),
    .B(_02960_),
    .Y(_02961_));
 NOR2x1_ASAP7_75t_R _32544_ (.A(net3171),
    .B(net3276),
    .Y(_02962_));
 NOR2x1_ASAP7_75t_R _32545_ (.A(net3170),
    .B(net3332),
    .Y(_02963_));
 NOR2x1_ASAP7_75t_R _32546_ (.A(net1157),
    .B(net3171),
    .Y(_02964_));
 OR3x1_ASAP7_75t_R _32547_ (.A(_02962_),
    .B(_02963_),
    .C(_02964_),
    .Y(_02965_));
 AO21x1_ASAP7_75t_R _32548_ (.A1(_01819_),
    .A2(net3169),
    .B(net2549),
    .Y(_02966_));
 NAND2x1_ASAP7_75t_R _32549_ (.A(_01930_),
    .B(_02114_),
    .Y(_02967_));
 NAND3x1_ASAP7_75t_R _32550_ (.A(_02966_),
    .B(_02186_),
    .C(_02967_),
    .Y(_02968_));
 AO21x1_ASAP7_75t_R _32551_ (.A1(_01832_),
    .A2(_01877_),
    .B(net2193),
    .Y(_02969_));
 AO21x1_ASAP7_75t_R _32552_ (.A1(_01799_),
    .A2(_01908_),
    .B(net2193),
    .Y(_02970_));
 NAND2x1_ASAP7_75t_R _32553_ (.A(_02969_),
    .B(_02970_),
    .Y(_02971_));
 NOR3x1_ASAP7_75t_R _32554_ (.A(_02965_),
    .B(_02968_),
    .C(_02971_),
    .Y(_02972_));
 AND2x2_ASAP7_75t_R _32555_ (.A(_02961_),
    .B(_02972_),
    .Y(_02973_));
 INVx2_ASAP7_75t_R _32556_ (.A(_02973_),
    .Y(_02974_));
 NAND2x1_ASAP7_75t_R _32557_ (.A(_02190_),
    .B(_02498_),
    .Y(_02975_));
 AO21x1_ASAP7_75t_R _32558_ (.A1(_02500_),
    .A2(_01825_),
    .B(net3125),
    .Y(_02976_));
 NAND2x1_ASAP7_75t_R _32559_ (.A(_02975_),
    .B(_02976_),
    .Y(_02977_));
 NOR2x1_ASAP7_75t_R _32560_ (.A(net2369),
    .B(net2262),
    .Y(_02978_));
 AOI211x1_ASAP7_75t_R _32561_ (.A1(_01770_),
    .A2(_01776_),
    .B(net2262),
    .C(_01870_),
    .Y(_02979_));
 OR3x1_ASAP7_75t_R _32562_ (.A(_02977_),
    .B(_02978_),
    .C(_02979_),
    .Y(_02980_));
 AO21x1_ASAP7_75t_R _32563_ (.A1(_01795_),
    .A2(_02559_),
    .B(_01955_),
    .Y(_02981_));
 INVx1_ASAP7_75t_R _32564_ (.A(_02221_),
    .Y(_02982_));
 OA21x2_ASAP7_75t_R _32565_ (.A1(_02981_),
    .A2(net1448),
    .B(_02982_),
    .Y(_02983_));
 AO21x1_ASAP7_75t_R _32566_ (.A1(_02110_),
    .A2(net3276),
    .B(_01955_),
    .Y(_02984_));
 AO21x1_ASAP7_75t_R _32567_ (.A1(net1413),
    .A2(_01824_),
    .B(_01955_),
    .Y(_02985_));
 NAND3x1_ASAP7_75t_R _32568_ (.A(_02983_),
    .B(_02984_),
    .C(_02985_),
    .Y(_02986_));
 NOR2x1_ASAP7_75t_R _32569_ (.A(_02980_),
    .B(_02986_),
    .Y(_02987_));
 AO21x1_ASAP7_75t_R _32570_ (.A1(_01869_),
    .A2(_01786_),
    .B(net1302),
    .Y(_02988_));
 AO21x1_ASAP7_75t_R _32571_ (.A1(_01824_),
    .A2(net1458),
    .B(_01967_),
    .Y(_02989_));
 OA21x2_ASAP7_75t_R _32572_ (.A1(_01967_),
    .A2(_02988_),
    .B(_02989_),
    .Y(_02990_));
 OA211x2_ASAP7_75t_R _32573_ (.A1(net1116),
    .A2(_01776_),
    .B(_01970_),
    .C(net1131),
    .Y(_02991_));
 AOI21x1_ASAP7_75t_R _32574_ (.A1(net2654),
    .A2(_01970_),
    .B(_02991_),
    .Y(_02992_));
 NAND2x1_ASAP7_75t_R _32575_ (.A(_02990_),
    .B(_02992_),
    .Y(_02993_));
 OA211x2_ASAP7_75t_R _32576_ (.A1(net1116),
    .A2(_01776_),
    .B(_01974_),
    .C(net1461),
    .Y(_02994_));
 NOR2x1_ASAP7_75t_R _32577_ (.A(_01795_),
    .B(_01977_),
    .Y(_02995_));
 OA21x2_ASAP7_75t_R _32578_ (.A1(_01806_),
    .A2(_01890_),
    .B(_01974_),
    .Y(_02996_));
 OR3x1_ASAP7_75t_R _32579_ (.A(_02994_),
    .B(_02995_),
    .C(_02996_),
    .Y(_02997_));
 NOR2x1_ASAP7_75t_R _32580_ (.A(_02993_),
    .B(_02997_),
    .Y(_02998_));
 NAND2x1_ASAP7_75t_R _32581_ (.A(_02987_),
    .B(_02998_),
    .Y(_02999_));
 NOR2x2_ASAP7_75t_R _32582_ (.A(_02974_),
    .B(_02999_),
    .Y(_03000_));
 NAND2x2_ASAP7_75t_R _32583_ (.A(_02951_),
    .B(_03000_),
    .Y(_03001_));
 TAPCELL_ASAP7_75t_R PHY_540 ();
 NAND2x2_ASAP7_75t_R _32585_ (.A(_01987_),
    .B(_03001_),
    .Y(_03003_));
 INVx4_ASAP7_75t_R _32586_ (.A(_03001_),
    .Y(_03004_));
 NAND2x1_ASAP7_75t_R _32587_ (.A(_02240_),
    .B(_03004_),
    .Y(_03005_));
 AO21x1_ASAP7_75t_R _32588_ (.A1(net2120),
    .A2(net2361),
    .B(_01334_),
    .Y(_03006_));
 AND2x2_ASAP7_75t_R _32589_ (.A(_03006_),
    .B(_02688_),
    .Y(_03007_));
 AO21x1_ASAP7_75t_R _32590_ (.A1(net1866),
    .A2(net1803),
    .B(_01334_),
    .Y(_03008_));
 OA21x2_ASAP7_75t_R _32591_ (.A1(_01334_),
    .A2(net1076),
    .B(_03008_),
    .Y(_03009_));
 NAND2x1_ASAP7_75t_R _32592_ (.A(_03007_),
    .B(_03009_),
    .Y(_03010_));
 NOR2x2_ASAP7_75t_R _32593_ (.A(net2361),
    .B(_01345_),
    .Y(_03011_));
 NOR2x2_ASAP7_75t_R _32594_ (.A(_03011_),
    .B(_02066_),
    .Y(_03012_));
 AO21x2_ASAP7_75t_R _32595_ (.A1(net2522),
    .A2(net1698),
    .B(_01345_),
    .Y(_03013_));
 AO21x1_ASAP7_75t_R _32596_ (.A1(net1076),
    .A2(_01259_),
    .B(net3240),
    .Y(_03014_));
 NAND3x2_ASAP7_75t_R _32597_ (.B(net3288),
    .C(_03014_),
    .Y(_03015_),
    .A(_03012_));
 NOR2x2_ASAP7_75t_R _32598_ (.A(_03010_),
    .B(_03015_),
    .Y(_03016_));
 AO21x2_ASAP7_75t_R _32599_ (.A1(net2361),
    .A2(net1142),
    .B(_01322_),
    .Y(_03017_));
 OAI21x1_ASAP7_75t_R _32600_ (.A1(net2460),
    .A2(_01226_),
    .B(_03017_),
    .Y(_03018_));
 AO21x2_ASAP7_75t_R _32601_ (.A1(net1802),
    .A2(net1698),
    .B(_01322_),
    .Y(_03019_));
 NAND2x1_ASAP7_75t_R _32602_ (.A(_02061_),
    .B(_01329_),
    .Y(_03020_));
 NAND2x1_ASAP7_75t_R _32603_ (.A(net1331),
    .B(_01329_),
    .Y(_03021_));
 NAND3x1_ASAP7_75t_R _32604_ (.A(_03019_),
    .B(_03020_),
    .C(_03021_),
    .Y(_03022_));
 NOR2x1_ASAP7_75t_R _32605_ (.A(_03018_),
    .B(_03022_),
    .Y(_03023_));
 AO21x1_ASAP7_75t_R _32606_ (.A1(_01113_),
    .A2(_02032_),
    .B(_01308_),
    .Y(_03024_));
 AO21x1_ASAP7_75t_R _32607_ (.A1(net1752),
    .A2(_01453_),
    .B(_01308_),
    .Y(_03025_));
 AND3x1_ASAP7_75t_R _32608_ (.A(_03024_),
    .B(_03025_),
    .C(_02080_),
    .Y(_03026_));
 AND2x2_ASAP7_75t_R _32609_ (.A(_03023_),
    .B(_03026_),
    .Y(_03027_));
 NAND2x2_ASAP7_75t_R _32610_ (.A(_03016_),
    .B(_03027_),
    .Y(_03028_));
 AO21x1_ASAP7_75t_R _32611_ (.A1(net1266),
    .A2(net938),
    .B(net3315),
    .Y(_03029_));
 NAND2x1_ASAP7_75t_R _32612_ (.A(_01405_),
    .B(_01265_),
    .Y(_03030_));
 INVx1_ASAP7_75t_R _32613_ (.A(_01410_),
    .Y(_03031_));
 AND3x1_ASAP7_75t_R _32614_ (.A(_03029_),
    .B(_03030_),
    .C(_03031_),
    .Y(_03032_));
 AND3x1_ASAP7_75t_R _32615_ (.A(_02623_),
    .B(_01251_),
    .C(_01187_),
    .Y(_03033_));
 AOI21x1_ASAP7_75t_R _32616_ (.A1(_01112_),
    .A2(_01244_),
    .B(_03033_),
    .Y(_03034_));
 AND2x2_ASAP7_75t_R _32617_ (.A(_03032_),
    .B(_03034_),
    .Y(_03035_));
 AO21x1_ASAP7_75t_R _32618_ (.A1(_01416_),
    .A2(_01173_),
    .B(_01283_),
    .Y(_03036_));
 AO21x1_ASAP7_75t_R _32619_ (.A1(_01416_),
    .A2(_01474_),
    .B(_01281_),
    .Y(_03037_));
 AOI211x1_ASAP7_75t_R _32620_ (.A1(_01416_),
    .A2(_01180_),
    .B(_03036_),
    .C(_03037_),
    .Y(_03038_));
 AO21x1_ASAP7_75t_R _32621_ (.A1(net2723),
    .A2(net1572),
    .B(net3145),
    .Y(_03039_));
 OAI21x1_ASAP7_75t_R _32622_ (.A1(net3145),
    .A2(net940),
    .B(_03039_),
    .Y(_03040_));
 AND3x1_ASAP7_75t_R _32623_ (.A(_01288_),
    .B(_01187_),
    .C(_01279_),
    .Y(_03041_));
 AOI211x1_ASAP7_75t_R _32624_ (.A1(_01288_),
    .A2(_01374_),
    .B(_03040_),
    .C(_03041_),
    .Y(_03042_));
 NAND3x2_ASAP7_75t_R _32625_ (.B(_03038_),
    .C(_03042_),
    .Y(_03043_),
    .A(_03035_));
 NOR2x2_ASAP7_75t_R _32626_ (.A(_03028_),
    .B(_03043_),
    .Y(_03044_));
 AOI211x1_ASAP7_75t_R _32627_ (.A1(net1341),
    .A2(_01096_),
    .B(_01229_),
    .C(_01204_),
    .Y(_03045_));
 OA21x2_ASAP7_75t_R _32628_ (.A1(_01327_),
    .A2(_02061_),
    .B(_01234_),
    .Y(_03046_));
 NOR2x1_ASAP7_75t_R _32629_ (.A(_03045_),
    .B(_03046_),
    .Y(_03047_));
 AO221x1_ASAP7_75t_R _32630_ (.A1(net2872),
    .A2(net3289),
    .B1(_01159_),
    .B2(_01248_),
    .C(_01229_),
    .Y(_03048_));
 NAND2x1_ASAP7_75t_R _32631_ (.A(_03047_),
    .B(_03048_),
    .Y(_03049_));
 NAND2x1_ASAP7_75t_R _32632_ (.A(_01218_),
    .B(_02600_),
    .Y(_03050_));
 NAND2x1_ASAP7_75t_R _32633_ (.A(_01328_),
    .B(_01218_),
    .Y(_03051_));
 AND3x1_ASAP7_75t_R _32634_ (.A(_03050_),
    .B(_02620_),
    .C(_03051_),
    .Y(_03052_));
 AOI211x1_ASAP7_75t_R _32635_ (.A1(net1341),
    .A2(net3289),
    .B(_01215_),
    .C(net1429),
    .Y(_03053_));
 NOR2x2_ASAP7_75t_R _32636_ (.A(_01215_),
    .B(net2731),
    .Y(_03054_));
 AOI211x1_ASAP7_75t_R _32637_ (.A1(_01218_),
    .A2(_01160_),
    .B(_03053_),
    .C(_03054_),
    .Y(_03055_));
 NAND2x1_ASAP7_75t_R _32638_ (.A(_03052_),
    .B(_03055_),
    .Y(_03056_));
 NOR2x1_ASAP7_75t_R _32639_ (.A(_03049_),
    .B(_03056_),
    .Y(_03057_));
 NAND2x1_ASAP7_75t_R _32640_ (.A(_01109_),
    .B(_01210_),
    .Y(_03058_));
 AO21x1_ASAP7_75t_R _32641_ (.A1(net2872),
    .A2(net1277),
    .B(_03058_),
    .Y(_03059_));
 OAI21x1_ASAP7_75t_R _32642_ (.A1(net3154),
    .A2(_01303_),
    .B(_03059_),
    .Y(_03060_));
 NAND2x1_ASAP7_75t_R _32643_ (.A(net1333),
    .B(_01210_),
    .Y(_03061_));
 NAND2x1_ASAP7_75t_R _32644_ (.A(_01327_),
    .B(_01210_),
    .Y(_03062_));
 NAND3x1_ASAP7_75t_R _32645_ (.A(_01433_),
    .B(_03061_),
    .C(_03062_),
    .Y(_03063_));
 AO21x1_ASAP7_75t_R _32646_ (.A1(_01303_),
    .A2(net938),
    .B(net3144),
    .Y(_03064_));
 AO21x1_ASAP7_75t_R _32647_ (.A1(net940),
    .A2(_01259_),
    .B(net3144),
    .Y(_03065_));
 NAND3x1_ASAP7_75t_R _32648_ (.A(_03064_),
    .B(_03065_),
    .C(_02632_),
    .Y(_03066_));
 NOR3x1_ASAP7_75t_R _32649_ (.A(_03060_),
    .B(_03063_),
    .C(_03066_),
    .Y(_03067_));
 NAND2x1_ASAP7_75t_R _32650_ (.A(_03057_),
    .B(_03067_),
    .Y(_03068_));
 AO21x1_ASAP7_75t_R _32651_ (.A1(_01303_),
    .A2(_01321_),
    .B(_01120_),
    .Y(_03069_));
 NAND2x1_ASAP7_75t_R _32652_ (.A(_01103_),
    .B(_01286_),
    .Y(_03070_));
 NAND2x2_ASAP7_75t_R _32653_ (.A(_01103_),
    .B(_02619_),
    .Y(_03071_));
 AND3x1_ASAP7_75t_R _32654_ (.A(_03069_),
    .B(_03070_),
    .C(_03071_),
    .Y(_03072_));
 NAND2x1_ASAP7_75t_R _32655_ (.A(_01187_),
    .B(_02593_),
    .Y(_03073_));
 OA21x2_ASAP7_75t_R _32656_ (.A1(net1277),
    .A2(_03073_),
    .B(_02590_),
    .Y(_03074_));
 OA21x2_ASAP7_75t_R _32657_ (.A1(_01204_),
    .A2(_01133_),
    .B(_01465_),
    .Y(_03075_));
 AND3x1_ASAP7_75t_R _32658_ (.A(_03072_),
    .B(_03074_),
    .C(_03075_),
    .Y(_03076_));
 AO21x1_ASAP7_75t_R _32659_ (.A1(net2125),
    .A2(net1141),
    .B(_01170_),
    .Y(_03077_));
 AO21x1_ASAP7_75t_R _32660_ (.A1(_01138_),
    .A2(_01226_),
    .B(_01170_),
    .Y(_03078_));
 NAND2x1_ASAP7_75t_R _32661_ (.A(_01160_),
    .B(_01171_),
    .Y(_03079_));
 AND3x1_ASAP7_75t_R _32662_ (.A(_03077_),
    .B(_03078_),
    .C(_03079_),
    .Y(_03080_));
 OA21x2_ASAP7_75t_R _32663_ (.A1(_01166_),
    .A2(_02023_),
    .B(_01163_),
    .Y(_03081_));
 OA21x2_ASAP7_75t_R _32664_ (.A1(net2443),
    .A2(_01160_),
    .B(_01163_),
    .Y(_03082_));
 NOR2x1_ASAP7_75t_R _32665_ (.A(_02032_),
    .B(_01156_),
    .Y(_03083_));
 NOR3x1_ASAP7_75t_R _32666_ (.A(_03081_),
    .B(_03082_),
    .C(_03083_),
    .Y(_03084_));
 AO21x1_ASAP7_75t_R _32667_ (.A1(net1884),
    .A2(net940),
    .B(_01170_),
    .Y(_03085_));
 OA21x2_ASAP7_75t_R _32668_ (.A1(_01143_),
    .A2(_01170_),
    .B(_03085_),
    .Y(_03086_));
 AND3x1_ASAP7_75t_R _32669_ (.A(_03080_),
    .B(_03084_),
    .C(_03086_),
    .Y(_03087_));
 NAND2x1_ASAP7_75t_R _32670_ (.A(_03076_),
    .B(_03087_),
    .Y(_03088_));
 NOR2x1_ASAP7_75t_R _32671_ (.A(_03068_),
    .B(_03088_),
    .Y(_03089_));
 NAND2x2_ASAP7_75t_R _32672_ (.A(_03044_),
    .B(_03089_),
    .Y(_03090_));
 INVx1_ASAP7_75t_R _32673_ (.A(_03090_),
    .Y(_03091_));
 AOI21x1_ASAP7_75t_R _32674_ (.A1(_03003_),
    .A2(_03005_),
    .B(_03091_),
    .Y(_03092_));
 AO21x1_ASAP7_75t_R _32675_ (.A1(_03000_),
    .A2(_02951_),
    .B(_01987_),
    .Y(_03093_));
 NAND2x1_ASAP7_75t_R _32676_ (.A(_01987_),
    .B(_03004_),
    .Y(_03094_));
 AOI21x1_ASAP7_75t_R _32677_ (.A1(_03093_),
    .A2(_03094_),
    .B(net2793),
    .Y(_03095_));
 NOR2x1_ASAP7_75t_R _32678_ (.A(_03092_),
    .B(_03095_),
    .Y(_03096_));
 AO21x2_ASAP7_75t_R _32679_ (.A1(_22045_),
    .A2(net996),
    .B(net1851),
    .Y(_03097_));
 AO21x1_ASAP7_75t_R _32680_ (.A1(_03097_),
    .A2(net2752),
    .B(_21976_),
    .Y(_03098_));
 NOR2x1_ASAP7_75t_R _32681_ (.A(_22024_),
    .B(_21962_),
    .Y(_03099_));
 INVx1_ASAP7_75t_R _32682_ (.A(_03099_),
    .Y(_03100_));
 NAND2x1_ASAP7_75t_R _32683_ (.A(_21957_),
    .B(_01087_),
    .Y(_03101_));
 AO21x1_ASAP7_75t_R _32684_ (.A1(_21920_),
    .A2(net1792),
    .B(_21962_),
    .Y(_03102_));
 AND4x1_ASAP7_75t_R _32685_ (.A(_03098_),
    .B(_03100_),
    .C(_03101_),
    .D(_03102_),
    .Y(_03103_));
 AO21x1_ASAP7_75t_R _32686_ (.A1(_21983_),
    .A2(_22018_),
    .B(_21901_),
    .Y(_03104_));
 NAND2x1_ASAP7_75t_R _32687_ (.A(_21877_),
    .B(_21926_),
    .Y(_03105_));
 AO21x1_ASAP7_75t_R _32688_ (.A1(_03105_),
    .A2(_22080_),
    .B(_21901_),
    .Y(_03106_));
 NOR2x2_ASAP7_75t_R _32689_ (.A(net2295),
    .B(_21895_),
    .Y(_03107_));
 NAND2x1_ASAP7_75t_R _32690_ (.A(_03107_),
    .B(_02323_),
    .Y(_03108_));
 NAND3x1_ASAP7_75t_R _32691_ (.A(_03104_),
    .B(_03106_),
    .C(_03108_),
    .Y(_03109_));
 INVx1_ASAP7_75t_R _32692_ (.A(_03109_),
    .Y(_03110_));
 OA21x2_ASAP7_75t_R _32693_ (.A1(_22046_),
    .A2(_21909_),
    .B(_21885_),
    .Y(_03111_));
 INVx1_ASAP7_75t_R _32694_ (.A(_03111_),
    .Y(_03112_));
 AO21x1_ASAP7_75t_R _32695_ (.A1(_21920_),
    .A2(net1632),
    .B(net2496),
    .Y(_03113_));
 AND2x2_ASAP7_75t_R _32696_ (.A(_03112_),
    .B(_03113_),
    .Y(_03114_));
 AO21x1_ASAP7_75t_R _32697_ (.A1(net2752),
    .A2(_21940_),
    .B(net2496),
    .Y(_03115_));
 OA21x2_ASAP7_75t_R _32698_ (.A1(net2510),
    .A2(net2496),
    .B(_03115_),
    .Y(_03116_));
 AND3x1_ASAP7_75t_R _32699_ (.A(_03110_),
    .B(_03114_),
    .C(_03116_),
    .Y(_03117_));
 NAND2x1_ASAP7_75t_R _32700_ (.A(_03103_),
    .B(_03117_),
    .Y(_03118_));
 AO21x1_ASAP7_75t_R _32701_ (.A1(net3172),
    .A2(net1834),
    .B(_21992_),
    .Y(_03119_));
 NAND2x1_ASAP7_75t_R _32702_ (.A(net2802),
    .B(_02758_),
    .Y(_03120_));
 NAND2x1_ASAP7_75t_R _32703_ (.A(_21872_),
    .B(_02758_),
    .Y(_03121_));
 AND3x1_ASAP7_75t_R _32704_ (.A(_03119_),
    .B(_03120_),
    .C(_03121_),
    .Y(_03122_));
 AO21x1_ASAP7_75t_R _32705_ (.A1(_02305_),
    .A2(_03105_),
    .B(_22004_),
    .Y(_03123_));
 AO21x1_ASAP7_75t_R _32706_ (.A1(net2752),
    .A2(_21940_),
    .B(_22004_),
    .Y(_03124_));
 OA21x2_ASAP7_75t_R _32707_ (.A1(_22004_),
    .A2(net2365),
    .B(_03124_),
    .Y(_03125_));
 AND3x1_ASAP7_75t_R _32708_ (.A(_03122_),
    .B(_03123_),
    .C(_03125_),
    .Y(_03126_));
 AO21x1_ASAP7_75t_R _32709_ (.A1(net3172),
    .A2(net1634),
    .B(net3156),
    .Y(_03127_));
 AND2x2_ASAP7_75t_R _32710_ (.A(_03127_),
    .B(_02747_),
    .Y(_03128_));
 AO21x2_ASAP7_75t_R _32711_ (.A1(_21934_),
    .A2(_22018_),
    .B(_22015_),
    .Y(_03129_));
 AO21x1_ASAP7_75t_R _32712_ (.A1(net2258),
    .A2(_21969_),
    .B(net3075),
    .Y(_03130_));
 AND2x2_ASAP7_75t_R _32713_ (.A(_03129_),
    .B(_03130_),
    .Y(_03131_));
 AOI22x1_ASAP7_75t_R _32714_ (.A1(_02340_),
    .A2(net994),
    .B1(_01085_),
    .B2(_22016_),
    .Y(_03132_));
 NAND2x1_ASAP7_75t_R _32715_ (.A(net1172),
    .B(net1649),
    .Y(_03133_));
 AO21x1_ASAP7_75t_R _32716_ (.A1(_03133_),
    .A2(net2258),
    .B(net2556),
    .Y(_03134_));
 AND4x1_ASAP7_75t_R _32717_ (.A(_03128_),
    .B(_03131_),
    .C(_03132_),
    .D(_03134_),
    .Y(_03135_));
 NAND2x1_ASAP7_75t_R _32718_ (.A(_03126_),
    .B(_03135_),
    .Y(_03136_));
 NOR2x2_ASAP7_75t_R _32719_ (.A(_03118_),
    .B(_03136_),
    .Y(_03137_));
 AO21x1_ASAP7_75t_R _32720_ (.A1(_21929_),
    .A2(net2801),
    .B(_22061_),
    .Y(_03138_));
 AO21x2_ASAP7_75t_R _32721_ (.A1(net2293),
    .A2(net1833),
    .B(_22061_),
    .Y(_03139_));
 AO21x1_ASAP7_75t_R _32722_ (.A1(_02259_),
    .A2(_02273_),
    .B(_22061_),
    .Y(_03140_));
 AND3x1_ASAP7_75t_R _32723_ (.A(_03138_),
    .B(_03139_),
    .C(_03140_),
    .Y(_03141_));
 AO21x1_ASAP7_75t_R _32724_ (.A1(_22024_),
    .A2(net2801),
    .B(_22064_),
    .Y(_03142_));
 AO21x1_ASAP7_75t_R _32725_ (.A1(net1629),
    .A2(net1833),
    .B(_22064_),
    .Y(_03143_));
 NAND2x1_ASAP7_75t_R _32726_ (.A(_22049_),
    .B(_22003_),
    .Y(_03144_));
 AND3x1_ASAP7_75t_R _32727_ (.A(_03142_),
    .B(_03143_),
    .C(_03144_),
    .Y(_03145_));
 NOR2x1_ASAP7_75t_R _32728_ (.A(net1711),
    .B(_22064_),
    .Y(_03146_));
 INVx1_ASAP7_75t_R _32729_ (.A(_21969_),
    .Y(_03147_));
 OA21x2_ASAP7_75t_R _32730_ (.A1(_01087_),
    .A2(_03147_),
    .B(_22049_),
    .Y(_03148_));
 AOI21x1_ASAP7_75t_R _32731_ (.A1(_21918_),
    .A2(_03146_),
    .B(_03148_),
    .Y(_03149_));
 AND3x1_ASAP7_75t_R _32732_ (.A(_03141_),
    .B(_03145_),
    .C(_03149_),
    .Y(_03150_));
 AO21x1_ASAP7_75t_R _32733_ (.A1(_02259_),
    .A2(_22018_),
    .B(_22077_),
    .Y(_03151_));
 AO21x1_ASAP7_75t_R _32734_ (.A1(net2260),
    .A2(_21940_),
    .B(_22077_),
    .Y(_03152_));
 AND2x2_ASAP7_75t_R _32735_ (.A(_03151_),
    .B(_03152_),
    .Y(_03153_));
 AO21x2_ASAP7_75t_R _32736_ (.A1(_02259_),
    .A2(net3236),
    .B(_22070_),
    .Y(_03154_));
 NAND2x1_ASAP7_75t_R _32737_ (.A(net1259),
    .B(_02292_),
    .Y(_03155_));
 AND2x2_ASAP7_75t_R _32738_ (.A(_03154_),
    .B(_03155_),
    .Y(_03156_));
 AO21x1_ASAP7_75t_R _32739_ (.A1(_21920_),
    .A2(net1833),
    .B(_22070_),
    .Y(_03157_));
 AND2x2_ASAP7_75t_R _32740_ (.A(_03157_),
    .B(_02728_),
    .Y(_03158_));
 NOR2x1_ASAP7_75t_R _32741_ (.A(net2293),
    .B(_22077_),
    .Y(_03159_));
 INVx1_ASAP7_75t_R _32742_ (.A(_02723_),
    .Y(_03160_));
 NOR2x1_ASAP7_75t_R _32743_ (.A(_03159_),
    .B(_03160_),
    .Y(_03161_));
 AND4x1_ASAP7_75t_R _32744_ (.A(_03153_),
    .B(_03156_),
    .C(_03158_),
    .D(_03161_),
    .Y(_03162_));
 NAND2x1_ASAP7_75t_R _32745_ (.A(_03150_),
    .B(_03162_),
    .Y(_03163_));
 NAND2x2_ASAP7_75t_R _32746_ (.A(_01079_),
    .B(net3167),
    .Y(_03164_));
 NAND2x1_ASAP7_75t_R _32747_ (.A(_03147_),
    .B(_01079_),
    .Y(_03165_));
 NAND2x1_ASAP7_75t_R _32748_ (.A(_03164_),
    .B(_03165_),
    .Y(_03166_));
 OA21x2_ASAP7_75t_R _32749_ (.A1(_22003_),
    .A2(_22053_),
    .B(_01079_),
    .Y(_03167_));
 NOR2x1_ASAP7_75t_R _32750_ (.A(net3152),
    .B(_22024_),
    .Y(_03168_));
 OR3x1_ASAP7_75t_R _32751_ (.A(_03166_),
    .B(_03167_),
    .C(_03168_),
    .Y(_03169_));
 NOR2x1_ASAP7_75t_R _32752_ (.A(_01072_),
    .B(_21995_),
    .Y(_03170_));
 AO21x1_ASAP7_75t_R _32753_ (.A1(net2802),
    .A2(_01073_),
    .B(_03170_),
    .Y(_03171_));
 NAND2x1_ASAP7_75t_R _32754_ (.A(net1259),
    .B(_01073_),
    .Y(_03172_));
 AO21x1_ASAP7_75t_R _32755_ (.A1(_22018_),
    .A2(_22019_),
    .B(_01072_),
    .Y(_03173_));
 NAND2x1_ASAP7_75t_R _32756_ (.A(_03172_),
    .B(_03173_),
    .Y(_03174_));
 NOR2x1_ASAP7_75t_R _32757_ (.A(_01072_),
    .B(net2294),
    .Y(_03175_));
 OR3x1_ASAP7_75t_R _32758_ (.A(_03171_),
    .B(_03174_),
    .C(_03175_),
    .Y(_03176_));
 NOR2x1_ASAP7_75t_R _32759_ (.A(_03176_),
    .B(_03169_),
    .Y(_03177_));
 AO21x1_ASAP7_75t_R _32760_ (.A1(net3155),
    .A2(_21890_),
    .B(_22091_),
    .Y(_03178_));
 OA21x2_ASAP7_75t_R _32761_ (.A1(net2420),
    .A2(_22091_),
    .B(_03178_),
    .Y(_03179_));
 AO21x1_ASAP7_75t_R _32762_ (.A1(net2298),
    .A2(_21997_),
    .B(_22091_),
    .Y(_03180_));
 INVx1_ASAP7_75t_R _32763_ (.A(_03180_),
    .Y(_03181_));
 OA211x2_ASAP7_75t_R _32764_ (.A1(_21887_),
    .A2(net1049),
    .B(_22092_),
    .C(_21926_),
    .Y(_03182_));
 NOR2x1_ASAP7_75t_R _32765_ (.A(_03181_),
    .B(_03182_),
    .Y(_03183_));
 NAND2x1_ASAP7_75t_R _32766_ (.A(_03179_),
    .B(_03183_),
    .Y(_03184_));
 OA21x2_ASAP7_75t_R _32767_ (.A1(_21909_),
    .A2(_21955_),
    .B(_02266_),
    .Y(_03185_));
 OA21x2_ASAP7_75t_R _32768_ (.A1(_22054_),
    .A2(_02269_),
    .B(_02266_),
    .Y(_03186_));
 OA21x2_ASAP7_75t_R _32769_ (.A1(_22083_),
    .A2(_02286_),
    .B(_02266_),
    .Y(_03187_));
 AOI211x1_ASAP7_75t_R _32770_ (.A1(net1139),
    .A2(_21876_),
    .B(_21895_),
    .C(_22100_),
    .Y(_03188_));
 OR4x1_ASAP7_75t_R _32771_ (.A(_03185_),
    .B(_03186_),
    .C(_03187_),
    .D(_03188_),
    .Y(_03189_));
 NOR2x1_ASAP7_75t_R _32772_ (.A(_03184_),
    .B(_03189_),
    .Y(_03190_));
 NAND2x1_ASAP7_75t_R _32773_ (.A(_03177_),
    .B(_03190_),
    .Y(_03191_));
 NOR2x1_ASAP7_75t_R _32774_ (.A(_03163_),
    .B(_03191_),
    .Y(_03192_));
 NAND2x2_ASAP7_75t_R _32775_ (.A(_03137_),
    .B(_03192_),
    .Y(_03193_));
 AO21x1_ASAP7_75t_R _32776_ (.A1(net2368),
    .A2(net2062),
    .B(_01505_),
    .Y(_03194_));
 AO21x1_ASAP7_75t_R _32777_ (.A1(_01699_),
    .A2(_01600_),
    .B(_01505_),
    .Y(_03195_));
 NAND2x2_ASAP7_75t_R _32778_ (.A(net1898),
    .B(net1576),
    .Y(_03196_));
 AO21x1_ASAP7_75t_R _32779_ (.A1(_03196_),
    .A2(_01590_),
    .B(_01505_),
    .Y(_03197_));
 AND3x1_ASAP7_75t_R _32780_ (.A(_03194_),
    .B(_03195_),
    .C(_03197_),
    .Y(_03198_));
 INVx1_ASAP7_75t_R _32781_ (.A(_01661_),
    .Y(_03199_));
 AO21x1_ASAP7_75t_R _32782_ (.A1(_01678_),
    .A2(_01674_),
    .B(net2334),
    .Y(_03200_));
 NAND2x1_ASAP7_75t_R _32783_ (.A(_01680_),
    .B(_01657_),
    .Y(_03201_));
 AND3x1_ASAP7_75t_R _32784_ (.A(_03199_),
    .B(_03200_),
    .C(_03201_),
    .Y(_03202_));
 AND2x2_ASAP7_75t_R _32785_ (.A(_03198_),
    .B(_03202_),
    .Y(_03203_));
 AO21x1_ASAP7_75t_R _32786_ (.A1(net3267),
    .A2(net1612),
    .B(_01624_),
    .Y(_03204_));
 NOR2x1_ASAP7_75t_R _32787_ (.A(_01624_),
    .B(_01699_),
    .Y(_03205_));
 INVx1_ASAP7_75t_R _32788_ (.A(_03205_),
    .Y(_03206_));
 AND2x2_ASAP7_75t_R _32789_ (.A(_03204_),
    .B(_03206_),
    .Y(_03207_));
 OA21x2_ASAP7_75t_R _32790_ (.A1(_01624_),
    .A2(net1457),
    .B(_03207_),
    .Y(_03208_));
 NAND2x1_ASAP7_75t_R _32791_ (.A(_02447_),
    .B(_01637_),
    .Y(_03209_));
 NAND2x1_ASAP7_75t_R _32792_ (.A(_01680_),
    .B(_01637_),
    .Y(_03210_));
 OA211x2_ASAP7_75t_R _32793_ (.A1(net2746),
    .A2(net2572),
    .B(_03209_),
    .C(_03210_),
    .Y(_03211_));
 NAND3x2_ASAP7_75t_R _32794_ (.B(_03208_),
    .C(_03211_),
    .Y(_03212_),
    .A(_03203_));
 AO21x1_ASAP7_75t_R _32795_ (.A1(_01670_),
    .A2(_01590_),
    .B(_01586_),
    .Y(_03213_));
 AO21x1_ASAP7_75t_R _32796_ (.A1(_01612_),
    .A2(_01540_),
    .B(net2348),
    .Y(_03214_));
 AND2x2_ASAP7_75t_R _32797_ (.A(_03213_),
    .B(_03214_),
    .Y(_03215_));
 NAND2x1_ASAP7_75t_R _32798_ (.A(_02425_),
    .B(_02829_),
    .Y(_03216_));
 NAND3x1_ASAP7_75t_R _32799_ (.A(_03215_),
    .B(_03216_),
    .C(_02438_),
    .Y(_03217_));
 AO21x1_ASAP7_75t_R _32800_ (.A1(net3261),
    .A2(net1605),
    .B(net2275),
    .Y(_03218_));
 OA21x2_ASAP7_75t_R _32801_ (.A1(net1457),
    .A2(net2275),
    .B(_03218_),
    .Y(_03219_));
 AO21x1_ASAP7_75t_R _32802_ (.A1(net2368),
    .A2(net1613),
    .B(net2275),
    .Y(_03220_));
 NAND3x1_ASAP7_75t_R _32803_ (.A(_03219_),
    .B(_02826_),
    .C(_03220_),
    .Y(_03221_));
 NOR2x1_ASAP7_75t_R _32804_ (.A(_03217_),
    .B(_03221_),
    .Y(_03222_));
 AO21x1_ASAP7_75t_R _32805_ (.A1(net3255),
    .A2(_01644_),
    .B(_01543_),
    .Y(_03223_));
 OA21x2_ASAP7_75t_R _32806_ (.A1(_02419_),
    .A2(_01543_),
    .B(_03223_),
    .Y(_03224_));
 AO21x1_ASAP7_75t_R _32807_ (.A1(net2368),
    .A2(net1612),
    .B(_01543_),
    .Y(_03225_));
 NAND3x1_ASAP7_75t_R _32808_ (.A(_03224_),
    .B(_02816_),
    .C(_03225_),
    .Y(_03226_));
 AO21x1_ASAP7_75t_R _32809_ (.A1(_01689_),
    .A2(_02372_),
    .B(_01571_),
    .Y(_03227_));
 NAND2x1_ASAP7_75t_R _32810_ (.A(_02456_),
    .B(_03227_),
    .Y(_03228_));
 NOR2x1_ASAP7_75t_R _32811_ (.A(net2524),
    .B(_01571_),
    .Y(_03229_));
 OA21x2_ASAP7_75t_R _32812_ (.A1(_02460_),
    .A2(_01680_),
    .B(_01565_),
    .Y(_03230_));
 OR3x1_ASAP7_75t_R _32813_ (.A(_03228_),
    .B(_03229_),
    .C(_03230_),
    .Y(_03231_));
 NOR2x1_ASAP7_75t_R _32814_ (.A(_03226_),
    .B(_03231_),
    .Y(_03232_));
 NAND2x1_ASAP7_75t_R _32815_ (.A(_03222_),
    .B(_03232_),
    .Y(_03233_));
 NOR2x2_ASAP7_75t_R _32816_ (.A(_03212_),
    .B(_03233_),
    .Y(_03234_));
 AO21x1_ASAP7_75t_R _32817_ (.A1(net2572),
    .A2(_02804_),
    .B(_01685_),
    .Y(_03235_));
 AO21x1_ASAP7_75t_R _32818_ (.A1(net1104),
    .A2(_01612_),
    .B(_01685_),
    .Y(_03236_));
 NAND2x1_ASAP7_75t_R _32819_ (.A(_01511_),
    .B(_01696_),
    .Y(_03237_));
 NAND3x1_ASAP7_75t_R _32820_ (.A(_03235_),
    .B(_03236_),
    .C(_03237_),
    .Y(_03238_));
 INVx1_ASAP7_75t_R _32821_ (.A(_03238_),
    .Y(_03239_));
 AO21x1_ASAP7_75t_R _32822_ (.A1(net2367),
    .A2(net1612),
    .B(_01701_),
    .Y(_03240_));
 AND2x2_ASAP7_75t_R _32823_ (.A(_03240_),
    .B(_02841_),
    .Y(_03241_));
 AO21x1_ASAP7_75t_R _32824_ (.A1(_01670_),
    .A2(_02361_),
    .B(_01701_),
    .Y(_03242_));
 OA21x2_ASAP7_75t_R _32825_ (.A1(_01644_),
    .A2(_01701_),
    .B(_03242_),
    .Y(_03243_));
 AND3x1_ASAP7_75t_R _32826_ (.A(_03239_),
    .B(_03241_),
    .C(_03243_),
    .Y(_03244_));
 AO21x1_ASAP7_75t_R _32827_ (.A1(net2572),
    .A2(net2254),
    .B(_01668_),
    .Y(_03245_));
 AO21x1_ASAP7_75t_R _32828_ (.A1(net2818),
    .A2(net2539),
    .B(_01668_),
    .Y(_03246_));
 NOR2x1_ASAP7_75t_R _32829_ (.A(_02372_),
    .B(_01668_),
    .Y(_03247_));
 INVx1_ASAP7_75t_R _32830_ (.A(_03247_),
    .Y(_03248_));
 AND3x1_ASAP7_75t_R _32831_ (.A(_03245_),
    .B(_03246_),
    .C(_03248_),
    .Y(_03249_));
 AO21x1_ASAP7_75t_R _32832_ (.A1(net3261),
    .A2(_01590_),
    .B(_01675_),
    .Y(_03250_));
 AO21x1_ASAP7_75t_R _32833_ (.A1(net1104),
    .A2(net2539),
    .B(_01675_),
    .Y(_03251_));
 NAND2x2_ASAP7_75t_R _32834_ (.A(_02461_),
    .B(_01681_),
    .Y(_03252_));
 AND3x1_ASAP7_75t_R _32835_ (.A(_03250_),
    .B(_03251_),
    .C(_03252_),
    .Y(_03253_));
 AOI211x1_ASAP7_75t_R _32836_ (.A1(net1120),
    .A2(_01494_),
    .B(net2733),
    .C(net2378),
    .Y(_03254_));
 OA21x2_ASAP7_75t_R _32837_ (.A1(_02457_),
    .A2(_01526_),
    .B(_01681_),
    .Y(_03255_));
 NOR2x1_ASAP7_75t_R _32838_ (.A(_03254_),
    .B(_03255_),
    .Y(_03256_));
 AND3x1_ASAP7_75t_R _32839_ (.A(_03249_),
    .B(_03253_),
    .C(_03256_),
    .Y(_03257_));
 NAND2x1_ASAP7_75t_R _32840_ (.A(_03244_),
    .B(_03257_),
    .Y(_03258_));
 INVx2_ASAP7_75t_R _32841_ (.A(_01540_),
    .Y(_03259_));
 NOR2x1_ASAP7_75t_R _32842_ (.A(_01590_),
    .B(_01707_),
    .Y(_03260_));
 AO21x1_ASAP7_75t_R _32843_ (.A1(_03259_),
    .A2(_01711_),
    .B(_03260_),
    .Y(_03261_));
 NAND2x1_ASAP7_75t_R _32844_ (.A(_01526_),
    .B(_01711_),
    .Y(_03262_));
 INVx1_ASAP7_75t_R _32845_ (.A(_03262_),
    .Y(_03263_));
 OA21x2_ASAP7_75t_R _32846_ (.A1(_02447_),
    .A2(_02424_),
    .B(_01711_),
    .Y(_03264_));
 OR3x1_ASAP7_75t_R _32847_ (.A(_03261_),
    .B(_03263_),
    .C(_03264_),
    .Y(_03265_));
 AO21x1_ASAP7_75t_R _32848_ (.A1(_01598_),
    .A2(_01600_),
    .B(_01715_),
    .Y(_03266_));
 OA21x2_ASAP7_75t_R _32849_ (.A1(net2570),
    .A2(_01715_),
    .B(_03266_),
    .Y(_03267_));
 NOR2x1_ASAP7_75t_R _32850_ (.A(net2777),
    .B(_01501_),
    .Y(_03268_));
 INVx1_ASAP7_75t_R _32851_ (.A(_01592_),
    .Y(_03269_));
 NAND2x1_ASAP7_75t_R _32852_ (.A(_03268_),
    .B(_03269_),
    .Y(_03270_));
 NOR2x1_ASAP7_75t_R _32853_ (.A(_00634_),
    .B(_03270_),
    .Y(_03271_));
 AOI211x1_ASAP7_75t_R _32854_ (.A1(_01491_),
    .A2(_01720_),
    .B(_03271_),
    .C(_02394_),
    .Y(_03272_));
 NAND2x1_ASAP7_75t_R _32855_ (.A(_03267_),
    .B(_03272_),
    .Y(_03273_));
 NOR2x2_ASAP7_75t_R _32856_ (.A(_03265_),
    .B(_03273_),
    .Y(_03274_));
 AO21x1_ASAP7_75t_R _32857_ (.A1(net1613),
    .A2(_01674_),
    .B(_01728_),
    .Y(_03275_));
 AO21x1_ASAP7_75t_R _32858_ (.A1(_01691_),
    .A2(_01699_),
    .B(_01728_),
    .Y(_03276_));
 NAND2x1_ASAP7_75t_R _32859_ (.A(_03275_),
    .B(_03276_),
    .Y(_03277_));
 INVx1_ASAP7_75t_R _32860_ (.A(_03277_),
    .Y(_03278_));
 OA21x2_ASAP7_75t_R _32861_ (.A1(_01562_),
    .A2(_03269_),
    .B(_02388_),
    .Y(_03279_));
 OA211x2_ASAP7_75t_R _32862_ (.A1(_01498_),
    .A2(net1263),
    .B(_02388_),
    .C(net1576),
    .Y(_03280_));
 NOR2x1_ASAP7_75t_R _32863_ (.A(_03279_),
    .B(_03280_),
    .Y(_03281_));
 NAND2x1_ASAP7_75t_R _32864_ (.A(_03278_),
    .B(_03281_),
    .Y(_03282_));
 OAI21x1_ASAP7_75t_R _32865_ (.A1(_01689_),
    .A2(_01735_),
    .B(_01736_),
    .Y(_03283_));
 AO21x1_ASAP7_75t_R _32866_ (.A1(net3136),
    .A2(_02419_),
    .B(_01735_),
    .Y(_03284_));
 NAND2x1_ASAP7_75t_R _32867_ (.A(_01746_),
    .B(_03284_),
    .Y(_03285_));
 AO21x1_ASAP7_75t_R _32868_ (.A1(_02447_),
    .A2(_01737_),
    .B(_01739_),
    .Y(_03286_));
 OR3x1_ASAP7_75t_R _32869_ (.A(_03283_),
    .B(_03285_),
    .C(_03286_),
    .Y(_03287_));
 NOR2x1_ASAP7_75t_R _32870_ (.A(_03282_),
    .B(_03287_),
    .Y(_03288_));
 NAND2x2_ASAP7_75t_R _32871_ (.A(_03274_),
    .B(_03288_),
    .Y(_03289_));
 NOR2x2_ASAP7_75t_R _32872_ (.A(_03258_),
    .B(_03289_),
    .Y(_03290_));
 NAND2x2_ASAP7_75t_R _32873_ (.A(_03234_),
    .B(_03290_),
    .Y(_03291_));
 XNOR2x2_ASAP7_75t_R _32874_ (.A(_03193_),
    .B(_03291_),
    .Y(_03292_));
 OAI22x1_ASAP7_75t_R _32875_ (.A1(_01138_),
    .A2(_01308_),
    .B1(net1266),
    .B2(net3154),
    .Y(_03293_));
 AOI211x1_ASAP7_75t_R _32876_ (.A1(_01233_),
    .A2(_01315_),
    .B(_03293_),
    .C(_01429_),
    .Y(_03294_));
 NAND2x1_ASAP7_75t_R _32877_ (.A(_01327_),
    .B(_01234_),
    .Y(_03295_));
 OAI21x1_ASAP7_75t_R _32878_ (.A1(net1266),
    .A2(_01170_),
    .B(_03295_),
    .Y(_03296_));
 NAND2x1_ASAP7_75t_R _32879_ (.A(net1684),
    .B(net1971),
    .Y(_03297_));
 AO21x1_ASAP7_75t_R _32880_ (.A1(_01303_),
    .A2(net938),
    .B(_01170_),
    .Y(_03298_));
 OAI21x1_ASAP7_75t_R _32881_ (.A1(_01229_),
    .A2(_03297_),
    .B(_03298_),
    .Y(_03299_));
 NOR2x1_ASAP7_75t_R _32882_ (.A(_03296_),
    .B(_03299_),
    .Y(_03300_));
 NAND2x1_ASAP7_75t_R _32883_ (.A(_03294_),
    .B(_03300_),
    .Y(_03301_));
 AO21x1_ASAP7_75t_R _32884_ (.A1(_01474_),
    .A2(_01163_),
    .B(_01410_),
    .Y(_03302_));
 OAI21x1_ASAP7_75t_R _32885_ (.A1(_01178_),
    .A2(_03073_),
    .B(_01386_),
    .Y(_03303_));
 NOR2x1_ASAP7_75t_R _32886_ (.A(_03302_),
    .B(_03303_),
    .Y(_03304_));
 INVx1_ASAP7_75t_R _32887_ (.A(_01465_),
    .Y(_03305_));
 AOI211x1_ASAP7_75t_R _32888_ (.A1(_01244_),
    .A2(net1277),
    .B(_03305_),
    .C(_01439_),
    .Y(_03306_));
 NAND2x1_ASAP7_75t_R _32889_ (.A(_03304_),
    .B(_03306_),
    .Y(_03307_));
 NOR2x1_ASAP7_75t_R _32890_ (.A(_03301_),
    .B(_03307_),
    .Y(_03308_));
 OAI22x1_ASAP7_75t_R _32891_ (.A1(net3145),
    .A2(_01153_),
    .B1(_01215_),
    .B2(_01453_),
    .Y(_03309_));
 NAND2x1_ASAP7_75t_R _32892_ (.A(_01418_),
    .B(_01472_),
    .Y(_03310_));
 NOR2x1_ASAP7_75t_R _32893_ (.A(_03309_),
    .B(_03310_),
    .Y(_03311_));
 NAND2x1_ASAP7_75t_R _32894_ (.A(_01423_),
    .B(_01389_),
    .Y(_03312_));
 NAND2x1_ASAP7_75t_R _32895_ (.A(_01327_),
    .B(_01197_),
    .Y(_03313_));
 OAI21x1_ASAP7_75t_R _32896_ (.A1(net1277),
    .A2(_02590_),
    .B(_03313_),
    .Y(_03314_));
 NOR2x1_ASAP7_75t_R _32897_ (.A(_03312_),
    .B(_03314_),
    .Y(_03315_));
 NAND2x1_ASAP7_75t_R _32898_ (.A(_03311_),
    .B(_03315_),
    .Y(_03316_));
 NOR2x1_ASAP7_75t_R _32899_ (.A(net2325),
    .B(net2872),
    .Y(_03317_));
 AOI22x1_ASAP7_75t_R _32900_ (.A1(_01337_),
    .A2(_01374_),
    .B1(_01163_),
    .B2(_03317_),
    .Y(_03318_));
 AOI22x1_ASAP7_75t_R _32901_ (.A1(_01251_),
    .A2(_01374_),
    .B1(_01337_),
    .B2(_01180_),
    .Y(_03319_));
 NAND2x1_ASAP7_75t_R _32902_ (.A(_03318_),
    .B(_03319_),
    .Y(_03320_));
 NOR2x1_ASAP7_75t_R _32903_ (.A(_00585_),
    .B(_01099_),
    .Y(_03321_));
 AOI22x1_ASAP7_75t_R _32904_ (.A1(_01351_),
    .A2(_01109_),
    .B1(_02061_),
    .B2(_03321_),
    .Y(_03322_));
 AOI22x1_ASAP7_75t_R _32905_ (.A1(_01416_),
    .A2(net1968),
    .B1(_02593_),
    .B2(_01405_),
    .Y(_03323_));
 NAND2x1_ASAP7_75t_R _32906_ (.A(_03322_),
    .B(_03323_),
    .Y(_03324_));
 NOR2x1_ASAP7_75t_R _32907_ (.A(_03320_),
    .B(_03324_),
    .Y(_03325_));
 AO21x1_ASAP7_75t_R _32908_ (.A1(_01306_),
    .A2(_01153_),
    .B(net3417),
    .Y(_03326_));
 NAND2x1_ASAP7_75t_R _32909_ (.A(_03326_),
    .B(_01412_),
    .Y(_03327_));
 AOI21x1_ASAP7_75t_R _32910_ (.A1(_01218_),
    .A2(_01305_),
    .B(_01402_),
    .Y(_03328_));
 OR3x1_ASAP7_75t_R _32911_ (.A(_01308_),
    .B(net2649),
    .C(_01178_),
    .Y(_03329_));
 NAND2x1_ASAP7_75t_R _32912_ (.A(_03328_),
    .B(_03329_),
    .Y(_03330_));
 NOR2x1_ASAP7_75t_R _32913_ (.A(_03327_),
    .B(_03330_),
    .Y(_03331_));
 NAND2x1_ASAP7_75t_R _32914_ (.A(_03325_),
    .B(_03331_),
    .Y(_03332_));
 NOR2x1_ASAP7_75t_R _32915_ (.A(_03316_),
    .B(_03332_),
    .Y(_03333_));
 NAND2x1_ASAP7_75t_R _32916_ (.A(_03308_),
    .B(_03333_),
    .Y(_03334_));
 NOR2x2_ASAP7_75t_R _32917_ (.A(_01404_),
    .B(_01451_),
    .Y(_03335_));
 AO21x1_ASAP7_75t_R _32918_ (.A1(net1572),
    .A2(net1122),
    .B(net3154),
    .Y(_03336_));
 NAND3x2_ASAP7_75t_R _32919_ (.B(_02013_),
    .C(_03336_),
    .Y(_03337_),
    .A(_03335_));
 NAND2x1_ASAP7_75t_R _32920_ (.A(_01186_),
    .B(_01097_),
    .Y(_03338_));
 NAND2x1_ASAP7_75t_R _32921_ (.A(net2443),
    .B(_01351_),
    .Y(_03339_));
 OAI21x1_ASAP7_75t_R _32922_ (.A1(_01156_),
    .A2(_03338_),
    .B(_03339_),
    .Y(_03340_));
 INVx1_ASAP7_75t_R _32923_ (.A(_01257_),
    .Y(_03341_));
 OAI21x1_ASAP7_75t_R _32924_ (.A1(_01112_),
    .A2(_03341_),
    .B(_01266_),
    .Y(_03342_));
 NOR2x1_ASAP7_75t_R _32925_ (.A(_03340_),
    .B(_03342_),
    .Y(_03343_));
 INVx1_ASAP7_75t_R _32926_ (.A(_01438_),
    .Y(_03344_));
 NAND2x1_ASAP7_75t_R _32927_ (.A(_01471_),
    .B(_01458_),
    .Y(_03345_));
 NOR2x1_ASAP7_75t_R _32928_ (.A(_03344_),
    .B(_03345_),
    .Y(_03346_));
 NAND2x1_ASAP7_75t_R _32929_ (.A(_03343_),
    .B(_03346_),
    .Y(_03347_));
 NOR2x2_ASAP7_75t_R _32930_ (.A(_03337_),
    .B(_03347_),
    .Y(_03348_));
 OAI22x1_ASAP7_75t_R _32931_ (.A1(net938),
    .A2(_01334_),
    .B1(net3240),
    .B2(_01259_),
    .Y(_03349_));
 OAI22x1_ASAP7_75t_R _32932_ (.A1(net3320),
    .A2(net3240),
    .B1(net1266),
    .B2(_01229_),
    .Y(_03350_));
 NOR2x1_ASAP7_75t_R _32933_ (.A(_03349_),
    .B(_03350_),
    .Y(_03351_));
 OAI22x1_ASAP7_75t_R _32934_ (.A1(net938),
    .A2(net3154),
    .B1(_01306_),
    .B2(_01229_),
    .Y(_03352_));
 OA21x2_ASAP7_75t_R _32935_ (.A1(_01268_),
    .A2(_01374_),
    .B(_01329_),
    .Y(_03353_));
 NOR2x1_ASAP7_75t_R _32936_ (.A(_03352_),
    .B(_03353_),
    .Y(_03354_));
 NAND2x1_ASAP7_75t_R _32937_ (.A(_03351_),
    .B(_03354_),
    .Y(_03355_));
 OAI22x1_ASAP7_75t_R _32938_ (.A1(net3145),
    .A2(_01303_),
    .B1(_01133_),
    .B2(net2723),
    .Y(_03356_));
 OAI21x1_ASAP7_75t_R _32939_ (.A1(net1122),
    .A2(_01133_),
    .B(_01460_),
    .Y(_03357_));
 NOR2x1_ASAP7_75t_R _32940_ (.A(_03356_),
    .B(_03357_),
    .Y(_03358_));
 OAI22x1_ASAP7_75t_R _32941_ (.A1(net2651),
    .A2(net3417),
    .B1(net1158),
    .B2(_01133_),
    .Y(_03359_));
 NAND2x1_ASAP7_75t_R _32942_ (.A(_01383_),
    .B(_02635_),
    .Y(_03360_));
 NOR2x1_ASAP7_75t_R _32943_ (.A(_03359_),
    .B(_03360_),
    .Y(_03361_));
 NAND2x1_ASAP7_75t_R _32944_ (.A(_03358_),
    .B(_03361_),
    .Y(_03362_));
 NOR2x2_ASAP7_75t_R _32945_ (.A(_03355_),
    .B(_03362_),
    .Y(_03363_));
 OA21x2_ASAP7_75t_R _32946_ (.A1(_01328_),
    .A2(_01209_),
    .B(_01218_),
    .Y(_03364_));
 OAI22x1_ASAP7_75t_R _32947_ (.A1(net1158),
    .A2(net3154),
    .B1(net3145),
    .B2(net938),
    .Y(_03365_));
 NOR2x1_ASAP7_75t_R _32948_ (.A(_03364_),
    .B(_03365_),
    .Y(_03366_));
 NOR2x1_ASAP7_75t_R _32949_ (.A(_01229_),
    .B(net2651),
    .Y(_03367_));
 AOI211x1_ASAP7_75t_R _32950_ (.A1(_01288_),
    .A2(_02600_),
    .B(_01440_),
    .C(_03367_),
    .Y(_03368_));
 NAND2x1_ASAP7_75t_R _32951_ (.A(_03366_),
    .B(_03368_),
    .Y(_03369_));
 AND2x2_ASAP7_75t_R _32952_ (.A(_02683_),
    .B(_02015_),
    .Y(_03370_));
 AOI21x1_ASAP7_75t_R _32953_ (.A1(_01234_),
    .A2(net2443),
    .B(_01395_),
    .Y(_03371_));
 AO21x1_ASAP7_75t_R _32954_ (.A1(net3320),
    .A2(net1122),
    .B(net2460),
    .Y(_03372_));
 NAND3x2_ASAP7_75t_R _32955_ (.B(_03371_),
    .C(_03372_),
    .Y(_03373_),
    .A(_03370_));
 NOR2x2_ASAP7_75t_R _32956_ (.A(_03369_),
    .B(_03373_),
    .Y(_03374_));
 NAND3x2_ASAP7_75t_R _32957_ (.B(_03363_),
    .C(_03374_),
    .Y(_03375_),
    .A(_03348_));
 NOR2x2_ASAP7_75t_R _32958_ (.A(_03334_),
    .B(_03375_),
    .Y(_03376_));
 XOR2x2_ASAP7_75t_R _32959_ (.A(_02692_),
    .B(_03376_),
    .Y(_03377_));
 XOR2x1_ASAP7_75t_R _32960_ (.A(_03292_),
    .Y(_03378_),
    .B(_03377_));
 NAND2x1_ASAP7_75t_R _32961_ (.A(_03096_),
    .B(_03378_),
    .Y(_03379_));
 XOR2x2_ASAP7_75t_R _32962_ (.A(_03001_),
    .B(_01987_),
    .Y(_03380_));
 XOR2x1_ASAP7_75t_R _32963_ (.A(_03380_),
    .Y(_03381_),
    .B(net2793));
 XOR2x2_ASAP7_75t_R _32964_ (.A(_02692_),
    .B(_01480_),
    .Y(_03382_));
 XOR2x1_ASAP7_75t_R _32965_ (.A(_03292_),
    .Y(_03383_),
    .B(_03382_));
 NAND2x1_ASAP7_75t_R _32966_ (.A(_03381_),
    .B(_03383_),
    .Y(_03384_));
 AOI21x1_ASAP7_75t_R _32967_ (.A1(_03379_),
    .A2(_03384_),
    .B(_18753_),
    .Y(_03385_));
 OAI21x1_ASAP7_75t_R _32968_ (.A1(_02904_),
    .A2(_03385_),
    .B(_00481_),
    .Y(_03386_));
 AND2x2_ASAP7_75t_R _32969_ (.A(_18753_),
    .B(_00880_),
    .Y(_03387_));
 XOR2x1_ASAP7_75t_R _32970_ (.A(_03377_),
    .Y(_03388_),
    .B(net2793));
 XOR2x1_ASAP7_75t_R _32971_ (.A(_03292_),
    .Y(_03389_),
    .B(_03380_));
 NAND2x1_ASAP7_75t_R _32972_ (.A(_03388_),
    .B(_03389_),
    .Y(_03390_));
 XOR2x1_ASAP7_75t_R _32973_ (.A(_03377_),
    .Y(_03391_),
    .B(_03091_));
 XNOR2x1_ASAP7_75t_R _32974_ (.B(_03292_),
    .Y(_03392_),
    .A(_03380_));
 NAND2x1_ASAP7_75t_R _32975_ (.A(_03391_),
    .B(_03392_),
    .Y(_03393_));
 TAPCELL_ASAP7_75t_R PHY_539 ();
 AOI21x1_ASAP7_75t_R _32977_ (.A1(_03390_),
    .A2(_03393_),
    .B(_18753_),
    .Y(_03395_));
 INVx1_ASAP7_75t_R _32978_ (.A(_00481_),
    .Y(_03396_));
 OAI21x1_ASAP7_75t_R _32979_ (.A1(_03387_),
    .A2(_03395_),
    .B(_03396_),
    .Y(_03397_));
 NAND2x2_ASAP7_75t_R _32980_ (.A(_03386_),
    .B(_03397_),
    .Y(_00116_));
 AND2x2_ASAP7_75t_R _32981_ (.A(net390),
    .B(_00879_),
    .Y(_03398_));
 XOR2x2_ASAP7_75t_R _32982_ (.A(_03090_),
    .B(_01480_),
    .Y(_03399_));
 AO21x1_ASAP7_75t_R _32983_ (.A1(_01630_),
    .A2(net3149),
    .B(net2794),
    .Y(_03400_));
 AND3x1_ASAP7_75t_R _32984_ (.A(_03213_),
    .B(_03400_),
    .C(_01596_),
    .Y(_03401_));
 OA21x2_ASAP7_75t_R _32985_ (.A1(net3147),
    .A2(_01688_),
    .B(_02825_),
    .Y(_03402_));
 AOI21x1_ASAP7_75t_R _32986_ (.A1(net3255),
    .A2(net3265),
    .B(_01603_),
    .Y(_03403_));
 NOR3x1_ASAP7_75t_R _32987_ (.A(_03402_),
    .B(_03403_),
    .C(_02441_),
    .Y(_03404_));
 AO21x1_ASAP7_75t_R _32988_ (.A1(_01689_),
    .A2(_01600_),
    .B(net2348),
    .Y(_03405_));
 OA21x2_ASAP7_75t_R _32989_ (.A1(net1613),
    .A2(net2348),
    .B(_03405_),
    .Y(_03406_));
 NAND3x1_ASAP7_75t_R _32990_ (.A(_03401_),
    .B(_03404_),
    .C(_03406_),
    .Y(_03407_));
 AO21x1_ASAP7_75t_R _32991_ (.A1(_02419_),
    .A2(net2728),
    .B(_01543_),
    .Y(_03408_));
 NAND2x1_ASAP7_75t_R _32992_ (.A(_01575_),
    .B(_01550_),
    .Y(_03409_));
 AND4x1_ASAP7_75t_R _32993_ (.A(_01558_),
    .B(_03408_),
    .C(_03409_),
    .D(_02817_),
    .Y(_03410_));
 AO21x1_ASAP7_75t_R _32994_ (.A1(_01565_),
    .A2(_01635_),
    .B(_01578_),
    .Y(_03411_));
 AOI211x1_ASAP7_75t_R _32995_ (.A1(_01565_),
    .A2(_02457_),
    .B(_03411_),
    .C(_02455_),
    .Y(_03412_));
 NAND2x1_ASAP7_75t_R _32996_ (.A(_03410_),
    .B(_03412_),
    .Y(_03413_));
 NOR2x1_ASAP7_75t_R _32997_ (.A(_03407_),
    .B(_03413_),
    .Y(_03414_));
 INVx2_ASAP7_75t_R _32998_ (.A(_01527_),
    .Y(_03415_));
 NOR2x1_ASAP7_75t_R _32999_ (.A(net2572),
    .B(_01505_),
    .Y(_03416_));
 AOI21x1_ASAP7_75t_R _33000_ (.A1(_01641_),
    .A2(_01500_),
    .B(_01505_),
    .Y(_03417_));
 OR3x1_ASAP7_75t_R _33001_ (.A(_03415_),
    .B(_03416_),
    .C(_03417_),
    .Y(_03418_));
 OA21x2_ASAP7_75t_R _33002_ (.A1(_02460_),
    .A2(_01680_),
    .B(_01657_),
    .Y(_03419_));
 NOR2x1_ASAP7_75t_R _33003_ (.A(net2524),
    .B(net2334),
    .Y(_03420_));
 AOI21x1_ASAP7_75t_R _33004_ (.A1(_01600_),
    .A2(_01687_),
    .B(net2334),
    .Y(_03421_));
 OR3x1_ASAP7_75t_R _33005_ (.A(_03419_),
    .B(_03420_),
    .C(_03421_),
    .Y(_03422_));
 NOR2x1_ASAP7_75t_R _33006_ (.A(_03418_),
    .B(_03422_),
    .Y(_03423_));
 AO21x1_ASAP7_75t_R _33007_ (.A1(net3267),
    .A2(net2572),
    .B(_01636_),
    .Y(_03424_));
 AO21x1_ASAP7_75t_R _33008_ (.A1(_01670_),
    .A2(_01540_),
    .B(_01636_),
    .Y(_03425_));
 AND3x1_ASAP7_75t_R _33009_ (.A(_03424_),
    .B(_03425_),
    .C(_03209_),
    .Y(_03426_));
 AO21x1_ASAP7_75t_R _33010_ (.A1(_01641_),
    .A2(_01590_),
    .B(_01624_),
    .Y(_03427_));
 AO21x1_ASAP7_75t_R _33011_ (.A1(_01569_),
    .A2(_01540_),
    .B(_01624_),
    .Y(_03428_));
 OAI21x1_ASAP7_75t_R _33012_ (.A1(_01619_),
    .A2(_02414_),
    .B(_01621_),
    .Y(_03429_));
 NAND3x1_ASAP7_75t_R _33013_ (.A(_03427_),
    .B(_03428_),
    .C(_03429_),
    .Y(_03430_));
 INVx1_ASAP7_75t_R _33014_ (.A(_03430_),
    .Y(_03431_));
 AND2x2_ASAP7_75t_R _33015_ (.A(_03426_),
    .B(_03431_),
    .Y(_03432_));
 AND2x2_ASAP7_75t_R _33016_ (.A(_03423_),
    .B(_03432_),
    .Y(_03433_));
 NAND2x2_ASAP7_75t_R _33017_ (.A(_03414_),
    .B(_03433_),
    .Y(_03434_));
 AOI211x1_ASAP7_75t_R _33018_ (.A1(net1120),
    .A2(net1263),
    .B(net3175),
    .C(net1238),
    .Y(_03435_));
 OA21x2_ASAP7_75t_R _33019_ (.A1(_02425_),
    .A2(_02447_),
    .B(_02388_),
    .Y(_03436_));
 NOR2x2_ASAP7_75t_R _33020_ (.A(_03435_),
    .B(_03436_),
    .Y(_03437_));
 AO21x1_ASAP7_75t_R _33021_ (.A1(_01515_),
    .A2(net3130),
    .B(net2625),
    .Y(_03438_));
 AO21x1_ASAP7_75t_R _33022_ (.A1(_03438_),
    .A2(net2571),
    .B(_01735_),
    .Y(_03439_));
 AO21x1_ASAP7_75t_R _33023_ (.A1(_01592_),
    .A2(_01732_),
    .B(net3175),
    .Y(_03440_));
 NAND3x2_ASAP7_75t_R _33024_ (.B(_03439_),
    .C(_03440_),
    .Y(_03441_),
    .A(_03437_));
 NAND2x1_ASAP7_75t_R _33025_ (.A(net1263),
    .B(net3146),
    .Y(_03442_));
 AOI21x1_ASAP7_75t_R _33026_ (.A1(_03442_),
    .A2(_01598_),
    .B(_01715_),
    .Y(_03443_));
 OR2x2_ASAP7_75t_R _33027_ (.A(_03443_),
    .B(_02874_),
    .Y(_03444_));
 AOI211x1_ASAP7_75t_R _33028_ (.A1(_01498_),
    .A2(_01494_),
    .B(net3256),
    .C(net1239),
    .Y(_03445_));
 AOI21x1_ASAP7_75t_R _33029_ (.A1(net3257),
    .A2(_01711_),
    .B(_03445_),
    .Y(_03446_));
 AOI211x1_ASAP7_75t_R _33030_ (.A1(net1120),
    .A2(net1263),
    .B(_01707_),
    .C(net2071),
    .Y(_03447_));
 AOI21x1_ASAP7_75t_R _33031_ (.A1(_03259_),
    .A2(_01711_),
    .B(_03447_),
    .Y(_03448_));
 NAND2x2_ASAP7_75t_R _33032_ (.A(_03446_),
    .B(_03448_),
    .Y(_03449_));
 NOR3x2_ASAP7_75t_R _33033_ (.B(_03444_),
    .C(_03449_),
    .Y(_03450_),
    .A(_03441_));
 AO21x1_ASAP7_75t_R _33034_ (.A1(net1605),
    .A2(net1597),
    .B(_01701_),
    .Y(_03451_));
 AO21x1_ASAP7_75t_R _33035_ (.A1(net1613),
    .A2(_01600_),
    .B(_01701_),
    .Y(_03452_));
 OA211x2_ASAP7_75t_R _33036_ (.A1(_01500_),
    .A2(_01701_),
    .B(_03451_),
    .C(_03452_),
    .Y(_03453_));
 AO21x1_ASAP7_75t_R _33037_ (.A1(_01691_),
    .A2(_01699_),
    .B(_01668_),
    .Y(_03454_));
 NAND2x2_ASAP7_75t_R _33038_ (.A(_02447_),
    .B(_02368_),
    .Y(_03455_));
 NAND3x2_ASAP7_75t_R _33039_ (.B(_01672_),
    .C(_03455_),
    .Y(_03456_),
    .A(_03454_));
 AO21x1_ASAP7_75t_R _33040_ (.A1(net3135),
    .A2(net2818),
    .B(_01675_),
    .Y(_03457_));
 AO21x1_ASAP7_75t_R _33041_ (.A1(net2368),
    .A2(_01691_),
    .B(_01675_),
    .Y(_03458_));
 NAND3x2_ASAP7_75t_R _33042_ (.B(_03458_),
    .C(_03252_),
    .Y(_03459_),
    .A(_03457_));
 NOR2x2_ASAP7_75t_R _33043_ (.A(_03456_),
    .B(_03459_),
    .Y(_03460_));
 INVx1_ASAP7_75t_R _33044_ (.A(_01695_),
    .Y(_03461_));
 AND3x2_ASAP7_75t_R _33045_ (.A(_03461_),
    .B(_03237_),
    .C(_02366_),
    .Y(_03462_));
 NAND3x2_ASAP7_75t_R _33046_ (.B(_03460_),
    .C(_03462_),
    .Y(_03463_),
    .A(_03453_));
 INVx1_ASAP7_75t_R _33047_ (.A(_03463_),
    .Y(_03464_));
 NAND2x2_ASAP7_75t_R _33048_ (.A(_03450_),
    .B(_03464_),
    .Y(_03465_));
 NOR2x2_ASAP7_75t_R _33049_ (.A(_03434_),
    .B(_03465_),
    .Y(_03466_));
 XOR2x1_ASAP7_75t_R _33050_ (.A(_03399_),
    .Y(_03467_),
    .B(net3150));
 AO21x1_ASAP7_75t_R _33051_ (.A1(_01113_),
    .A2(_01138_),
    .B(net3154),
    .Y(_03468_));
 AO21x1_ASAP7_75t_R _33052_ (.A1(net1158),
    .A2(_01303_),
    .B(_01202_),
    .Y(_03469_));
 AND4x1_ASAP7_75t_R _33053_ (.A(_03468_),
    .B(_03469_),
    .C(_02636_),
    .D(_02635_),
    .Y(_03470_));
 INVx1_ASAP7_75t_R _33054_ (.A(_01259_),
    .Y(_03471_));
 AOI211x1_ASAP7_75t_R _33055_ (.A1(net1341),
    .A2(net1277),
    .B(_01221_),
    .C(net3144),
    .Y(_03472_));
 AO21x1_ASAP7_75t_R _33056_ (.A1(net1275),
    .A2(_01306_),
    .B(_01191_),
    .Y(_03473_));
 OAI21x1_ASAP7_75t_R _33057_ (.A1(net3144),
    .A2(net1158),
    .B(_03473_),
    .Y(_03474_));
 AOI211x1_ASAP7_75t_R _33058_ (.A1(_01197_),
    .A2(_03471_),
    .B(_03472_),
    .C(_03474_),
    .Y(_03475_));
 NAND2x1_ASAP7_75t_R _33059_ (.A(_03470_),
    .B(_03475_),
    .Y(_03476_));
 OA21x2_ASAP7_75t_R _33060_ (.A1(_01179_),
    .A2(_01270_),
    .B(_01234_),
    .Y(_03477_));
 OA211x2_ASAP7_75t_R _33061_ (.A1(net3142),
    .A2(net3289),
    .B(_01234_),
    .C(_01109_),
    .Y(_03478_));
 NOR2x1_ASAP7_75t_R _33062_ (.A(_03477_),
    .B(_03478_),
    .Y(_03479_));
 OA211x2_ASAP7_75t_R _33063_ (.A1(_01204_),
    .A2(_01215_),
    .B(_03051_),
    .C(_01220_),
    .Y(_03480_));
 AOI21x1_ASAP7_75t_R _33064_ (.A1(_01234_),
    .A2(_02061_),
    .B(_01235_),
    .Y(_03481_));
 NAND3x1_ASAP7_75t_R _33065_ (.A(_03479_),
    .B(_03480_),
    .C(_03481_),
    .Y(_03482_));
 NOR2x1_ASAP7_75t_R _33066_ (.A(_03482_),
    .B(_03476_),
    .Y(_03483_));
 NAND2x1_ASAP7_75t_R _33067_ (.A(_03071_),
    .B(_01144_),
    .Y(_03484_));
 AO21x1_ASAP7_75t_R _33068_ (.A1(net1828),
    .A2(_01447_),
    .B(_01133_),
    .Y(_03485_));
 AO21x1_ASAP7_75t_R _33069_ (.A1(net1158),
    .A2(_01226_),
    .B(_01133_),
    .Y(_03486_));
 NAND2x1_ASAP7_75t_R _33070_ (.A(_03485_),
    .B(_03486_),
    .Y(_03487_));
 OR3x1_ASAP7_75t_R _33071_ (.A(_02027_),
    .B(_03484_),
    .C(_03487_),
    .Y(_03488_));
 AO21x1_ASAP7_75t_R _33072_ (.A1(_01115_),
    .A2(_01138_),
    .B(_01156_),
    .Y(_03489_));
 NOR2x1_ASAP7_75t_R _33073_ (.A(net1141),
    .B(_01156_),
    .Y(_03490_));
 INVx1_ASAP7_75t_R _33074_ (.A(_03490_),
    .Y(_03491_));
 AND4x1_ASAP7_75t_R _33075_ (.A(_03489_),
    .B(_01158_),
    .C(_01167_),
    .D(_03491_),
    .Y(_03492_));
 INVx1_ASAP7_75t_R _33076_ (.A(_03492_),
    .Y(_03493_));
 OA21x2_ASAP7_75t_R _33077_ (.A1(_01328_),
    .A2(_02023_),
    .B(_01171_),
    .Y(_03494_));
 OA21x2_ASAP7_75t_R _33078_ (.A1(_01209_),
    .A2(_01270_),
    .B(_01171_),
    .Y(_03495_));
 NOR2x1_ASAP7_75t_R _33079_ (.A(net1076),
    .B(_01170_),
    .Y(_03496_));
 OR3x1_ASAP7_75t_R _33080_ (.A(_03494_),
    .B(_03495_),
    .C(_03496_),
    .Y(_03497_));
 NOR3x1_ASAP7_75t_R _33081_ (.A(_03488_),
    .B(_03493_),
    .C(_03497_),
    .Y(_03498_));
 NAND2x1_ASAP7_75t_R _33082_ (.A(_03483_),
    .B(_03498_),
    .Y(_03499_));
 AO21x1_ASAP7_75t_R _33083_ (.A1(net2717),
    .A2(net1572),
    .B(_01276_),
    .Y(_03500_));
 OA21x2_ASAP7_75t_R _33084_ (.A1(net3320),
    .A2(net3417),
    .B(_03500_),
    .Y(_03501_));
 AO21x1_ASAP7_75t_R _33085_ (.A1(net1865),
    .A2(_01447_),
    .B(_01287_),
    .Y(_03502_));
 AO21x1_ASAP7_75t_R _33086_ (.A1(_01303_),
    .A2(_01248_),
    .B(_01287_),
    .Y(_03503_));
 AND2x2_ASAP7_75t_R _33087_ (.A(_03502_),
    .B(_03503_),
    .Y(_03504_));
 AO21x1_ASAP7_75t_R _33088_ (.A1(_01228_),
    .A2(net938),
    .B(_01276_),
    .Y(_03505_));
 NAND2x1_ASAP7_75t_R _33089_ (.A(_01406_),
    .B(_01416_),
    .Y(_03506_));
 AND2x2_ASAP7_75t_R _33090_ (.A(_03505_),
    .B(_03506_),
    .Y(_03507_));
 NAND3x2_ASAP7_75t_R _33091_ (.B(_03504_),
    .C(_03507_),
    .Y(_03508_),
    .A(_03501_));
 AO21x1_ASAP7_75t_R _33092_ (.A1(net1266),
    .A2(_01303_),
    .B(_01243_),
    .Y(_03509_));
 AO21x1_ASAP7_75t_R _33093_ (.A1(net2522),
    .A2(_01259_),
    .B(_01243_),
    .Y(_03510_));
 NAND2x1_ASAP7_75t_R _33094_ (.A(net2443),
    .B(_01251_),
    .Y(_03511_));
 AND3x1_ASAP7_75t_R _33095_ (.A(_03509_),
    .B(_03510_),
    .C(_03511_),
    .Y(_03512_));
 NAND2x1_ASAP7_75t_R _33096_ (.A(_01266_),
    .B(_02056_),
    .Y(_03513_));
 OA211x2_ASAP7_75t_R _33097_ (.A1(_01106_),
    .A2(_02623_),
    .B(_01265_),
    .C(_01186_),
    .Y(_03514_));
 NOR2x1_ASAP7_75t_R _33098_ (.A(_03513_),
    .B(_03514_),
    .Y(_03515_));
 NAND2x1_ASAP7_75t_R _33099_ (.A(_03515_),
    .B(_03512_),
    .Y(_03516_));
 NOR2x2_ASAP7_75t_R _33100_ (.A(_03508_),
    .B(_03516_),
    .Y(_03517_));
 OA21x2_ASAP7_75t_R _33101_ (.A1(_01268_),
    .A2(_01160_),
    .B(_01315_),
    .Y(_03518_));
 NOR2x1_ASAP7_75t_R _33102_ (.A(_01226_),
    .B(_01308_),
    .Y(_03519_));
 OR3x2_ASAP7_75t_R _33103_ (.A(_03518_),
    .B(_02083_),
    .C(_03519_),
    .Y(_03520_));
 AO21x1_ASAP7_75t_R _33104_ (.A1(net1158),
    .A2(net938),
    .B(net2460),
    .Y(_03521_));
 INVx1_ASAP7_75t_R _33105_ (.A(_01395_),
    .Y(_03522_));
 NAND2x2_ASAP7_75t_R _33106_ (.A(_01305_),
    .B(_01329_),
    .Y(_03523_));
 NAND3x2_ASAP7_75t_R _33107_ (.B(_03522_),
    .C(_03523_),
    .Y(_03524_),
    .A(_03521_));
 OAI21x1_ASAP7_75t_R _33108_ (.A1(net1572),
    .A2(net2460),
    .B(_03019_),
    .Y(_03525_));
 NOR3x2_ASAP7_75t_R _33109_ (.B(_03524_),
    .C(_03525_),
    .Y(_03526_),
    .A(_03520_));
 OA21x2_ASAP7_75t_R _33110_ (.A1(_01204_),
    .A2(_01334_),
    .B(_01386_),
    .Y(_03527_));
 AO21x1_ASAP7_75t_R _33111_ (.A1(net2120),
    .A2(_01318_),
    .B(_01334_),
    .Y(_03528_));
 NAND2x1_ASAP7_75t_R _33112_ (.A(_01474_),
    .B(_01337_),
    .Y(_03529_));
 AND3x1_ASAP7_75t_R _33113_ (.A(_03528_),
    .B(_01372_),
    .C(_03529_),
    .Y(_03530_));
 NAND2x1_ASAP7_75t_R _33114_ (.A(_03527_),
    .B(_03530_),
    .Y(_03531_));
 AO21x1_ASAP7_75t_R _33115_ (.A1(_01113_),
    .A2(_01226_),
    .B(net3240),
    .Y(_03532_));
 OA21x2_ASAP7_75t_R _33116_ (.A1(net1158),
    .A2(net3240),
    .B(_03532_),
    .Y(_03533_));
 AO21x1_ASAP7_75t_R _33117_ (.A1(net2544),
    .A2(net1076),
    .B(_01345_),
    .Y(_03534_));
 AND3x1_ASAP7_75t_R _33118_ (.A(_03013_),
    .B(_03534_),
    .C(_01347_),
    .Y(_03535_));
 NAND2x1_ASAP7_75t_R _33119_ (.A(_03533_),
    .B(_03535_),
    .Y(_03536_));
 NOR2x2_ASAP7_75t_R _33120_ (.A(_03531_),
    .B(_03536_),
    .Y(_03537_));
 NAND3x2_ASAP7_75t_R _33121_ (.B(_03526_),
    .C(_03537_),
    .Y(_03538_),
    .A(_03517_));
 NOR2x2_ASAP7_75t_R _33122_ (.A(_03499_),
    .B(_03538_),
    .Y(_03539_));
 AO21x1_ASAP7_75t_R _33123_ (.A1(net2293),
    .A2(net1048),
    .B(_01072_),
    .Y(_03540_));
 INVx1_ASAP7_75t_R _33124_ (.A(_03170_),
    .Y(_03541_));
 NAND3x1_ASAP7_75t_R _33125_ (.A(_03540_),
    .B(_03541_),
    .C(_02715_),
    .Y(_03542_));
 INVx1_ASAP7_75t_R _33126_ (.A(_03542_),
    .Y(_03543_));
 AO21x1_ASAP7_75t_R _33127_ (.A1(_21929_),
    .A2(_21995_),
    .B(net3152),
    .Y(_03544_));
 NAND2x1_ASAP7_75t_R _33128_ (.A(_02269_),
    .B(_01079_),
    .Y(_03545_));
 AND2x2_ASAP7_75t_R _33129_ (.A(_03544_),
    .B(_03545_),
    .Y(_03546_));
 NAND2x1_ASAP7_75t_R _33130_ (.A(_21878_),
    .B(_01079_),
    .Y(_03547_));
 AND3x2_ASAP7_75t_R _33131_ (.A(_01083_),
    .B(_03547_),
    .C(_03165_),
    .Y(_03548_));
 NAND3x2_ASAP7_75t_R _33132_ (.B(_03546_),
    .C(_03548_),
    .Y(_03549_),
    .A(_03543_));
 AO21x1_ASAP7_75t_R _33133_ (.A1(_21929_),
    .A2(net3280),
    .B(net3081),
    .Y(_03550_));
 AO21x1_ASAP7_75t_R _33134_ (.A1(net3173),
    .A2(net1792),
    .B(_22100_),
    .Y(_03551_));
 NAND2x1_ASAP7_75t_R _33135_ (.A(_21909_),
    .B(_02266_),
    .Y(_03552_));
 AND3x2_ASAP7_75t_R _33136_ (.A(_03550_),
    .B(_03551_),
    .C(_03552_),
    .Y(_03553_));
 AO21x1_ASAP7_75t_R _33137_ (.A1(_21877_),
    .A2(_00550_),
    .B(net2006),
    .Y(_03554_));
 AO21x1_ASAP7_75t_R _33138_ (.A1(_03554_),
    .A2(net1829),
    .B(_22091_),
    .Y(_03555_));
 AO21x1_ASAP7_75t_R _33139_ (.A1(_22019_),
    .A2(_22098_),
    .B(_22100_),
    .Y(_03556_));
 NAND3x2_ASAP7_75t_R _33140_ (.B(_03555_),
    .C(_03556_),
    .Y(_03557_),
    .A(_03553_));
 NOR2x2_ASAP7_75t_R _33141_ (.A(_03549_),
    .B(_03557_),
    .Y(_03558_));
 AO21x1_ASAP7_75t_R _33142_ (.A1(_22024_),
    .A2(_21929_),
    .B(_22061_),
    .Y(_03559_));
 AO21x1_ASAP7_75t_R _33143_ (.A1(net2365),
    .A2(_22057_),
    .B(_22061_),
    .Y(_03560_));
 NAND2x1_ASAP7_75t_R _33144_ (.A(_22053_),
    .B(_22062_),
    .Y(_03561_));
 AND3x1_ASAP7_75t_R _33145_ (.A(_03559_),
    .B(_03560_),
    .C(_03561_),
    .Y(_03562_));
 AO21x1_ASAP7_75t_R _33146_ (.A1(_21920_),
    .A2(_21929_),
    .B(_22064_),
    .Y(_03563_));
 AO21x1_ASAP7_75t_R _33147_ (.A1(net2266),
    .A2(net2365),
    .B(_22064_),
    .Y(_03564_));
 NAND2x1_ASAP7_75t_R _33148_ (.A(_22049_),
    .B(_01087_),
    .Y(_03565_));
 AND3x1_ASAP7_75t_R _33149_ (.A(_03563_),
    .B(_03564_),
    .C(_03565_),
    .Y(_03566_));
 NAND2x2_ASAP7_75t_R _33150_ (.A(_03562_),
    .B(_03566_),
    .Y(_03567_));
 INVx1_ASAP7_75t_R _33151_ (.A(_03151_),
    .Y(_03568_));
 OR3x2_ASAP7_75t_R _33152_ (.A(_02297_),
    .B(_03568_),
    .C(_22086_),
    .Y(_03569_));
 AO21x1_ASAP7_75t_R _33153_ (.A1(net1038),
    .A2(net2510),
    .B(_22070_),
    .Y(_03570_));
 AO21x1_ASAP7_75t_R _33154_ (.A1(net1048),
    .A2(net2801),
    .B(_22070_),
    .Y(_03571_));
 NOR2x1_ASAP7_75t_R _33155_ (.A(_22057_),
    .B(_22070_),
    .Y(_03572_));
 INVx1_ASAP7_75t_R _33156_ (.A(_03572_),
    .Y(_03573_));
 NAND3x2_ASAP7_75t_R _33157_ (.B(_03571_),
    .C(_03573_),
    .Y(_03574_),
    .A(_03570_));
 NOR3x2_ASAP7_75t_R _33158_ (.B(_03569_),
    .C(_03574_),
    .Y(_03575_),
    .A(_03567_));
 NAND2x2_ASAP7_75t_R _33159_ (.A(_03558_),
    .B(_03575_),
    .Y(_03576_));
 AO21x1_ASAP7_75t_R _33160_ (.A1(net2296),
    .A2(net1630),
    .B(_22004_),
    .Y(_03577_));
 NAND2x1_ASAP7_75t_R _33161_ (.A(net2802),
    .B(_22005_),
    .Y(_03578_));
 AND3x1_ASAP7_75t_R _33162_ (.A(_03577_),
    .B(_22007_),
    .C(_03578_),
    .Y(_03579_));
 NAND2x1_ASAP7_75t_R _33163_ (.A(_21953_),
    .B(_02758_),
    .Y(_03580_));
 NAND2x1_ASAP7_75t_R _33164_ (.A(_01085_),
    .B(_02758_),
    .Y(_03581_));
 AND3x1_ASAP7_75t_R _33165_ (.A(_21999_),
    .B(_03580_),
    .C(_03581_),
    .Y(_03582_));
 AO21x1_ASAP7_75t_R _33166_ (.A1(_21890_),
    .A2(net2420),
    .B(net3151),
    .Y(_03583_));
 AND3x4_ASAP7_75t_R _33167_ (.A(_03579_),
    .B(_03582_),
    .C(_03583_),
    .Y(_03584_));
 AO21x1_ASAP7_75t_R _33168_ (.A1(_21983_),
    .A2(_22057_),
    .B(_21893_),
    .Y(_03585_));
 NAND2x1_ASAP7_75t_R _33169_ (.A(_21885_),
    .B(_22003_),
    .Y(_03586_));
 AND3x1_ASAP7_75t_R _33170_ (.A(_03585_),
    .B(_21910_),
    .C(_03586_),
    .Y(_03587_));
 AO21x1_ASAP7_75t_R _33171_ (.A1(_22080_),
    .A2(net1834),
    .B(_21901_),
    .Y(_03588_));
 OAI21x1_ASAP7_75t_R _33172_ (.A1(net3280),
    .A2(net1751),
    .B(_03588_),
    .Y(_03589_));
 AO21x1_ASAP7_75t_R _33173_ (.A1(_21967_),
    .A2(net2420),
    .B(_21901_),
    .Y(_03590_));
 OAI21x1_ASAP7_75t_R _33174_ (.A1(net2365),
    .A2(net1751),
    .B(_03590_),
    .Y(_03591_));
 NOR2x1_ASAP7_75t_R _33175_ (.A(_03589_),
    .B(_03591_),
    .Y(_03592_));
 NAND2x1_ASAP7_75t_R _33176_ (.A(_03587_),
    .B(_03592_),
    .Y(_03593_));
 OAI21x1_ASAP7_75t_R _33177_ (.A1(_21962_),
    .A2(_02305_),
    .B(_21958_),
    .Y(_03594_));
 OA211x2_ASAP7_75t_R _33178_ (.A1(_21888_),
    .A2(_21918_),
    .B(_21957_),
    .C(_21872_),
    .Y(_03595_));
 NOR2x1_ASAP7_75t_R _33179_ (.A(_03594_),
    .B(_03595_),
    .Y(_03596_));
 AO21x1_ASAP7_75t_R _33180_ (.A1(net3155),
    .A2(_21969_),
    .B(_21976_),
    .Y(_03597_));
 INVx1_ASAP7_75t_R _33181_ (.A(_03597_),
    .Y(_03598_));
 OA211x2_ASAP7_75t_R _33182_ (.A1(net1139),
    .A2(_21876_),
    .B(_21980_),
    .C(net2589),
    .Y(_03599_));
 NOR2x1_ASAP7_75t_R _33183_ (.A(_03598_),
    .B(_03599_),
    .Y(_03600_));
 NAND2x1_ASAP7_75t_R _33184_ (.A(_03596_),
    .B(_03600_),
    .Y(_03601_));
 NOR2x2_ASAP7_75t_R _33185_ (.A(_03601_),
    .B(_03593_),
    .Y(_03602_));
 NOR2x2_ASAP7_75t_R _33186_ (.A(_22015_),
    .B(net1630),
    .Y(_03603_));
 OA21x2_ASAP7_75t_R _33187_ (.A1(_22075_),
    .A2(net2802),
    .B(_22016_),
    .Y(_03604_));
 NOR2x2_ASAP7_75t_R _33188_ (.A(_03603_),
    .B(_03604_),
    .Y(_03605_));
 AO21x1_ASAP7_75t_R _33189_ (.A1(net2420),
    .A2(_22008_),
    .B(net3075),
    .Y(_03606_));
 NAND3x2_ASAP7_75t_R _33190_ (.B(_03129_),
    .C(_03606_),
    .Y(_03607_),
    .A(_03605_));
 AOI21x1_ASAP7_75t_R _33191_ (.A1(_22019_),
    .A2(net2266),
    .B(net3156),
    .Y(_03608_));
 NOR2x1_ASAP7_75t_R _33192_ (.A(_02348_),
    .B(_03608_),
    .Y(_03609_));
 AO21x1_ASAP7_75t_R _33193_ (.A1(net1829),
    .A2(net3172),
    .B(net2556),
    .Y(_03610_));
 AO21x1_ASAP7_75t_R _33194_ (.A1(net1630),
    .A2(net1833),
    .B(net3156),
    .Y(_03611_));
 NAND2x1_ASAP7_75t_R _33195_ (.A(_22075_),
    .B(_22034_),
    .Y(_03612_));
 AND3x1_ASAP7_75t_R _33196_ (.A(_03610_),
    .B(_03611_),
    .C(_03612_),
    .Y(_03613_));
 NAND2x1_ASAP7_75t_R _33197_ (.A(_03609_),
    .B(_03613_),
    .Y(_03614_));
 NOR2x2_ASAP7_75t_R _33198_ (.A(_03614_),
    .B(_03607_),
    .Y(_03615_));
 NAND3x2_ASAP7_75t_R _33199_ (.B(_03602_),
    .C(_03615_),
    .Y(_03616_),
    .A(_03584_));
 NOR2x2_ASAP7_75t_R _33200_ (.A(_03576_),
    .B(_03616_),
    .Y(_03617_));
 XOR2x2_ASAP7_75t_R _33201_ (.A(_03539_),
    .B(_03617_),
    .Y(_03618_));
 OA211x2_ASAP7_75t_R _33202_ (.A1(_01770_),
    .A2(net1455),
    .B(_01904_),
    .C(_01830_),
    .Y(_03619_));
 NOR2x1_ASAP7_75t_R _33203_ (.A(_02521_),
    .B(_03619_),
    .Y(_03620_));
 AO21x1_ASAP7_75t_R _33204_ (.A1(_01832_),
    .A2(_01877_),
    .B(net2140),
    .Y(_03621_));
 INVx2_ASAP7_75t_R _33205_ (.A(_01916_),
    .Y(_03622_));
 NAND2x1_ASAP7_75t_R _33206_ (.A(_01787_),
    .B(_03622_),
    .Y(_03623_));
 AND2x2_ASAP7_75t_R _33207_ (.A(_03621_),
    .B(_03623_),
    .Y(_03624_));
 NAND3x1_ASAP7_75t_R _33208_ (.A(_03620_),
    .B(_02204_),
    .C(_03624_),
    .Y(_03625_));
 AO21x1_ASAP7_75t_R _33209_ (.A1(net1413),
    .A2(net1527),
    .B(net2195),
    .Y(_03626_));
 NAND2x1_ASAP7_75t_R _33210_ (.A(net1454),
    .B(net1464),
    .Y(_03627_));
 AO21x1_ASAP7_75t_R _33211_ (.A1(_03627_),
    .A2(_01908_),
    .B(net2195),
    .Y(_03628_));
 NAND2x1_ASAP7_75t_R _33212_ (.A(_01806_),
    .B(_01940_),
    .Y(_03629_));
 AND3x1_ASAP7_75t_R _33213_ (.A(_03626_),
    .B(_03628_),
    .C(_03629_),
    .Y(_03630_));
 NOR2x1_ASAP7_75t_R _33214_ (.A(_02149_),
    .B(net2549),
    .Y(_03631_));
 INVx1_ASAP7_75t_R _33215_ (.A(_03631_),
    .Y(_03632_));
 AND3x1_ASAP7_75t_R _33216_ (.A(_01927_),
    .B(_02967_),
    .C(_03632_),
    .Y(_03633_));
 AOI21x1_ASAP7_75t_R _33217_ (.A1(net950),
    .A2(_02535_),
    .B(_02963_),
    .Y(_03634_));
 NAND3x1_ASAP7_75t_R _33218_ (.A(_03630_),
    .B(_03633_),
    .C(_03634_),
    .Y(_03635_));
 NOR2x1_ASAP7_75t_R _33219_ (.A(_03625_),
    .B(_03635_),
    .Y(_03636_));
 AO21x1_ASAP7_75t_R _33220_ (.A1(net2563),
    .A2(net1138),
    .B(_01977_),
    .Y(_03637_));
 AO21x1_ASAP7_75t_R _33221_ (.A1(_02129_),
    .A2(_01934_),
    .B(_01977_),
    .Y(_03638_));
 NOR2x1_ASAP7_75t_R _33222_ (.A(_01836_),
    .B(_01977_),
    .Y(_03639_));
 INVx1_ASAP7_75t_R _33223_ (.A(_03639_),
    .Y(_03640_));
 AND3x1_ASAP7_75t_R _33224_ (.A(_03637_),
    .B(_03638_),
    .C(_03640_),
    .Y(_03641_));
 AO21x1_ASAP7_75t_R _33225_ (.A1(net1413),
    .A2(_01824_),
    .B(_01967_),
    .Y(_03642_));
 AO21x1_ASAP7_75t_R _33226_ (.A1(net2307),
    .A2(net3275),
    .B(_01967_),
    .Y(_03643_));
 NAND2x1_ASAP7_75t_R _33227_ (.A(_01970_),
    .B(_02177_),
    .Y(_03644_));
 INVx1_ASAP7_75t_R _33228_ (.A(_01935_),
    .Y(_03645_));
 NAND2x1_ASAP7_75t_R _33229_ (.A(_01970_),
    .B(_03645_),
    .Y(_03646_));
 AND4x1_ASAP7_75t_R _33230_ (.A(_03642_),
    .B(_03643_),
    .C(_03644_),
    .D(_03646_),
    .Y(_03647_));
 NAND2x1_ASAP7_75t_R _33231_ (.A(_03647_),
    .B(_03641_),
    .Y(_03648_));
 NOR2x1_ASAP7_75t_R _33232_ (.A(_01831_),
    .B(net2264),
    .Y(_03649_));
 INVx1_ASAP7_75t_R _33233_ (.A(_03649_),
    .Y(_03650_));
 AO21x1_ASAP7_75t_R _33234_ (.A1(net3131),
    .A2(net1157),
    .B(net2264),
    .Y(_03651_));
 NAND2x1_ASAP7_75t_R _33235_ (.A(_03650_),
    .B(_03651_),
    .Y(_03652_));
 NOR2x1_ASAP7_75t_R _33236_ (.A(_01908_),
    .B(net2263),
    .Y(_03653_));
 NOR2x1_ASAP7_75t_R _33237_ (.A(net2307),
    .B(net2352),
    .Y(_03654_));
 INVx1_ASAP7_75t_R _33238_ (.A(_01955_),
    .Y(_03655_));
 OA21x2_ASAP7_75t_R _33239_ (.A1(_02918_),
    .A2(_02117_),
    .B(_03655_),
    .Y(_03656_));
 OR4x1_ASAP7_75t_R _33240_ (.A(_03652_),
    .B(_03653_),
    .C(_03654_),
    .D(_03656_),
    .Y(_03657_));
 NOR2x1_ASAP7_75t_R _33241_ (.A(_03657_),
    .B(_03648_),
    .Y(_03658_));
 NAND2x2_ASAP7_75t_R _33242_ (.A(_03658_),
    .B(_03636_),
    .Y(_03659_));
 AO21x1_ASAP7_75t_R _33243_ (.A1(net3254),
    .A2(net1157),
    .B(net3128),
    .Y(_03660_));
 AO21x1_ASAP7_75t_R _33244_ (.A1(net1138),
    .A2(_02559_),
    .B(_01894_),
    .Y(_03661_));
 AND3x1_ASAP7_75t_R _33245_ (.A(_03660_),
    .B(_03661_),
    .C(_02914_),
    .Y(_03662_));
 NAND2x2_ASAP7_75t_R _33246_ (.A(_02117_),
    .B(_01876_),
    .Y(_03663_));
 AO21x1_ASAP7_75t_R _33247_ (.A1(_01785_),
    .A2(_01832_),
    .B(_01878_),
    .Y(_03664_));
 NAND2x1_ASAP7_75t_R _33248_ (.A(_03663_),
    .B(_03664_),
    .Y(_03665_));
 INVx1_ASAP7_75t_R _33249_ (.A(_03665_),
    .Y(_03666_));
 AO21x1_ASAP7_75t_R _33250_ (.A1(_01799_),
    .A2(net1138),
    .B(_01878_),
    .Y(_03667_));
 OA21x2_ASAP7_75t_R _33251_ (.A1(_01857_),
    .A2(_01878_),
    .B(_03667_),
    .Y(_03668_));
 NAND3x1_ASAP7_75t_R _33252_ (.A(_03662_),
    .B(_03666_),
    .C(_03668_),
    .Y(_03669_));
 AO21x1_ASAP7_75t_R _33253_ (.A1(net2175),
    .A2(_01946_),
    .B(_01851_),
    .Y(_03670_));
 AND3x1_ASAP7_75t_R _33254_ (.A(_03670_),
    .B(_02562_),
    .C(_02109_),
    .Y(_03671_));
 NAND2x1_ASAP7_75t_R _33255_ (.A(net2619),
    .B(net2218),
    .Y(_03672_));
 OA21x2_ASAP7_75t_R _33256_ (.A1(_03672_),
    .A2(_01911_),
    .B(_01864_),
    .Y(_03673_));
 AO21x1_ASAP7_75t_R _33257_ (.A1(net2560),
    .A2(net1245),
    .B(net2494),
    .Y(_03674_));
 AO21x1_ASAP7_75t_R _33258_ (.A1(_02110_),
    .A2(_02100_),
    .B(net2494),
    .Y(_03675_));
 NAND2x1_ASAP7_75t_R _33259_ (.A(_03674_),
    .B(_03675_),
    .Y(_03676_));
 NOR2x1_ASAP7_75t_R _33260_ (.A(_03673_),
    .B(_03676_),
    .Y(_03677_));
 AOI211x1_ASAP7_75t_R _33261_ (.A1(net1116),
    .A2(_01776_),
    .B(_01857_),
    .C(_01851_),
    .Y(_03678_));
 NAND2x1_ASAP7_75t_R _33262_ (.A(_01882_),
    .B(_01847_),
    .Y(_03679_));
 NAND2x1_ASAP7_75t_R _33263_ (.A(_01847_),
    .B(_02177_),
    .Y(_03680_));
 NAND2x1_ASAP7_75t_R _33264_ (.A(_03679_),
    .B(_03680_),
    .Y(_03681_));
 NOR2x1_ASAP7_75t_R _33265_ (.A(_03678_),
    .B(_03681_),
    .Y(_03682_));
 NAND3x1_ASAP7_75t_R _33266_ (.A(_03671_),
    .B(_03677_),
    .C(_03682_),
    .Y(_03683_));
 NOR2x1_ASAP7_75t_R _33267_ (.A(_03669_),
    .B(_03683_),
    .Y(_03684_));
 AO21x1_ASAP7_75t_R _33268_ (.A1(net2175),
    .A2(_01832_),
    .B(_01781_),
    .Y(_03685_));
 AO21x1_ASAP7_75t_R _33269_ (.A1(net1527),
    .A2(net1157),
    .B(_01781_),
    .Y(_03686_));
 NAND2x1_ASAP7_75t_R _33270_ (.A(net3274),
    .B(_02131_),
    .Y(_03687_));
 AND3x1_ASAP7_75t_R _33271_ (.A(_03685_),
    .B(_03686_),
    .C(_03687_),
    .Y(_03688_));
 AO21x1_ASAP7_75t_R _33272_ (.A1(net2563),
    .A2(net1138),
    .B(_01781_),
    .Y(_03689_));
 AO21x1_ASAP7_75t_R _33273_ (.A1(net2619),
    .A2(_01837_),
    .B(_01781_),
    .Y(_03690_));
 NOR2x1_ASAP7_75t_R _33274_ (.A(_01781_),
    .B(_01908_),
    .Y(_03691_));
 INVx1_ASAP7_75t_R _33275_ (.A(_03691_),
    .Y(_03692_));
 AND3x1_ASAP7_75t_R _33276_ (.A(_03689_),
    .B(_03690_),
    .C(_03692_),
    .Y(_03693_));
 OA21x2_ASAP7_75t_R _33277_ (.A1(_01855_),
    .A2(net2654),
    .B(_01762_),
    .Y(_03694_));
 OA21x2_ASAP7_75t_R _33278_ (.A1(_01976_),
    .A2(_02099_),
    .B(_01762_),
    .Y(_03695_));
 NOR2x1_ASAP7_75t_R _33279_ (.A(_03694_),
    .B(_03695_),
    .Y(_03696_));
 NAND3x1_ASAP7_75t_R _33280_ (.A(_03688_),
    .B(_03693_),
    .C(_03696_),
    .Y(_03697_));
 AO21x1_ASAP7_75t_R _33281_ (.A1(net3132),
    .A2(net1157),
    .B(_01828_),
    .Y(_03698_));
 NAND2x1_ASAP7_75t_R _33282_ (.A(_02936_),
    .B(_03698_),
    .Y(_03699_));
 NAND2x1_ASAP7_75t_R _33283_ (.A(_02142_),
    .B(_01835_),
    .Y(_03700_));
 OR2x2_ASAP7_75t_R _33284_ (.A(_03699_),
    .B(_03700_),
    .Y(_03701_));
 OA21x2_ASAP7_75t_R _33285_ (.A1(_02124_),
    .A2(_02114_),
    .B(_01810_),
    .Y(_03702_));
 OA21x2_ASAP7_75t_R _33286_ (.A1(_02190_),
    .A2(_02117_),
    .B(_01810_),
    .Y(_03703_));
 NAND2x1_ASAP7_75t_R _33287_ (.A(_01911_),
    .B(_01810_),
    .Y(_03704_));
 INVx1_ASAP7_75t_R _33288_ (.A(_03704_),
    .Y(_03705_));
 OR3x1_ASAP7_75t_R _33289_ (.A(_03702_),
    .B(_03703_),
    .C(_03705_),
    .Y(_03706_));
 OR2x2_ASAP7_75t_R _33290_ (.A(_03701_),
    .B(_03706_),
    .Y(_03707_));
 NOR2x1_ASAP7_75t_R _33291_ (.A(_03707_),
    .B(_03697_),
    .Y(_03708_));
 NAND2x1_ASAP7_75t_R _33292_ (.A(_03684_),
    .B(_03708_),
    .Y(_03709_));
 NOR2x2_ASAP7_75t_R _33293_ (.A(_03659_),
    .B(_03709_),
    .Y(_03710_));
 XOR2x2_ASAP7_75t_R _33294_ (.A(_03710_),
    .B(net2710),
    .Y(_03711_));
 XOR2x2_ASAP7_75t_R _33295_ (.A(_03618_),
    .B(_03711_),
    .Y(_03712_));
 NAND2x1_ASAP7_75t_R _33296_ (.A(_03467_),
    .B(_03712_),
    .Y(_03713_));
 XOR2x2_ASAP7_75t_R _33297_ (.A(_03090_),
    .B(_03376_),
    .Y(_03714_));
 XOR2x1_ASAP7_75t_R _33298_ (.A(_03714_),
    .Y(_03715_),
    .B(net3150));
 XNOR2x2_ASAP7_75t_R _33299_ (.A(_03711_),
    .B(_03618_),
    .Y(_03716_));
 NAND2x1_ASAP7_75t_R _33300_ (.A(_03715_),
    .B(_03716_),
    .Y(_03717_));
 AOI21x1_ASAP7_75t_R _33301_ (.A1(_03713_),
    .A2(_03717_),
    .B(_18753_),
    .Y(_03718_));
 INVx1_ASAP7_75t_R _33302_ (.A(_00480_),
    .Y(_03719_));
 OAI21x1_ASAP7_75t_R _33303_ (.A1(_03398_),
    .A2(_03718_),
    .B(_03719_),
    .Y(_03720_));
 NOR2x1_ASAP7_75t_R _33304_ (.A(net395),
    .B(_00879_),
    .Y(_03721_));
 NAND2x1_ASAP7_75t_R _33305_ (.A(_03715_),
    .B(_03712_),
    .Y(_03722_));
 NAND2x1_ASAP7_75t_R _33306_ (.A(_03716_),
    .B(_03467_),
    .Y(_03723_));
 AOI21x1_ASAP7_75t_R _33307_ (.A1(_03722_),
    .A2(_03723_),
    .B(_18753_),
    .Y(_03724_));
 OAI21x1_ASAP7_75t_R _33308_ (.A1(_03721_),
    .A2(_03724_),
    .B(_00480_),
    .Y(_03725_));
 NAND2x1_ASAP7_75t_R _33309_ (.A(_03725_),
    .B(_03720_),
    .Y(_00117_));
 NAND2x1_ASAP7_75t_R _33310_ (.A(_00878_),
    .B(net390),
    .Y(_03726_));
 INVx1_ASAP7_75t_R _33311_ (.A(_21911_),
    .Y(_03727_));
 AO21x1_ASAP7_75t_R _33312_ (.A1(net3155),
    .A2(_21983_),
    .B(_21893_),
    .Y(_03728_));
 INVx1_ASAP7_75t_R _33313_ (.A(_21894_),
    .Y(_03729_));
 INVx1_ASAP7_75t_R _33314_ (.A(_21897_),
    .Y(_03730_));
 NAND3x2_ASAP7_75t_R _33315_ (.B(_03729_),
    .C(_03730_),
    .Y(_03731_),
    .A(_03728_));
 NOR2x2_ASAP7_75t_R _33316_ (.A(_03727_),
    .B(_03731_),
    .Y(_03732_));
 NAND3x2_ASAP7_75t_R _33317_ (.B(net1751),
    .C(_21868_),
    .Y(_03733_),
    .A(_03732_));
 NOR3x2_ASAP7_75t_R _33318_ (.B(_21865_),
    .C(_21867_),
    .Y(_03734_),
    .A(_03733_));
 OR3x1_ASAP7_75t_R _33319_ (.A(_22061_),
    .B(net2005),
    .C(net1139),
    .Y(_03735_));
 NOR2x1_ASAP7_75t_R _33320_ (.A(net1629),
    .B(_22061_),
    .Y(_03736_));
 AOI211x1_ASAP7_75t_R _33321_ (.A1(_21887_),
    .A2(_21876_),
    .B(_22061_),
    .C(net1039),
    .Y(_03737_));
 NOR2x1_ASAP7_75t_R _33322_ (.A(_03736_),
    .B(_03737_),
    .Y(_03738_));
 NAND2x1_ASAP7_75t_R _33323_ (.A(_03735_),
    .B(_03738_),
    .Y(_03739_));
 OA21x2_ASAP7_75t_R _33324_ (.A1(_02316_),
    .A2(_21881_),
    .B(_22049_),
    .Y(_03740_));
 AOI211x1_ASAP7_75t_R _33325_ (.A1(_21887_),
    .A2(_21876_),
    .B(_22064_),
    .C(_21895_),
    .Y(_03741_));
 NOR2x1_ASAP7_75t_R _33326_ (.A(_03740_),
    .B(_03741_),
    .Y(_03742_));
 OA21x2_ASAP7_75t_R _33327_ (.A1(net1792),
    .A2(_22064_),
    .B(_22051_),
    .Y(_03743_));
 NAND2x1_ASAP7_75t_R _33328_ (.A(_03743_),
    .B(_03742_),
    .Y(_03744_));
 NOR2x1_ASAP7_75t_R _33329_ (.A(_03739_),
    .B(_03744_),
    .Y(_03745_));
 NAND2x1_ASAP7_75t_R _33330_ (.A(net3083),
    .B(_02292_),
    .Y(_03746_));
 NAND3x1_ASAP7_75t_R _33331_ (.A(_02290_),
    .B(_03154_),
    .C(_03746_),
    .Y(_03747_));
 AOI211x1_ASAP7_75t_R _33332_ (.A1(net1139),
    .A2(net1049),
    .B(net1711),
    .C(_22077_),
    .Y(_03748_));
 INVx1_ASAP7_75t_R _33333_ (.A(_03748_),
    .Y(_03749_));
 NAND2x1_ASAP7_75t_R _33334_ (.A(_22084_),
    .B(net2802),
    .Y(_03750_));
 AO21x1_ASAP7_75t_R _33335_ (.A1(net2752),
    .A2(_02273_),
    .B(_22077_),
    .Y(_03751_));
 NAND3x1_ASAP7_75t_R _33336_ (.A(_03749_),
    .B(_03750_),
    .C(_03751_),
    .Y(_03752_));
 NOR2x1_ASAP7_75t_R _33337_ (.A(_03747_),
    .B(_03752_),
    .Y(_03753_));
 NAND2x1_ASAP7_75t_R _33338_ (.A(_03745_),
    .B(_03753_),
    .Y(_03754_));
 AO31x2_ASAP7_75t_R _33339_ (.A1(_21907_),
    .A2(net3173),
    .A3(net1048),
    .B(_01072_),
    .Y(_03755_));
 AO31x2_ASAP7_75t_R _33340_ (.A1(net2261),
    .A2(net2265),
    .A3(net3225),
    .B(_01072_),
    .Y(_03756_));
 NAND2x1_ASAP7_75t_R _33341_ (.A(_03755_),
    .B(_03756_),
    .Y(_03757_));
 AOI211x1_ASAP7_75t_R _33342_ (.A1(_21887_),
    .A2(net1049),
    .B(net3152),
    .C(net1709),
    .Y(_03758_));
 INVx1_ASAP7_75t_R _33343_ (.A(_03758_),
    .Y(_03759_));
 AO21x1_ASAP7_75t_R _33344_ (.A1(_21995_),
    .A2(_21944_),
    .B(net3143),
    .Y(_03760_));
 NAND3x1_ASAP7_75t_R _33345_ (.A(_03759_),
    .B(_03760_),
    .C(_03545_),
    .Y(_03761_));
 NOR2x1_ASAP7_75t_R _33346_ (.A(_03757_),
    .B(_03761_),
    .Y(_03762_));
 AO21x1_ASAP7_75t_R _33347_ (.A1(net2510),
    .A2(net2420),
    .B(net3082),
    .Y(_03763_));
 AO21x1_ASAP7_75t_R _33348_ (.A1(net1829),
    .A2(_21995_),
    .B(net3082),
    .Y(_03764_));
 NAND2x1_ASAP7_75t_R _33349_ (.A(_03763_),
    .B(_03764_),
    .Y(_03765_));
 AO31x2_ASAP7_75t_R _33350_ (.A1(_22024_),
    .A2(net1792),
    .A3(_22080_),
    .B(_22091_),
    .Y(_03766_));
 OA21x2_ASAP7_75t_R _33351_ (.A1(_22014_),
    .A2(_03107_),
    .B(_22092_),
    .Y(_03767_));
 AOI21x1_ASAP7_75t_R _33352_ (.A1(_01082_),
    .A2(_22092_),
    .B(_03767_),
    .Y(_03768_));
 NAND2x1_ASAP7_75t_R _33353_ (.A(_03766_),
    .B(_03768_),
    .Y(_03769_));
 NOR2x1_ASAP7_75t_R _33354_ (.A(_03765_),
    .B(_03769_),
    .Y(_03770_));
 NAND2x2_ASAP7_75t_R _33355_ (.A(_03762_),
    .B(_03770_),
    .Y(_03771_));
 NOR2x2_ASAP7_75t_R _33356_ (.A(_03771_),
    .B(_03754_),
    .Y(_03772_));
 AO21x1_ASAP7_75t_R _33357_ (.A1(_21890_),
    .A2(_03133_),
    .B(net3151),
    .Y(_03773_));
 AO21x1_ASAP7_75t_R _33358_ (.A1(_02305_),
    .A2(net3280),
    .B(net3151),
    .Y(_03774_));
 NAND2x2_ASAP7_75t_R _33359_ (.A(_03773_),
    .B(_03774_),
    .Y(_03775_));
 AO21x1_ASAP7_75t_R _33360_ (.A1(net3172),
    .A2(net1792),
    .B(net3148),
    .Y(_03776_));
 OAI21x1_ASAP7_75t_R _33361_ (.A1(net3148),
    .A2(_21929_),
    .B(_03776_),
    .Y(_03777_));
 NOR3x2_ASAP7_75t_R _33362_ (.B(_03777_),
    .C(_22011_),
    .Y(_03778_),
    .A(_03775_));
 NAND2x1_ASAP7_75t_R _33363_ (.A(_21909_),
    .B(_22034_),
    .Y(_03779_));
 NAND2x1_ASAP7_75t_R _33364_ (.A(_03779_),
    .B(_03611_),
    .Y(_03780_));
 AO21x1_ASAP7_75t_R _33365_ (.A1(_22018_),
    .A2(_22019_),
    .B(net3156),
    .Y(_03781_));
 NAND2x1_ASAP7_75t_R _33366_ (.A(_22031_),
    .B(_03781_),
    .Y(_03782_));
 NOR2x1_ASAP7_75t_R _33367_ (.A(_03780_),
    .B(_03782_),
    .Y(_03783_));
 AO21x1_ASAP7_75t_R _33368_ (.A1(net2258),
    .A2(_02273_),
    .B(net3075),
    .Y(_03784_));
 NAND2x1_ASAP7_75t_R _33369_ (.A(_03784_),
    .B(_03129_),
    .Y(_03785_));
 AO21x1_ASAP7_75t_R _33370_ (.A1(_02340_),
    .A2(net993),
    .B(_03603_),
    .Y(_03786_));
 NOR2x1_ASAP7_75t_R _33371_ (.A(_03785_),
    .B(_03786_),
    .Y(_03787_));
 NAND2x1_ASAP7_75t_R _33372_ (.A(_03783_),
    .B(_03787_),
    .Y(_03788_));
 INVx1_ASAP7_75t_R _33373_ (.A(_03788_),
    .Y(_03789_));
 NAND2x1_ASAP7_75t_R _33374_ (.A(_03778_),
    .B(_03789_),
    .Y(_03790_));
 AOI221x1_ASAP7_75t_R _33375_ (.A1(net1139),
    .A2(_21876_),
    .B1(net1710),
    .B2(_21895_),
    .C(net2497),
    .Y(_03791_));
 INVx1_ASAP7_75t_R _33376_ (.A(_21910_),
    .Y(_03792_));
 NOR3x2_ASAP7_75t_R _33377_ (.B(_03792_),
    .C(_02315_),
    .Y(_03793_),
    .A(_03791_));
 AO21x1_ASAP7_75t_R _33378_ (.A1(net2510),
    .A2(_21895_),
    .B(_21976_),
    .Y(_03794_));
 OAI21x1_ASAP7_75t_R _33379_ (.A1(_21929_),
    .A2(_21976_),
    .B(_03794_),
    .Y(_03795_));
 AO21x1_ASAP7_75t_R _33380_ (.A1(net2752),
    .A2(_21940_),
    .B(_21962_),
    .Y(_03796_));
 NAND2x1_ASAP7_75t_R _33381_ (.A(net1650),
    .B(_21957_),
    .Y(_03797_));
 OAI21x1_ASAP7_75t_R _33382_ (.A1(_02304_),
    .A2(_02722_),
    .B(_21957_),
    .Y(_03798_));
 NAND3x1_ASAP7_75t_R _33383_ (.A(_03796_),
    .B(_03797_),
    .C(_03798_),
    .Y(_03799_));
 NOR2x1_ASAP7_75t_R _33384_ (.A(_03795_),
    .B(_03799_),
    .Y(_03800_));
 AOI21x1_ASAP7_75t_R _33385_ (.A1(net3077),
    .A2(_03097_),
    .B(net1751),
    .Y(_03801_));
 AO21x1_ASAP7_75t_R _33386_ (.A1(net2258),
    .A2(_21940_),
    .B(net1751),
    .Y(_03802_));
 AO21x1_ASAP7_75t_R _33387_ (.A1(_21983_),
    .A2(_21890_),
    .B(net1751),
    .Y(_03803_));
 NAND2x1_ASAP7_75t_R _33388_ (.A(_03802_),
    .B(_03803_),
    .Y(_03804_));
 NOR2x2_ASAP7_75t_R _33389_ (.A(_03801_),
    .B(_03804_),
    .Y(_03805_));
 NAND3x1_ASAP7_75t_R _33390_ (.A(_03793_),
    .B(_03800_),
    .C(_03805_),
    .Y(_03806_));
 NOR2x1_ASAP7_75t_R _33391_ (.A(_03790_),
    .B(_03806_),
    .Y(_03807_));
 NAND2x2_ASAP7_75t_R _33392_ (.A(_03807_),
    .B(_03772_),
    .Y(_03808_));
 NOR2x2_ASAP7_75t_R _33393_ (.A(_03734_),
    .B(_03808_),
    .Y(_03809_));
 NOR2x1_ASAP7_75t_R _33394_ (.A(_01307_),
    .B(_01370_),
    .Y(_03810_));
 NAND2x2_ASAP7_75t_R _33395_ (.A(_00585_),
    .B(_03810_),
    .Y(_03811_));
 AO21x1_ASAP7_75t_R _33396_ (.A1(_01228_),
    .A2(_01113_),
    .B(_01133_),
    .Y(_03812_));
 AND2x2_ASAP7_75t_R _33397_ (.A(_03812_),
    .B(_01465_),
    .Y(_03813_));
 AO21x1_ASAP7_75t_R _33398_ (.A1(net1752),
    .A2(_01292_),
    .B(_01120_),
    .Y(_03814_));
 AO21x1_ASAP7_75t_R _33399_ (.A1(_01172_),
    .A2(_01128_),
    .B(_01120_),
    .Y(_03815_));
 NAND2x1_ASAP7_75t_R _33400_ (.A(_01103_),
    .B(_01406_),
    .Y(_03816_));
 AND3x1_ASAP7_75t_R _33401_ (.A(_03814_),
    .B(_03815_),
    .C(_03816_),
    .Y(_03817_));
 NAND2x1_ASAP7_75t_R _33402_ (.A(_03813_),
    .B(_03817_),
    .Y(_03818_));
 OA21x2_ASAP7_75t_R _33403_ (.A1(_01209_),
    .A2(_01305_),
    .B(_01163_),
    .Y(_03819_));
 NAND2x1_ASAP7_75t_R _33404_ (.A(_01186_),
    .B(net3142),
    .Y(_03820_));
 NOR2x1_ASAP7_75t_R _33405_ (.A(_03820_),
    .B(_01156_),
    .Y(_03821_));
 NOR2x1_ASAP7_75t_R _33406_ (.A(net2125),
    .B(_01156_),
    .Y(_03822_));
 NOR3x1_ASAP7_75t_R _33407_ (.A(_03819_),
    .B(_03821_),
    .C(_03822_),
    .Y(_03823_));
 AOI211x1_ASAP7_75t_R _33408_ (.A1(net1341),
    .A2(_01096_),
    .B(_01170_),
    .C(_01221_),
    .Y(_03824_));
 OA21x2_ASAP7_75t_R _33409_ (.A1(_02600_),
    .A2(_02592_),
    .B(_01171_),
    .Y(_03825_));
 NOR2x1_ASAP7_75t_R _33410_ (.A(_03824_),
    .B(_03825_),
    .Y(_03826_));
 AOI21x1_ASAP7_75t_R _33411_ (.A1(net2443),
    .A2(_01171_),
    .B(_01177_),
    .Y(_03827_));
 NAND3x1_ASAP7_75t_R _33412_ (.A(_03823_),
    .B(_03826_),
    .C(_03827_),
    .Y(_03828_));
 NOR2x1_ASAP7_75t_R _33413_ (.A(_03818_),
    .B(_03828_),
    .Y(_03829_));
 AO21x1_ASAP7_75t_R _33414_ (.A1(net2121),
    .A2(net2361),
    .B(_01202_),
    .Y(_03830_));
 AO21x1_ASAP7_75t_R _33415_ (.A1(_03297_),
    .A2(net1294),
    .B(_01202_),
    .Y(_03831_));
 AND3x1_ASAP7_75t_R _33416_ (.A(_03830_),
    .B(_03831_),
    .C(_03058_),
    .Y(_03832_));
 AO21x1_ASAP7_75t_R _33417_ (.A1(net2316),
    .A2(_01252_),
    .B(_01191_),
    .Y(_03833_));
 AO21x1_ASAP7_75t_R _33418_ (.A1(net2121),
    .A2(net1428),
    .B(_01191_),
    .Y(_03834_));
 AND3x1_ASAP7_75t_R _33419_ (.A(_03833_),
    .B(_03834_),
    .C(_03313_),
    .Y(_03835_));
 NAND2x1_ASAP7_75t_R _33420_ (.A(_03832_),
    .B(_03835_),
    .Y(_03836_));
 NOR2x1_ASAP7_75t_R _33421_ (.A(_01215_),
    .B(_01138_),
    .Y(_03837_));
 NOR3x1_ASAP7_75t_R _33422_ (.A(_01451_),
    .B(_03837_),
    .C(_03054_),
    .Y(_03838_));
 OA21x2_ASAP7_75t_R _33423_ (.A1(_01160_),
    .A2(_01305_),
    .B(_01234_),
    .Y(_03839_));
 AOI21x1_ASAP7_75t_R _33424_ (.A1(_01234_),
    .A2(_01313_),
    .B(_03839_),
    .Y(_03840_));
 AO21x1_ASAP7_75t_R _33425_ (.A1(net1119),
    .A2(_01453_),
    .B(_01215_),
    .Y(_03841_));
 NAND3x1_ASAP7_75t_R _33426_ (.A(_03838_),
    .B(_03840_),
    .C(_03841_),
    .Y(_03842_));
 NOR2x1_ASAP7_75t_R _33427_ (.A(_03836_),
    .B(_03842_),
    .Y(_03843_));
 NAND2x1_ASAP7_75t_R _33428_ (.A(_03829_),
    .B(_03843_),
    .Y(_03844_));
 NOR2x1_ASAP7_75t_R _33429_ (.A(net1696),
    .B(_01243_),
    .Y(_03845_));
 AOI211x1_ASAP7_75t_R _33430_ (.A1(_01209_),
    .A2(_01251_),
    .B(_03845_),
    .C(_01244_),
    .Y(_03846_));
 INVx1_ASAP7_75t_R _33431_ (.A(_02051_),
    .Y(_03847_));
 AO21x1_ASAP7_75t_R _33432_ (.A1(_03847_),
    .A2(_01321_),
    .B(net3315),
    .Y(_03848_));
 AO21x1_ASAP7_75t_R _33433_ (.A1(_01172_),
    .A2(net1572),
    .B(net3315),
    .Y(_03849_));
 AND3x1_ASAP7_75t_R _33434_ (.A(_03848_),
    .B(_03849_),
    .C(_03341_),
    .Y(_03850_));
 NAND2x1_ASAP7_75t_R _33435_ (.A(_03846_),
    .B(_03850_),
    .Y(_03851_));
 AO21x1_ASAP7_75t_R _33436_ (.A1(_03847_),
    .A2(_01248_),
    .B(_01287_),
    .Y(_03852_));
 INVx1_ASAP7_75t_R _33437_ (.A(_03852_),
    .Y(_03853_));
 AOI221x1_ASAP7_75t_R _33438_ (.A1(net1341),
    .A2(_01096_),
    .B1(_01204_),
    .B2(_01221_),
    .C(_01287_),
    .Y(_03854_));
 NOR2x1_ASAP7_75t_R _33439_ (.A(_03853_),
    .B(_03854_),
    .Y(_03855_));
 AND2x2_ASAP7_75t_R _33440_ (.A(_01423_),
    .B(_03506_),
    .Y(_03856_));
 AO21x1_ASAP7_75t_R _33441_ (.A1(_01252_),
    .A2(_01292_),
    .B(_01276_),
    .Y(_03857_));
 AO21x1_ASAP7_75t_R _33442_ (.A1(_01125_),
    .A2(_01194_),
    .B(_01276_),
    .Y(_03858_));
 AND2x2_ASAP7_75t_R _33443_ (.A(_03857_),
    .B(_03858_),
    .Y(_03859_));
 NAND3x1_ASAP7_75t_R _33444_ (.A(_03855_),
    .B(_03856_),
    .C(_03859_),
    .Y(_03860_));
 NOR2x1_ASAP7_75t_R _33445_ (.A(_03851_),
    .B(_03860_),
    .Y(_03861_));
 INVx1_ASAP7_75t_R _33446_ (.A(_01316_),
    .Y(_03862_));
 AO21x1_ASAP7_75t_R _33447_ (.A1(net2361),
    .A2(net1142),
    .B(_01308_),
    .Y(_03863_));
 NAND2x1_ASAP7_75t_R _33448_ (.A(_02677_),
    .B(_03863_),
    .Y(_03864_));
 NOR2x1_ASAP7_75t_R _33449_ (.A(_03862_),
    .B(_03864_),
    .Y(_03865_));
 AO21x1_ASAP7_75t_R _33450_ (.A1(_03847_),
    .A2(_01226_),
    .B(_01322_),
    .Y(_03866_));
 NAND2x1_ASAP7_75t_R _33451_ (.A(_01253_),
    .B(_01329_),
    .Y(_03867_));
 AND3x1_ASAP7_75t_R _33452_ (.A(_03019_),
    .B(_03866_),
    .C(_03867_),
    .Y(_03868_));
 NAND2x1_ASAP7_75t_R _33453_ (.A(_03865_),
    .B(_03868_),
    .Y(_03869_));
 AO21x1_ASAP7_75t_R _33454_ (.A1(net2120),
    .A2(_01248_),
    .B(_01345_),
    .Y(_03870_));
 AO21x1_ASAP7_75t_R _33455_ (.A1(net1293),
    .A2(net3341),
    .B(_01345_),
    .Y(_03871_));
 AND3x4_ASAP7_75t_R _33456_ (.A(_03870_),
    .B(_03013_),
    .C(_03871_),
    .Y(_03872_));
 AO21x1_ASAP7_75t_R _33457_ (.A1(_01348_),
    .A2(net1698),
    .B(_01334_),
    .Y(_03873_));
 AND2x2_ASAP7_75t_R _33458_ (.A(_01341_),
    .B(_03873_),
    .Y(_03874_));
 AO31x2_ASAP7_75t_R _33459_ (.A1(net1142),
    .A2(net2123),
    .A3(_01138_),
    .B(_01334_),
    .Y(_03875_));
 AND2x4_ASAP7_75t_R _33460_ (.A(_03875_),
    .B(_03874_),
    .Y(_03876_));
 NAND2x2_ASAP7_75t_R _33461_ (.A(_03872_),
    .B(_03876_),
    .Y(_03877_));
 NOR2x2_ASAP7_75t_R _33462_ (.A(_03869_),
    .B(_03877_),
    .Y(_03878_));
 NAND2x2_ASAP7_75t_R _33463_ (.A(_03861_),
    .B(_03878_),
    .Y(_03879_));
 NOR2x2_ASAP7_75t_R _33464_ (.A(_03844_),
    .B(_03879_),
    .Y(_03880_));
 NAND2x2_ASAP7_75t_R _33465_ (.A(_03811_),
    .B(_03880_),
    .Y(_03881_));
 NOR2x2_ASAP7_75t_R _33466_ (.A(_03809_),
    .B(net2117),
    .Y(_03882_));
 NAND2x2_ASAP7_75t_R _33467_ (.A(_03809_),
    .B(net2117),
    .Y(_03883_));
 INVx2_ASAP7_75t_R _33468_ (.A(_03883_),
    .Y(_03884_));
 INVx4_ASAP7_75t_R _33469_ (.A(_01539_),
    .Y(_03885_));
 AO21x1_ASAP7_75t_R _33470_ (.A1(net1597),
    .A2(net1104),
    .B(net3175),
    .Y(_03886_));
 AO21x1_ASAP7_75t_R _33471_ (.A1(net2572),
    .A2(_01598_),
    .B(net3175),
    .Y(_03887_));
 NAND2x1_ASAP7_75t_R _33472_ (.A(_03886_),
    .B(_03887_),
    .Y(_03888_));
 AO21x1_ASAP7_75t_R _33473_ (.A1(net1605),
    .A2(_03196_),
    .B(_01735_),
    .Y(_03889_));
 AO21x1_ASAP7_75t_R _33474_ (.A1(net1612),
    .A2(_01674_),
    .B(_01735_),
    .Y(_03890_));
 NAND3x1_ASAP7_75t_R _33475_ (.A(_03889_),
    .B(_03890_),
    .C(_01738_),
    .Y(_03891_));
 NOR2x1_ASAP7_75t_R _33476_ (.A(_03888_),
    .B(_03891_),
    .Y(_03892_));
 AO21x1_ASAP7_75t_R _33477_ (.A1(net2366),
    .A2(net1613),
    .B(_01715_),
    .Y(_03893_));
 NAND2x1_ASAP7_75t_R _33478_ (.A(net1896),
    .B(net1888),
    .Y(_03894_));
 AO21x1_ASAP7_75t_R _33479_ (.A1(_03894_),
    .A2(net1457),
    .B(_01715_),
    .Y(_03895_));
 NAND2x1_ASAP7_75t_R _33480_ (.A(_01599_),
    .B(_01720_),
    .Y(_03896_));
 NAND3x1_ASAP7_75t_R _33481_ (.A(_03893_),
    .B(_03895_),
    .C(_03896_),
    .Y(_03897_));
 AO21x1_ASAP7_75t_R _33482_ (.A1(net2524),
    .A2(net3261),
    .B(net3256),
    .Y(_03898_));
 AO21x1_ASAP7_75t_R _33483_ (.A1(net1613),
    .A2(_01524_),
    .B(net3256),
    .Y(_03899_));
 INVx1_ASAP7_75t_R _33484_ (.A(_03260_),
    .Y(_03900_));
 NAND3x1_ASAP7_75t_R _33485_ (.A(_03898_),
    .B(_03899_),
    .C(_03900_),
    .Y(_03901_));
 NOR2x1_ASAP7_75t_R _33486_ (.A(_03897_),
    .B(_03901_),
    .Y(_03902_));
 NAND2x1_ASAP7_75t_R _33487_ (.A(_03892_),
    .B(_03902_),
    .Y(_03903_));
 AO21x1_ASAP7_75t_R _33488_ (.A1(_01689_),
    .A2(_01674_),
    .B(_01701_),
    .Y(_03904_));
 NAND2x1_ASAP7_75t_R _33489_ (.A(_03242_),
    .B(_03904_),
    .Y(_03905_));
 AO21x1_ASAP7_75t_R _33490_ (.A1(_01630_),
    .A2(_02363_),
    .B(_01685_),
    .Y(_03906_));
 OAI21x1_ASAP7_75t_R _33491_ (.A1(_01511_),
    .A2(_01516_),
    .B(_01696_),
    .Y(_03907_));
 NAND2x2_ASAP7_75t_R _33492_ (.A(_02457_),
    .B(_01696_),
    .Y(_03908_));
 NAND3x2_ASAP7_75t_R _33493_ (.B(_03907_),
    .C(_03908_),
    .Y(_03909_),
    .A(_03906_));
 NOR2x2_ASAP7_75t_R _33494_ (.A(_03905_),
    .B(_03909_),
    .Y(_03910_));
 NAND2x2_ASAP7_75t_R _33495_ (.A(_03259_),
    .B(_02368_),
    .Y(_03911_));
 NAND3x2_ASAP7_75t_R _33496_ (.B(_02855_),
    .C(_03911_),
    .Y(_03912_),
    .A(_02369_));
 OAI21x1_ASAP7_75t_R _33497_ (.A1(net2406),
    .A2(_01526_),
    .B(_02368_),
    .Y(_03913_));
 NAND2x2_ASAP7_75t_R _33498_ (.A(net3257),
    .B(_02368_),
    .Y(_03914_));
 NAND2x2_ASAP7_75t_R _33499_ (.A(_01719_),
    .B(_02368_),
    .Y(_03915_));
 NAND3x2_ASAP7_75t_R _33500_ (.B(_03914_),
    .C(_03915_),
    .Y(_03916_),
    .A(_03913_));
 NOR2x2_ASAP7_75t_R _33501_ (.A(_03912_),
    .B(_03916_),
    .Y(_03917_));
 AO21x1_ASAP7_75t_R _33502_ (.A1(net3261),
    .A2(_02419_),
    .B(net2733),
    .Y(_03918_));
 AO21x1_ASAP7_75t_R _33503_ (.A1(_01678_),
    .A2(net1612),
    .B(net2733),
    .Y(_03919_));
 AO21x1_ASAP7_75t_R _33504_ (.A1(net1104),
    .A2(_01569_),
    .B(net2733),
    .Y(_03920_));
 AND3x2_ASAP7_75t_R _33505_ (.A(_03918_),
    .B(_03919_),
    .C(_03920_),
    .Y(_03921_));
 NAND3x2_ASAP7_75t_R _33506_ (.B(_03917_),
    .C(_03921_),
    .Y(_03922_),
    .A(_03910_));
 NOR2x2_ASAP7_75t_R _33507_ (.A(_03903_),
    .B(_03922_),
    .Y(_03923_));
 AO21x1_ASAP7_75t_R _33508_ (.A1(net2368),
    .A2(net1612),
    .B(_01571_),
    .Y(_03924_));
 NAND2x1_ASAP7_75t_R _33509_ (.A(_02821_),
    .B(_03924_),
    .Y(_03925_));
 OAI21x1_ASAP7_75t_R _33510_ (.A1(_02457_),
    .A2(_02414_),
    .B(_01550_),
    .Y(_03926_));
 AO21x1_ASAP7_75t_R _33511_ (.A1(net3261),
    .A2(_02419_),
    .B(_01543_),
    .Y(_03927_));
 NAND2x1_ASAP7_75t_R _33512_ (.A(_03926_),
    .B(_03927_),
    .Y(_03928_));
 NOR3x1_ASAP7_75t_R _33513_ (.A(_03925_),
    .B(_03928_),
    .C(_01574_),
    .Y(_03929_));
 AO31x2_ASAP7_75t_R _33514_ (.A1(net2257),
    .A2(net2065),
    .A3(_01699_),
    .B(_01603_),
    .Y(_03930_));
 AO21x1_ASAP7_75t_R _33515_ (.A1(_01590_),
    .A2(net3255),
    .B(_01603_),
    .Y(_03931_));
 AND2x2_ASAP7_75t_R _33516_ (.A(_01614_),
    .B(_03931_),
    .Y(_03932_));
 NAND2x1_ASAP7_75t_R _33517_ (.A(_03930_),
    .B(_03932_),
    .Y(_03933_));
 AOI22x1_ASAP7_75t_R _33518_ (.A1(_02437_),
    .A2(net1026),
    .B1(net3257),
    .B2(_02829_),
    .Y(_03934_));
 NOR2x1_ASAP7_75t_R _33519_ (.A(_01732_),
    .B(_01586_),
    .Y(_03935_));
 INVx1_ASAP7_75t_R _33520_ (.A(_03935_),
    .Y(_03936_));
 AND2x2_ASAP7_75t_R _33521_ (.A(_03213_),
    .B(_03936_),
    .Y(_03937_));
 NAND2x1_ASAP7_75t_R _33522_ (.A(_03934_),
    .B(_03937_),
    .Y(_03938_));
 NOR2x1_ASAP7_75t_R _33523_ (.A(_03933_),
    .B(_03938_),
    .Y(_03939_));
 NAND2x1_ASAP7_75t_R _33524_ (.A(_03929_),
    .B(_03939_),
    .Y(_03940_));
 AOI221x1_ASAP7_75t_R _33525_ (.A1(net1120),
    .A2(_01494_),
    .B1(net2077),
    .B2(_01644_),
    .C(_01505_),
    .Y(_03941_));
 NAND2x2_ASAP7_75t_R _33526_ (.A(_02427_),
    .B(_02426_),
    .Y(_03942_));
 NOR3x2_ASAP7_75t_R _33527_ (.B(_03415_),
    .C(_03942_),
    .Y(_03943_),
    .A(_03941_));
 AO21x1_ASAP7_75t_R _33528_ (.A1(net1597),
    .A2(_01644_),
    .B(_01636_),
    .Y(_03944_));
 OAI21x1_ASAP7_75t_R _33529_ (.A1(net2746),
    .A2(_01691_),
    .B(_03944_),
    .Y(_03945_));
 AO21x1_ASAP7_75t_R _33530_ (.A1(_01630_),
    .A2(net1104),
    .B(_01624_),
    .Y(_03946_));
 OAI21x1_ASAP7_75t_R _33531_ (.A1(_02414_),
    .A2(_01549_),
    .B(_01621_),
    .Y(_03947_));
 NAND2x2_ASAP7_75t_R _33532_ (.A(net1889),
    .B(_01621_),
    .Y(_03948_));
 NAND3x2_ASAP7_75t_R _33533_ (.B(_03947_),
    .C(_03948_),
    .Y(_03949_),
    .A(_03946_));
 NOR2x2_ASAP7_75t_R _33534_ (.A(_03945_),
    .B(_03949_),
    .Y(_03950_));
 AO21x1_ASAP7_75t_R _33535_ (.A1(net1104),
    .A2(_01612_),
    .B(_01532_),
    .Y(_03951_));
 AO21x1_ASAP7_75t_R _33536_ (.A1(net3261),
    .A2(_02419_),
    .B(net2334),
    .Y(_03952_));
 NAND2x1_ASAP7_75t_R _33537_ (.A(_03951_),
    .B(_03952_),
    .Y(_03953_));
 AO21x2_ASAP7_75t_R _33538_ (.A1(net2572),
    .A2(net2254),
    .B(net2334),
    .Y(_03954_));
 OAI21x1_ASAP7_75t_R _33539_ (.A1(_01600_),
    .A2(net2335),
    .B(_03954_),
    .Y(_03955_));
 NOR2x2_ASAP7_75t_R _33540_ (.A(_03953_),
    .B(_03955_),
    .Y(_03956_));
 NAND3x2_ASAP7_75t_R _33541_ (.B(_03950_),
    .C(_03956_),
    .Y(_03957_),
    .A(_03943_));
 NOR2x2_ASAP7_75t_R _33542_ (.A(_03940_),
    .B(_03957_),
    .Y(_03958_));
 NAND2x2_ASAP7_75t_R _33543_ (.A(_03923_),
    .B(_03958_),
    .Y(_03959_));
 NOR2x2_ASAP7_75t_R _33544_ (.A(_03885_),
    .B(_03959_),
    .Y(_03960_));
 OAI21x1_ASAP7_75t_R _33545_ (.A1(_03882_),
    .A2(_03884_),
    .B(_03960_),
    .Y(_03961_));
 INVx1_ASAP7_75t_R _33546_ (.A(_03778_),
    .Y(_03962_));
 NOR2x1_ASAP7_75t_R _33547_ (.A(_03788_),
    .B(_03962_),
    .Y(_03963_));
 INVx1_ASAP7_75t_R _33548_ (.A(_03800_),
    .Y(_03964_));
 NAND2x1_ASAP7_75t_R _33549_ (.A(_03805_),
    .B(_03793_),
    .Y(_03965_));
 NOR2x1_ASAP7_75t_R _33550_ (.A(_03964_),
    .B(_03965_),
    .Y(_03966_));
 NAND2x1_ASAP7_75t_R _33551_ (.A(_03963_),
    .B(_03966_),
    .Y(_03967_));
 INVx2_ASAP7_75t_R _33552_ (.A(_03772_),
    .Y(_03968_));
 NOR2x2_ASAP7_75t_R _33553_ (.A(_03967_),
    .B(_03968_),
    .Y(_03969_));
 NAND2x2_ASAP7_75t_R _33554_ (.A(net2791),
    .B(_03969_),
    .Y(_03970_));
 NOR2x2_ASAP7_75t_R _33555_ (.A(_03970_),
    .B(net2117),
    .Y(_03971_));
 AOI21x1_ASAP7_75t_R _33556_ (.A1(_03811_),
    .A2(_03880_),
    .B(net3287),
    .Y(_03972_));
 NAND3x2_ASAP7_75t_R _33557_ (.B(_03958_),
    .C(_03923_),
    .Y(_03973_),
    .A(net3127));
 OAI21x1_ASAP7_75t_R _33558_ (.A1(_03971_),
    .A2(_03972_),
    .B(_03973_),
    .Y(_03974_));
 AO21x1_ASAP7_75t_R _33559_ (.A1(net1253),
    .A2(net2286),
    .B(_01916_),
    .Y(_03975_));
 OA21x2_ASAP7_75t_R _33560_ (.A1(_01761_),
    .A2(_02988_),
    .B(_03975_),
    .Y(_03976_));
 AO21x1_ASAP7_75t_R _33561_ (.A1(net3254),
    .A2(net1157),
    .B(_01955_),
    .Y(_03977_));
 AND4x1_ASAP7_75t_R _33562_ (.A(_03670_),
    .B(_03977_),
    .C(_03679_),
    .D(_03632_),
    .Y(_03978_));
 NAND2x1_ASAP7_75t_R _33563_ (.A(_03976_),
    .B(_03978_),
    .Y(_03979_));
 NOR2x1_ASAP7_75t_R _33564_ (.A(_01938_),
    .B(_01809_),
    .Y(_03980_));
 AOI21x1_ASAP7_75t_R _33565_ (.A1(_01762_),
    .A2(_02136_),
    .B(_03980_),
    .Y(_03981_));
 OA21x2_ASAP7_75t_R _33566_ (.A1(net2306),
    .A2(_01936_),
    .B(_01942_),
    .Y(_03982_));
 NAND2x1_ASAP7_75t_R _33567_ (.A(_03981_),
    .B(_03982_),
    .Y(_03983_));
 NOR2x1_ASAP7_75t_R _33568_ (.A(_03979_),
    .B(_03983_),
    .Y(_03984_));
 AND3x1_ASAP7_75t_R _33569_ (.A(_01888_),
    .B(_01787_),
    .C(_01770_),
    .Y(_03985_));
 INVx1_ASAP7_75t_R _33570_ (.A(_01877_),
    .Y(_03986_));
 NAND2x1_ASAP7_75t_R _33571_ (.A(_01847_),
    .B(_03986_),
    .Y(_03987_));
 OAI21x1_ASAP7_75t_R _33572_ (.A1(net2619),
    .A2(net2140),
    .B(_03987_),
    .Y(_03988_));
 AOI211x1_ASAP7_75t_R _33573_ (.A1(_02131_),
    .A2(_01816_),
    .B(_03985_),
    .C(_03988_),
    .Y(_03989_));
 AOI21x1_ASAP7_75t_R _33574_ (.A1(_01806_),
    .A2(_01974_),
    .B(_02991_),
    .Y(_03990_));
 AO21x1_ASAP7_75t_R _33575_ (.A1(_01905_),
    .A2(_01828_),
    .B(net1527),
    .Y(_03991_));
 AO21x1_ASAP7_75t_R _33576_ (.A1(_01977_),
    .A2(net2352),
    .B(_01821_),
    .Y(_03992_));
 AND2x2_ASAP7_75t_R _33577_ (.A(_03991_),
    .B(_03992_),
    .Y(_03993_));
 NAND3x1_ASAP7_75t_R _33578_ (.A(_03989_),
    .B(_03990_),
    .C(_03993_),
    .Y(_03994_));
 NAND2x1_ASAP7_75t_R _33579_ (.A(net2330),
    .B(_01930_),
    .Y(_03995_));
 NAND2x1_ASAP7_75t_R _33580_ (.A(_01847_),
    .B(_01806_),
    .Y(_03996_));
 AND4x1_ASAP7_75t_R _33581_ (.A(_02571_),
    .B(_01872_),
    .C(_03995_),
    .D(_03996_),
    .Y(_03997_));
 OA21x2_ASAP7_75t_R _33582_ (.A1(net2286),
    .A2(_01828_),
    .B(_03692_),
    .Y(_03998_));
 AND3x1_ASAP7_75t_R _33583_ (.A(_03998_),
    .B(_02910_),
    .C(_02906_),
    .Y(_03999_));
 NAND2x1_ASAP7_75t_R _33584_ (.A(_03997_),
    .B(_03999_),
    .Y(_04000_));
 NOR2x1_ASAP7_75t_R _33585_ (.A(_03994_),
    .B(_04000_),
    .Y(_04001_));
 NAND2x1_ASAP7_75t_R _33586_ (.A(_03984_),
    .B(_04001_),
    .Y(_04002_));
 NAND2x1_ASAP7_75t_R _33587_ (.A(_03655_),
    .B(_01816_),
    .Y(_04003_));
 NAND2x1_ASAP7_75t_R _33588_ (.A(_01784_),
    .B(_03622_),
    .Y(_04004_));
 AND4x1_ASAP7_75t_R _33589_ (.A(_03640_),
    .B(_04003_),
    .C(_03704_),
    .D(_04004_),
    .Y(_04005_));
 AOI22x1_ASAP7_75t_R _33590_ (.A1(_02151_),
    .A2(_01974_),
    .B1(net2654),
    .B2(_02141_),
    .Y(_04006_));
 OA21x2_ASAP7_75t_R _33591_ (.A1(_01828_),
    .A2(_02134_),
    .B(_04006_),
    .Y(_04007_));
 OR3x1_ASAP7_75t_R _33592_ (.A(_01851_),
    .B(net1451),
    .C(_01857_),
    .Y(_04008_));
 AND2x2_ASAP7_75t_R _33593_ (.A(_04008_),
    .B(_02118_),
    .Y(_04009_));
 NAND3x1_ASAP7_75t_R _33594_ (.A(_04005_),
    .B(_04007_),
    .C(_04009_),
    .Y(_04010_));
 AO21x1_ASAP7_75t_R _33595_ (.A1(_02498_),
    .A2(net2301),
    .B(_02535_),
    .Y(_04011_));
 AO21x1_ASAP7_75t_R _33596_ (.A1(net1253),
    .A2(_01821_),
    .B(_01781_),
    .Y(_04012_));
 INVx1_ASAP7_75t_R _33597_ (.A(_04012_),
    .Y(_04013_));
 AO221x1_ASAP7_75t_R _33598_ (.A1(_02131_),
    .A2(_01843_),
    .B1(_02211_),
    .B2(_04011_),
    .C(_04013_),
    .Y(_04014_));
 NOR2x1_ASAP7_75t_R _33599_ (.A(_04010_),
    .B(_04014_),
    .Y(_04015_));
 OA211x2_ASAP7_75t_R _33600_ (.A1(net2300),
    .A2(net1556),
    .B(_01970_),
    .C(_01818_),
    .Y(_04016_));
 AND3x1_ASAP7_75t_R _33601_ (.A(_01830_),
    .B(_00595_),
    .C(_01845_),
    .Y(_04017_));
 AO21x1_ASAP7_75t_R _33602_ (.A1(net1116),
    .A2(_04017_),
    .B(_01891_),
    .Y(_04018_));
 NOR2x1_ASAP7_75t_R _33603_ (.A(_04016_),
    .B(_04018_),
    .Y(_04019_));
 NOR2x1_ASAP7_75t_R _33604_ (.A(_01878_),
    .B(_01824_),
    .Y(_04020_));
 INVx1_ASAP7_75t_R _33605_ (.A(_04020_),
    .Y(_04021_));
 INVx1_ASAP7_75t_R _33606_ (.A(_02483_),
    .Y(_04022_));
 AND4x1_ASAP7_75t_R _33607_ (.A(_02101_),
    .B(_02186_),
    .C(_04021_),
    .D(_04022_),
    .Y(_04023_));
 NAND2x1_ASAP7_75t_R _33608_ (.A(_04019_),
    .B(_04023_),
    .Y(_04024_));
 NAND2x1_ASAP7_75t_R _33609_ (.A(_02918_),
    .B(_01762_),
    .Y(_04025_));
 AND4x1_ASAP7_75t_R _33610_ (.A(_04025_),
    .B(_02924_),
    .C(_02198_),
    .D(_02522_),
    .Y(_04026_));
 AOI22x1_ASAP7_75t_R _33611_ (.A1(_01816_),
    .A2(_03622_),
    .B1(_01806_),
    .B2(_02141_),
    .Y(_04027_));
 AO21x1_ASAP7_75t_R _33612_ (.A1(net1527),
    .A2(net1157),
    .B(net2140),
    .Y(_04028_));
 AND3x1_ASAP7_75t_R _33613_ (.A(_04027_),
    .B(_01950_),
    .C(_04028_),
    .Y(_04029_));
 NAND2x1_ASAP7_75t_R _33614_ (.A(_04026_),
    .B(_04029_),
    .Y(_04030_));
 AO21x1_ASAP7_75t_R _33615_ (.A1(_02500_),
    .A2(_01857_),
    .B(net2263),
    .Y(_04031_));
 NAND2x1_ASAP7_75t_R _33616_ (.A(_01930_),
    .B(_01886_),
    .Y(_04032_));
 AND3x1_ASAP7_75t_R _33617_ (.A(_04031_),
    .B(_04032_),
    .C(_03663_),
    .Y(_04033_));
 NAND2x1_ASAP7_75t_R _33618_ (.A(net1558),
    .B(_01940_),
    .Y(_04034_));
 OA21x2_ASAP7_75t_R _33619_ (.A1(_02559_),
    .A2(net2352),
    .B(_04034_),
    .Y(_04035_));
 OA21x2_ASAP7_75t_R _33620_ (.A1(_02110_),
    .A2(_01936_),
    .B(_02519_),
    .Y(_04036_));
 AND2x2_ASAP7_75t_R _33621_ (.A(_04035_),
    .B(_04036_),
    .Y(_04037_));
 NAND2x1_ASAP7_75t_R _33622_ (.A(_04033_),
    .B(_04037_),
    .Y(_04038_));
 NOR3x1_ASAP7_75t_R _33623_ (.A(_04024_),
    .B(_04030_),
    .C(_04038_),
    .Y(_04039_));
 NAND2x1_ASAP7_75t_R _33624_ (.A(_04015_),
    .B(_04039_),
    .Y(_04040_));
 NOR2x2_ASAP7_75t_R _33625_ (.A(_04002_),
    .B(_04040_),
    .Y(_04041_));
 XNOR2x2_ASAP7_75t_R _33626_ (.A(_03539_),
    .B(_04041_),
    .Y(_04042_));
 INVx1_ASAP7_75t_R _33627_ (.A(_04042_),
    .Y(_04043_));
 NAND3x2_ASAP7_75t_R _33628_ (.B(_03974_),
    .C(_04043_),
    .Y(_04044_),
    .A(_03961_));
 INVx2_ASAP7_75t_R _33629_ (.A(_03882_),
    .Y(_04045_));
 AOI21x1_ASAP7_75t_R _33630_ (.A1(_03883_),
    .A2(_04045_),
    .B(_03973_),
    .Y(_04046_));
 NAND2x2_ASAP7_75t_R _33631_ (.A(_03881_),
    .B(_03970_),
    .Y(_04047_));
 INVx2_ASAP7_75t_R _33632_ (.A(_03971_),
    .Y(_04048_));
 AOI21x1_ASAP7_75t_R _33633_ (.A1(_04047_),
    .A2(_04048_),
    .B(_03960_),
    .Y(_04049_));
 OAI21x1_ASAP7_75t_R _33634_ (.A1(_04046_),
    .A2(_04049_),
    .B(_04042_),
    .Y(_04050_));
 NAND3x1_ASAP7_75t_R _33635_ (.A(_04044_),
    .B(net395),
    .C(_04050_),
    .Y(_04051_));
 INVx1_ASAP7_75t_R _33636_ (.A(_00479_),
    .Y(_04052_));
 AOI21x1_ASAP7_75t_R _33637_ (.A1(_03726_),
    .A2(_04051_),
    .B(_04052_),
    .Y(_04053_));
 OR2x2_ASAP7_75t_R _33638_ (.A(net395),
    .B(_00878_),
    .Y(_04054_));
 AO21x1_ASAP7_75t_R _33639_ (.A1(_04044_),
    .A2(_04050_),
    .B(_18753_),
    .Y(_04055_));
 AOI21x1_ASAP7_75t_R _33640_ (.A1(_04054_),
    .A2(_04055_),
    .B(_00479_),
    .Y(_04056_));
 NOR2x1_ASAP7_75t_R _33641_ (.A(_04053_),
    .B(_04056_),
    .Y(_00118_));
 NOR2x1_ASAP7_75t_R _33642_ (.A(net395),
    .B(_00877_),
    .Y(_04057_));
 NOR2x1_ASAP7_75t_R _33643_ (.A(_01276_),
    .B(_01113_),
    .Y(_04058_));
 OR3x1_ASAP7_75t_R _33644_ (.A(_01281_),
    .B(_04058_),
    .C(_01278_),
    .Y(_04059_));
 NAND2x1_ASAP7_75t_R _33645_ (.A(_01361_),
    .B(_02665_),
    .Y(_04060_));
 AO21x1_ASAP7_75t_R _33646_ (.A1(net3320),
    .A2(_01259_),
    .B(net3417),
    .Y(_04061_));
 INVx1_ASAP7_75t_R _33647_ (.A(_04061_),
    .Y(_04062_));
 NOR3x1_ASAP7_75t_R _33648_ (.A(_04059_),
    .B(_04060_),
    .C(_04062_),
    .Y(_04063_));
 NAND2x1_ASAP7_75t_R _33649_ (.A(_03030_),
    .B(_01412_),
    .Y(_04064_));
 AO21x1_ASAP7_75t_R _33650_ (.A1(net1802),
    .A2(_01148_),
    .B(net3315),
    .Y(_04065_));
 OAI21x1_ASAP7_75t_R _33651_ (.A1(net3315),
    .A2(_01153_),
    .B(_04065_),
    .Y(_04066_));
 OR2x2_ASAP7_75t_R _33652_ (.A(_04064_),
    .B(_04066_),
    .Y(_04067_));
 OA21x2_ASAP7_75t_R _33653_ (.A1(_01173_),
    .A2(_01166_),
    .B(_01251_),
    .Y(_04068_));
 OR3x1_ASAP7_75t_R _33654_ (.A(_04068_),
    .B(_03845_),
    .C(_01407_),
    .Y(_04069_));
 NOR2x1_ASAP7_75t_R _33655_ (.A(_04067_),
    .B(_04069_),
    .Y(_04070_));
 NAND2x1_ASAP7_75t_R _33656_ (.A(_04063_),
    .B(_04070_),
    .Y(_04071_));
 AO21x1_ASAP7_75t_R _33657_ (.A1(_01113_),
    .A2(_01138_),
    .B(_01345_),
    .Y(_04072_));
 OAI21x1_ASAP7_75t_R _33658_ (.A1(net3240),
    .A2(_01226_),
    .B(_04072_),
    .Y(_04073_));
 OAI21x1_ASAP7_75t_R _33659_ (.A1(net2544),
    .A2(net3240),
    .B(_01349_),
    .Y(_04074_));
 AO21x1_ASAP7_75t_R _33660_ (.A1(_01160_),
    .A2(_01351_),
    .B(_03011_),
    .Y(_04075_));
 NOR3x2_ASAP7_75t_R _33661_ (.B(_04074_),
    .C(_04075_),
    .Y(_04076_),
    .A(_04073_));
 AO21x1_ASAP7_75t_R _33662_ (.A1(_01306_),
    .A2(_01226_),
    .B(net2460),
    .Y(_04077_));
 AO21x1_ASAP7_75t_R _33663_ (.A1(_01348_),
    .A2(_01204_),
    .B(net2460),
    .Y(_04078_));
 NAND3x2_ASAP7_75t_R _33664_ (.B(_04077_),
    .C(_04078_),
    .Y(_04079_),
    .A(_03017_));
 AO21x1_ASAP7_75t_R _33665_ (.A1(net1158),
    .A2(net1266),
    .B(_01308_),
    .Y(_04080_));
 AO21x1_ASAP7_75t_R _33666_ (.A1(net1884),
    .A2(net1119),
    .B(_01308_),
    .Y(_04081_));
 NAND2x2_ASAP7_75t_R _33667_ (.A(_01233_),
    .B(_01315_),
    .Y(_04082_));
 NAND3x2_ASAP7_75t_R _33668_ (.B(_04081_),
    .C(_04082_),
    .Y(_04083_),
    .A(_04080_));
 NOR2x2_ASAP7_75t_R _33669_ (.A(_04079_),
    .B(_04083_),
    .Y(_04084_));
 AO21x1_ASAP7_75t_R _33670_ (.A1(_01113_),
    .A2(net2651),
    .B(_01334_),
    .Y(_04085_));
 AO21x1_ASAP7_75t_R _33671_ (.A1(net1119),
    .A2(_01143_),
    .B(_01334_),
    .Y(_04086_));
 AND3x2_ASAP7_75t_R _33672_ (.A(_04085_),
    .B(_04086_),
    .C(_01373_),
    .Y(_04087_));
 NAND3x2_ASAP7_75t_R _33673_ (.B(_04084_),
    .C(_04087_),
    .Y(_04088_),
    .A(_04076_));
 NOR2x2_ASAP7_75t_R _33674_ (.A(_04071_),
    .B(_04088_),
    .Y(_04089_));
 AO21x1_ASAP7_75t_R _33675_ (.A1(_01113_),
    .A2(_01226_),
    .B(_01191_),
    .Y(_04090_));
 AO21x1_ASAP7_75t_R _33676_ (.A1(net1158),
    .A2(_01303_),
    .B(_01191_),
    .Y(_04091_));
 AO21x1_ASAP7_75t_R _33677_ (.A1(net1884),
    .A2(net1119),
    .B(_01191_),
    .Y(_04092_));
 NAND2x1_ASAP7_75t_R _33678_ (.A(_01233_),
    .B(_01197_),
    .Y(_04093_));
 AND4x2_ASAP7_75t_R _33679_ (.A(_04090_),
    .B(_04091_),
    .C(_04092_),
    .D(_04093_),
    .Y(_04094_));
 AO21x1_ASAP7_75t_R _33680_ (.A1(_01138_),
    .A2(net2731),
    .B(_01202_),
    .Y(_04095_));
 NAND2x1_ASAP7_75t_R _33681_ (.A(_01210_),
    .B(_01173_),
    .Y(_04096_));
 NAND2x1_ASAP7_75t_R _33682_ (.A(_02023_),
    .B(_01210_),
    .Y(_04097_));
 AND4x2_ASAP7_75t_R _33683_ (.A(_01433_),
    .B(_04095_),
    .C(_04096_),
    .D(_04097_),
    .Y(_04098_));
 AO21x1_ASAP7_75t_R _33684_ (.A1(net940),
    .A2(_01447_),
    .B(_01229_),
    .Y(_04099_));
 AO21x1_ASAP7_75t_R _33685_ (.A1(_01228_),
    .A2(_01306_),
    .B(_01229_),
    .Y(_04100_));
 NAND2x1_ASAP7_75t_R _33686_ (.A(_04099_),
    .B(_04100_),
    .Y(_04101_));
 AO21x1_ASAP7_75t_R _33687_ (.A1(net1158),
    .A2(net938),
    .B(_01215_),
    .Y(_04102_));
 AO21x1_ASAP7_75t_R _33688_ (.A1(net1884),
    .A2(net1076),
    .B(_01215_),
    .Y(_04103_));
 NAND2x2_ASAP7_75t_R _33689_ (.A(_01270_),
    .B(_01218_),
    .Y(_04104_));
 NAND3x2_ASAP7_75t_R _33690_ (.B(_04103_),
    .C(_04104_),
    .Y(_04105_),
    .A(_04102_));
 NOR2x2_ASAP7_75t_R _33691_ (.A(_04101_),
    .B(_04105_),
    .Y(_04106_));
 NAND3x2_ASAP7_75t_R _33692_ (.B(_04098_),
    .C(_04106_),
    .Y(_04107_),
    .A(_04094_));
 OAI21x1_ASAP7_75t_R _33693_ (.A1(_01259_),
    .A2(_01156_),
    .B(_02034_),
    .Y(_04108_));
 AOI211x1_ASAP7_75t_R _33694_ (.A1(_01474_),
    .A2(_01163_),
    .B(_04108_),
    .C(_03082_),
    .Y(_04109_));
 AO21x1_ASAP7_75t_R _33695_ (.A1(net1158),
    .A2(_01303_),
    .B(_01120_),
    .Y(_04110_));
 NAND2x2_ASAP7_75t_R _33696_ (.A(_04110_),
    .B(_01458_),
    .Y(_04111_));
 AO21x1_ASAP7_75t_R _33697_ (.A1(_01348_),
    .A2(_01447_),
    .B(_01133_),
    .Y(_04112_));
 AO21x1_ASAP7_75t_R _33698_ (.A1(_01113_),
    .A2(_02032_),
    .B(_01133_),
    .Y(_04113_));
 NAND2x2_ASAP7_75t_R _33699_ (.A(_04112_),
    .B(_04113_),
    .Y(_04114_));
 AO21x1_ASAP7_75t_R _33700_ (.A1(_01153_),
    .A2(net1122),
    .B(_01120_),
    .Y(_04115_));
 AO21x1_ASAP7_75t_R _33701_ (.A1(net1884),
    .A2(net1119),
    .B(_01120_),
    .Y(_04116_));
 NAND2x2_ASAP7_75t_R _33702_ (.A(_04115_),
    .B(_04116_),
    .Y(_04117_));
 NOR3x2_ASAP7_75t_R _33703_ (.B(_04114_),
    .C(_04117_),
    .Y(_04118_),
    .A(_04111_));
 AO21x1_ASAP7_75t_R _33704_ (.A1(net1158),
    .A2(net1266),
    .B(_01170_),
    .Y(_04119_));
 AO21x1_ASAP7_75t_R _33705_ (.A1(_01306_),
    .A2(_01226_),
    .B(_01170_),
    .Y(_04120_));
 AO21x1_ASAP7_75t_R _33706_ (.A1(_01153_),
    .A2(_01221_),
    .B(_01170_),
    .Y(_04121_));
 AND3x2_ASAP7_75t_R _33707_ (.A(_04119_),
    .B(_04120_),
    .C(_04121_),
    .Y(_04122_));
 NAND3x2_ASAP7_75t_R _33708_ (.B(_04118_),
    .C(_04122_),
    .Y(_04123_),
    .A(_04109_));
 NOR2x2_ASAP7_75t_R _33709_ (.A(_04107_),
    .B(_04123_),
    .Y(_04124_));
 NAND2x2_ASAP7_75t_R _33710_ (.A(_04089_),
    .B(_04124_),
    .Y(_04125_));
 NOR2x2_ASAP7_75t_R _33711_ (.A(_01371_),
    .B(_04125_),
    .Y(_04126_));
 AO21x1_ASAP7_75t_R _33712_ (.A1(_22019_),
    .A2(_21895_),
    .B(net3151),
    .Y(_04127_));
 AND3x1_ASAP7_75t_R _33713_ (.A(_03119_),
    .B(_21996_),
    .C(_04127_),
    .Y(_04128_));
 AO21x1_ASAP7_75t_R _33714_ (.A1(net3172),
    .A2(net1048),
    .B(net3148),
    .Y(_04129_));
 AO21x1_ASAP7_75t_R _33715_ (.A1(net991),
    .A2(_03133_),
    .B(net3148),
    .Y(_04130_));
 NAND3x1_ASAP7_75t_R _33716_ (.A(_04128_),
    .B(_04129_),
    .C(_04130_),
    .Y(_04131_));
 AO21x1_ASAP7_75t_R _33717_ (.A1(net1829),
    .A2(net3172),
    .B(net3075),
    .Y(_04132_));
 AO21x1_ASAP7_75t_R _33718_ (.A1(_21995_),
    .A2(net3280),
    .B(net3075),
    .Y(_04133_));
 NAND2x1_ASAP7_75t_R _33719_ (.A(_03107_),
    .B(_22016_),
    .Y(_04134_));
 AND4x1_ASAP7_75t_R _33720_ (.A(_04132_),
    .B(_04133_),
    .C(_22022_),
    .D(_04134_),
    .Y(_04135_));
 AOI22x1_ASAP7_75t_R _33721_ (.A1(_02348_),
    .A2(_21879_),
    .B1(_22034_),
    .B2(_01082_),
    .Y(_04136_));
 NAND2x1_ASAP7_75t_R _33722_ (.A(_22053_),
    .B(_22034_),
    .Y(_04137_));
 AO21x1_ASAP7_75t_R _33723_ (.A1(_22076_),
    .A2(_21929_),
    .B(net2556),
    .Y(_04138_));
 AND3x1_ASAP7_75t_R _33724_ (.A(_04136_),
    .B(_04137_),
    .C(_04138_),
    .Y(_04139_));
 NAND2x1_ASAP7_75t_R _33725_ (.A(_04135_),
    .B(_04139_),
    .Y(_04140_));
 NOR2x1_ASAP7_75t_R _33726_ (.A(_04131_),
    .B(_04140_),
    .Y(_04141_));
 AND2x2_ASAP7_75t_R _33727_ (.A(_21911_),
    .B(_02774_),
    .Y(_04142_));
 AO21x1_ASAP7_75t_R _33728_ (.A1(_22076_),
    .A2(_21944_),
    .B(net1751),
    .Y(_04143_));
 AO21x1_ASAP7_75t_R _33729_ (.A1(net1048),
    .A2(_22080_),
    .B(net1751),
    .Y(_04144_));
 AO21x1_ASAP7_75t_R _33730_ (.A1(net2365),
    .A2(_21969_),
    .B(net1751),
    .Y(_04145_));
 NAND2x1_ASAP7_75t_R _33731_ (.A(_22053_),
    .B(_02323_),
    .Y(_04146_));
 AND4x1_ASAP7_75t_R _33732_ (.A(_04143_),
    .B(_04144_),
    .C(_04145_),
    .D(_04146_),
    .Y(_04147_));
 NAND2x1_ASAP7_75t_R _33733_ (.A(_04142_),
    .B(_04147_),
    .Y(_04148_));
 OA21x2_ASAP7_75t_R _33734_ (.A1(_02765_),
    .A2(_03107_),
    .B(_21980_),
    .Y(_04149_));
 INVx2_ASAP7_75t_R _33735_ (.A(_21978_),
    .Y(_04150_));
 NOR2x1_ASAP7_75t_R _33736_ (.A(_21976_),
    .B(_04150_),
    .Y(_04151_));
 NOR2x1_ASAP7_75t_R _33737_ (.A(net2510),
    .B(_21976_),
    .Y(_04152_));
 OR3x1_ASAP7_75t_R _33738_ (.A(_04149_),
    .B(_04151_),
    .C(_04152_),
    .Y(_04153_));
 INVx1_ASAP7_75t_R _33739_ (.A(_04153_),
    .Y(_04154_));
 OA21x2_ASAP7_75t_R _33740_ (.A1(_22053_),
    .A2(_02269_),
    .B(_21957_),
    .Y(_04155_));
 NOR2x1_ASAP7_75t_R _33741_ (.A(_03099_),
    .B(_04155_),
    .Y(_04156_));
 NAND2x1_ASAP7_75t_R _33742_ (.A(_21957_),
    .B(_02316_),
    .Y(_04157_));
 AO21x1_ASAP7_75t_R _33743_ (.A1(net2752),
    .A2(net991),
    .B(_21962_),
    .Y(_04158_));
 AND3x1_ASAP7_75t_R _33744_ (.A(_04156_),
    .B(_04157_),
    .C(_04158_),
    .Y(_04159_));
 NAND2x1_ASAP7_75t_R _33745_ (.A(_04154_),
    .B(_04159_),
    .Y(_04160_));
 NOR2x2_ASAP7_75t_R _33746_ (.A(_04148_),
    .B(_04160_),
    .Y(_04161_));
 NAND2x2_ASAP7_75t_R _33747_ (.A(_04141_),
    .B(_04161_),
    .Y(_04162_));
 AO21x1_ASAP7_75t_R _33748_ (.A1(_22024_),
    .A2(net1792),
    .B(_01072_),
    .Y(_04163_));
 AO21x1_ASAP7_75t_R _33749_ (.A1(net1038),
    .A2(_22019_),
    .B(_01072_),
    .Y(_04164_));
 NAND2x1_ASAP7_75t_R _33750_ (.A(_03107_),
    .B(_01073_),
    .Y(_04165_));
 AND3x1_ASAP7_75t_R _33751_ (.A(_04163_),
    .B(_04164_),
    .C(_04165_),
    .Y(_04166_));
 OAI21x1_ASAP7_75t_R _33752_ (.A1(net3083),
    .A2(net2039),
    .B(_01079_),
    .Y(_04167_));
 AO21x1_ASAP7_75t_R _33753_ (.A1(net1829),
    .A2(net1048),
    .B(net2424),
    .Y(_04168_));
 NAND2x1_ASAP7_75t_R _33754_ (.A(_04167_),
    .B(_04168_),
    .Y(_04169_));
 AO21x1_ASAP7_75t_R _33755_ (.A1(net1038),
    .A2(net3225),
    .B(net2424),
    .Y(_04170_));
 OAI21x1_ASAP7_75t_R _33756_ (.A1(net991),
    .A2(net2424),
    .B(_04170_),
    .Y(_04171_));
 NOR2x1_ASAP7_75t_R _33757_ (.A(_04171_),
    .B(_04169_),
    .Y(_04172_));
 NAND2x1_ASAP7_75t_R _33758_ (.A(_04166_),
    .B(_04172_),
    .Y(_04173_));
 OA211x2_ASAP7_75t_R _33759_ (.A1(_21887_),
    .A2(_21876_),
    .B(_22092_),
    .C(net2589),
    .Y(_04174_));
 INVx1_ASAP7_75t_R _33760_ (.A(_04174_),
    .Y(_04175_));
 AO21x1_ASAP7_75t_R _33761_ (.A1(_21995_),
    .A2(_22080_),
    .B(net3081),
    .Y(_04176_));
 AO21x1_ASAP7_75t_R _33762_ (.A1(net2510),
    .A2(_22057_),
    .B(net3081),
    .Y(_04177_));
 AND2x2_ASAP7_75t_R _33763_ (.A(_04176_),
    .B(_04177_),
    .Y(_04178_));
 AO21x1_ASAP7_75t_R _33764_ (.A1(net3225),
    .A2(net991),
    .B(_22091_),
    .Y(_04179_));
 NAND3x2_ASAP7_75t_R _33765_ (.B(_04178_),
    .C(_04179_),
    .Y(_04180_),
    .A(_04175_));
 NOR2x2_ASAP7_75t_R _33766_ (.A(_04180_),
    .B(_04173_),
    .Y(_04181_));
 AO21x1_ASAP7_75t_R _33767_ (.A1(_22019_),
    .A2(_22057_),
    .B(_22070_),
    .Y(_04182_));
 AND3x1_ASAP7_75t_R _33768_ (.A(_04182_),
    .B(_02728_),
    .C(_03746_),
    .Y(_04183_));
 OAI21x1_ASAP7_75t_R _33769_ (.A1(net3083),
    .A2(net2040),
    .B(_22084_),
    .Y(_04184_));
 OA21x2_ASAP7_75t_R _33770_ (.A1(_21876_),
    .A2(_02295_),
    .B(_04184_),
    .Y(_04185_));
 AO21x1_ASAP7_75t_R _33771_ (.A1(net1038),
    .A2(_21983_),
    .B(_22077_),
    .Y(_04186_));
 AO21x1_ASAP7_75t_R _33772_ (.A1(_22008_),
    .A2(_02273_),
    .B(_22077_),
    .Y(_04187_));
 AND2x2_ASAP7_75t_R _33773_ (.A(_04186_),
    .B(_04187_),
    .Y(_04188_));
 AND3x2_ASAP7_75t_R _33774_ (.A(_04183_),
    .B(_04185_),
    .C(_04188_),
    .Y(_04189_));
 OA21x2_ASAP7_75t_R _33775_ (.A1(_02765_),
    .A2(_22014_),
    .B(_22062_),
    .Y(_04190_));
 NOR2x2_ASAP7_75t_R _33776_ (.A(_04190_),
    .B(_02287_),
    .Y(_04191_));
 NAND2x2_ASAP7_75t_R _33777_ (.A(net3083),
    .B(_22062_),
    .Y(_04192_));
 NAND3x2_ASAP7_75t_R _33778_ (.B(_04192_),
    .C(_03139_),
    .Y(_04193_),
    .A(_04191_));
 AOI211x1_ASAP7_75t_R _33779_ (.A1(_01087_),
    .A2(_22049_),
    .B(_03146_),
    .C(_22067_),
    .Y(_04194_));
 OA21x2_ASAP7_75t_R _33780_ (.A1(_01085_),
    .A2(_02269_),
    .B(_22049_),
    .Y(_04195_));
 OA21x2_ASAP7_75t_R _33781_ (.A1(_21909_),
    .A2(net3083),
    .B(_22049_),
    .Y(_04196_));
 AOI211x1_ASAP7_75t_R _33782_ (.A1(net2040),
    .A2(_22049_),
    .B(_04195_),
    .C(_04196_),
    .Y(_04197_));
 NAND2x1_ASAP7_75t_R _33783_ (.A(_04194_),
    .B(_04197_),
    .Y(_04198_));
 NOR2x2_ASAP7_75t_R _33784_ (.A(_04193_),
    .B(_04198_),
    .Y(_04199_));
 NAND3x2_ASAP7_75t_R _33785_ (.B(_04189_),
    .C(_04199_),
    .Y(_04200_),
    .A(_04181_));
 NOR3x2_ASAP7_75t_R _33786_ (.B(_03734_),
    .C(_04200_),
    .Y(_04201_),
    .A(_04162_));
 NOR2x2_ASAP7_75t_R _33787_ (.A(_04201_),
    .B(_04126_),
    .Y(_04202_));
 NAND3x2_ASAP7_75t_R _33788_ (.B(_04089_),
    .C(_04124_),
    .Y(_04203_),
    .A(_03811_));
 NOR2x1_ASAP7_75t_R _33789_ (.A(_04162_),
    .B(_04200_),
    .Y(_04204_));
 NAND2x2_ASAP7_75t_R _33790_ (.A(net2791),
    .B(_04204_),
    .Y(_04205_));
 NOR2x2_ASAP7_75t_R _33791_ (.A(_04203_),
    .B(_04205_),
    .Y(_04206_));
 AO21x1_ASAP7_75t_R _33792_ (.A1(_01727_),
    .A2(_03442_),
    .B(net3256),
    .Y(_04207_));
 NAND2x1_ASAP7_75t_R _33793_ (.A(_02461_),
    .B(_01711_),
    .Y(_04208_));
 AO21x1_ASAP7_75t_R _33794_ (.A1(net3261),
    .A2(net1605),
    .B(net3256),
    .Y(_04209_));
 AND3x1_ASAP7_75t_R _33795_ (.A(_04207_),
    .B(_04208_),
    .C(_04209_),
    .Y(_04210_));
 OAI22x1_ASAP7_75t_R _33796_ (.A1(_03270_),
    .A2(_00634_),
    .B1(net1605),
    .B2(_01715_),
    .Y(_04211_));
 NOR2x1_ASAP7_75t_R _33797_ (.A(_01630_),
    .B(_01715_),
    .Y(_04212_));
 AO21x1_ASAP7_75t_R _33798_ (.A1(_01699_),
    .A2(net1612),
    .B(_01715_),
    .Y(_04213_));
 INVx1_ASAP7_75t_R _33799_ (.A(_04213_),
    .Y(_04214_));
 NOR3x1_ASAP7_75t_R _33800_ (.A(_04211_),
    .B(_04212_),
    .C(_04214_),
    .Y(_04215_));
 NAND2x1_ASAP7_75t_R _33801_ (.A(_04210_),
    .B(_04215_),
    .Y(_04216_));
 AO21x1_ASAP7_75t_R _33802_ (.A1(_01598_),
    .A2(_01674_),
    .B(net3175),
    .Y(_04217_));
 AO21x1_ASAP7_75t_R _33803_ (.A1(net1597),
    .A2(_01500_),
    .B(net3175),
    .Y(_04218_));
 AND2x2_ASAP7_75t_R _33804_ (.A(_04217_),
    .B(_04218_),
    .Y(_04219_));
 INVx1_ASAP7_75t_R _33805_ (.A(_04219_),
    .Y(_04220_));
 OA211x2_ASAP7_75t_R _33806_ (.A1(_01498_),
    .A2(_01494_),
    .B(_01737_),
    .C(net3146),
    .Y(_04221_));
 OA21x2_ASAP7_75t_R _33807_ (.A1(_02461_),
    .A2(_01514_),
    .B(_01737_),
    .Y(_04222_));
 OR3x1_ASAP7_75t_R _33808_ (.A(_04220_),
    .B(_04221_),
    .C(_04222_),
    .Y(_04223_));
 NOR2x2_ASAP7_75t_R _33809_ (.A(_04216_),
    .B(_04223_),
    .Y(_04224_));
 AO21x1_ASAP7_75t_R _33810_ (.A1(net2366),
    .A2(net1613),
    .B(net2733),
    .Y(_04225_));
 AO21x1_ASAP7_75t_R _33811_ (.A1(_01598_),
    .A2(_01600_),
    .B(net2733),
    .Y(_04226_));
 AO21x1_ASAP7_75t_R _33812_ (.A1(net2075),
    .A2(_01569_),
    .B(net2733),
    .Y(_04227_));
 AND3x1_ASAP7_75t_R _33813_ (.A(_04225_),
    .B(_04226_),
    .C(_04227_),
    .Y(_04228_));
 AND3x1_ASAP7_75t_R _33814_ (.A(_02370_),
    .B(_02369_),
    .C(_03911_),
    .Y(_04229_));
 OA21x2_ASAP7_75t_R _33815_ (.A1(_01689_),
    .A2(_01668_),
    .B(_03245_),
    .Y(_04230_));
 NAND3x1_ASAP7_75t_R _33816_ (.A(_04228_),
    .B(_04229_),
    .C(_04230_),
    .Y(_04231_));
 AO21x1_ASAP7_75t_R _33817_ (.A1(net2572),
    .A2(net1613),
    .B(_01685_),
    .Y(_04232_));
 OAI21x1_ASAP7_75t_R _33818_ (.A1(_01685_),
    .A2(_01727_),
    .B(_04232_),
    .Y(_04233_));
 AO21x1_ASAP7_75t_R _33819_ (.A1(_01592_),
    .A2(_01500_),
    .B(_01701_),
    .Y(_04234_));
 AO21x1_ASAP7_75t_R _33820_ (.A1(_01689_),
    .A2(_02372_),
    .B(_01701_),
    .Y(_04235_));
 NAND2x1_ASAP7_75t_R _33821_ (.A(_04234_),
    .B(_04235_),
    .Y(_04236_));
 NAND2x1_ASAP7_75t_R _33822_ (.A(_02449_),
    .B(_01696_),
    .Y(_04237_));
 AO21x1_ASAP7_75t_R _33823_ (.A1(_01630_),
    .A2(net1457),
    .B(_01685_),
    .Y(_04238_));
 NAND2x1_ASAP7_75t_R _33824_ (.A(_04237_),
    .B(_04238_),
    .Y(_04239_));
 OA21x2_ASAP7_75t_R _33825_ (.A1(_02453_),
    .A2(_01514_),
    .B(_01696_),
    .Y(_04240_));
 OR4x1_ASAP7_75t_R _33826_ (.A(_04233_),
    .B(_04236_),
    .C(_04239_),
    .D(_04240_),
    .Y(_04241_));
 NOR2x1_ASAP7_75t_R _33827_ (.A(_04231_),
    .B(_04241_),
    .Y(_04242_));
 NAND2x2_ASAP7_75t_R _33828_ (.A(_04224_),
    .B(_04242_),
    .Y(_04243_));
 AO21x1_ASAP7_75t_R _33829_ (.A1(net2062),
    .A2(net2254),
    .B(_01624_),
    .Y(_04244_));
 NAND2x1_ASAP7_75t_R _33830_ (.A(_03206_),
    .B(_04244_),
    .Y(_04245_));
 NOR2x1_ASAP7_75t_R _33831_ (.A(_01569_),
    .B(_01624_),
    .Y(_04246_));
 AO21x1_ASAP7_75t_R _33832_ (.A1(net1605),
    .A2(net1597),
    .B(_01624_),
    .Y(_04247_));
 INVx1_ASAP7_75t_R _33833_ (.A(_04247_),
    .Y(_04248_));
 OR3x2_ASAP7_75t_R _33834_ (.A(_04245_),
    .B(_04246_),
    .C(_04248_),
    .Y(_04249_));
 AO21x1_ASAP7_75t_R _33835_ (.A1(net2524),
    .A2(_01540_),
    .B(net2334),
    .Y(_04250_));
 AO21x1_ASAP7_75t_R _33836_ (.A1(_01678_),
    .A2(net2379),
    .B(net2334),
    .Y(_04251_));
 AND2x2_ASAP7_75t_R _33837_ (.A(_04250_),
    .B(_04251_),
    .Y(_04252_));
 NAND3x2_ASAP7_75t_R _33838_ (.B(_01528_),
    .C(_02794_),
    .Y(_04253_),
    .A(_04252_));
 NAND2x2_ASAP7_75t_R _33839_ (.A(_01582_),
    .B(_01637_),
    .Y(_04254_));
 AO21x1_ASAP7_75t_R _33840_ (.A1(_01630_),
    .A2(_02363_),
    .B(net2746),
    .Y(_04255_));
 OA21x2_ASAP7_75t_R _33841_ (.A1(net1597),
    .A2(net2746),
    .B(_04255_),
    .Y(_04256_));
 NAND2x2_ASAP7_75t_R _33842_ (.A(_04254_),
    .B(_04256_),
    .Y(_04257_));
 NOR3x2_ASAP7_75t_R _33843_ (.B(_04253_),
    .C(_04257_),
    .Y(_04258_),
    .A(_04249_));
 AO21x1_ASAP7_75t_R _33844_ (.A1(_01689_),
    .A2(_01691_),
    .B(net2275),
    .Y(_04259_));
 OA21x2_ASAP7_75t_R _33845_ (.A1(net1612),
    .A2(net2275),
    .B(_04259_),
    .Y(_04260_));
 OA21x2_ASAP7_75t_R _33846_ (.A1(net1605),
    .A2(net2275),
    .B(_02442_),
    .Y(_04261_));
 NAND2x1_ASAP7_75t_R _33847_ (.A(_04260_),
    .B(_04261_),
    .Y(_04262_));
 NAND2x1_ASAP7_75t_R _33848_ (.A(_01680_),
    .B(_02829_),
    .Y(_04263_));
 AND2x2_ASAP7_75t_R _33849_ (.A(_01594_),
    .B(_04263_),
    .Y(_04264_));
 AO21x1_ASAP7_75t_R _33850_ (.A1(net2366),
    .A2(net2572),
    .B(net2348),
    .Y(_04265_));
 AOI211x1_ASAP7_75t_R _33851_ (.A1(_01498_),
    .A2(net1263),
    .B(net2348),
    .C(net1243),
    .Y(_04266_));
 INVx1_ASAP7_75t_R _33852_ (.A(_04266_),
    .Y(_04267_));
 NAND3x1_ASAP7_75t_R _33853_ (.A(_04264_),
    .B(_04265_),
    .C(_04267_),
    .Y(_04268_));
 NOR2x1_ASAP7_75t_R _33854_ (.A(_04262_),
    .B(_04268_),
    .Y(_04269_));
 AND3x1_ASAP7_75t_R _33855_ (.A(_03225_),
    .B(_03223_),
    .C(_01551_),
    .Y(_04270_));
 AO21x1_ASAP7_75t_R _33856_ (.A1(net2366),
    .A2(net1613),
    .B(_01571_),
    .Y(_04271_));
 AO21x1_ASAP7_75t_R _33857_ (.A1(_03894_),
    .A2(net1457),
    .B(_01571_),
    .Y(_04272_));
 AND2x2_ASAP7_75t_R _33858_ (.A(_04271_),
    .B(_04272_),
    .Y(_04273_));
 AND2x2_ASAP7_75t_R _33859_ (.A(_04270_),
    .B(_04273_),
    .Y(_04274_));
 AND2x2_ASAP7_75t_R _33860_ (.A(_04269_),
    .B(_04274_),
    .Y(_04275_));
 NAND2x2_ASAP7_75t_R _33861_ (.A(_04258_),
    .B(_04275_),
    .Y(_04276_));
 NOR2x1_ASAP7_75t_R _33862_ (.A(_04243_),
    .B(_04276_),
    .Y(_04277_));
 NAND2x2_ASAP7_75t_R _33863_ (.A(net3127),
    .B(_04277_),
    .Y(_04278_));
 OAI21x1_ASAP7_75t_R _33864_ (.A1(_04202_),
    .A2(_04206_),
    .B(_04278_),
    .Y(_04279_));
 NOR2x2_ASAP7_75t_R _33865_ (.A(_04203_),
    .B(_04201_),
    .Y(_04280_));
 NOR2x2_ASAP7_75t_R _33866_ (.A(_04126_),
    .B(_04205_),
    .Y(_04281_));
 NOR3x2_ASAP7_75t_R _33867_ (.B(_04243_),
    .C(_03885_),
    .Y(_04282_),
    .A(_04276_));
 OAI21x1_ASAP7_75t_R _33868_ (.A1(_04280_),
    .A2(_04281_),
    .B(_04282_),
    .Y(_04283_));
 AOI21x1_ASAP7_75t_R _33869_ (.A1(net953),
    .A2(_02535_),
    .B(_02536_),
    .Y(_04284_));
 AO21x1_ASAP7_75t_R _33870_ (.A1(_01908_),
    .A2(net2371),
    .B(net2384),
    .Y(_04285_));
 AND3x1_ASAP7_75t_R _33871_ (.A(_04284_),
    .B(_03632_),
    .C(_04285_),
    .Y(_04286_));
 AO21x1_ASAP7_75t_R _33872_ (.A1(_01824_),
    .A2(net1157),
    .B(net2194),
    .Y(_04287_));
 AO21x1_ASAP7_75t_R _33873_ (.A1(_01799_),
    .A2(net2286),
    .B(net2194),
    .Y(_04288_));
 NAND2x1_ASAP7_75t_R _33874_ (.A(_01940_),
    .B(_02176_),
    .Y(_04289_));
 NOR2x1_ASAP7_75t_R _33875_ (.A(net2194),
    .B(net3276),
    .Y(_04290_));
 INVx1_ASAP7_75t_R _33876_ (.A(_04290_),
    .Y(_04291_));
 AND4x1_ASAP7_75t_R _33877_ (.A(_04287_),
    .B(_04288_),
    .C(_04289_),
    .D(_04291_),
    .Y(_04292_));
 NAND2x2_ASAP7_75t_R _33878_ (.A(_04286_),
    .B(_04292_),
    .Y(_04293_));
 AO21x1_ASAP7_75t_R _33879_ (.A1(net1413),
    .A2(net1157),
    .B(_01905_),
    .Y(_04294_));
 OAI21x1_ASAP7_75t_R _33880_ (.A1(_01905_),
    .A2(_01946_),
    .B(_04294_),
    .Y(_04295_));
 NOR2x1_ASAP7_75t_R _33881_ (.A(_04295_),
    .B(_02205_),
    .Y(_04296_));
 AO21x1_ASAP7_75t_R _33882_ (.A1(_02500_),
    .A2(_01832_),
    .B(_01916_),
    .Y(_04297_));
 OA211x2_ASAP7_75t_R _33883_ (.A1(net2563),
    .A2(net2140),
    .B(_03975_),
    .C(_04297_),
    .Y(_04298_));
 NAND2x1_ASAP7_75t_R _33884_ (.A(_04296_),
    .B(_04298_),
    .Y(_04299_));
 NOR2x2_ASAP7_75t_R _33885_ (.A(_04293_),
    .B(_04299_),
    .Y(_04300_));
 AO21x1_ASAP7_75t_R _33886_ (.A1(net2307),
    .A2(net3275),
    .B(net2262),
    .Y(_04301_));
 INVx1_ASAP7_75t_R _33887_ (.A(_02229_),
    .Y(_04302_));
 AND4x1_ASAP7_75t_R _33888_ (.A(_04301_),
    .B(_04302_),
    .C(_02502_),
    .D(_02975_),
    .Y(_04303_));
 NAND2x1_ASAP7_75t_R _33889_ (.A(_02177_),
    .B(_03655_),
    .Y(_04304_));
 OA211x2_ASAP7_75t_R _33890_ (.A1(_01946_),
    .A2(net2352),
    .B(_02981_),
    .C(_04304_),
    .Y(_04305_));
 NAND2x1_ASAP7_75t_R _33891_ (.A(_04303_),
    .B(_04305_),
    .Y(_04306_));
 AO221x1_ASAP7_75t_R _33892_ (.A1(net1116),
    .A2(_01776_),
    .B1(_01870_),
    .B2(_01857_),
    .C(_01967_),
    .Y(_04307_));
 INVx1_ASAP7_75t_R _33893_ (.A(_02101_),
    .Y(_04308_));
 NOR2x1_ASAP7_75t_R _33894_ (.A(_02491_),
    .B(_04308_),
    .Y(_04309_));
 AND2x2_ASAP7_75t_R _33895_ (.A(_04307_),
    .B(_04309_),
    .Y(_04310_));
 NOR2x2_ASAP7_75t_R _33896_ (.A(net951),
    .B(_01870_),
    .Y(_04311_));
 AO21x1_ASAP7_75t_R _33897_ (.A1(_04311_),
    .A2(_01974_),
    .B(_02484_),
    .Y(_04312_));
 OA21x2_ASAP7_75t_R _33898_ (.A1(_01976_),
    .A2(_01806_),
    .B(_01974_),
    .Y(_04313_));
 AO21x1_ASAP7_75t_R _33899_ (.A1(_02114_),
    .A2(_01974_),
    .B(_02483_),
    .Y(_04314_));
 NOR3x1_ASAP7_75t_R _33900_ (.A(_04312_),
    .B(_04313_),
    .C(_04314_),
    .Y(_04315_));
 NAND2x1_ASAP7_75t_R _33901_ (.A(_04310_),
    .B(_04315_),
    .Y(_04316_));
 NOR2x1_ASAP7_75t_R _33902_ (.A(_04306_),
    .B(_04316_),
    .Y(_04317_));
 NAND2x2_ASAP7_75t_R _33903_ (.A(_04300_),
    .B(_04317_),
    .Y(_04318_));
 OA21x2_ASAP7_75t_R _33904_ (.A1(net1253),
    .A2(net2494),
    .B(_01868_),
    .Y(_04319_));
 AO21x1_ASAP7_75t_R _33905_ (.A1(net3254),
    .A2(_01785_),
    .B(_01851_),
    .Y(_04320_));
 AO21x1_ASAP7_75t_R _33906_ (.A1(net1138),
    .A2(net2619),
    .B(_01851_),
    .Y(_04321_));
 AND2x2_ASAP7_75t_R _33907_ (.A(_04320_),
    .B(_04321_),
    .Y(_04322_));
 AO31x2_ASAP7_75t_R _33908_ (.A1(net2175),
    .A2(net1157),
    .A3(_01934_),
    .B(net2494),
    .Y(_04323_));
 NAND3x2_ASAP7_75t_R _33909_ (.B(_04322_),
    .C(_04323_),
    .Y(_04324_),
    .A(_04319_));
 OA211x2_ASAP7_75t_R _33910_ (.A1(net1116),
    .A2(_01776_),
    .B(_01888_),
    .C(net1466),
    .Y(_04325_));
 INVx1_ASAP7_75t_R _33911_ (.A(_04325_),
    .Y(_04326_));
 AO21x1_ASAP7_75t_R _33912_ (.A1(_02110_),
    .A2(net3276),
    .B(net2459),
    .Y(_04327_));
 NAND2x1_ASAP7_75t_R _33913_ (.A(_01890_),
    .B(_01888_),
    .Y(_04328_));
 AND3x1_ASAP7_75t_R _33914_ (.A(_04327_),
    .B(_02913_),
    .C(_04328_),
    .Y(_04329_));
 NAND2x2_ASAP7_75t_R _33915_ (.A(_04326_),
    .B(_04329_),
    .Y(_04330_));
 AO31x2_ASAP7_75t_R _33916_ (.A1(net1253),
    .A2(net2395),
    .A3(_01908_),
    .B(_01878_),
    .Y(_04331_));
 AO21x1_ASAP7_75t_R _33917_ (.A1(net1317),
    .A2(net3277),
    .B(_01878_),
    .Y(_04332_));
 NAND2x1_ASAP7_75t_R _33918_ (.A(_01784_),
    .B(_01876_),
    .Y(_04333_));
 AND3x1_ASAP7_75t_R _33919_ (.A(_04332_),
    .B(_02907_),
    .C(_04333_),
    .Y(_04334_));
 NAND2x2_ASAP7_75t_R _33920_ (.A(_04331_),
    .B(_04334_),
    .Y(_04335_));
 NOR3x2_ASAP7_75t_R _33921_ (.B(_04330_),
    .C(_04335_),
    .Y(_04336_),
    .A(_04324_));
 AO21x1_ASAP7_75t_R _33922_ (.A1(_02110_),
    .A2(_01934_),
    .B(_01828_),
    .Y(_04337_));
 NAND2x1_ASAP7_75t_R _33923_ (.A(_04337_),
    .B(_01835_),
    .Y(_04338_));
 AO21x1_ASAP7_75t_R _33924_ (.A1(_01836_),
    .A2(_01837_),
    .B(_01809_),
    .Y(_04339_));
 AO21x1_ASAP7_75t_R _33925_ (.A1(_01821_),
    .A2(_01774_),
    .B(_01809_),
    .Y(_04340_));
 NAND2x1_ASAP7_75t_R _33926_ (.A(_04339_),
    .B(_04340_),
    .Y(_04341_));
 AOI211x1_ASAP7_75t_R _33927_ (.A1(_01806_),
    .A2(_01810_),
    .B(_04338_),
    .C(_04341_),
    .Y(_04342_));
 INVx1_ASAP7_75t_R _33928_ (.A(_04342_),
    .Y(_04343_));
 AO21x1_ASAP7_75t_R _33929_ (.A1(net2619),
    .A2(_01837_),
    .B(_01761_),
    .Y(_04344_));
 AO21x1_ASAP7_75t_R _33930_ (.A1(net1253),
    .A2(net2286),
    .B(_01761_),
    .Y(_04345_));
 NAND2x1_ASAP7_75t_R _33931_ (.A(_04344_),
    .B(_04345_),
    .Y(_04346_));
 AO21x1_ASAP7_75t_R _33932_ (.A1(_02110_),
    .A2(net3276),
    .B(_01761_),
    .Y(_04347_));
 OAI21x1_ASAP7_75t_R _33933_ (.A1(_01761_),
    .A2(_01946_),
    .B(_04347_),
    .Y(_04348_));
 AOI211x1_ASAP7_75t_R _33934_ (.A1(_01762_),
    .A2(net2330),
    .B(_04346_),
    .C(_04348_),
    .Y(_04349_));
 OA211x2_ASAP7_75t_R _33935_ (.A1(_01770_),
    .A2(net1452),
    .B(_02131_),
    .C(net1459),
    .Y(_04350_));
 AO21x1_ASAP7_75t_R _33936_ (.A1(_02918_),
    .A2(_02131_),
    .B(_02947_),
    .Y(_04351_));
 OA21x2_ASAP7_75t_R _33937_ (.A1(_02124_),
    .A2(_01886_),
    .B(_02131_),
    .Y(_04352_));
 NOR3x1_ASAP7_75t_R _33938_ (.A(_04350_),
    .B(_04351_),
    .C(_04352_),
    .Y(_04353_));
 NAND2x1_ASAP7_75t_R _33939_ (.A(_04349_),
    .B(_04353_),
    .Y(_04354_));
 NOR2x1_ASAP7_75t_R _33940_ (.A(_04343_),
    .B(_04354_),
    .Y(_04355_));
 NAND2x1_ASAP7_75t_R _33941_ (.A(_04336_),
    .B(_04355_),
    .Y(_04356_));
 NOR2x2_ASAP7_75t_R _33942_ (.A(_04318_),
    .B(_04356_),
    .Y(_04357_));
 NAND2x2_ASAP7_75t_R _33943_ (.A(_02247_),
    .B(_04357_),
    .Y(_04358_));
 INVx2_ASAP7_75t_R _33944_ (.A(_03881_),
    .Y(_04359_));
 XOR2x1_ASAP7_75t_R _33945_ (.A(net3139),
    .Y(_04360_),
    .B(_04359_));
 INVx1_ASAP7_75t_R _33946_ (.A(_04360_),
    .Y(_04361_));
 AOI21x1_ASAP7_75t_R _33947_ (.A1(_04279_),
    .A2(_04283_),
    .B(_04361_),
    .Y(_04362_));
 NOR2x2_ASAP7_75t_R _33948_ (.A(net3237),
    .B(_04282_),
    .Y(_04363_));
 NOR2x2_ASAP7_75t_R _33949_ (.A(_04205_),
    .B(_04278_),
    .Y(_04364_));
 OAI21x1_ASAP7_75t_R _33950_ (.A1(_04363_),
    .A2(_04364_),
    .B(_04126_),
    .Y(_04365_));
 NOR2x1_ASAP7_75t_R _33951_ (.A(_04205_),
    .B(_04282_),
    .Y(_04366_));
 NOR2x1_ASAP7_75t_R _33952_ (.A(net3237),
    .B(_04278_),
    .Y(_04367_));
 OAI21x1_ASAP7_75t_R _33953_ (.A1(_04366_),
    .A2(_04367_),
    .B(_04203_),
    .Y(_04368_));
 AOI21x1_ASAP7_75t_R _33954_ (.A1(_04365_),
    .A2(_04368_),
    .B(_04360_),
    .Y(_04369_));
 TAPCELL_ASAP7_75t_R PHY_538 ();
 OAI21x1_ASAP7_75t_R _33956_ (.A1(_04362_),
    .A2(_04369_),
    .B(net395),
    .Y(_04371_));
 INVx1_ASAP7_75t_R _33957_ (.A(_04371_),
    .Y(_04372_));
 OAI21x1_ASAP7_75t_R _33958_ (.A1(_04057_),
    .A2(_04372_),
    .B(_00478_),
    .Y(_04373_));
 INVx1_ASAP7_75t_R _33959_ (.A(_04057_),
    .Y(_04374_));
 NAND3x1_ASAP7_75t_R _33960_ (.A(_04371_),
    .B(_14358_),
    .C(_04374_),
    .Y(_04375_));
 NAND2x1_ASAP7_75t_R _33961_ (.A(_04375_),
    .B(_04373_),
    .Y(_00119_));
 AO21x1_ASAP7_75t_R _33962_ (.A1(net2266),
    .A2(_22019_),
    .B(_22061_),
    .Y(_04376_));
 AO21x1_ASAP7_75t_R _33963_ (.A1(net2420),
    .A2(_22008_),
    .B(_22061_),
    .Y(_04377_));
 NAND3x1_ASAP7_75t_R _33964_ (.A(_04376_),
    .B(_04377_),
    .C(_04192_),
    .Y(_04378_));
 AO21x1_ASAP7_75t_R _33965_ (.A1(_21890_),
    .A2(net2420),
    .B(_22064_),
    .Y(_04379_));
 NOR2x1_ASAP7_75t_R _33966_ (.A(_04196_),
    .B(_22055_),
    .Y(_04380_));
 NAND2x1_ASAP7_75t_R _33967_ (.A(_04379_),
    .B(_04380_),
    .Y(_04381_));
 NOR2x1_ASAP7_75t_R _33968_ (.A(_04378_),
    .B(_04381_),
    .Y(_04382_));
 NAND2x1_ASAP7_75t_R _33969_ (.A(_22084_),
    .B(_01085_),
    .Y(_04383_));
 NAND3x1_ASAP7_75t_R _33970_ (.A(_04184_),
    .B(_02721_),
    .C(_04383_),
    .Y(_04384_));
 OAI21x1_ASAP7_75t_R _33971_ (.A1(_22070_),
    .A2(_02261_),
    .B(_03154_),
    .Y(_04385_));
 AO21x1_ASAP7_75t_R _33972_ (.A1(_22024_),
    .A2(net2801),
    .B(_22070_),
    .Y(_04386_));
 AO21x1_ASAP7_75t_R _33973_ (.A1(net1629),
    .A2(net1833),
    .B(_22070_),
    .Y(_04387_));
 NAND2x1_ASAP7_75t_R _33974_ (.A(_04386_),
    .B(_04387_),
    .Y(_04388_));
 NOR3x1_ASAP7_75t_R _33975_ (.A(_04384_),
    .B(_04385_),
    .C(_04388_),
    .Y(_04389_));
 NAND2x1_ASAP7_75t_R _33976_ (.A(_04382_),
    .B(_04389_),
    .Y(_04390_));
 INVx1_ASAP7_75t_R _33977_ (.A(_02696_),
    .Y(_04391_));
 AOI211x1_ASAP7_75t_R _33978_ (.A1(_21887_),
    .A2(_21876_),
    .B(_22091_),
    .C(net1040),
    .Y(_04392_));
 NOR2x1_ASAP7_75t_R _33979_ (.A(_04391_),
    .B(_04392_),
    .Y(_04393_));
 NOR2x1_ASAP7_75t_R _33980_ (.A(_22091_),
    .B(net3236),
    .Y(_04394_));
 NOR2x1_ASAP7_75t_R _33981_ (.A(_04394_),
    .B(_03767_),
    .Y(_04395_));
 NAND2x1_ASAP7_75t_R _33982_ (.A(_04393_),
    .B(_04395_),
    .Y(_04396_));
 AO21x1_ASAP7_75t_R _33983_ (.A1(_22099_),
    .A2(_02261_),
    .B(_22100_),
    .Y(_04397_));
 AOI211x1_ASAP7_75t_R _33984_ (.A1(net1407),
    .A2(net1170),
    .B(net3080),
    .C(net1845),
    .Y(_04398_));
 OA21x2_ASAP7_75t_R _33985_ (.A1(_21953_),
    .A2(_21955_),
    .B(_02266_),
    .Y(_04399_));
 NOR2x1_ASAP7_75t_R _33986_ (.A(_04398_),
    .B(_04399_),
    .Y(_04400_));
 NAND2x1_ASAP7_75t_R _33987_ (.A(_04397_),
    .B(_04400_),
    .Y(_04401_));
 NOR2x1_ASAP7_75t_R _33988_ (.A(_04396_),
    .B(_04401_),
    .Y(_04402_));
 AO31x2_ASAP7_75t_R _33989_ (.A1(net2261),
    .A2(_21969_),
    .A3(_22019_),
    .B(_01072_),
    .Y(_04403_));
 NOR2x1_ASAP7_75t_R _33990_ (.A(_01072_),
    .B(_22076_),
    .Y(_04404_));
 AOI211x1_ASAP7_75t_R _33991_ (.A1(net1139),
    .A2(net1169),
    .B(_01072_),
    .C(net1846),
    .Y(_04405_));
 NOR2x1_ASAP7_75t_R _33992_ (.A(_04404_),
    .B(_04405_),
    .Y(_04406_));
 NAND2x1_ASAP7_75t_R _33993_ (.A(_04403_),
    .B(_04406_),
    .Y(_04407_));
 AOI211x1_ASAP7_75t_R _33994_ (.A1(_21887_),
    .A2(net1169),
    .B(_01078_),
    .C(_21895_),
    .Y(_04408_));
 INVx1_ASAP7_75t_R _33995_ (.A(_04408_),
    .Y(_04409_));
 AO21x1_ASAP7_75t_R _33996_ (.A1(_21929_),
    .A2(net1629),
    .B(_01078_),
    .Y(_04410_));
 NAND3x1_ASAP7_75t_R _33997_ (.A(_04409_),
    .B(_03164_),
    .C(_04410_),
    .Y(_04411_));
 NOR2x1_ASAP7_75t_R _33998_ (.A(_04407_),
    .B(_04411_),
    .Y(_04412_));
 NAND2x1_ASAP7_75t_R _33999_ (.A(_04402_),
    .B(_04412_),
    .Y(_04413_));
 NOR2x1_ASAP7_75t_R _34000_ (.A(_04413_),
    .B(_04390_),
    .Y(_04414_));
 AO21x1_ASAP7_75t_R _34001_ (.A1(net1834),
    .A2(net1045),
    .B(net2513),
    .Y(_04415_));
 AO21x1_ASAP7_75t_R _34002_ (.A1(net2365),
    .A2(_21969_),
    .B(net2513),
    .Y(_04416_));
 NAND2x1_ASAP7_75t_R _34003_ (.A(_04415_),
    .B(_04416_),
    .Y(_04417_));
 AOI21x1_ASAP7_75t_R _34004_ (.A1(net993),
    .A2(_02348_),
    .B(_03608_),
    .Y(_04418_));
 AOI211x1_ASAP7_75t_R _34005_ (.A1(_21887_),
    .A2(net1171),
    .B(net3156),
    .C(net1853),
    .Y(_04419_));
 OA21x2_ASAP7_75t_R _34006_ (.A1(net2038),
    .A2(_21909_),
    .B(_22034_),
    .Y(_04420_));
 NOR2x1_ASAP7_75t_R _34007_ (.A(_04419_),
    .B(_04420_),
    .Y(_04421_));
 NAND2x1_ASAP7_75t_R _34008_ (.A(_04418_),
    .B(_04421_),
    .Y(_04422_));
 NOR2x1_ASAP7_75t_R _34009_ (.A(_04417_),
    .B(_04422_),
    .Y(_04423_));
 AO21x1_ASAP7_75t_R _34010_ (.A1(net2267),
    .A2(net2337),
    .B(net3148),
    .Y(_04424_));
 AO21x1_ASAP7_75t_R _34011_ (.A1(_22024_),
    .A2(net1834),
    .B(net3148),
    .Y(_04425_));
 AO21x1_ASAP7_75t_R _34012_ (.A1(net2259),
    .A2(_02273_),
    .B(net3148),
    .Y(_04426_));
 NAND3x1_ASAP7_75t_R _34013_ (.A(_04424_),
    .B(_04425_),
    .C(_04426_),
    .Y(_04427_));
 AO31x2_ASAP7_75t_R _34014_ (.A1(net3172),
    .A2(_04150_),
    .A3(net1631),
    .B(_21992_),
    .Y(_04428_));
 AOI211x1_ASAP7_75t_R _34015_ (.A1(_21878_),
    .A2(_02758_),
    .B(_02759_),
    .C(_02760_),
    .Y(_04429_));
 NAND2x1_ASAP7_75t_R _34016_ (.A(_04428_),
    .B(_04429_),
    .Y(_04430_));
 NOR2x1_ASAP7_75t_R _34017_ (.A(_04427_),
    .B(_04430_),
    .Y(_04431_));
 NAND2x1_ASAP7_75t_R _34018_ (.A(_04423_),
    .B(_04431_),
    .Y(_04432_));
 AO21x1_ASAP7_75t_R _34019_ (.A1(_02312_),
    .A2(_04150_),
    .B(_21976_),
    .Y(_04433_));
 AO21x1_ASAP7_75t_R _34020_ (.A1(_21967_),
    .A2(net2420),
    .B(_21976_),
    .Y(_04434_));
 NAND2x1_ASAP7_75t_R _34021_ (.A(_02316_),
    .B(_21980_),
    .Y(_04435_));
 NAND3x1_ASAP7_75t_R _34022_ (.A(_04433_),
    .B(_04434_),
    .C(_04435_),
    .Y(_04436_));
 INVx1_ASAP7_75t_R _34023_ (.A(_21958_),
    .Y(_04437_));
 NOR2x1_ASAP7_75t_R _34024_ (.A(_04437_),
    .B(_04155_),
    .Y(_04438_));
 AND2x2_ASAP7_75t_R _34025_ (.A(_21972_),
    .B(_03101_),
    .Y(_04439_));
 NAND2x1_ASAP7_75t_R _34026_ (.A(_04438_),
    .B(_04439_),
    .Y(_04440_));
 NOR2x1_ASAP7_75t_R _34027_ (.A(_04436_),
    .B(_04440_),
    .Y(_04441_));
 AO21x1_ASAP7_75t_R _34028_ (.A1(net2297),
    .A2(net1834),
    .B(net2497),
    .Y(_04442_));
 AOI211x1_ASAP7_75t_R _34029_ (.A1(_21887_),
    .A2(_21876_),
    .B(_21895_),
    .C(net2497),
    .Y(_04443_));
 INVx1_ASAP7_75t_R _34030_ (.A(_04443_),
    .Y(_04444_));
 NAND2x1_ASAP7_75t_R _34031_ (.A(_04442_),
    .B(_04444_),
    .Y(_04445_));
 AOI211x1_ASAP7_75t_R _34032_ (.A1(_21887_),
    .A2(net1173),
    .B(_21901_),
    .C(_21895_),
    .Y(_04446_));
 NOR2x1_ASAP7_75t_R _34033_ (.A(_21915_),
    .B(_04446_),
    .Y(_04447_));
 AO31x2_ASAP7_75t_R _34034_ (.A1(_03097_),
    .A2(_21995_),
    .A3(_21929_),
    .B(_21901_),
    .Y(_04448_));
 NAND2x1_ASAP7_75t_R _34035_ (.A(_04447_),
    .B(_04448_),
    .Y(_04449_));
 NOR2x2_ASAP7_75t_R _34036_ (.A(_04445_),
    .B(_04449_),
    .Y(_04450_));
 NAND2x2_ASAP7_75t_R _34037_ (.A(_04441_),
    .B(_04450_),
    .Y(_04451_));
 NOR2x2_ASAP7_75t_R _34038_ (.A(_04432_),
    .B(_04451_),
    .Y(_04452_));
 NAND2x2_ASAP7_75t_R _34039_ (.A(_04414_),
    .B(_04452_),
    .Y(_04453_));
 XOR2x2_ASAP7_75t_R _34040_ (.A(_01480_),
    .B(_04453_),
    .Y(_04454_));
 AO21x1_ASAP7_75t_R _34041_ (.A1(_02110_),
    .A2(_02100_),
    .B(_01828_),
    .Y(_04455_));
 AO21x1_ASAP7_75t_R _34042_ (.A1(_01799_),
    .A2(_02134_),
    .B(_01828_),
    .Y(_04456_));
 AND2x2_ASAP7_75t_R _34043_ (.A(_04455_),
    .B(_04456_),
    .Y(_04457_));
 OA21x2_ASAP7_75t_R _34044_ (.A1(net2330),
    .A2(net3274),
    .B(_01810_),
    .Y(_04458_));
 NOR2x1_ASAP7_75t_R _34045_ (.A(_04458_),
    .B(_01812_),
    .Y(_04459_));
 OA21x2_ASAP7_75t_R _34046_ (.A1(net2654),
    .A2(_04311_),
    .B(_01810_),
    .Y(_04460_));
 OA21x2_ASAP7_75t_R _34047_ (.A1(_01855_),
    .A2(_01886_),
    .B(_01810_),
    .Y(_04461_));
 NOR2x1_ASAP7_75t_R _34048_ (.A(_04460_),
    .B(_04461_),
    .Y(_04462_));
 NAND3x1_ASAP7_75t_R _34049_ (.A(_04457_),
    .B(_04459_),
    .C(_04462_),
    .Y(_04463_));
 AO21x1_ASAP7_75t_R _34050_ (.A1(net1413),
    .A2(net1527),
    .B(_01781_),
    .Y(_04464_));
 AO21x1_ASAP7_75t_R _34051_ (.A1(_01785_),
    .A2(_01832_),
    .B(_01781_),
    .Y(_04465_));
 AO21x1_ASAP7_75t_R _34052_ (.A1(_01795_),
    .A2(_01870_),
    .B(_01781_),
    .Y(_04466_));
 AND3x1_ASAP7_75t_R _34053_ (.A(_04464_),
    .B(_04465_),
    .C(_04466_),
    .Y(_04467_));
 OAI21x1_ASAP7_75t_R _34054_ (.A1(net3272),
    .A2(_01976_),
    .B(_01762_),
    .Y(_04468_));
 AND3x1_ASAP7_75t_R _34055_ (.A(_04468_),
    .B(_02576_),
    .C(_04344_),
    .Y(_04469_));
 NAND2x1_ASAP7_75t_R _34056_ (.A(_04467_),
    .B(_04469_),
    .Y(_04470_));
 NOR2x1_ASAP7_75t_R _34057_ (.A(_04463_),
    .B(_04470_),
    .Y(_04471_));
 AO21x1_ASAP7_75t_R _34058_ (.A1(net2175),
    .A2(net1157),
    .B(_01878_),
    .Y(_04472_));
 AO21x1_ASAP7_75t_R _34059_ (.A1(net1253),
    .A2(_01799_),
    .B(_01878_),
    .Y(_04473_));
 NAND2x1_ASAP7_75t_R _34060_ (.A(_01858_),
    .B(_01876_),
    .Y(_04474_));
 AND3x1_ASAP7_75t_R _34061_ (.A(_04472_),
    .B(_04473_),
    .C(_04474_),
    .Y(_04475_));
 AO21x1_ASAP7_75t_R _34062_ (.A1(net2560),
    .A2(net1527),
    .B(net2459),
    .Y(_04476_));
 AO21x1_ASAP7_75t_R _34063_ (.A1(_02110_),
    .A2(_01832_),
    .B(net2459),
    .Y(_04477_));
 NAND2x1_ASAP7_75t_R _34064_ (.A(_04476_),
    .B(_04477_),
    .Y(_04478_));
 OA21x2_ASAP7_75t_R _34065_ (.A1(_02544_),
    .A2(_04311_),
    .B(_01888_),
    .Y(_04479_));
 AO21x1_ASAP7_75t_R _34066_ (.A1(_02114_),
    .A2(_01888_),
    .B(_04479_),
    .Y(_04480_));
 NOR2x1_ASAP7_75t_R _34067_ (.A(_04478_),
    .B(_04480_),
    .Y(_04481_));
 NAND2x1_ASAP7_75t_R _34068_ (.A(_04475_),
    .B(_04481_),
    .Y(_04482_));
 AO21x1_ASAP7_75t_R _34069_ (.A1(_01785_),
    .A2(_01934_),
    .B(_01851_),
    .Y(_04483_));
 INVx1_ASAP7_75t_R _34070_ (.A(_02920_),
    .Y(_04484_));
 AND3x1_ASAP7_75t_R _34071_ (.A(_04483_),
    .B(_03680_),
    .C(_04484_),
    .Y(_04485_));
 OA211x2_ASAP7_75t_R _34072_ (.A1(_01770_),
    .A2(_01776_),
    .B(_01864_),
    .C(net1559),
    .Y(_04486_));
 INVx1_ASAP7_75t_R _34073_ (.A(_04486_),
    .Y(_04487_));
 AO21x1_ASAP7_75t_R _34074_ (.A1(net2395),
    .A2(_01908_),
    .B(net2494),
    .Y(_04488_));
 NAND3x1_ASAP7_75t_R _34075_ (.A(_04485_),
    .B(_04487_),
    .C(_04488_),
    .Y(_04489_));
 NOR2x1_ASAP7_75t_R _34076_ (.A(_04482_),
    .B(_04489_),
    .Y(_04490_));
 NAND2x1_ASAP7_75t_R _34077_ (.A(_04471_),
    .B(_04490_),
    .Y(_04491_));
 OA21x2_ASAP7_75t_R _34078_ (.A1(_01816_),
    .A2(net2330),
    .B(_01904_),
    .Y(_04492_));
 OAI21x1_ASAP7_75t_R _34079_ (.A1(_04311_),
    .A2(_02544_),
    .B(_01904_),
    .Y(_04493_));
 NAND2x1_ASAP7_75t_R _34080_ (.A(_02517_),
    .B(_04493_),
    .Y(_04494_));
 NOR2x1_ASAP7_75t_R _34081_ (.A(_04492_),
    .B(_04494_),
    .Y(_04495_));
 AO21x1_ASAP7_75t_R _34082_ (.A1(net3134),
    .A2(_01770_),
    .B(_03623_),
    .Y(_04496_));
 AO21x1_ASAP7_75t_R _34083_ (.A1(_02191_),
    .A2(_01877_),
    .B(net2140),
    .Y(_04497_));
 NAND3x1_ASAP7_75t_R _34084_ (.A(_04495_),
    .B(_04496_),
    .C(_04497_),
    .Y(_04498_));
 AO21x1_ASAP7_75t_R _34085_ (.A1(_02110_),
    .A2(_01946_),
    .B(net2193),
    .Y(_04499_));
 NAND2x1_ASAP7_75t_R _34086_ (.A(_02918_),
    .B(_01940_),
    .Y(_04500_));
 AND3x1_ASAP7_75t_R _34087_ (.A(_04499_),
    .B(_01939_),
    .C(_04500_),
    .Y(_04501_));
 AO21x1_ASAP7_75t_R _34088_ (.A1(net2560),
    .A2(net1316),
    .B(net2549),
    .Y(_04502_));
 AO21x1_ASAP7_75t_R _34089_ (.A1(_01785_),
    .A2(_01832_),
    .B(net2549),
    .Y(_04503_));
 AND2x2_ASAP7_75t_R _34090_ (.A(_04502_),
    .B(_04503_),
    .Y(_04504_));
 AOI22x1_ASAP7_75t_R _34091_ (.A1(_02183_),
    .A2(net3259),
    .B1(_01930_),
    .B2(_01858_),
    .Y(_04505_));
 AND2x2_ASAP7_75t_R _34092_ (.A(_04504_),
    .B(_04505_),
    .Y(_04506_));
 NAND2x1_ASAP7_75t_R _34093_ (.A(_04501_),
    .B(_04506_),
    .Y(_04507_));
 NOR2x1_ASAP7_75t_R _34094_ (.A(_04498_),
    .B(_04507_),
    .Y(_04508_));
 AO21x1_ASAP7_75t_R _34095_ (.A1(_02129_),
    .A2(_01850_),
    .B(_01977_),
    .Y(_04509_));
 AO21x1_ASAP7_75t_R _34096_ (.A1(net2619),
    .A2(_01837_),
    .B(_01977_),
    .Y(_04510_));
 NAND2x1_ASAP7_75t_R _34097_ (.A(_01974_),
    .B(_01871_),
    .Y(_04511_));
 AND3x1_ASAP7_75t_R _34098_ (.A(_04509_),
    .B(_04510_),
    .C(_04511_),
    .Y(_04512_));
 AOI211x1_ASAP7_75t_R _34099_ (.A1(net2655),
    .A2(_01970_),
    .B(_02102_),
    .C(_02991_),
    .Y(_04513_));
 NAND2x1_ASAP7_75t_R _34100_ (.A(_04512_),
    .B(_04513_),
    .Y(_04514_));
 AO21x1_ASAP7_75t_R _34101_ (.A1(net2307),
    .A2(_01837_),
    .B(net2352),
    .Y(_04515_));
 INVx1_ASAP7_75t_R _34102_ (.A(_01957_),
    .Y(_04516_));
 AND3x1_ASAP7_75t_R _34103_ (.A(_04515_),
    .B(_04516_),
    .C(_04304_),
    .Y(_04517_));
 AO21x1_ASAP7_75t_R _34104_ (.A1(net1253),
    .A2(net1138),
    .B(net3125),
    .Y(_04518_));
 AO21x1_ASAP7_75t_R _34105_ (.A1(net2307),
    .A2(_01908_),
    .B(net2264),
    .Y(_04519_));
 AND4x1_ASAP7_75t_R _34106_ (.A(_04518_),
    .B(_01951_),
    .C(_04519_),
    .D(_03650_),
    .Y(_04520_));
 NAND2x1_ASAP7_75t_R _34107_ (.A(_04517_),
    .B(_04520_),
    .Y(_04521_));
 NOR2x1_ASAP7_75t_R _34108_ (.A(_04514_),
    .B(_04521_),
    .Y(_04522_));
 NAND2x2_ASAP7_75t_R _34109_ (.A(_04508_),
    .B(_04522_),
    .Y(_04523_));
 NOR2x2_ASAP7_75t_R _34110_ (.A(_04491_),
    .B(_04523_),
    .Y(_04524_));
 NAND2x2_ASAP7_75t_R _34111_ (.A(_02247_),
    .B(_04524_),
    .Y(_04525_));
 XOR2x2_ASAP7_75t_R _34112_ (.A(_04454_),
    .B(_04525_),
    .Y(_04526_));
 AO21x1_ASAP7_75t_R _34113_ (.A1(net1026),
    .A2(_02441_),
    .B(_03403_),
    .Y(_04527_));
 AO21x1_ASAP7_75t_R _34114_ (.A1(net1612),
    .A2(_01674_),
    .B(net2275),
    .Y(_04528_));
 OAI21x1_ASAP7_75t_R _34115_ (.A1(net2275),
    .A2(_01583_),
    .B(_04528_),
    .Y(_04529_));
 AO21x1_ASAP7_75t_R _34116_ (.A1(net1612),
    .A2(net1242),
    .B(net2348),
    .Y(_04530_));
 AO21x1_ASAP7_75t_R _34117_ (.A1(_01670_),
    .A2(_01540_),
    .B(net2348),
    .Y(_04531_));
 NAND2x2_ASAP7_75t_R _34118_ (.A(_04530_),
    .B(_04531_),
    .Y(_04532_));
 NOR3x2_ASAP7_75t_R _34119_ (.B(_04529_),
    .C(_04532_),
    .Y(_04533_),
    .A(_04527_));
 AO21x1_ASAP7_75t_R _34120_ (.A1(net1605),
    .A2(net1597),
    .B(_01571_),
    .Y(_04534_));
 AO21x1_ASAP7_75t_R _34121_ (.A1(_01699_),
    .A2(net1612),
    .B(_01571_),
    .Y(_04535_));
 AO21x1_ASAP7_75t_R _34122_ (.A1(net1457),
    .A2(net2538),
    .B(_01571_),
    .Y(_04536_));
 NAND3x1_ASAP7_75t_R _34123_ (.A(_04534_),
    .B(_04535_),
    .C(_04536_),
    .Y(_04537_));
 AO21x1_ASAP7_75t_R _34124_ (.A1(net2818),
    .A2(net2538),
    .B(net3264),
    .Y(_04538_));
 NAND2x1_ASAP7_75t_R _34125_ (.A(_01516_),
    .B(_01550_),
    .Y(_04539_));
 AND2x2_ASAP7_75t_R _34126_ (.A(_04538_),
    .B(_04539_),
    .Y(_04540_));
 AO21x1_ASAP7_75t_R _34127_ (.A1(_01699_),
    .A2(_01600_),
    .B(net3264),
    .Y(_04541_));
 AO21x1_ASAP7_75t_R _34128_ (.A1(net2368),
    .A2(net2062),
    .B(net3264),
    .Y(_04542_));
 NAND2x1_ASAP7_75t_R _34129_ (.A(_04541_),
    .B(_04542_),
    .Y(_04543_));
 INVx1_ASAP7_75t_R _34130_ (.A(_04543_),
    .Y(_04544_));
 NAND2x1_ASAP7_75t_R _34131_ (.A(_04540_),
    .B(_04544_),
    .Y(_04545_));
 NOR2x1_ASAP7_75t_R _34132_ (.A(_04537_),
    .B(_04545_),
    .Y(_04546_));
 NAND2x1_ASAP7_75t_R _34133_ (.A(_04533_),
    .B(_04546_),
    .Y(_04547_));
 AO21x1_ASAP7_75t_R _34134_ (.A1(_01629_),
    .A2(net1457),
    .B(_01624_),
    .Y(_04548_));
 NAND3x1_ASAP7_75t_R _34135_ (.A(_04548_),
    .B(_01622_),
    .C(_04244_),
    .Y(_04549_));
 NAND2x1_ASAP7_75t_R _34136_ (.A(_01511_),
    .B(_01637_),
    .Y(_04550_));
 AO21x1_ASAP7_75t_R _34137_ (.A1(_01630_),
    .A2(net2795),
    .B(_01636_),
    .Y(_04551_));
 NAND2x1_ASAP7_75t_R _34138_ (.A(_04550_),
    .B(_04551_),
    .Y(_04552_));
 NAND2x1_ASAP7_75t_R _34139_ (.A(_04254_),
    .B(_02409_),
    .Y(_04553_));
 NOR2x1_ASAP7_75t_R _34140_ (.A(_04552_),
    .B(_04553_),
    .Y(_04554_));
 INVx1_ASAP7_75t_R _34141_ (.A(_04554_),
    .Y(_04555_));
 NOR2x1_ASAP7_75t_R _34142_ (.A(_04549_),
    .B(_04555_),
    .Y(_04556_));
 NAND2x2_ASAP7_75t_R _34143_ (.A(_01719_),
    .B(_01657_),
    .Y(_04557_));
 NAND3x2_ASAP7_75t_R _34144_ (.B(_04557_),
    .C(_02421_),
    .Y(_04558_),
    .A(_03954_));
 AO21x1_ASAP7_75t_R _34145_ (.A1(_01569_),
    .A2(net1104),
    .B(_01505_),
    .Y(_04559_));
 AO21x1_ASAP7_75t_R _34146_ (.A1(net2572),
    .A2(net1612),
    .B(_01505_),
    .Y(_04560_));
 NAND2x2_ASAP7_75t_R _34147_ (.A(_04559_),
    .B(_04560_),
    .Y(_04561_));
 AO21x1_ASAP7_75t_R _34148_ (.A1(_01569_),
    .A2(_02363_),
    .B(net2334),
    .Y(_04562_));
 OAI21x1_ASAP7_75t_R _34149_ (.A1(net2079),
    .A2(net2336),
    .B(_04562_),
    .Y(_04563_));
 NOR3x2_ASAP7_75t_R _34150_ (.B(_04561_),
    .C(_04563_),
    .Y(_04564_),
    .A(_04558_));
 NAND2x2_ASAP7_75t_R _34151_ (.A(_04556_),
    .B(_04564_),
    .Y(_04565_));
 NOR2x2_ASAP7_75t_R _34152_ (.A(_04547_),
    .B(_04565_),
    .Y(_04566_));
 NOR2x1_ASAP7_75t_R _34153_ (.A(_01668_),
    .B(_01689_),
    .Y(_04567_));
 AOI221x1_ASAP7_75t_R _34154_ (.A1(_01498_),
    .A2(_01494_),
    .B1(net2074),
    .B2(_01644_),
    .C(_01668_),
    .Y(_04568_));
 NOR2x1_ASAP7_75t_R _34155_ (.A(_04567_),
    .B(_04568_),
    .Y(_04569_));
 AO21x1_ASAP7_75t_R _34156_ (.A1(_02419_),
    .A2(net2728),
    .B(_01675_),
    .Y(_04570_));
 NAND2x1_ASAP7_75t_R _34157_ (.A(_01575_),
    .B(_01681_),
    .Y(_04571_));
 AND3x1_ASAP7_75t_R _34158_ (.A(_01677_),
    .B(_04570_),
    .C(_04571_),
    .Y(_04572_));
 NAND2x1_ASAP7_75t_R _34159_ (.A(_04569_),
    .B(_04572_),
    .Y(_04573_));
 AO21x1_ASAP7_75t_R _34160_ (.A1(_01630_),
    .A2(_02363_),
    .B(_01701_),
    .Y(_04574_));
 NAND2x1_ASAP7_75t_R _34161_ (.A(_04574_),
    .B(_03242_),
    .Y(_04575_));
 AO21x1_ASAP7_75t_R _34162_ (.A1(net2062),
    .A2(net2254),
    .B(_01701_),
    .Y(_04576_));
 AO21x1_ASAP7_75t_R _34163_ (.A1(_01699_),
    .A2(_01600_),
    .B(_01701_),
    .Y(_04577_));
 NAND2x1_ASAP7_75t_R _34164_ (.A(_04576_),
    .B(_04577_),
    .Y(_04578_));
 NOR2x1_ASAP7_75t_R _34165_ (.A(_04575_),
    .B(_04578_),
    .Y(_04579_));
 AO21x1_ASAP7_75t_R _34166_ (.A1(_01727_),
    .A2(net2367),
    .B(_01685_),
    .Y(_04580_));
 AO21x1_ASAP7_75t_R _34167_ (.A1(net3135),
    .A2(_01641_),
    .B(_01685_),
    .Y(_04581_));
 AND2x2_ASAP7_75t_R _34168_ (.A(_04580_),
    .B(_04581_),
    .Y(_04582_));
 NAND2x1_ASAP7_75t_R _34169_ (.A(_04579_),
    .B(_04582_),
    .Y(_04583_));
 NOR2x2_ASAP7_75t_R _34170_ (.A(_04573_),
    .B(_04583_),
    .Y(_04584_));
 INVx1_ASAP7_75t_R _34171_ (.A(_04584_),
    .Y(_04585_));
 NOR2x1_ASAP7_75t_R _34172_ (.A(_02391_),
    .B(_01731_),
    .Y(_04586_));
 AOI211x1_ASAP7_75t_R _34173_ (.A1(net1120),
    .A2(net1895),
    .B(_01728_),
    .C(net2377),
    .Y(_04587_));
 OA21x2_ASAP7_75t_R _34174_ (.A1(_01719_),
    .A2(_01575_),
    .B(_02388_),
    .Y(_04588_));
 NOR2x1_ASAP7_75t_R _34175_ (.A(_04587_),
    .B(_04588_),
    .Y(_04589_));
 NAND2x1_ASAP7_75t_R _34176_ (.A(_04586_),
    .B(_04589_),
    .Y(_04590_));
 AOI211x1_ASAP7_75t_R _34177_ (.A1(_01498_),
    .A2(_01494_),
    .B(_01735_),
    .C(net1238),
    .Y(_04591_));
 AOI21x1_ASAP7_75t_R _34178_ (.A1(_03196_),
    .A2(net2524),
    .B(_01735_),
    .Y(_04592_));
 OR3x1_ASAP7_75t_R _34179_ (.A(_04591_),
    .B(_02868_),
    .C(_04592_),
    .Y(_04593_));
 NOR2x2_ASAP7_75t_R _34180_ (.A(_04590_),
    .B(_04593_),
    .Y(_04594_));
 AOI211x1_ASAP7_75t_R _34181_ (.A1(net1120),
    .A2(net1263),
    .B(_01715_),
    .C(_01644_),
    .Y(_04595_));
 NOR2x1_ASAP7_75t_R _34182_ (.A(_04595_),
    .B(_03271_),
    .Y(_04596_));
 AOI211x1_ASAP7_75t_R _34183_ (.A1(net1120),
    .A2(net1896),
    .B(_01715_),
    .C(net2379),
    .Y(_04597_));
 AOI21x1_ASAP7_75t_R _34184_ (.A1(_01720_),
    .A2(net2406),
    .B(_04597_),
    .Y(_04598_));
 NAND2x1_ASAP7_75t_R _34185_ (.A(_04596_),
    .B(_04598_),
    .Y(_04599_));
 OA21x2_ASAP7_75t_R _34186_ (.A1(_01635_),
    .A2(_01719_),
    .B(_01711_),
    .Y(_04600_));
 OA21x2_ASAP7_75t_R _34187_ (.A1(_02449_),
    .A2(_02798_),
    .B(_01711_),
    .Y(_04601_));
 OR3x1_ASAP7_75t_R _34188_ (.A(_04600_),
    .B(_04601_),
    .C(_03260_),
    .Y(_04602_));
 NOR2x2_ASAP7_75t_R _34189_ (.A(_04599_),
    .B(_04602_),
    .Y(_04603_));
 NAND2x1_ASAP7_75t_R _34190_ (.A(_04594_),
    .B(_04603_),
    .Y(_04604_));
 NOR2x1_ASAP7_75t_R _34191_ (.A(_04585_),
    .B(_04604_),
    .Y(_04605_));
 NAND2x2_ASAP7_75t_R _34192_ (.A(_04566_),
    .B(_04605_),
    .Y(_04606_));
 XOR2x1_ASAP7_75t_R _34193_ (.A(_04126_),
    .Y(_04607_),
    .B(_04606_));
 XOR2x1_ASAP7_75t_R _34194_ (.A(_04526_),
    .Y(_04608_),
    .B(_04607_));
 AND2x2_ASAP7_75t_R _34195_ (.A(_18753_),
    .B(_00876_),
    .Y(_04609_));
 AO21x1_ASAP7_75t_R _34196_ (.A1(_04608_),
    .A2(net395),
    .B(_04609_),
    .Y(_04610_));
 XOR2x1_ASAP7_75t_R _34197_ (.A(_04610_),
    .Y(_00120_),
    .B(_00477_));
 AND2x2_ASAP7_75t_R _34198_ (.A(_18753_),
    .B(_00875_),
    .Y(_04611_));
 NOR2x2_ASAP7_75t_R _34199_ (.A(_01371_),
    .B(_01360_),
    .Y(_04612_));
 INVx2_ASAP7_75t_R _34200_ (.A(_04612_),
    .Y(_04613_));
 NAND2x1_ASAP7_75t_R _34201_ (.A(_04613_),
    .B(_01991_),
    .Y(_04614_));
 NAND2x1_ASAP7_75t_R _34202_ (.A(_04612_),
    .B(_01094_),
    .Y(_04615_));
 INVx1_ASAP7_75t_R _34203_ (.A(_04566_),
    .Y(_04616_));
 NAND3x2_ASAP7_75t_R _34204_ (.B(_04594_),
    .C(_04603_),
    .Y(_04617_),
    .A(_04584_));
 NOR2x2_ASAP7_75t_R _34205_ (.A(_04616_),
    .B(_04617_),
    .Y(_04618_));
 AO21x2_ASAP7_75t_R _34206_ (.A1(_04614_),
    .A2(_04615_),
    .B(_04618_),
    .Y(_04619_));
 XOR2x1_ASAP7_75t_R _34207_ (.A(_01094_),
    .Y(_04620_),
    .B(_04612_));
 NAND2x2_ASAP7_75t_R _34208_ (.A(_04620_),
    .B(_04618_),
    .Y(_04621_));
 NAND3x1_ASAP7_75t_R _34209_ (.A(_04619_),
    .B(_04621_),
    .C(_02249_),
    .Y(_04622_));
 AO21x1_ASAP7_75t_R _34210_ (.A1(_04619_),
    .A2(_04621_),
    .B(_02249_),
    .Y(_04623_));
 AOI21x1_ASAP7_75t_R _34211_ (.A1(_04622_),
    .A2(_04623_),
    .B(_18753_),
    .Y(_04624_));
 OAI21x1_ASAP7_75t_R _34212_ (.A1(_04611_),
    .A2(_04624_),
    .B(_14601_),
    .Y(_04625_));
 TAPCELL_ASAP7_75t_R PHY_537 ();
 NOR2x1_ASAP7_75t_R _34214_ (.A(net395),
    .B(_00875_),
    .Y(_04627_));
 INVx1_ASAP7_75t_R _34215_ (.A(_02249_),
    .Y(_04628_));
 NAND3x1_ASAP7_75t_R _34216_ (.A(_04619_),
    .B(_04621_),
    .C(_04628_),
    .Y(_04629_));
 AO21x1_ASAP7_75t_R _34217_ (.A1(_04619_),
    .A2(_04621_),
    .B(_04628_),
    .Y(_04630_));
 AOI21x1_ASAP7_75t_R _34218_ (.A1(_04629_),
    .A2(_04630_),
    .B(_18753_),
    .Y(_04631_));
 OAI21x1_ASAP7_75t_R _34219_ (.A1(_04627_),
    .A2(_04631_),
    .B(_00476_),
    .Y(_04632_));
 NAND2x2_ASAP7_75t_R _34220_ (.A(_04632_),
    .B(_04625_),
    .Y(_00081_));
 OAI21x1_ASAP7_75t_R _34221_ (.A1(_01371_),
    .A2(_02090_),
    .B(_02357_),
    .Y(_04633_));
 INVx2_ASAP7_75t_R _34222_ (.A(_02357_),
    .Y(_04634_));
 NAND2x2_ASAP7_75t_R _34223_ (.A(_04634_),
    .B(_02091_),
    .Y(_04635_));
 NAND2x2_ASAP7_75t_R _34224_ (.A(_04633_),
    .B(_04635_),
    .Y(_04636_));
 XOR2x2_ASAP7_75t_R _34225_ (.A(_01754_),
    .B(_04618_),
    .Y(_04637_));
 XOR2x1_ASAP7_75t_R _34226_ (.A(_04636_),
    .Y(_04638_),
    .B(_04637_));
 XOR2x1_ASAP7_75t_R _34227_ (.A(_02249_),
    .Y(_04639_),
    .B(_02589_));
 INVx1_ASAP7_75t_R _34228_ (.A(_04639_),
    .Y(_04640_));
 NAND2x1_ASAP7_75t_R _34229_ (.A(_04638_),
    .B(_04640_),
    .Y(_04641_));
 INVx1_ASAP7_75t_R _34230_ (.A(_01753_),
    .Y(_04642_));
 OAI21x1_ASAP7_75t_R _34231_ (.A1(_03885_),
    .A2(_04642_),
    .B(_04618_),
    .Y(_04643_));
 NAND3x2_ASAP7_75t_R _34232_ (.B(_04606_),
    .C(net3126),
    .Y(_04644_),
    .A(_01753_));
 NAND2x2_ASAP7_75t_R _34233_ (.A(_04643_),
    .B(_04644_),
    .Y(_04645_));
 XOR2x1_ASAP7_75t_R _34234_ (.A(_04636_),
    .Y(_04646_),
    .B(_04645_));
 AOI21x1_ASAP7_75t_R _34235_ (.A1(_04639_),
    .A2(_04646_),
    .B(_18753_),
    .Y(_04647_));
 AND2x2_ASAP7_75t_R _34236_ (.A(_18753_),
    .B(_00874_),
    .Y(_04648_));
 AOI21x1_ASAP7_75t_R _34237_ (.A1(_04641_),
    .A2(_04647_),
    .B(_04648_),
    .Y(_04649_));
 XNOR2x1_ASAP7_75t_R _34238_ (.B(_04649_),
    .Y(_00082_),
    .A(_00475_));
 AND2x2_ASAP7_75t_R _34239_ (.A(_18753_),
    .B(_00873_),
    .Y(_04650_));
 INVx1_ASAP7_75t_R _34240_ (.A(_02719_),
    .Y(_04651_));
 NAND2x1_ASAP7_75t_R _34241_ (.A(_02744_),
    .B(_02730_),
    .Y(_04652_));
 NOR2x2_ASAP7_75t_R _34242_ (.A(_04651_),
    .B(_04652_),
    .Y(_04653_));
 INVx1_ASAP7_75t_R _34243_ (.A(_02764_),
    .Y(_04654_));
 NOR2x2_ASAP7_75t_R _34244_ (.A(_02783_),
    .B(_04654_),
    .Y(_04655_));
 NAND2x2_ASAP7_75t_R _34245_ (.A(_04653_),
    .B(_04655_),
    .Y(_04656_));
 NOR2x2_ASAP7_75t_R _34246_ (.A(_04656_),
    .B(net2523),
    .Y(_04657_));
 AOI21x1_ASAP7_75t_R _34247_ (.A1(_02645_),
    .A2(_02691_),
    .B(_02786_),
    .Y(_04658_));
 OAI21x1_ASAP7_75t_R _34248_ (.A1(_04657_),
    .A2(_04658_),
    .B(_03004_),
    .Y(_04659_));
 NOR2x2_ASAP7_75t_R _34249_ (.A(_02786_),
    .B(net2523),
    .Y(_04660_));
 AND2x2_ASAP7_75t_R _34250_ (.A(_02692_),
    .B(_02786_),
    .Y(_04661_));
 OAI21x1_ASAP7_75t_R _34251_ (.A1(_04660_),
    .A2(_04661_),
    .B(net2672),
    .Y(_04662_));
 XOR2x2_ASAP7_75t_R _34252_ (.A(_02588_),
    .B(net2574),
    .Y(_04663_));
 AOI21x1_ASAP7_75t_R _34253_ (.A1(_04659_),
    .A2(_04662_),
    .B(_04663_),
    .Y(_04664_));
 XNOR2x2_ASAP7_75t_R _34254_ (.A(net2574),
    .B(_02588_),
    .Y(_04665_));
 NAND2x1_ASAP7_75t_R _34255_ (.A(_04659_),
    .B(_04662_),
    .Y(_04666_));
 NOR2x1_ASAP7_75t_R _34256_ (.A(_04665_),
    .B(_04666_),
    .Y(_04667_));
 OAI21x1_ASAP7_75t_R _34257_ (.A1(_04664_),
    .A2(_04667_),
    .B(net396),
    .Y(_04668_));
 INVx1_ASAP7_75t_R _34258_ (.A(_04668_),
    .Y(_04669_));
 INVx1_ASAP7_75t_R _34259_ (.A(_00474_),
    .Y(_04670_));
 OAI21x1_ASAP7_75t_R _34260_ (.A1(_04650_),
    .A2(_04669_),
    .B(_04670_),
    .Y(_04671_));
 INVx1_ASAP7_75t_R _34261_ (.A(_04650_),
    .Y(_04672_));
 NAND3x1_ASAP7_75t_R _34262_ (.A(_04668_),
    .B(_00474_),
    .C(_04672_),
    .Y(_04673_));
 NAND2x1_ASAP7_75t_R _34263_ (.A(_04673_),
    .B(_04671_),
    .Y(_00083_));
 NOR2x1_ASAP7_75t_R _34264_ (.A(net396),
    .B(_00872_),
    .Y(_04674_));
 XOR2x2_ASAP7_75t_R _34265_ (.A(_03090_),
    .B(_03710_),
    .Y(_04675_));
 XOR2x2_ASAP7_75t_R _34266_ (.A(_02888_),
    .B(_04606_),
    .Y(_04676_));
 XNOR2x1_ASAP7_75t_R _34267_ (.B(_04676_),
    .Y(_04677_),
    .A(_04675_));
 INVx2_ASAP7_75t_R _34268_ (.A(_03193_),
    .Y(_04678_));
 AOI21x1_ASAP7_75t_R _34269_ (.A1(_03003_),
    .A2(_03005_),
    .B(_04678_),
    .Y(_04679_));
 AOI21x1_ASAP7_75t_R _34270_ (.A1(_03093_),
    .A2(_03094_),
    .B(net2700),
    .Y(_04680_));
 NOR2x1_ASAP7_75t_R _34271_ (.A(_04679_),
    .B(_04680_),
    .Y(_04681_));
 NAND2x1_ASAP7_75t_R _34272_ (.A(_04677_),
    .B(_04681_),
    .Y(_04682_));
 XOR2x2_ASAP7_75t_R _34273_ (.A(_04676_),
    .B(_04675_),
    .Y(_04683_));
 OAI21x1_ASAP7_75t_R _34274_ (.A1(_04679_),
    .A2(_04680_),
    .B(net3270),
    .Y(_04684_));
 AOI21x1_ASAP7_75t_R _34275_ (.A1(_04682_),
    .A2(_04684_),
    .B(_18753_),
    .Y(_04685_));
 OAI21x1_ASAP7_75t_R _34276_ (.A1(_04674_),
    .A2(_04685_),
    .B(_00473_),
    .Y(_04686_));
 AND2x2_ASAP7_75t_R _34277_ (.A(_18753_),
    .B(_00872_),
    .Y(_04687_));
 XOR2x2_ASAP7_75t_R _34278_ (.A(_03193_),
    .B(_03090_),
    .Y(_04688_));
 INVx3_ASAP7_75t_R _34279_ (.A(_03710_),
    .Y(_04689_));
 XOR2x1_ASAP7_75t_R _34280_ (.A(_04688_),
    .Y(_04690_),
    .B(_04689_));
 XOR2x1_ASAP7_75t_R _34281_ (.A(_03380_),
    .Y(_04691_),
    .B(_04676_));
 NAND2x1_ASAP7_75t_R _34282_ (.A(_04690_),
    .B(_04691_),
    .Y(_04692_));
 XOR2x1_ASAP7_75t_R _34283_ (.A(_04688_),
    .Y(_04693_),
    .B(_03710_));
 XNOR2x1_ASAP7_75t_R _34284_ (.B(_03380_),
    .Y(_04694_),
    .A(_04676_));
 NAND2x1_ASAP7_75t_R _34285_ (.A(_04693_),
    .B(_04694_),
    .Y(_04695_));
 AOI21x1_ASAP7_75t_R _34286_ (.A1(_04692_),
    .A2(_04695_),
    .B(_18753_),
    .Y(_04696_));
 INVx1_ASAP7_75t_R _34287_ (.A(_00473_),
    .Y(_04697_));
 OAI21x1_ASAP7_75t_R _34288_ (.A1(_04687_),
    .A2(_04696_),
    .B(_04697_),
    .Y(_04698_));
 NAND2x1_ASAP7_75t_R _34289_ (.A(_04698_),
    .B(_04686_),
    .Y(_00084_));
 AND2x2_ASAP7_75t_R _34290_ (.A(_18753_),
    .B(_00871_),
    .Y(_04699_));
 XOR2x1_ASAP7_75t_R _34291_ (.A(net2646),
    .Y(_04700_),
    .B(_04041_));
 XOR2x2_ASAP7_75t_R _34292_ (.A(_03291_),
    .B(_04606_),
    .Y(_04701_));
 XOR2x1_ASAP7_75t_R _34293_ (.A(_04701_),
    .Y(_04702_),
    .B(net2827));
 NAND2x1_ASAP7_75t_R _34294_ (.A(_04700_),
    .B(_04702_),
    .Y(_04703_));
 NOR2x1_ASAP7_75t_R _34295_ (.A(_03711_),
    .B(_04701_),
    .Y(_04704_));
 AND2x2_ASAP7_75t_R _34296_ (.A(_04701_),
    .B(_03711_),
    .Y(_04705_));
 INVx3_ASAP7_75t_R _34297_ (.A(_04041_),
    .Y(_04706_));
 XOR2x1_ASAP7_75t_R _34298_ (.A(_03618_),
    .Y(_04707_),
    .B(_04706_));
 OAI21x1_ASAP7_75t_R _34299_ (.A1(_04704_),
    .A2(_04705_),
    .B(_04707_),
    .Y(_04708_));
 AOI21x1_ASAP7_75t_R _34300_ (.A1(_04703_),
    .A2(_04708_),
    .B(net388),
    .Y(_04709_));
 INVx1_ASAP7_75t_R _34301_ (.A(_00472_),
    .Y(_04710_));
 OAI21x1_ASAP7_75t_R _34302_ (.A1(_04699_),
    .A2(_04709_),
    .B(_04710_),
    .Y(_04711_));
 NOR2x1_ASAP7_75t_R _34303_ (.A(net396),
    .B(_00871_),
    .Y(_04712_));
 XOR2x1_ASAP7_75t_R _34304_ (.A(_04701_),
    .Y(_04713_),
    .B(_04041_));
 NAND2x1_ASAP7_75t_R _34305_ (.A(_04713_),
    .B(_03716_),
    .Y(_04714_));
 XOR2x1_ASAP7_75t_R _34306_ (.A(_04701_),
    .Y(_04715_),
    .B(_04706_));
 NAND2x1_ASAP7_75t_R _34307_ (.A(_03712_),
    .B(_04715_),
    .Y(_04716_));
 AOI21x1_ASAP7_75t_R _34308_ (.A1(_04714_),
    .A2(_04716_),
    .B(_18753_),
    .Y(_04717_));
 OAI21x1_ASAP7_75t_R _34309_ (.A1(_04712_),
    .A2(_04717_),
    .B(_00472_),
    .Y(_04718_));
 NAND2x1_ASAP7_75t_R _34310_ (.A(_04718_),
    .B(_04711_),
    .Y(_00085_));
 INVx1_ASAP7_75t_R _34311_ (.A(net3139),
    .Y(_04719_));
 AOI21x1_ASAP7_75t_R _34312_ (.A1(_04047_),
    .A2(_04048_),
    .B(_04719_),
    .Y(_04720_));
 AOI21x1_ASAP7_75t_R _34313_ (.A1(_03883_),
    .A2(_04045_),
    .B(net3140),
    .Y(_04721_));
 XOR2x2_ASAP7_75t_R _34314_ (.A(_04041_),
    .B(_03466_),
    .Y(_04722_));
 NOR3x1_ASAP7_75t_R _34315_ (.A(_04720_),
    .B(_04721_),
    .C(_04722_),
    .Y(_04723_));
 OAI21x1_ASAP7_75t_R _34316_ (.A1(_04721_),
    .A2(_04720_),
    .B(_04722_),
    .Y(_04724_));
 NAND2x1_ASAP7_75t_R _34317_ (.A(_04724_),
    .B(net395),
    .Y(_04725_));
 OR2x2_ASAP7_75t_R _34318_ (.A(net395),
    .B(_00870_),
    .Y(_04726_));
 OAI21x1_ASAP7_75t_R _34319_ (.A1(_04723_),
    .A2(_04725_),
    .B(_04726_),
    .Y(_04727_));
 XNOR2x1_ASAP7_75t_R _34320_ (.B(_04727_),
    .Y(_00086_),
    .A(_00471_));
 OAI21x1_ASAP7_75t_R _34321_ (.A1(_04202_),
    .A2(_04206_),
    .B(_04525_),
    .Y(_04728_));
 INVx2_ASAP7_75t_R _34322_ (.A(_04525_),
    .Y(_04729_));
 OAI21x1_ASAP7_75t_R _34323_ (.A1(_04280_),
    .A2(_04281_),
    .B(_04729_),
    .Y(_04730_));
 XOR2x1_ASAP7_75t_R _34324_ (.A(net3139),
    .Y(_04731_),
    .B(_03960_));
 INVx1_ASAP7_75t_R _34325_ (.A(_04731_),
    .Y(_04732_));
 AOI21x1_ASAP7_75t_R _34326_ (.A1(_04728_),
    .A2(_04730_),
    .B(_04732_),
    .Y(_04733_));
 OAI21x1_ASAP7_75t_R _34327_ (.A1(_04202_),
    .A2(_04206_),
    .B(_04729_),
    .Y(_04734_));
 OAI21x1_ASAP7_75t_R _34328_ (.A1(_04280_),
    .A2(_04281_),
    .B(_04525_),
    .Y(_04735_));
 AOI21x1_ASAP7_75t_R _34329_ (.A1(_04734_),
    .A2(_04735_),
    .B(_04731_),
    .Y(_04736_));
 OAI21x1_ASAP7_75t_R _34330_ (.A1(_04733_),
    .A2(_04736_),
    .B(net395),
    .Y(_04737_));
 INVx1_ASAP7_75t_R _34331_ (.A(_00470_),
    .Y(_04738_));
 NOR2x1_ASAP7_75t_R _34332_ (.A(net392),
    .B(_00869_),
    .Y(_04739_));
 INVx1_ASAP7_75t_R _34333_ (.A(_04739_),
    .Y(_04740_));
 NAND3x1_ASAP7_75t_R _34334_ (.A(_04737_),
    .B(_04738_),
    .C(_04740_),
    .Y(_04741_));
 AO21x1_ASAP7_75t_R _34335_ (.A1(_04737_),
    .A2(_04740_),
    .B(_04738_),
    .Y(_04742_));
 NAND2x1_ASAP7_75t_R _34336_ (.A(_04741_),
    .B(_04742_),
    .Y(_00087_));
 XOR2x2_ASAP7_75t_R _34337_ (.A(_04282_),
    .B(net2710),
    .Y(_04743_));
 XOR2x1_ASAP7_75t_R _34338_ (.A(_04526_),
    .Y(_04744_),
    .B(_04743_));
 AND2x2_ASAP7_75t_R _34339_ (.A(net389),
    .B(_00868_),
    .Y(_04745_));
 AO21x1_ASAP7_75t_R _34340_ (.A1(_04744_),
    .A2(net395),
    .B(_04745_),
    .Y(_04746_));
 XOR2x1_ASAP7_75t_R _34341_ (.A(_04746_),
    .Y(_00088_),
    .B(_00469_));
 INVx8_ASAP7_75t_R _34342_ (.A(_04453_),
    .Y(_04747_));
 TAPCELL_ASAP7_75t_R PHY_536 ();
 NOR2x1_ASAP7_75t_R _34344_ (.A(_04747_),
    .B(_04612_),
    .Y(_04749_));
 NOR2x1_ASAP7_75t_R _34345_ (.A(_04453_),
    .B(_04613_),
    .Y(_04750_));
 NOR2x2_ASAP7_75t_R _34346_ (.A(_02107_),
    .B(_02239_),
    .Y(_04751_));
 OAI21x1_ASAP7_75t_R _34347_ (.A1(_04749_),
    .A2(_04750_),
    .B(_04751_),
    .Y(_04752_));
 NAND2x2_ASAP7_75t_R _34348_ (.A(_02247_),
    .B(_02245_),
    .Y(_04753_));
 NOR2x1_ASAP7_75t_R _34349_ (.A(_04749_),
    .B(_04750_),
    .Y(_04754_));
 NAND2x1_ASAP7_75t_R _34350_ (.A(_04754_),
    .B(_04753_),
    .Y(_04755_));
 AOI21x1_ASAP7_75t_R _34351_ (.A1(_04752_),
    .A2(_04755_),
    .B(_04637_),
    .Y(_04756_));
 NAND2x1_ASAP7_75t_R _34352_ (.A(_04612_),
    .B(_04751_),
    .Y(_04757_));
 NAND2x1_ASAP7_75t_R _34353_ (.A(_04613_),
    .B(_04753_),
    .Y(_04758_));
 NAND3x1_ASAP7_75t_R _34354_ (.A(_04757_),
    .B(_04758_),
    .C(net3269),
    .Y(_04759_));
 AO21x1_ASAP7_75t_R _34355_ (.A1(_04757_),
    .A2(_04758_),
    .B(net3269),
    .Y(_04760_));
 AOI21x1_ASAP7_75t_R _34356_ (.A1(_04759_),
    .A2(_04760_),
    .B(_04645_),
    .Y(_04761_));
 OAI21x1_ASAP7_75t_R _34357_ (.A1(_04756_),
    .A2(_04761_),
    .B(net396),
    .Y(_04762_));
 NOR2x1_ASAP7_75t_R _34358_ (.A(net396),
    .B(_00867_),
    .Y(_04763_));
 INVx1_ASAP7_75t_R _34359_ (.A(_04763_),
    .Y(_04764_));
 NAND3x1_ASAP7_75t_R _34360_ (.A(_04762_),
    .B(_15661_),
    .C(_04764_),
    .Y(_04765_));
 AO21x1_ASAP7_75t_R _34361_ (.A1(_04762_),
    .A2(_04764_),
    .B(_15661_),
    .Y(_04766_));
 NAND2x1_ASAP7_75t_R _34362_ (.A(_04765_),
    .B(_04766_),
    .Y(_00049_));
 AND2x2_ASAP7_75t_R _34363_ (.A(_18753_),
    .B(_00866_),
    .Y(_04767_));
 NAND2x2_ASAP7_75t_R _34364_ (.A(_04645_),
    .B(_04665_),
    .Y(_04768_));
 INVx1_ASAP7_75t_R _34365_ (.A(_04768_),
    .Y(_04769_));
 NAND2x2_ASAP7_75t_R _34366_ (.A(_04663_),
    .B(_04637_),
    .Y(_04770_));
 INVx1_ASAP7_75t_R _34367_ (.A(_04770_),
    .Y(_04771_));
 INVx1_ASAP7_75t_R _34368_ (.A(_01093_),
    .Y(_04772_));
 OAI21x1_ASAP7_75t_R _34369_ (.A1(_03734_),
    .A2(_04772_),
    .B(_04747_),
    .Y(_04773_));
 NAND3x2_ASAP7_75t_R _34370_ (.B(net2031),
    .C(net2789),
    .Y(_04774_),
    .A(_01093_));
 AOI21x1_ASAP7_75t_R _34371_ (.A1(_04773_),
    .A2(_04774_),
    .B(net2042),
    .Y(_04775_));
 NAND3x2_ASAP7_75t_R _34372_ (.B(_01093_),
    .C(net2789),
    .Y(_04776_),
    .A(net3269));
 AO21x1_ASAP7_75t_R _34373_ (.A1(_01093_),
    .A2(net2790),
    .B(_04747_),
    .Y(_04777_));
 AOI21x1_ASAP7_75t_R _34374_ (.A1(_04776_),
    .A2(_04777_),
    .B(_02092_),
    .Y(_04778_));
 NOR2x2_ASAP7_75t_R _34375_ (.A(_04775_),
    .B(_04778_),
    .Y(_04779_));
 OAI21x1_ASAP7_75t_R _34376_ (.A1(_04769_),
    .A2(_04771_),
    .B(_04779_),
    .Y(_04780_));
 AOI21x1_ASAP7_75t_R _34377_ (.A1(_04773_),
    .A2(_04774_),
    .B(_02092_),
    .Y(_04781_));
 AOI21x1_ASAP7_75t_R _34378_ (.A1(_04776_),
    .A2(_04777_),
    .B(net2042),
    .Y(_04782_));
 NOR2x1_ASAP7_75t_R _34379_ (.A(_04781_),
    .B(_04782_),
    .Y(_04783_));
 NAND3x1_ASAP7_75t_R _34380_ (.A(_04783_),
    .B(_04770_),
    .C(_04768_),
    .Y(_04784_));
 TAPCELL_ASAP7_75t_R PHY_535 ();
 AOI21x1_ASAP7_75t_R _34382_ (.A1(_04780_),
    .A2(_04784_),
    .B(_18753_),
    .Y(_04786_));
 OAI21x1_ASAP7_75t_R _34383_ (.A1(_04767_),
    .A2(_04786_),
    .B(_15784_),
    .Y(_04787_));
 NOR2x1_ASAP7_75t_R _34384_ (.A(net396),
    .B(_00866_),
    .Y(_04788_));
 NAND3x1_ASAP7_75t_R _34385_ (.A(_04779_),
    .B(_04770_),
    .C(_04768_),
    .Y(_04789_));
 AO21x1_ASAP7_75t_R _34386_ (.A1(_04768_),
    .A2(_04770_),
    .B(_04779_),
    .Y(_04790_));
 AOI21x1_ASAP7_75t_R _34387_ (.A1(_04789_),
    .A2(_04790_),
    .B(_18753_),
    .Y(_04791_));
 OAI21x1_ASAP7_75t_R _34388_ (.A1(_04788_),
    .A2(_04791_),
    .B(_00467_),
    .Y(_04792_));
 NAND2x2_ASAP7_75t_R _34389_ (.A(_04792_),
    .B(_04787_),
    .Y(_00050_));
 NOR2x1_ASAP7_75t_R _34390_ (.A(net396),
    .B(_00865_),
    .Y(_04793_));
 NOR2x2_ASAP7_75t_R _34391_ (.A(_02888_),
    .B(net2523),
    .Y(_04794_));
 AOI22x1_ASAP7_75t_R _34392_ (.A1(_02691_),
    .A2(_02645_),
    .B1(_02887_),
    .B2(_02837_),
    .Y(_04795_));
 OA21x2_ASAP7_75t_R _34393_ (.A1(_04794_),
    .A2(_04795_),
    .B(net2674),
    .Y(_04796_));
 NOR3x1_ASAP7_75t_R _34394_ (.A(_04794_),
    .B(_04795_),
    .C(net2674),
    .Y(_04797_));
 OAI21x1_ASAP7_75t_R _34395_ (.A1(_04796_),
    .A2(_04797_),
    .B(_02472_),
    .Y(_04798_));
 XOR2x1_ASAP7_75t_R _34396_ (.A(net2672),
    .Y(_04799_),
    .B(_02692_));
 NOR2x1_ASAP7_75t_R _34397_ (.A(_02888_),
    .B(_04799_),
    .Y(_04800_));
 XNOR2x1_ASAP7_75t_R _34398_ (.B(net2672),
    .Y(_04801_),
    .A(net2523));
 NOR2x1_ASAP7_75t_R _34399_ (.A(_02896_),
    .B(_04801_),
    .Y(_04802_));
 OAI21x1_ASAP7_75t_R _34400_ (.A1(_04800_),
    .A2(_04802_),
    .B(_02468_),
    .Y(_04803_));
 AOI21x1_ASAP7_75t_R _34401_ (.A1(_04798_),
    .A2(_04803_),
    .B(_18753_),
    .Y(_04804_));
 NOR2x2_ASAP7_75t_R _34402_ (.A(_04793_),
    .B(_04804_),
    .Y(_04805_));
 XOR2x1_ASAP7_75t_R _34403_ (.A(_04805_),
    .Y(_00051_),
    .B(_00466_));
 NAND2x1_ASAP7_75t_R _34404_ (.A(_00864_),
    .B(net388),
    .Y(_04806_));
 NOR2x1_ASAP7_75t_R _34405_ (.A(_04675_),
    .B(_04676_),
    .Y(_04807_));
 AND2x2_ASAP7_75t_R _34406_ (.A(_04676_),
    .B(_04675_),
    .Y(_04808_));
 NOR2x2_ASAP7_75t_R _34407_ (.A(_04453_),
    .B(_04656_),
    .Y(_04809_));
 NOR2x2_ASAP7_75t_R _34408_ (.A(_04747_),
    .B(_02786_),
    .Y(_04810_));
 OAI21x1_ASAP7_75t_R _34409_ (.A1(_04809_),
    .A2(_04810_),
    .B(_03291_),
    .Y(_04811_));
 NOR2x1_ASAP7_75t_R _34410_ (.A(_04747_),
    .B(_04656_),
    .Y(_04812_));
 AO21x1_ASAP7_75t_R _34411_ (.A1(_04653_),
    .A2(_04655_),
    .B(_04453_),
    .Y(_04813_));
 INVx1_ASAP7_75t_R _34412_ (.A(_04813_),
    .Y(_04814_));
 INVx2_ASAP7_75t_R _34413_ (.A(_03291_),
    .Y(_04815_));
 OAI21x1_ASAP7_75t_R _34414_ (.A1(_04812_),
    .A2(_04814_),
    .B(_04815_),
    .Y(_04816_));
 NAND2x1_ASAP7_75t_R _34415_ (.A(_04816_),
    .B(_04811_),
    .Y(_04817_));
 OAI21x1_ASAP7_75t_R _34416_ (.A1(_04807_),
    .A2(_04808_),
    .B(_04817_),
    .Y(_04818_));
 INVx1_ASAP7_75t_R _34417_ (.A(_04818_),
    .Y(_04819_));
 INVx1_ASAP7_75t_R _34418_ (.A(_04817_),
    .Y(_04820_));
 NAND2x2_ASAP7_75t_R _34419_ (.A(_04683_),
    .B(_04820_),
    .Y(_04821_));
 INVx1_ASAP7_75t_R _34420_ (.A(_04821_),
    .Y(_04822_));
 OAI21x1_ASAP7_75t_R _34421_ (.A1(_04819_),
    .A2(_04822_),
    .B(net396),
    .Y(_04823_));
 INVx2_ASAP7_75t_R _34422_ (.A(_00465_),
    .Y(_04824_));
 AOI21x1_ASAP7_75t_R _34423_ (.A1(_04806_),
    .A2(_04823_),
    .B(_04824_),
    .Y(_04825_));
 OR2x2_ASAP7_75t_R _34424_ (.A(net396),
    .B(_00864_),
    .Y(_04826_));
 NAND3x1_ASAP7_75t_R _34425_ (.A(_04821_),
    .B(_04818_),
    .C(net396),
    .Y(_04827_));
 AOI21x1_ASAP7_75t_R _34426_ (.A1(_04826_),
    .A2(_04827_),
    .B(_00465_),
    .Y(_04828_));
 NOR2x1_ASAP7_75t_R _34427_ (.A(_04825_),
    .B(_04828_),
    .Y(_00052_));
 AND2x2_ASAP7_75t_R _34428_ (.A(net388),
    .B(_00863_),
    .Y(_04829_));
 XOR2x2_ASAP7_75t_R _34429_ (.A(_03193_),
    .B(_04747_),
    .Y(_04830_));
 INVx3_ASAP7_75t_R _34430_ (.A(_03539_),
    .Y(_04831_));
 XOR2x1_ASAP7_75t_R _34431_ (.A(_04830_),
    .Y(_04832_),
    .B(_04831_));
 INVx1_ASAP7_75t_R _34432_ (.A(_03450_),
    .Y(_04833_));
 NOR2x1_ASAP7_75t_R _34433_ (.A(_03463_),
    .B(_04833_),
    .Y(_04834_));
 INVx1_ASAP7_75t_R _34434_ (.A(_03434_),
    .Y(_04835_));
 NAND2x2_ASAP7_75t_R _34435_ (.A(_04834_),
    .B(_04835_),
    .Y(_04836_));
 XOR2x2_ASAP7_75t_R _34436_ (.A(_04041_),
    .B(_04836_),
    .Y(_04837_));
 XOR2x1_ASAP7_75t_R _34437_ (.A(_04837_),
    .Y(_04838_),
    .B(_04701_));
 NAND2x1_ASAP7_75t_R _34438_ (.A(_04832_),
    .B(_04838_),
    .Y(_04839_));
 XOR2x1_ASAP7_75t_R _34439_ (.A(_04830_),
    .Y(_04840_),
    .B(_03539_));
 XOR2x1_ASAP7_75t_R _34440_ (.A(_04722_),
    .Y(_04841_),
    .B(_04701_));
 NAND2x1_ASAP7_75t_R _34441_ (.A(_04840_),
    .B(_04841_),
    .Y(_04842_));
 AOI21x1_ASAP7_75t_R _34442_ (.A1(_04839_),
    .A2(_04842_),
    .B(net388),
    .Y(_04843_));
 INVx1_ASAP7_75t_R _34443_ (.A(_00464_),
    .Y(_04844_));
 OAI21x1_ASAP7_75t_R _34444_ (.A1(_04829_),
    .A2(_04843_),
    .B(_04844_),
    .Y(_04845_));
 NOR2x1_ASAP7_75t_R _34445_ (.A(net396),
    .B(_00863_),
    .Y(_04846_));
 XOR2x2_ASAP7_75t_R _34446_ (.A(_03193_),
    .B(net2031),
    .Y(_04847_));
 NOR2x2_ASAP7_75t_R _34447_ (.A(_04847_),
    .B(_04837_),
    .Y(_04848_));
 NOR2x1_ASAP7_75t_R _34448_ (.A(_04722_),
    .B(_04830_),
    .Y(_04849_));
 AOI21x1_ASAP7_75t_R _34449_ (.A1(_03290_),
    .A2(_03234_),
    .B(_04618_),
    .Y(_04850_));
 NOR2x1_ASAP7_75t_R _34450_ (.A(net3260),
    .B(net3176),
    .Y(_04851_));
 OAI21x1_ASAP7_75t_R _34451_ (.A1(_04850_),
    .A2(_04851_),
    .B(_03539_),
    .Y(_04852_));
 NOR2x1_ASAP7_75t_R _34452_ (.A(_04618_),
    .B(net3176),
    .Y(_04853_));
 NOR2x1_ASAP7_75t_R _34453_ (.A(net3260),
    .B(_04815_),
    .Y(_04854_));
 OAI21x1_ASAP7_75t_R _34454_ (.A1(_04853_),
    .A2(_04854_),
    .B(_04831_),
    .Y(_04855_));
 NAND2x1_ASAP7_75t_R _34455_ (.A(_04852_),
    .B(_04855_),
    .Y(_04856_));
 OAI21x1_ASAP7_75t_R _34456_ (.A1(_04848_),
    .A2(_04849_),
    .B(_04856_),
    .Y(_04857_));
 XOR2x1_ASAP7_75t_R _34457_ (.A(_04701_),
    .Y(_04858_),
    .B(_04831_));
 NOR2x1_ASAP7_75t_R _34458_ (.A(_04848_),
    .B(_04849_),
    .Y(_04859_));
 NAND2x1_ASAP7_75t_R _34459_ (.A(_04859_),
    .B(_04858_),
    .Y(_04860_));
 AOI21x1_ASAP7_75t_R _34460_ (.A1(_04857_),
    .A2(_04860_),
    .B(net388),
    .Y(_04861_));
 OAI21x1_ASAP7_75t_R _34461_ (.A1(_04846_),
    .A2(_04861_),
    .B(_00464_),
    .Y(_04862_));
 NAND2x1_ASAP7_75t_R _34462_ (.A(_04862_),
    .B(_04845_),
    .Y(_00053_));
 NOR2x1_ASAP7_75t_R _34463_ (.A(net394),
    .B(_00862_),
    .Y(_04863_));
 NAND2x2_ASAP7_75t_R _34464_ (.A(_03466_),
    .B(_03617_),
    .Y(_04864_));
 OAI22x1_ASAP7_75t_R _34465_ (.A1(_03465_),
    .A2(_03434_),
    .B1(_03616_),
    .B2(_03576_),
    .Y(_04865_));
 AO21x1_ASAP7_75t_R _34466_ (.A1(_04864_),
    .A2(_04865_),
    .B(_04358_),
    .Y(_04866_));
 NAND3x2_ASAP7_75t_R _34467_ (.B(_04864_),
    .C(_04865_),
    .Y(_04867_),
    .A(net3139));
 XOR2x2_ASAP7_75t_R _34468_ (.A(_03881_),
    .B(_03960_),
    .Y(_04868_));
 AOI21x1_ASAP7_75t_R _34469_ (.A1(_04866_),
    .A2(_04867_),
    .B(_04868_),
    .Y(_04869_));
 INVx2_ASAP7_75t_R _34470_ (.A(_04868_),
    .Y(_04870_));
 NAND2x1_ASAP7_75t_R _34471_ (.A(_04866_),
    .B(_04867_),
    .Y(_04871_));
 NOR2x1_ASAP7_75t_R _34472_ (.A(_04871_),
    .B(_04870_),
    .Y(_04872_));
 OAI21x1_ASAP7_75t_R _34473_ (.A1(_04869_),
    .A2(_04872_),
    .B(net396),
    .Y(_04873_));
 INVx1_ASAP7_75t_R _34474_ (.A(_04873_),
    .Y(_04874_));
 OAI21x1_ASAP7_75t_R _34475_ (.A1(_04863_),
    .A2(_04874_),
    .B(_00463_),
    .Y(_04875_));
 INVx1_ASAP7_75t_R _34476_ (.A(_04863_),
    .Y(_04876_));
 NAND3x1_ASAP7_75t_R _34477_ (.A(_04873_),
    .B(_16060_),
    .C(_04876_),
    .Y(_04877_));
 NAND2x1_ASAP7_75t_R _34478_ (.A(_04875_),
    .B(_04877_),
    .Y(_00054_));
 NAND2x1_ASAP7_75t_R _34479_ (.A(_03809_),
    .B(_04126_),
    .Y(_04878_));
 NAND2x1_ASAP7_75t_R _34480_ (.A(_03970_),
    .B(_04203_),
    .Y(_04879_));
 AOI21x1_ASAP7_75t_R _34481_ (.A1(_04878_),
    .A2(_04879_),
    .B(_04729_),
    .Y(_04880_));
 NAND2x1_ASAP7_75t_R _34482_ (.A(_03970_),
    .B(_04126_),
    .Y(_04881_));
 NAND2x1_ASAP7_75t_R _34483_ (.A(_03809_),
    .B(_04203_),
    .Y(_04882_));
 AOI21x1_ASAP7_75t_R _34484_ (.A1(_04881_),
    .A2(_04882_),
    .B(net3340),
    .Y(_04883_));
 XOR2x2_ASAP7_75t_R _34485_ (.A(_04282_),
    .B(_03960_),
    .Y(_04884_));
 NOR3x1_ASAP7_75t_R _34486_ (.A(_04880_),
    .B(_04883_),
    .C(_04884_),
    .Y(_04885_));
 OAI21x1_ASAP7_75t_R _34487_ (.A1(_04880_),
    .A2(_04883_),
    .B(_04884_),
    .Y(_04886_));
 NAND2x1_ASAP7_75t_R _34488_ (.A(_04886_),
    .B(net396),
    .Y(_04887_));
 OR2x2_ASAP7_75t_R _34489_ (.A(net396),
    .B(_00861_),
    .Y(_04888_));
 OAI21x1_ASAP7_75t_R _34490_ (.A1(_04885_),
    .A2(_04887_),
    .B(_04888_),
    .Y(_04889_));
 XOR2x1_ASAP7_75t_R _34491_ (.A(_04889_),
    .Y(_00055_),
    .B(_16130_));
 NOR2x2_ASAP7_75t_R _34492_ (.A(net2392),
    .B(net3237),
    .Y(_04890_));
 NOR2x1_ASAP7_75t_R _34493_ (.A(_03376_),
    .B(_04205_),
    .Y(_04891_));
 OAI21x1_ASAP7_75t_R _34494_ (.A1(_04890_),
    .A2(_04891_),
    .B(net3260),
    .Y(_04892_));
 NOR2x2_ASAP7_75t_R _34495_ (.A(_03376_),
    .B(_04201_),
    .Y(_04893_));
 NOR2x1_ASAP7_75t_R _34496_ (.A(net2392),
    .B(_04205_),
    .Y(_04894_));
 OAI21x1_ASAP7_75t_R _34497_ (.A1(_04893_),
    .A2(_04894_),
    .B(_04618_),
    .Y(_04895_));
 AOI21x1_ASAP7_75t_R _34498_ (.A1(_04892_),
    .A2(_04895_),
    .B(_04743_),
    .Y(_04896_));
 OAI21x1_ASAP7_75t_R _34499_ (.A1(_04890_),
    .A2(_04891_),
    .B(_04618_),
    .Y(_04897_));
 OAI21x1_ASAP7_75t_R _34500_ (.A1(_04893_),
    .A2(_04894_),
    .B(net3260),
    .Y(_04898_));
 INVx1_ASAP7_75t_R _34501_ (.A(_04743_),
    .Y(_04899_));
 AOI21x1_ASAP7_75t_R _34502_ (.A1(_04897_),
    .A2(_04898_),
    .B(_04899_),
    .Y(_04900_));
 OAI21x1_ASAP7_75t_R _34503_ (.A1(_04896_),
    .A2(_04900_),
    .B(net395),
    .Y(_04901_));
 INVx2_ASAP7_75t_R _34504_ (.A(_00461_),
    .Y(_04902_));
 NOR2x1_ASAP7_75t_R _34505_ (.A(net394),
    .B(_00860_),
    .Y(_04903_));
 INVx1_ASAP7_75t_R _34506_ (.A(_04903_),
    .Y(_04904_));
 NAND3x1_ASAP7_75t_R _34507_ (.A(_04901_),
    .B(_04902_),
    .C(_04904_),
    .Y(_04905_));
 AO21x1_ASAP7_75t_R _34508_ (.A1(_04901_),
    .A2(_04904_),
    .B(_04902_),
    .Y(_04906_));
 NAND2x1_ASAP7_75t_R _34509_ (.A(_04906_),
    .B(_04905_),
    .Y(_00056_));
 XOR2x1_ASAP7_75t_R _34510_ (.A(_04454_),
    .Y(_04907_),
    .B(_04751_));
 XNOR2x1_ASAP7_75t_R _34511_ (.B(_01754_),
    .Y(_04908_),
    .A(_01094_));
 XOR2x1_ASAP7_75t_R _34512_ (.A(_04907_),
    .Y(_04909_),
    .B(_04908_));
 NOR2x1_ASAP7_75t_R _34513_ (.A(net395),
    .B(_00859_),
    .Y(_04910_));
 AO21x1_ASAP7_75t_R _34514_ (.A1(_04909_),
    .A2(net395),
    .B(_04910_),
    .Y(_04911_));
 XNOR2x1_ASAP7_75t_R _34515_ (.B(_04911_),
    .Y(_00017_),
    .A(_00460_));
 NOR2x1_ASAP7_75t_R _34516_ (.A(net395),
    .B(_00858_),
    .Y(_04912_));
 OAI21x1_ASAP7_75t_R _34517_ (.A1(_01481_),
    .A2(_01482_),
    .B(_02588_),
    .Y(_04913_));
 NOR2x1_ASAP7_75t_R _34518_ (.A(net2392),
    .B(_04612_),
    .Y(_04914_));
 NOR3x1_ASAP7_75t_R _34519_ (.A(_03376_),
    .B(_01360_),
    .C(_01371_),
    .Y(_04915_));
 OAI21x1_ASAP7_75t_R _34520_ (.A1(_04914_),
    .A2(_04915_),
    .B(_02589_),
    .Y(_04916_));
 NAND2x2_ASAP7_75t_R _34521_ (.A(_04913_),
    .B(_04916_),
    .Y(_04917_));
 INVx1_ASAP7_75t_R _34522_ (.A(_04917_),
    .Y(_04918_));
 NAND2x2_ASAP7_75t_R _34523_ (.A(_04774_),
    .B(_04773_),
    .Y(_04919_));
 XOR2x1_ASAP7_75t_R _34524_ (.A(_02472_),
    .Y(_04920_),
    .B(_04919_));
 NAND2x1_ASAP7_75t_R _34525_ (.A(_04918_),
    .B(_04920_),
    .Y(_04921_));
 INVx1_ASAP7_75t_R _34526_ (.A(_04919_),
    .Y(_04922_));
 NAND2x1_ASAP7_75t_R _34527_ (.A(_02472_),
    .B(_04922_),
    .Y(_04923_));
 NAND2x2_ASAP7_75t_R _34528_ (.A(_04919_),
    .B(_02468_),
    .Y(_04924_));
 NAND3x1_ASAP7_75t_R _34529_ (.A(net3314),
    .B(_04923_),
    .C(_04924_),
    .Y(_04925_));
 AOI21x1_ASAP7_75t_R _34530_ (.A1(_04921_),
    .A2(_04925_),
    .B(_18753_),
    .Y(_04926_));
 OAI21x1_ASAP7_75t_R _34531_ (.A1(_04912_),
    .A2(_04926_),
    .B(_00459_),
    .Y(_04927_));
 AOI21x1_ASAP7_75t_R _34532_ (.A1(_04924_),
    .A2(_04923_),
    .B(net3314),
    .Y(_04928_));
 NOR2x1_ASAP7_75t_R _34533_ (.A(_04918_),
    .B(_04920_),
    .Y(_04929_));
 OAI21x1_ASAP7_75t_R _34534_ (.A1(_04928_),
    .A2(_04929_),
    .B(net395),
    .Y(_04930_));
 INVx1_ASAP7_75t_R _34535_ (.A(_00459_),
    .Y(_04931_));
 INVx1_ASAP7_75t_R _34536_ (.A(_04912_),
    .Y(_04932_));
 NAND3x1_ASAP7_75t_R _34537_ (.A(_04930_),
    .B(_04931_),
    .C(_04932_),
    .Y(_04933_));
 NAND2x1_ASAP7_75t_R _34538_ (.A(_04933_),
    .B(_04927_),
    .Y(_00018_));
 AND2x2_ASAP7_75t_R _34539_ (.A(_18753_),
    .B(_00857_),
    .Y(_04934_));
 AOI21x1_ASAP7_75t_R _34540_ (.A1(_04633_),
    .A2(_04635_),
    .B(net2673),
    .Y(_04935_));
 INVx1_ASAP7_75t_R _34541_ (.A(_04935_),
    .Y(_04936_));
 NAND3x1_ASAP7_75t_R _34542_ (.A(_04635_),
    .B(_04633_),
    .C(net2673),
    .Y(_04937_));
 XOR2x1_ASAP7_75t_R _34543_ (.A(_02888_),
    .Y(_04938_),
    .B(_02786_));
 INVx1_ASAP7_75t_R _34544_ (.A(_04938_),
    .Y(_04939_));
 AOI21x1_ASAP7_75t_R _34545_ (.A1(_04936_),
    .A2(_04937_),
    .B(_04939_),
    .Y(_04940_));
 NAND2x1_ASAP7_75t_R _34546_ (.A(_02357_),
    .B(net2042),
    .Y(_04941_));
 NAND2x1_ASAP7_75t_R _34547_ (.A(_04634_),
    .B(_02092_),
    .Y(_04942_));
 AOI21x1_ASAP7_75t_R _34548_ (.A1(_04941_),
    .A2(_04942_),
    .B(_03004_),
    .Y(_04943_));
 NOR3x1_ASAP7_75t_R _34549_ (.A(_04943_),
    .B(_04935_),
    .C(_04938_),
    .Y(_04944_));
 OAI21x1_ASAP7_75t_R _34550_ (.A1(_04940_),
    .A2(_04944_),
    .B(net396),
    .Y(_04945_));
 INVx1_ASAP7_75t_R _34551_ (.A(_04945_),
    .Y(_04946_));
 INVx1_ASAP7_75t_R _34552_ (.A(_00458_),
    .Y(_04947_));
 OAI21x1_ASAP7_75t_R _34553_ (.A1(_04934_),
    .A2(_04946_),
    .B(_04947_),
    .Y(_04948_));
 INVx1_ASAP7_75t_R _34554_ (.A(_04934_),
    .Y(_04949_));
 NAND3x1_ASAP7_75t_R _34555_ (.A(_04945_),
    .B(_00458_),
    .C(_04949_),
    .Y(_04950_));
 NAND2x1_ASAP7_75t_R _34556_ (.A(_04948_),
    .B(_04950_),
    .Y(_00019_));
 AND2x2_ASAP7_75t_R _34557_ (.A(_18753_),
    .B(_00856_),
    .Y(_04951_));
 NOR2x1_ASAP7_75t_R _34558_ (.A(net2700),
    .B(net3176),
    .Y(_04952_));
 NOR2x1_ASAP7_75t_R _34559_ (.A(_04678_),
    .B(_04815_),
    .Y(_04953_));
 OAI21x1_ASAP7_75t_R _34560_ (.A1(_04952_),
    .A2(_04953_),
    .B(_04689_),
    .Y(_04954_));
 NOR2x1_ASAP7_75t_R _34561_ (.A(_03291_),
    .B(_04678_),
    .Y(_04955_));
 NOR2x1_ASAP7_75t_R _34562_ (.A(net2700),
    .B(_04815_),
    .Y(_04956_));
 OAI21x1_ASAP7_75t_R _34563_ (.A1(_04955_),
    .A2(_04956_),
    .B(_03710_),
    .Y(_04957_));
 NAND2x1_ASAP7_75t_R _34564_ (.A(_04954_),
    .B(_04957_),
    .Y(_04958_));
 NOR2x2_ASAP7_75t_R _34565_ (.A(_04809_),
    .B(_04810_),
    .Y(_04959_));
 XOR2x1_ASAP7_75t_R _34566_ (.A(_03382_),
    .Y(_04960_),
    .B(_04959_));
 NAND2x1_ASAP7_75t_R _34567_ (.A(_04960_),
    .B(_04958_),
    .Y(_04961_));
 XOR2x1_ASAP7_75t_R _34568_ (.A(_03377_),
    .Y(_04962_),
    .B(_04959_));
 XOR2x1_ASAP7_75t_R _34569_ (.A(_03292_),
    .Y(_04963_),
    .B(_04689_));
 NAND2x1_ASAP7_75t_R _34570_ (.A(_04963_),
    .B(_04962_),
    .Y(_04964_));
 AOI21x1_ASAP7_75t_R _34571_ (.A1(_04961_),
    .A2(_04964_),
    .B(_18753_),
    .Y(_04965_));
 INVx2_ASAP7_75t_R _34572_ (.A(_00457_),
    .Y(_04966_));
 OAI21x1_ASAP7_75t_R _34573_ (.A1(_04951_),
    .A2(_04965_),
    .B(_04966_),
    .Y(_04967_));
 NOR2x1_ASAP7_75t_R _34574_ (.A(net396),
    .B(_00856_),
    .Y(_04968_));
 XOR2x1_ASAP7_75t_R _34575_ (.A(_04959_),
    .Y(_04969_),
    .B(_03710_));
 NAND2x1_ASAP7_75t_R _34576_ (.A(_03378_),
    .B(_04969_),
    .Y(_04970_));
 XOR2x1_ASAP7_75t_R _34577_ (.A(_04959_),
    .Y(_04971_),
    .B(_04689_));
 NAND2x1_ASAP7_75t_R _34578_ (.A(_04971_),
    .B(_03383_),
    .Y(_04972_));
 AOI21x1_ASAP7_75t_R _34579_ (.A1(_04970_),
    .A2(_04972_),
    .B(_18753_),
    .Y(_04973_));
 OAI21x1_ASAP7_75t_R _34580_ (.A1(_04968_),
    .A2(_04973_),
    .B(_00457_),
    .Y(_04974_));
 NAND2x1_ASAP7_75t_R _34581_ (.A(_04974_),
    .B(_04967_),
    .Y(_00020_));
 AND2x2_ASAP7_75t_R _34582_ (.A(_18753_),
    .B(_00855_),
    .Y(_04975_));
 INVx1_ASAP7_75t_R _34583_ (.A(_04975_),
    .Y(_04976_));
 NOR2x1_ASAP7_75t_R _34584_ (.A(_03399_),
    .B(_04830_),
    .Y(_04977_));
 NOR2x1_ASAP7_75t_R _34585_ (.A(_03714_),
    .B(_04847_),
    .Y(_04978_));
 AOI21x1_ASAP7_75t_R _34586_ (.A1(_04865_),
    .A2(_04864_),
    .B(_04706_),
    .Y(_04979_));
 OAI21x1_ASAP7_75t_R _34587_ (.A1(_03576_),
    .A2(_03616_),
    .B(_03466_),
    .Y(_04980_));
 NAND2x1_ASAP7_75t_R _34588_ (.A(_03617_),
    .B(_04836_),
    .Y(_04981_));
 AOI21x1_ASAP7_75t_R _34589_ (.A1(_04980_),
    .A2(_04981_),
    .B(_04041_),
    .Y(_04982_));
 NOR2x1_ASAP7_75t_R _34590_ (.A(_04979_),
    .B(_04982_),
    .Y(_04983_));
 OAI21x1_ASAP7_75t_R _34591_ (.A1(_04977_),
    .A2(_04978_),
    .B(_04983_),
    .Y(_04984_));
 NOR2x1_ASAP7_75t_R _34592_ (.A(_03399_),
    .B(_04847_),
    .Y(_04985_));
 NOR2x1_ASAP7_75t_R _34593_ (.A(_03714_),
    .B(_04830_),
    .Y(_04986_));
 AOI21x1_ASAP7_75t_R _34594_ (.A1(_04865_),
    .A2(_04864_),
    .B(_04041_),
    .Y(_04987_));
 AOI21x1_ASAP7_75t_R _34595_ (.A1(_04980_),
    .A2(_04981_),
    .B(_04706_),
    .Y(_04988_));
 NOR2x1_ASAP7_75t_R _34596_ (.A(_04987_),
    .B(_04988_),
    .Y(_04989_));
 OAI21x1_ASAP7_75t_R _34597_ (.A1(_04985_),
    .A2(_04986_),
    .B(_04989_),
    .Y(_04990_));
 AOI21x1_ASAP7_75t_R _34598_ (.A1(_04984_),
    .A2(_04990_),
    .B(net388),
    .Y(_04991_));
 INVx1_ASAP7_75t_R _34599_ (.A(_04991_),
    .Y(_04992_));
 INVx1_ASAP7_75t_R _34600_ (.A(_00456_),
    .Y(_04993_));
 AOI21x1_ASAP7_75t_R _34601_ (.A1(_04976_),
    .A2(_04992_),
    .B(_04993_),
    .Y(_04994_));
 NOR3x1_ASAP7_75t_R _34602_ (.A(_04991_),
    .B(_00456_),
    .C(_04975_),
    .Y(_04995_));
 NOR2x1_ASAP7_75t_R _34603_ (.A(_04994_),
    .B(_04995_),
    .Y(_00021_));
 NOR2x2_ASAP7_75t_R _34604_ (.A(net395),
    .B(_00854_),
    .Y(_04996_));
 INVx1_ASAP7_75t_R _34605_ (.A(_04996_),
    .Y(_04997_));
 NOR2x2_ASAP7_75t_R _34606_ (.A(_03960_),
    .B(net3287),
    .Y(_04998_));
 NOR2x1_ASAP7_75t_R _34607_ (.A(_03973_),
    .B(_03970_),
    .Y(_04999_));
 OAI21x1_ASAP7_75t_R _34608_ (.A1(_04998_),
    .A2(_04999_),
    .B(_04719_),
    .Y(_05000_));
 INVx1_ASAP7_75t_R _34609_ (.A(_05000_),
    .Y(_05001_));
 NAND2x2_ASAP7_75t_R _34610_ (.A(_03960_),
    .B(_03809_),
    .Y(_05002_));
 OAI22x1_ASAP7_75t_R _34611_ (.A1(_03808_),
    .A2(_03734_),
    .B1(_03959_),
    .B2(_03885_),
    .Y(_05003_));
 NAND3x2_ASAP7_75t_R _34612_ (.B(_05003_),
    .C(net3140),
    .Y(_05004_),
    .A(_05002_));
 INVx1_ASAP7_75t_R _34613_ (.A(_05004_),
    .Y(_05005_));
 OAI21x1_ASAP7_75t_R _34614_ (.A1(_05001_),
    .A2(_05005_),
    .B(net2396),
    .Y(_05006_));
 INVx2_ASAP7_75t_R _34615_ (.A(net2396),
    .Y(_05007_));
 NAND3x1_ASAP7_75t_R _34616_ (.A(_05004_),
    .B(_05000_),
    .C(_05007_),
    .Y(_05008_));
 AOI21x1_ASAP7_75t_R _34617_ (.A1(_05006_),
    .A2(_05008_),
    .B(_18753_),
    .Y(_05009_));
 INVx1_ASAP7_75t_R _34618_ (.A(_05009_),
    .Y(_05010_));
 AOI21x1_ASAP7_75t_R _34619_ (.A1(_04997_),
    .A2(_05010_),
    .B(_00455_),
    .Y(_05011_));
 INVx1_ASAP7_75t_R _34620_ (.A(_00455_),
    .Y(_05012_));
 NOR3x1_ASAP7_75t_R _34621_ (.A(_05009_),
    .B(_05012_),
    .C(_04996_),
    .Y(_05013_));
 NOR2x1_ASAP7_75t_R _34622_ (.A(_05011_),
    .B(_05013_),
    .Y(_00022_));
 NOR2x1_ASAP7_75t_R _34623_ (.A(net395),
    .B(_00853_),
    .Y(_05014_));
 OAI21x1_ASAP7_75t_R _34624_ (.A1(_03971_),
    .A2(_03972_),
    .B(net3340),
    .Y(_05015_));
 AO21x2_ASAP7_75t_R _34625_ (.A1(_04045_),
    .A2(_03883_),
    .B(net3340),
    .Y(_05016_));
 NOR2x2_ASAP7_75t_R _34626_ (.A(_04363_),
    .B(_04364_),
    .Y(_05017_));
 AOI21x1_ASAP7_75t_R _34627_ (.A1(_05015_),
    .A2(_05016_),
    .B(_05017_),
    .Y(_05018_));
 INVx1_ASAP7_75t_R _34628_ (.A(_05018_),
    .Y(_05019_));
 NAND3x1_ASAP7_75t_R _34629_ (.A(_05016_),
    .B(_05017_),
    .C(_05015_),
    .Y(_05020_));
 AOI21x1_ASAP7_75t_R _34630_ (.A1(_05019_),
    .A2(_05020_),
    .B(_18753_),
    .Y(_05021_));
 OAI21x1_ASAP7_75t_R _34631_ (.A1(_05014_),
    .A2(_05021_),
    .B(_00454_),
    .Y(_05022_));
 NOR2x1_ASAP7_75t_R _34632_ (.A(net3287),
    .B(net3340),
    .Y(_05023_));
 NOR2x1_ASAP7_75t_R _34633_ (.A(_03970_),
    .B(_04729_),
    .Y(_05024_));
 OAI21x1_ASAP7_75t_R _34634_ (.A1(_05023_),
    .A2(_05024_),
    .B(_03881_),
    .Y(_05025_));
 XOR2x1_ASAP7_75t_R _34635_ (.A(_04525_),
    .Y(_05026_),
    .B(net3287));
 NAND2x1_ASAP7_75t_R _34636_ (.A(_04359_),
    .B(_05026_),
    .Y(_05027_));
 INVx1_ASAP7_75t_R _34637_ (.A(_05017_),
    .Y(_05028_));
 AOI21x1_ASAP7_75t_R _34638_ (.A1(_05025_),
    .A2(_05027_),
    .B(_05028_),
    .Y(_05029_));
 OAI21x1_ASAP7_75t_R _34639_ (.A1(_05018_),
    .A2(_05029_),
    .B(net395),
    .Y(_05030_));
 INVx1_ASAP7_75t_R _34640_ (.A(_00454_),
    .Y(_05031_));
 INVx1_ASAP7_75t_R _34641_ (.A(_05014_),
    .Y(_05032_));
 NAND3x1_ASAP7_75t_R _34642_ (.A(_05030_),
    .B(_05031_),
    .C(_05032_),
    .Y(_05033_));
 NAND2x1_ASAP7_75t_R _34643_ (.A(_05033_),
    .B(_05022_),
    .Y(_00023_));
 AND2x2_ASAP7_75t_R _34644_ (.A(_18753_),
    .B(_00852_),
    .Y(_05034_));
 OA21x2_ASAP7_75t_R _34645_ (.A1(_04281_),
    .A2(_04280_),
    .B(net3269),
    .Y(_05035_));
 OA21x2_ASAP7_75t_R _34646_ (.A1(_04206_),
    .A2(_04202_),
    .B(net2031),
    .Y(_05036_));
 XNOR2x2_ASAP7_75t_R _34647_ (.A(net2710),
    .B(_04606_),
    .Y(_05037_));
 INVx1_ASAP7_75t_R _34648_ (.A(_05037_),
    .Y(_05038_));
 OAI21x1_ASAP7_75t_R _34649_ (.A1(_05035_),
    .A2(_05036_),
    .B(_05038_),
    .Y(_05039_));
 OA21x2_ASAP7_75t_R _34650_ (.A1(_04206_),
    .A2(_04202_),
    .B(net3269),
    .Y(_05040_));
 OA21x2_ASAP7_75t_R _34651_ (.A1(_04281_),
    .A2(_04280_),
    .B(net2031),
    .Y(_05041_));
 OAI21x1_ASAP7_75t_R _34652_ (.A1(_05040_),
    .A2(_05041_),
    .B(_05037_),
    .Y(_05042_));
 AOI21x1_ASAP7_75t_R _34653_ (.A1(_05039_),
    .A2(_05042_),
    .B(_18753_),
    .Y(_05043_));
 INVx1_ASAP7_75t_R _34654_ (.A(_00453_),
    .Y(_05044_));
 OAI21x1_ASAP7_75t_R _34655_ (.A1(_05034_),
    .A2(_05043_),
    .B(_05044_),
    .Y(_05045_));
 NOR2x1_ASAP7_75t_R _34656_ (.A(net396),
    .B(_00852_),
    .Y(_05046_));
 OAI21x1_ASAP7_75t_R _34657_ (.A1(_05035_),
    .A2(_05036_),
    .B(_05037_),
    .Y(_05047_));
 OAI21x1_ASAP7_75t_R _34658_ (.A1(_05040_),
    .A2(_05041_),
    .B(_05038_),
    .Y(_05048_));
 AOI21x1_ASAP7_75t_R _34659_ (.A1(_05047_),
    .A2(_05048_),
    .B(_18753_),
    .Y(_05049_));
 OAI21x1_ASAP7_75t_R _34660_ (.A1(_05046_),
    .A2(_05049_),
    .B(_00453_),
    .Y(_05050_));
 NAND2x1_ASAP7_75t_R _34661_ (.A(_05050_),
    .B(_05045_),
    .Y(_00024_));
 NOR2x1_ASAP7_75t_R _34662_ (.A(net394),
    .B(_00851_),
    .Y(_05051_));
 INVx1_ASAP7_75t_R _34663_ (.A(_05051_),
    .Y(_05052_));
 TAPCELL_ASAP7_75t_R PHY_534 ();
 TAPCELL_ASAP7_75t_R PHY_533 ();
 TAPCELL_ASAP7_75t_R PHY_532 ();
 NOR2x2_ASAP7_75t_R _34667_ (.A(_00621_),
    .B(net3099),
    .Y(_05056_));
 TAPCELL_ASAP7_75t_R PHY_531 ();
 NAND2x2_ASAP7_75t_R _34669_ (.A(net3438),
    .B(net1491),
    .Y(_05058_));
 INVx2_ASAP7_75t_R _34670_ (.A(_05058_),
    .Y(_05059_));
 NOR2x2_ASAP7_75t_R _34671_ (.A(_00617_),
    .B(_00618_),
    .Y(_05060_));
 AND2x6_ASAP7_75t_R _34672_ (.A(_00619_),
    .B(_00620_),
    .Y(_05061_));
 NAND2x2_ASAP7_75t_R _34673_ (.A(_05060_),
    .B(_05061_),
    .Y(_05062_));
 INVx3_ASAP7_75t_R _34674_ (.A(_05062_),
    .Y(_05063_));
 NAND2x1_ASAP7_75t_R _34675_ (.A(_05059_),
    .B(_05063_),
    .Y(_05064_));
 INVx5_ASAP7_75t_R _34676_ (.A(net2468),
    .Y(_05065_));
 NOR2x2_ASAP7_75t_R _34677_ (.A(net2782),
    .B(_05065_),
    .Y(_05066_));
 TAPCELL_ASAP7_75t_R PHY_530 ();
 INVx11_ASAP7_75t_R _34679_ (.A(net1147),
    .Y(_05068_));
 NOR2x2_ASAP7_75t_R _34680_ (.A(net1319),
    .B(_05068_),
    .Y(_05069_));
 NAND2x2_ASAP7_75t_R _34681_ (.A(net2171),
    .B(_05069_),
    .Y(_05070_));
 TAPCELL_ASAP7_75t_R PHY_529 ();
 NOR2x2_ASAP7_75t_R _34683_ (.A(net1319),
    .B(net1147),
    .Y(_05072_));
 NAND2x2_ASAP7_75t_R _34684_ (.A(_05072_),
    .B(net2169),
    .Y(_05073_));
 TAPCELL_ASAP7_75t_R PHY_528 ();
 INVx2_ASAP7_75t_R _34686_ (.A(_00619_),
    .Y(_05075_));
 NOR2x2_ASAP7_75t_R _34687_ (.A(_00620_),
    .B(_05075_),
    .Y(_05076_));
 INVx3_ASAP7_75t_R _34688_ (.A(_00617_),
    .Y(_05077_));
 NOR2x2_ASAP7_75t_R _34689_ (.A(_00618_),
    .B(_05077_),
    .Y(_05078_));
 NAND2x2_ASAP7_75t_R _34690_ (.A(_05076_),
    .B(_05078_),
    .Y(_05079_));
 TAPCELL_ASAP7_75t_R PHY_527 ();
 AO21x1_ASAP7_75t_R _34692_ (.A1(net1764),
    .A2(_05073_),
    .B(net2493),
    .Y(_05081_));
 NAND2x2_ASAP7_75t_R _34693_ (.A(_05064_),
    .B(_05081_),
    .Y(_05082_));
 NAND2x2_ASAP7_75t_R _34694_ (.A(_00621_),
    .B(_00622_),
    .Y(_05083_));
 NOR2x2_ASAP7_75t_R _34695_ (.A(net1156),
    .B(net1522),
    .Y(_05084_));
 NOR2x2_ASAP7_75t_R _34696_ (.A(_00619_),
    .B(_00620_),
    .Y(_05085_));
 NAND2x2_ASAP7_75t_R _34697_ (.A(_05085_),
    .B(_05078_),
    .Y(_05086_));
 CKINVDCx6p67_ASAP7_75t_R _34698_ (.A(_05086_),
    .Y(_05087_));
 NAND2x2_ASAP7_75t_R _34699_ (.A(_05084_),
    .B(_05087_),
    .Y(_05088_));
 NAND2x2_ASAP7_75t_R _34700_ (.A(net1319),
    .B(net1147),
    .Y(_05089_));
 NAND2x2_ASAP7_75t_R _34701_ (.A(net2782),
    .B(_05065_),
    .Y(_05090_));
 TAPCELL_ASAP7_75t_R PHY_526 ();
 NOR2x2_ASAP7_75t_R _34703_ (.A(_05089_),
    .B(_05090_),
    .Y(_05092_));
 INVx2_ASAP7_75t_R _34704_ (.A(_00622_),
    .Y(_05093_));
 NOR2x2_ASAP7_75t_R _34705_ (.A(net3094),
    .B(_05093_),
    .Y(_05094_));
 NAND2x2_ASAP7_75t_R _34706_ (.A(_05072_),
    .B(net2223),
    .Y(_05095_));
 INVx3_ASAP7_75t_R _34707_ (.A(_05095_),
    .Y(_05096_));
 NAND2x2_ASAP7_75t_R _34708_ (.A(_00617_),
    .B(_00618_),
    .Y(_05097_));
 INVx2_ASAP7_75t_R _34709_ (.A(_00620_),
    .Y(_05098_));
 NAND2x1_ASAP7_75t_R _34710_ (.A(_00619_),
    .B(_05098_),
    .Y(_05099_));
 NOR2x2_ASAP7_75t_R _34711_ (.A(_05097_),
    .B(_05099_),
    .Y(_05100_));
 OAI21x1_ASAP7_75t_R _34712_ (.A1(_05092_),
    .A2(_05096_),
    .B(_05100_),
    .Y(_05101_));
 NAND2x2_ASAP7_75t_R _34713_ (.A(_05088_),
    .B(_05101_),
    .Y(_05102_));
 CKINVDCx16_ASAP7_75t_R _34714_ (.A(net1326),
    .Y(_05103_));
 NOR2x2_ASAP7_75t_R _34715_ (.A(net1151),
    .B(_05103_),
    .Y(_05104_));
 NAND2x2_ASAP7_75t_R _34716_ (.A(net1485),
    .B(_05104_),
    .Y(_05105_));
 INVx5_ASAP7_75t_R _34717_ (.A(_05105_),
    .Y(_05106_));
 NAND2x2_ASAP7_75t_R _34718_ (.A(_05078_),
    .B(_05061_),
    .Y(_05107_));
 CKINVDCx5p33_ASAP7_75t_R _34719_ (.A(_05107_),
    .Y(_05108_));
 NAND2x2_ASAP7_75t_R _34720_ (.A(_05106_),
    .B(_05108_),
    .Y(_05109_));
 NOR2x2_ASAP7_75t_R _34721_ (.A(net1148),
    .B(_05090_),
    .Y(_05110_));
 TAPCELL_ASAP7_75t_R PHY_525 ();
 NAND2x1_ASAP7_75t_R _34723_ (.A(net1148),
    .B(net1487),
    .Y(_05112_));
 INVx1_ASAP7_75t_R _34724_ (.A(_05112_),
    .Y(_05113_));
 OAI21x1_ASAP7_75t_R _34725_ (.A1(_05110_),
    .A2(_05113_),
    .B(_05108_),
    .Y(_05114_));
 NAND2x2_ASAP7_75t_R _34726_ (.A(_05109_),
    .B(_05114_),
    .Y(_05115_));
 NOR3x2_ASAP7_75t_R _34727_ (.B(_05102_),
    .C(_05115_),
    .Y(_05116_),
    .A(_05082_));
 NOR2x2_ASAP7_75t_R _34728_ (.A(_00619_),
    .B(_05098_),
    .Y(_05117_));
 NAND2x2_ASAP7_75t_R _34729_ (.A(_05060_),
    .B(_05117_),
    .Y(_05118_));
 NAND2x2_ASAP7_75t_R _34730_ (.A(net1323),
    .B(net2169),
    .Y(_05119_));
 NOR2x1_ASAP7_75t_R _34731_ (.A(_05118_),
    .B(_05119_),
    .Y(_05120_));
 INVx2_ASAP7_75t_R _34732_ (.A(_05120_),
    .Y(_05121_));
 NAND2x2_ASAP7_75t_R _34733_ (.A(_05068_),
    .B(net2169),
    .Y(_05122_));
 INVx2_ASAP7_75t_R _34734_ (.A(_05122_),
    .Y(_05123_));
 NAND2x2_ASAP7_75t_R _34735_ (.A(_05123_),
    .B(_05087_),
    .Y(_05124_));
 TAPCELL_ASAP7_75t_R PHY_524 ();
 NAND2x2_ASAP7_75t_R _34737_ (.A(_05060_),
    .B(_05076_),
    .Y(_05126_));
 CKINVDCx6p67_ASAP7_75t_R _34738_ (.A(_05126_),
    .Y(_05127_));
 NAND2x2_ASAP7_75t_R _34739_ (.A(net2223),
    .B(_05127_),
    .Y(_05128_));
 NAND3x2_ASAP7_75t_R _34740_ (.B(_05124_),
    .C(_05128_),
    .Y(_05129_),
    .A(_05121_));
 TAPCELL_ASAP7_75t_R PHY_523 ();
 NAND2x2_ASAP7_75t_R _34742_ (.A(_05072_),
    .B(net1485),
    .Y(_05131_));
 TAPCELL_ASAP7_75t_R PHY_522 ();
 TAPCELL_ASAP7_75t_R PHY_521 ();
 AO21x2_ASAP7_75t_R _34745_ (.A1(_05105_),
    .A2(net2643),
    .B(_05118_),
    .Y(_05134_));
 NAND2x2_ASAP7_75t_R _34746_ (.A(net1490),
    .B(_05069_),
    .Y(_05135_));
 TAPCELL_ASAP7_75t_R PHY_520 ();
 TAPCELL_ASAP7_75t_R PHY_519 ();
 NAND2x2_ASAP7_75t_R _34749_ (.A(_05060_),
    .B(_05085_),
    .Y(_05138_));
 TAPCELL_ASAP7_75t_R PHY_518 ();
 AO21x1_ASAP7_75t_R _34751_ (.A1(net990),
    .A2(_05090_),
    .B(_05138_),
    .Y(_05140_));
 TAPCELL_ASAP7_75t_R PHY_517 ();
 NOR2x2_ASAP7_75t_R _34753_ (.A(net1320),
    .B(net1520),
    .Y(_05142_));
 INVx4_ASAP7_75t_R _34754_ (.A(_05142_),
    .Y(_05143_));
 NOR2x1_ASAP7_75t_R _34755_ (.A(_05138_),
    .B(_05143_),
    .Y(_05144_));
 INVx1_ASAP7_75t_R _34756_ (.A(_05144_),
    .Y(_05145_));
 NAND3x2_ASAP7_75t_R _34757_ (.B(_05140_),
    .C(_05145_),
    .Y(_05146_),
    .A(_05134_));
 NOR2x2_ASAP7_75t_R _34758_ (.A(_05129_),
    .B(_05146_),
    .Y(_05147_));
 NAND2x2_ASAP7_75t_R _34759_ (.A(_05116_),
    .B(_05147_),
    .Y(_05148_));
 INVx1_ASAP7_75t_R _34760_ (.A(_05148_),
    .Y(_05149_));
 NAND2x2_ASAP7_75t_R _34761_ (.A(_05103_),
    .B(net2226),
    .Y(_05150_));
 INVx4_ASAP7_75t_R _34762_ (.A(_05150_),
    .Y(_05151_));
 INVx4_ASAP7_75t_R _34763_ (.A(_05097_),
    .Y(_05152_));
 NAND2x2_ASAP7_75t_R _34764_ (.A(_05061_),
    .B(_05152_),
    .Y(_05153_));
 INVx5_ASAP7_75t_R _34765_ (.A(_05153_),
    .Y(_05154_));
 NAND2x2_ASAP7_75t_R _34766_ (.A(_05151_),
    .B(_05154_),
    .Y(_05155_));
 NAND2x2_ASAP7_75t_R _34767_ (.A(net2169),
    .B(net3456),
    .Y(_05156_));
 NAND2x2_ASAP7_75t_R _34768_ (.A(net3456),
    .B(net2223),
    .Y(_05157_));
 TAPCELL_ASAP7_75t_R PHY_516 ();
 TAPCELL_ASAP7_75t_R PHY_515 ();
 AO21x1_ASAP7_75t_R _34771_ (.A1(net1867),
    .A2(net2056),
    .B(_05153_),
    .Y(_05160_));
 NAND2x1_ASAP7_75t_R _34772_ (.A(_05155_),
    .B(_05160_),
    .Y(_05161_));
 INVx5_ASAP7_75t_R _34773_ (.A(_05083_),
    .Y(_05162_));
 NAND2x2_ASAP7_75t_R _34774_ (.A(_05069_),
    .B(_05162_),
    .Y(_05163_));
 TAPCELL_ASAP7_75t_R PHY_514 ();
 NAND2x2_ASAP7_75t_R _34776_ (.A(_05072_),
    .B(_05162_),
    .Y(_05165_));
 TAPCELL_ASAP7_75t_R PHY_513 ();
 AO21x1_ASAP7_75t_R _34778_ (.A1(net3440),
    .A2(net2315),
    .B(_05153_),
    .Y(_05167_));
 AO21x2_ASAP7_75t_R _34779_ (.A1(_05070_),
    .A2(_05073_),
    .B(_05153_),
    .Y(_05168_));
 NAND2x1_ASAP7_75t_R _34780_ (.A(_05167_),
    .B(_05168_),
    .Y(_05169_));
 NOR2x2_ASAP7_75t_R _34781_ (.A(_05161_),
    .B(_05169_),
    .Y(_05170_));
 INVx3_ASAP7_75t_R _34782_ (.A(net3108),
    .Y(_05171_));
 NAND2x1_ASAP7_75t_R _34783_ (.A(_05110_),
    .B(_05171_),
    .Y(_05172_));
 INVx3_ASAP7_75t_R _34784_ (.A(net1945),
    .Y(_05173_));
 NAND2x2_ASAP7_75t_R _34785_ (.A(_05078_),
    .B(_05117_),
    .Y(_05174_));
 INVx3_ASAP7_75t_R _34786_ (.A(_05174_),
    .Y(_05175_));
 NAND2x1_ASAP7_75t_R _34787_ (.A(_05173_),
    .B(_05175_),
    .Y(_05176_));
 NAND2x2_ASAP7_75t_R _34788_ (.A(net2467),
    .B(_05093_),
    .Y(_05177_));
 NOR2x2_ASAP7_75t_R _34789_ (.A(net1305),
    .B(_05177_),
    .Y(_05178_));
 NAND2x2_ASAP7_75t_R _34790_ (.A(_00620_),
    .B(_05075_),
    .Y(_05179_));
 NAND2x1_ASAP7_75t_R _34791_ (.A(_00618_),
    .B(_05077_),
    .Y(_05180_));
 NOR2x2_ASAP7_75t_R _34792_ (.A(_05179_),
    .B(_05180_),
    .Y(_05181_));
 NAND2x1_ASAP7_75t_R _34793_ (.A(_05178_),
    .B(_05181_),
    .Y(_05182_));
 NAND3x1_ASAP7_75t_R _34794_ (.A(_05172_),
    .B(_05176_),
    .C(_05182_),
    .Y(_05183_));
 INVx6_ASAP7_75t_R _34795_ (.A(_05089_),
    .Y(_05184_));
 NAND2x2_ASAP7_75t_R _34796_ (.A(net1485),
    .B(_05184_),
    .Y(_05185_));
 NAND2x2_ASAP7_75t_R _34797_ (.A(_05117_),
    .B(_05152_),
    .Y(_05186_));
 TAPCELL_ASAP7_75t_R PHY_512 ();
 AO21x1_ASAP7_75t_R _34799_ (.A1(net1767),
    .A2(net3451),
    .B(_05186_),
    .Y(_05188_));
 TAPCELL_ASAP7_75t_R PHY_511 ();
 NAND2x2_ASAP7_75t_R _34801_ (.A(net1152),
    .B(_05103_),
    .Y(_05190_));
 NOR2x2_ASAP7_75t_R _34802_ (.A(_05177_),
    .B(_05190_),
    .Y(_05191_));
 AOI22x1_ASAP7_75t_R _34803_ (.A1(_05154_),
    .A2(_05106_),
    .B1(_05100_),
    .B2(net3409),
    .Y(_05192_));
 NAND2x1_ASAP7_75t_R _34804_ (.A(_05188_),
    .B(_05192_),
    .Y(_05193_));
 NOR2x1_ASAP7_75t_R _34805_ (.A(_05183_),
    .B(_05193_),
    .Y(_05194_));
 NAND2x2_ASAP7_75t_R _34806_ (.A(_05170_),
    .B(_05194_),
    .Y(_05195_));
 INVx3_ASAP7_75t_R _34807_ (.A(_00618_),
    .Y(_05196_));
 NOR2x2_ASAP7_75t_R _34808_ (.A(_00617_),
    .B(_05196_),
    .Y(_05197_));
 NAND2x2_ASAP7_75t_R _34809_ (.A(_05076_),
    .B(_05197_),
    .Y(_05198_));
 INVx5_ASAP7_75t_R _34810_ (.A(_05198_),
    .Y(_05199_));
 NOR2x2_ASAP7_75t_R _34811_ (.A(net1524),
    .B(_05190_),
    .Y(_05200_));
 INVx4_ASAP7_75t_R _34812_ (.A(_05118_),
    .Y(_05201_));
 INVx3_ASAP7_75t_R _34813_ (.A(_05072_),
    .Y(_05202_));
 NOR2x2_ASAP7_75t_R _34814_ (.A(_05083_),
    .B(_05202_),
    .Y(_05203_));
 AOI22x1_ASAP7_75t_R _34815_ (.A1(_05199_),
    .A2(_05200_),
    .B1(_05201_),
    .B2(_05203_),
    .Y(_05204_));
 NOR2x2_ASAP7_75t_R _34816_ (.A(_05089_),
    .B(_05083_),
    .Y(_05205_));
 INVx11_ASAP7_75t_R _34817_ (.A(_05205_),
    .Y(_05206_));
 NOR2x1_ASAP7_75t_R _34818_ (.A(net3103),
    .B(_05206_),
    .Y(_05207_));
 NAND2x2_ASAP7_75t_R _34819_ (.A(_05197_),
    .B(_05061_),
    .Y(_05208_));
 NOR2x1_ASAP7_75t_R _34820_ (.A(_05208_),
    .B(_05163_),
    .Y(_05209_));
 NOR2x1_ASAP7_75t_R _34821_ (.A(_05207_),
    .B(_05209_),
    .Y(_05210_));
 NAND2x2_ASAP7_75t_R _34822_ (.A(net2223),
    .B(_05184_),
    .Y(_05211_));
 AO21x1_ASAP7_75t_R _34823_ (.A1(_05211_),
    .A2(net1836),
    .B(net3444),
    .Y(_05212_));
 AND3x1_ASAP7_75t_R _34824_ (.A(_05204_),
    .B(_05210_),
    .C(_05212_),
    .Y(_05213_));
 TAPCELL_ASAP7_75t_R PHY_510 ();
 NAND2x2_ASAP7_75t_R _34826_ (.A(_05085_),
    .B(_05152_),
    .Y(_05215_));
 AO21x1_ASAP7_75t_R _34827_ (.A1(_05211_),
    .A2(net1764),
    .B(_05215_),
    .Y(_05216_));
 NAND2x2_ASAP7_75t_R _34828_ (.A(net1319),
    .B(_05068_),
    .Y(_05217_));
 NOR2x2_ASAP7_75t_R _34829_ (.A(_05083_),
    .B(_05217_),
    .Y(_05218_));
 NOR2x1_ASAP7_75t_R _34830_ (.A(net3410),
    .B(net2418),
    .Y(_05219_));
 AOI21x1_ASAP7_75t_R _34831_ (.A1(_05199_),
    .A2(_05218_),
    .B(_05219_),
    .Y(_05220_));
 NAND2x1_ASAP7_75t_R _34832_ (.A(_05216_),
    .B(_05220_),
    .Y(_05221_));
 NAND2x2_ASAP7_75t_R _34833_ (.A(net2169),
    .B(_05184_),
    .Y(_05222_));
 NOR2x1_ASAP7_75t_R _34834_ (.A(_05138_),
    .B(net2126),
    .Y(_05223_));
 AOI21x1_ASAP7_75t_R _34835_ (.A1(_05127_),
    .A2(_05200_),
    .B(_05223_),
    .Y(_05224_));
 NAND2x2_ASAP7_75t_R _34836_ (.A(net3443),
    .B(_05162_),
    .Y(_05225_));
 NOR2x1_ASAP7_75t_R _34837_ (.A(_05138_),
    .B(_05225_),
    .Y(_05226_));
 AOI21x1_ASAP7_75t_R _34838_ (.A1(_05201_),
    .A2(_05205_),
    .B(_05226_),
    .Y(_05227_));
 NAND2x1_ASAP7_75t_R _34839_ (.A(_05224_),
    .B(_05227_),
    .Y(_05228_));
 NOR2x1_ASAP7_75t_R _34840_ (.A(_05221_),
    .B(_05228_),
    .Y(_05229_));
 NAND2x2_ASAP7_75t_R _34841_ (.A(_05213_),
    .B(_05229_),
    .Y(_05230_));
 NOR2x1_ASAP7_75t_R _34842_ (.A(_05195_),
    .B(_05230_),
    .Y(_05231_));
 NAND2x1_ASAP7_75t_R _34843_ (.A(_05149_),
    .B(_05231_),
    .Y(_05232_));
 INVx3_ASAP7_75t_R _34844_ (.A(_05084_),
    .Y(_05233_));
 AO21x1_ASAP7_75t_R _34845_ (.A1(net3440),
    .A2(_05233_),
    .B(_05215_),
    .Y(_05234_));
 NAND2x1_ASAP7_75t_R _34846_ (.A(net1401),
    .B(net1945),
    .Y(_05235_));
 OAI21x1_ASAP7_75t_R _34847_ (.A1(_05096_),
    .A2(_05235_),
    .B(_05087_),
    .Y(_05236_));
 NAND2x1_ASAP7_75t_R _34848_ (.A(_05234_),
    .B(_05236_),
    .Y(_05237_));
 NOR2x2_ASAP7_75t_R _34849_ (.A(net3439),
    .B(net2272),
    .Y(_05238_));
 NOR2x2_ASAP7_75t_R _34850_ (.A(_05177_),
    .B(_05202_),
    .Y(_05239_));
 NAND2x2_ASAP7_75t_R _34851_ (.A(_05085_),
    .B(_05197_),
    .Y(_05240_));
 INVx4_ASAP7_75t_R _34852_ (.A(_05240_),
    .Y(_05241_));
 OAI21x1_ASAP7_75t_R _34853_ (.A1(_05238_),
    .A2(_05239_),
    .B(_05241_),
    .Y(_05242_));
 NOR2x1_ASAP7_75t_R _34854_ (.A(net1525),
    .B(_05072_),
    .Y(_05243_));
 INVx2_ASAP7_75t_R _34855_ (.A(_05243_),
    .Y(_05244_));
 NOR2x2_ASAP7_75t_R _34856_ (.A(_05186_),
    .B(_05244_),
    .Y(_05245_));
 INVx3_ASAP7_75t_R _34857_ (.A(_05245_),
    .Y(_05246_));
 NOR2x2_ASAP7_75t_R _34858_ (.A(_05097_),
    .B(_05179_),
    .Y(_05247_));
 TAPCELL_ASAP7_75t_R PHY_509 ();
 NOR2x2_ASAP7_75t_R _34860_ (.A(_05090_),
    .B(_05184_),
    .Y(_05249_));
 NAND2x2_ASAP7_75t_R _34861_ (.A(_05247_),
    .B(_05249_),
    .Y(_05250_));
 NAND3x2_ASAP7_75t_R _34862_ (.B(_05246_),
    .C(_05250_),
    .Y(_05251_),
    .A(_05242_));
 NOR2x2_ASAP7_75t_R _34863_ (.A(_05237_),
    .B(_05251_),
    .Y(_05252_));
 TAPCELL_ASAP7_75t_R PHY_508 ();
 AO21x1_ASAP7_75t_R _34865_ (.A1(_05206_),
    .A2(_05143_),
    .B(_05240_),
    .Y(_05254_));
 NAND2x1_ASAP7_75t_R _34866_ (.A(net1485),
    .B(_05190_),
    .Y(_05255_));
 NAND2x2_ASAP7_75t_R _34867_ (.A(_05117_),
    .B(_05197_),
    .Y(_05256_));
 TAPCELL_ASAP7_75t_R PHY_507 ();
 AO21x1_ASAP7_75t_R _34869_ (.A1(net2056),
    .A2(_05255_),
    .B(_05256_),
    .Y(_05258_));
 NAND2x2_ASAP7_75t_R _34870_ (.A(_05103_),
    .B(net1488),
    .Y(_05259_));
 TAPCELL_ASAP7_75t_R PHY_506 ();
 AO21x1_ASAP7_75t_R _34872_ (.A1(_05105_),
    .A2(_05259_),
    .B(_05208_),
    .Y(_05261_));
 AND3x2_ASAP7_75t_R _34873_ (.A(_05254_),
    .B(_05258_),
    .C(_05261_),
    .Y(_05262_));
 AO21x1_ASAP7_75t_R _34874_ (.A1(_05222_),
    .A2(_05122_),
    .B(_05208_),
    .Y(_05263_));
 NOR2x2_ASAP7_75t_R _34875_ (.A(_05103_),
    .B(net1524),
    .Y(_05264_));
 INVx3_ASAP7_75t_R _34876_ (.A(_05264_),
    .Y(_05265_));
 AO21x1_ASAP7_75t_R _34877_ (.A1(_05265_),
    .A2(_05165_),
    .B(net2493),
    .Y(_05266_));
 OAI21x1_ASAP7_75t_R _34878_ (.A1(_05092_),
    .A2(_05110_),
    .B(_05175_),
    .Y(_05267_));
 AND3x1_ASAP7_75t_R _34879_ (.A(_05263_),
    .B(_05266_),
    .C(_05267_),
    .Y(_05268_));
 NAND3x2_ASAP7_75t_R _34880_ (.B(_05262_),
    .C(_05268_),
    .Y(_05269_),
    .A(_05252_));
 INVx1_ASAP7_75t_R _34881_ (.A(_05269_),
    .Y(_05270_));
 NAND2x2_ASAP7_75t_R _34882_ (.A(net1150),
    .B(net2170),
    .Y(_05271_));
 NOR2x2_ASAP7_75t_R _34883_ (.A(_05271_),
    .B(_05174_),
    .Y(_05272_));
 INVx1_ASAP7_75t_R _34884_ (.A(_05272_),
    .Y(_05273_));
 AO21x1_ASAP7_75t_R _34885_ (.A1(net3449),
    .A2(_05073_),
    .B(_05174_),
    .Y(_05274_));
 NAND2x1_ASAP7_75t_R _34886_ (.A(_05273_),
    .B(_05274_),
    .Y(_05275_));
 AO21x1_ASAP7_75t_R _34887_ (.A1(net3369),
    .A2(net1945),
    .B(_05126_),
    .Y(_05276_));
 NOR2x1_ASAP7_75t_R _34888_ (.A(_05095_),
    .B(_05208_),
    .Y(_05277_));
 NOR2x1_ASAP7_75t_R _34889_ (.A(_05222_),
    .B(_05107_),
    .Y(_05278_));
 NOR2x1_ASAP7_75t_R _34890_ (.A(_05277_),
    .B(_05278_),
    .Y(_05279_));
 NAND2x1_ASAP7_75t_R _34891_ (.A(_05276_),
    .B(_05279_),
    .Y(_05280_));
 NOR2x1_ASAP7_75t_R _34892_ (.A(_05275_),
    .B(_05280_),
    .Y(_05281_));
 NAND2x1_ASAP7_75t_R _34893_ (.A(net1945),
    .B(net3440),
    .Y(_05282_));
 OAI21x1_ASAP7_75t_R _34894_ (.A1(_05110_),
    .A2(_05282_),
    .B(_05063_),
    .Y(_05283_));
 TAPCELL_ASAP7_75t_R PHY_505 ();
 TAPCELL_ASAP7_75t_R PHY_504 ();
 AO21x1_ASAP7_75t_R _34897_ (.A1(_05206_),
    .A2(net3446),
    .B(net2621),
    .Y(_05286_));
 AO21x1_ASAP7_75t_R _34898_ (.A1(_05206_),
    .A2(net2056),
    .B(_05208_),
    .Y(_05287_));
 NAND3x1_ASAP7_75t_R _34899_ (.A(_05283_),
    .B(_05286_),
    .C(_05287_),
    .Y(_05288_));
 INVx1_ASAP7_75t_R _34900_ (.A(_05288_),
    .Y(_05289_));
 NAND2x1_ASAP7_75t_R _34901_ (.A(_05281_),
    .B(_05289_),
    .Y(_05290_));
 NOR2x2_ASAP7_75t_R _34902_ (.A(_05058_),
    .B(_05215_),
    .Y(_05291_));
 AOI21x1_ASAP7_75t_R _34903_ (.A1(_05131_),
    .A2(net1945),
    .B(_05186_),
    .Y(_05292_));
 NOR2x2_ASAP7_75t_R _34904_ (.A(_05291_),
    .B(_05292_),
    .Y(_05293_));
 NAND2x2_ASAP7_75t_R _34905_ (.A(_05142_),
    .B(_05100_),
    .Y(_05294_));
 TAPCELL_ASAP7_75t_R PHY_503 ();
 AO21x1_ASAP7_75t_R _34907_ (.A1(net990),
    .A2(net964),
    .B(_05198_),
    .Y(_05296_));
 NAND3x2_ASAP7_75t_R _34908_ (.B(_05294_),
    .C(_05296_),
    .Y(_05297_),
    .A(_05293_));
 INVx1_ASAP7_75t_R _34909_ (.A(_05297_),
    .Y(_05298_));
 NOR2x1_ASAP7_75t_R _34910_ (.A(_05240_),
    .B(_05185_),
    .Y(_05299_));
 NOR2x1_ASAP7_75t_R _34911_ (.A(_05165_),
    .B(_05174_),
    .Y(_05300_));
 NOR2x1_ASAP7_75t_R _34912_ (.A(_05299_),
    .B(_05300_),
    .Y(_05301_));
 NOR2x1_ASAP7_75t_R _34913_ (.A(_05131_),
    .B(_05079_),
    .Y(_05302_));
 NOR2x1_ASAP7_75t_R _34914_ (.A(_05225_),
    .B(_05174_),
    .Y(_05303_));
 NOR2x1_ASAP7_75t_R _34915_ (.A(_05302_),
    .B(_05303_),
    .Y(_05304_));
 NAND2x1_ASAP7_75t_R _34916_ (.A(_05301_),
    .B(_05304_),
    .Y(_05305_));
 NAND2x2_ASAP7_75t_R _34917_ (.A(_05076_),
    .B(_05152_),
    .Y(_05306_));
 OAI22x1_ASAP7_75t_R _34918_ (.A1(net3369),
    .A2(_05306_),
    .B1(_05153_),
    .B2(net990),
    .Y(_05307_));
 NOR2x2_ASAP7_75t_R _34919_ (.A(_05177_),
    .B(_05217_),
    .Y(_05308_));
 NAND2x1_ASAP7_75t_R _34920_ (.A(_05247_),
    .B(_05308_),
    .Y(_05309_));
 OAI21x1_ASAP7_75t_R _34921_ (.A1(net964),
    .A2(_05215_),
    .B(_05309_),
    .Y(_05310_));
 NOR2x1_ASAP7_75t_R _34922_ (.A(_05307_),
    .B(_05310_),
    .Y(_05311_));
 INVx1_ASAP7_75t_R _34923_ (.A(_05311_),
    .Y(_05312_));
 NOR2x1_ASAP7_75t_R _34924_ (.A(_05305_),
    .B(_05312_),
    .Y(_05313_));
 NAND2x1_ASAP7_75t_R _34925_ (.A(_05298_),
    .B(_05313_),
    .Y(_05314_));
 NOR2x1_ASAP7_75t_R _34926_ (.A(_05290_),
    .B(_05314_),
    .Y(_05315_));
 NAND2x2_ASAP7_75t_R _34927_ (.A(_05270_),
    .B(_05315_),
    .Y(_05316_));
 NOR2x2_ASAP7_75t_R _34928_ (.A(_05232_),
    .B(_05316_),
    .Y(_05317_));
 AO21x2_ASAP7_75t_R _34929_ (.A1(net3427),
    .A2(_05211_),
    .B(_05153_),
    .Y(_05318_));
 NAND2x2_ASAP7_75t_R _34930_ (.A(net1488),
    .B(_05154_),
    .Y(_05319_));
 NAND3x2_ASAP7_75t_R _34931_ (.B(_05319_),
    .C(_05155_),
    .Y(_05320_),
    .A(_05318_));
 AO21x2_ASAP7_75t_R _34932_ (.A1(_05163_),
    .A2(_05233_),
    .B(_05153_),
    .Y(_05321_));
 AO21x1_ASAP7_75t_R _34933_ (.A1(_05222_),
    .A2(net3449),
    .B(_05153_),
    .Y(_05322_));
 NAND3x2_ASAP7_75t_R _34934_ (.B(_05322_),
    .C(_05168_),
    .Y(_05323_),
    .A(_05321_));
 NOR2x2_ASAP7_75t_R _34935_ (.A(_05320_),
    .B(_05323_),
    .Y(_05324_));
 TAPCELL_ASAP7_75t_R PHY_502 ();
 OR3x2_ASAP7_75t_R _34937_ (.A(_05077_),
    .B(_05196_),
    .C(_00619_),
    .Y(_05326_));
 NAND3x2_ASAP7_75t_R _34938_ (.B(_05306_),
    .C(_05326_),
    .Y(_05327_),
    .A(_05324_));
 NOR2x1_ASAP7_75t_R _34939_ (.A(_05078_),
    .B(_05327_),
    .Y(_05328_));
 NAND2x2_ASAP7_75t_R _34940_ (.A(_00617_),
    .B(_05328_),
    .Y(_05329_));
 AO21x1_ASAP7_75t_R _34941_ (.A1(_05206_),
    .A2(net2314),
    .B(_05208_),
    .Y(_05330_));
 AO21x1_ASAP7_75t_R _34942_ (.A1(net3427),
    .A2(net2137),
    .B(_05208_),
    .Y(_05331_));
 INVx4_ASAP7_75t_R _34943_ (.A(_05208_),
    .Y(_05332_));
 NAND2x1_ASAP7_75t_R _34944_ (.A(_05308_),
    .B(_05332_),
    .Y(_05333_));
 NAND3x1_ASAP7_75t_R _34945_ (.A(_05330_),
    .B(_05331_),
    .C(_05333_),
    .Y(_05334_));
 NAND2x1_ASAP7_75t_R _34946_ (.A(_05073_),
    .B(_05233_),
    .Y(_05335_));
 OAI21x1_ASAP7_75t_R _34947_ (.A1(net3409),
    .A2(_05335_),
    .B(_05199_),
    .Y(_05336_));
 NAND2x2_ASAP7_75t_R _34948_ (.A(net2223),
    .B(_05069_),
    .Y(_05337_));
 AO21x2_ASAP7_75t_R _34949_ (.A1(net3427),
    .A2(net1877),
    .B(_05198_),
    .Y(_05338_));
 AO21x1_ASAP7_75t_R _34950_ (.A1(net3451),
    .A2(net2643),
    .B(_05198_),
    .Y(_05339_));
 NAND3x1_ASAP7_75t_R _34951_ (.A(_05336_),
    .B(_05338_),
    .C(_05339_),
    .Y(_05340_));
 NOR2x1_ASAP7_75t_R _34952_ (.A(_05334_),
    .B(_05340_),
    .Y(_05341_));
 NOR2x1_ASAP7_75t_R _34953_ (.A(_05256_),
    .B(_05206_),
    .Y(_05342_));
 TAPCELL_ASAP7_75t_R PHY_501 ();
 TAPCELL_ASAP7_75t_R PHY_500 ();
 CKINVDCx10_ASAP7_75t_R _34956_ (.A(net1485),
    .Y(_05345_));
 AOI221x1_ASAP7_75t_R _34957_ (.A1(net3436),
    .A2(net3442),
    .B1(_05345_),
    .B2(_05090_),
    .C(_05256_),
    .Y(_05346_));
 NOR2x1_ASAP7_75t_R _34958_ (.A(_05342_),
    .B(_05346_),
    .Y(_05347_));
 OAI21x1_ASAP7_75t_R _34959_ (.A1(_05173_),
    .A2(_05151_),
    .B(_05241_),
    .Y(_05348_));
 NAND2x1_ASAP7_75t_R _34960_ (.A(_05264_),
    .B(_05241_),
    .Y(_05349_));
 AND3x1_ASAP7_75t_R _34961_ (.A(_05348_),
    .B(_05242_),
    .C(_05349_),
    .Y(_05350_));
 NAND2x1_ASAP7_75t_R _34962_ (.A(_05347_),
    .B(_05350_),
    .Y(_05351_));
 INVx1_ASAP7_75t_R _34963_ (.A(_05351_),
    .Y(_05352_));
 NAND2x1_ASAP7_75t_R _34964_ (.A(_05341_),
    .B(_05352_),
    .Y(_05353_));
 TAPCELL_ASAP7_75t_R PHY_499 ();
 AO21x1_ASAP7_75t_R _34966_ (.A1(net1765),
    .A2(net3440),
    .B(net3412),
    .Y(_05355_));
 NOR2x1_ASAP7_75t_R _34967_ (.A(net3412),
    .B(_05095_),
    .Y(_05356_));
 AOI211x1_ASAP7_75t_R _34968_ (.A1(net3436),
    .A2(net1153),
    .B(net3412),
    .C(_05345_),
    .Y(_05357_));
 NOR2x1_ASAP7_75t_R _34969_ (.A(_05356_),
    .B(_05357_),
    .Y(_05358_));
 NAND2x1_ASAP7_75t_R _34970_ (.A(_05355_),
    .B(_05358_),
    .Y(_05359_));
 NAND2x2_ASAP7_75t_R _34971_ (.A(net3438),
    .B(net2226),
    .Y(_05360_));
 TAPCELL_ASAP7_75t_R PHY_498 ();
 AO31x2_ASAP7_75t_R _34973_ (.A1(_05259_),
    .A2(_05360_),
    .A3(net2417),
    .B(_05062_),
    .Y(_05362_));
 NOR2x1_ASAP7_75t_R _34974_ (.A(_05062_),
    .B(_05206_),
    .Y(_05363_));
 TAPCELL_ASAP7_75t_R PHY_497 ();
 AOI211x1_ASAP7_75t_R _34976_ (.A1(net1325),
    .A2(net1153),
    .B(_05062_),
    .C(net2274),
    .Y(_05365_));
 NOR2x1_ASAP7_75t_R _34977_ (.A(_05363_),
    .B(_05365_),
    .Y(_05366_));
 NAND2x1_ASAP7_75t_R _34978_ (.A(_05362_),
    .B(_05366_),
    .Y(_05367_));
 NOR2x2_ASAP7_75t_R _34979_ (.A(_05359_),
    .B(_05367_),
    .Y(_05368_));
 AO21x1_ASAP7_75t_R _34980_ (.A1(_05163_),
    .A2(_05265_),
    .B(net3444),
    .Y(_05369_));
 AOI211x1_ASAP7_75t_R _34981_ (.A1(net1323),
    .A2(net1155),
    .B(net3444),
    .C(net2274),
    .Y(_05370_));
 INVx1_ASAP7_75t_R _34982_ (.A(_05370_),
    .Y(_05371_));
 NAND2x2_ASAP7_75t_R _34983_ (.A(_05369_),
    .B(_05371_),
    .Y(_05372_));
 NOR2x1_ASAP7_75t_R _34984_ (.A(_05345_),
    .B(_05118_),
    .Y(_05373_));
 NAND2x2_ASAP7_75t_R _34985_ (.A(net3445),
    .B(_05373_),
    .Y(_05374_));
 OAI21x1_ASAP7_75t_R _34986_ (.A1(net3457),
    .A2(_05374_),
    .B(_05212_),
    .Y(_05375_));
 AO21x1_ASAP7_75t_R _34987_ (.A1(net2056),
    .A2(_05112_),
    .B(_05138_),
    .Y(_05376_));
 AO21x1_ASAP7_75t_R _34988_ (.A1(_05244_),
    .A2(_05119_),
    .B(_05138_),
    .Y(_05377_));
 NAND2x2_ASAP7_75t_R _34989_ (.A(_05376_),
    .B(_05377_),
    .Y(_05378_));
 NOR3x2_ASAP7_75t_R _34990_ (.B(_05375_),
    .C(_05378_),
    .Y(_05379_),
    .A(_05372_));
 NAND2x2_ASAP7_75t_R _34991_ (.A(_05368_),
    .B(_05379_),
    .Y(_05380_));
 NOR2x2_ASAP7_75t_R _34992_ (.A(_05353_),
    .B(_05380_),
    .Y(_05381_));
 AO21x1_ASAP7_75t_R _34993_ (.A1(net1237),
    .A2(net1523),
    .B(net2529),
    .Y(_05382_));
 AO21x1_ASAP7_75t_R _34994_ (.A1(net2056),
    .A2(_05259_),
    .B(net3455),
    .Y(_05383_));
 NAND2x2_ASAP7_75t_R _34995_ (.A(_05382_),
    .B(_05383_),
    .Y(_05384_));
 AO21x1_ASAP7_75t_R _34996_ (.A1(_05119_),
    .A2(net1894),
    .B(_05086_),
    .Y(_05385_));
 NAND2x2_ASAP7_75t_R _34997_ (.A(_05088_),
    .B(_05385_),
    .Y(_05386_));
 NAND2x1_ASAP7_75t_R _34998_ (.A(net1486),
    .B(_05087_),
    .Y(_05387_));
 NOR2x1_ASAP7_75t_R _34999_ (.A(_05072_),
    .B(_05090_),
    .Y(_05388_));
 NAND2x1_ASAP7_75t_R _35000_ (.A(_05388_),
    .B(_05087_),
    .Y(_05389_));
 OAI21x1_ASAP7_75t_R _35001_ (.A1(_05184_),
    .A2(_05387_),
    .B(_05389_),
    .Y(_05390_));
 NOR3x2_ASAP7_75t_R _35002_ (.B(_05386_),
    .C(_05390_),
    .Y(_05391_),
    .A(_05384_));
 AO21x1_ASAP7_75t_R _35003_ (.A1(net3096),
    .A2(net2027),
    .B(_05107_),
    .Y(_05392_));
 AO21x1_ASAP7_75t_R _35004_ (.A1(net3446),
    .A2(net1894),
    .B(_05107_),
    .Y(_05393_));
 AO21x1_ASAP7_75t_R _35005_ (.A1(net1403),
    .A2(net2645),
    .B(_05107_),
    .Y(_05394_));
 NAND3x1_ASAP7_75t_R _35006_ (.A(_05392_),
    .B(_05393_),
    .C(_05394_),
    .Y(_05395_));
 INVx1_ASAP7_75t_R _35007_ (.A(_05302_),
    .Y(_05396_));
 AO21x1_ASAP7_75t_R _35008_ (.A1(_05157_),
    .A2(net3096),
    .B(_05079_),
    .Y(_05397_));
 NAND2x1_ASAP7_75t_R _35009_ (.A(_05396_),
    .B(_05397_),
    .Y(_05398_));
 AO21x1_ASAP7_75t_R _35010_ (.A1(_05225_),
    .A2(_05165_),
    .B(_05079_),
    .Y(_05399_));
 AO21x1_ASAP7_75t_R _35011_ (.A1(net3369),
    .A2(net1767),
    .B(_05079_),
    .Y(_05400_));
 NAND2x1_ASAP7_75t_R _35012_ (.A(_05400_),
    .B(_05399_),
    .Y(_05401_));
 NOR2x1_ASAP7_75t_R _35013_ (.A(_05398_),
    .B(_05401_),
    .Y(_05402_));
 INVx1_ASAP7_75t_R _35014_ (.A(_05402_),
    .Y(_05403_));
 NOR2x1_ASAP7_75t_R _35015_ (.A(_05403_),
    .B(_05395_),
    .Y(_05404_));
 NAND2x1_ASAP7_75t_R _35016_ (.A(_05391_),
    .B(_05404_),
    .Y(_05405_));
 TAPCELL_ASAP7_75t_R PHY_496 ();
 AOI211x1_ASAP7_75t_R _35018_ (.A1(net3436),
    .A2(_05068_),
    .B(_05153_),
    .C(_05345_),
    .Y(_05407_));
 TAPCELL_ASAP7_75t_R PHY_495 ();
 OA21x2_ASAP7_75t_R _35020_ (.A1(_05178_),
    .A2(_05239_),
    .B(_05154_),
    .Y(_05409_));
 NOR2x2_ASAP7_75t_R _35021_ (.A(_05407_),
    .B(_05409_),
    .Y(_05410_));
 OA21x2_ASAP7_75t_R _35022_ (.A1(_05239_),
    .A2(_05178_),
    .B(_05100_),
    .Y(_05411_));
 AOI211x1_ASAP7_75t_R _35023_ (.A1(net3439),
    .A2(_05068_),
    .B(_05306_),
    .C(net1521),
    .Y(_05412_));
 NOR2x2_ASAP7_75t_R _35024_ (.A(_05411_),
    .B(_05412_),
    .Y(_05413_));
 AO31x2_ASAP7_75t_R _35025_ (.A1(_05131_),
    .A2(_05090_),
    .A3(_05058_),
    .B(_05306_),
    .Y(_05414_));
 NAND3x2_ASAP7_75t_R _35026_ (.B(_05413_),
    .C(_05414_),
    .Y(_05415_),
    .A(_05410_));
 INVx1_ASAP7_75t_R _35027_ (.A(_05415_),
    .Y(_05416_));
 AO21x2_ASAP7_75t_R _35028_ (.A1(net1767),
    .A2(_05073_),
    .B(_05186_),
    .Y(_05417_));
 OAI21x1_ASAP7_75t_R _35029_ (.A1(_05249_),
    .A2(_05106_),
    .B(_05247_),
    .Y(_05418_));
 NAND3x2_ASAP7_75t_R _35030_ (.B(_05418_),
    .C(_05246_),
    .Y(_05419_),
    .A(_05417_));
 INVx3_ASAP7_75t_R _35031_ (.A(_05215_),
    .Y(_05420_));
 OA21x2_ASAP7_75t_R _35032_ (.A1(_05123_),
    .A2(_05084_),
    .B(_05420_),
    .Y(_05421_));
 NOR2x2_ASAP7_75t_R _35033_ (.A(net1303),
    .B(_05345_),
    .Y(_05422_));
 OA31x2_ASAP7_75t_R _35034_ (.A1(_05422_),
    .A2(_05173_),
    .A3(_05151_),
    .B1(_05420_),
    .Y(_05423_));
 NOR3x1_ASAP7_75t_R _35035_ (.A(_05419_),
    .B(_05421_),
    .C(_05423_),
    .Y(_05424_));
 NAND2x1_ASAP7_75t_R _35036_ (.A(_05416_),
    .B(_05424_),
    .Y(_05425_));
 NOR2x2_ASAP7_75t_R _35037_ (.A(_05425_),
    .B(_05405_),
    .Y(_05426_));
 NAND2x2_ASAP7_75t_R _35038_ (.A(_05381_),
    .B(_05426_),
    .Y(_05427_));
 NAND3x2_ASAP7_75t_R _35039_ (.B(net3428),
    .C(net3114),
    .Y(_05428_),
    .A(_05317_));
 AOI21x1_ASAP7_75t_R _35040_ (.A1(net3428),
    .A2(_05317_),
    .B(net3114),
    .Y(_05429_));
 INVx2_ASAP7_75t_R _35041_ (.A(_05429_),
    .Y(_05430_));
 TAPCELL_ASAP7_75t_R PHY_494 ();
 NAND2x2_ASAP7_75t_R _35043_ (.A(_00579_),
    .B(net3112),
    .Y(_05432_));
 TAPCELL_ASAP7_75t_R PHY_493 ();
 NAND2x2_ASAP7_75t_R _35045_ (.A(net2114),
    .B(_00578_),
    .Y(_05434_));
 NOR2x2_ASAP7_75t_R _35046_ (.A(_05432_),
    .B(_05434_),
    .Y(_05435_));
 TAPCELL_ASAP7_75t_R PHY_492 ();
 TAPCELL_ASAP7_75t_R PHY_491 ();
 TAPCELL_ASAP7_75t_R PHY_490 ();
 INVx4_ASAP7_75t_R _35050_ (.A(net2726),
    .Y(_05439_));
 NAND2x2_ASAP7_75t_R _35051_ (.A(net2711),
    .B(_05439_),
    .Y(_05440_));
 NOR2x2_ASAP7_75t_R _35052_ (.A(net1314),
    .B(_05440_),
    .Y(_05441_));
 TAPCELL_ASAP7_75t_R PHY_489 ();
 CKINVDCx20_ASAP7_75t_R _35054_ (.A(net1310),
    .Y(_05443_));
 NOR2x2_ASAP7_75t_R _35055_ (.A(net1200),
    .B(_05443_),
    .Y(_05444_));
 INVx2_ASAP7_75t_R _35056_ (.A(_00582_),
    .Y(_05445_));
 NOR2x2_ASAP7_75t_R _35057_ (.A(net2726),
    .B(_05445_),
    .Y(_05446_));
 NAND2x2_ASAP7_75t_R _35058_ (.A(_05444_),
    .B(_05446_),
    .Y(_05447_));
 TAPCELL_ASAP7_75t_R PHY_488 ();
 NAND2x2_ASAP7_75t_R _35060_ (.A(net1310),
    .B(net1203),
    .Y(_05449_));
 INVx5_ASAP7_75t_R _35061_ (.A(_05449_),
    .Y(_05450_));
 NAND2x2_ASAP7_75t_R _35062_ (.A(_05446_),
    .B(_05450_),
    .Y(_05451_));
 TAPCELL_ASAP7_75t_R PHY_487 ();
 INVx8_ASAP7_75t_R _35064_ (.A(_05435_),
    .Y(_05453_));
 AOI21x1_ASAP7_75t_R _35065_ (.A1(_05447_),
    .A2(net3113),
    .B(_05453_),
    .Y(_05454_));
 NOR2x2_ASAP7_75t_R _35066_ (.A(net2726),
    .B(net2711),
    .Y(_05455_));
 TAPCELL_ASAP7_75t_R PHY_486 ();
 CKINVDCx20_ASAP7_75t_R _35068_ (.A(net1034),
    .Y(_05457_));
 NOR2x2_ASAP7_75t_R _35069_ (.A(_05457_),
    .B(_05453_),
    .Y(_05458_));
 AOI211x1_ASAP7_75t_R _35070_ (.A1(_05435_),
    .A2(_05441_),
    .B(_05454_),
    .C(_05458_),
    .Y(_05459_));
 NAND2x2_ASAP7_75t_R _35071_ (.A(net2726),
    .B(_00582_),
    .Y(_05460_));
 CKINVDCx6p67_ASAP7_75t_R _35072_ (.A(net1205),
    .Y(_05461_));
 NAND2x2_ASAP7_75t_R _35073_ (.A(_05444_),
    .B(_05461_),
    .Y(_05462_));
 NOR2x2_ASAP7_75t_R _35074_ (.A(net1311),
    .B(net1208),
    .Y(_05463_));
 INVx4_ASAP7_75t_R _35075_ (.A(_05463_),
    .Y(_05464_));
 AO21x1_ASAP7_75t_R _35076_ (.A1(_05462_),
    .A2(_05464_),
    .B(_05453_),
    .Y(_05465_));
 NOR2x2_ASAP7_75t_R _35077_ (.A(net2711),
    .B(_05439_),
    .Y(_05466_));
 NAND2x2_ASAP7_75t_R _35078_ (.A(net2016),
    .B(_05435_),
    .Y(_05467_));
 AND2x2_ASAP7_75t_R _35079_ (.A(_05465_),
    .B(_05467_),
    .Y(_05468_));
 INVx2_ASAP7_75t_R _35080_ (.A(_00579_),
    .Y(_05469_));
 NOR2x2_ASAP7_75t_R _35081_ (.A(net3112),
    .B(_05469_),
    .Y(_05470_));
 INVx3_ASAP7_75t_R _35082_ (.A(_05434_),
    .Y(_05471_));
 NAND2x2_ASAP7_75t_R _35083_ (.A(_05470_),
    .B(_05471_),
    .Y(_05472_));
 TAPCELL_ASAP7_75t_R PHY_485 ();
 NAND3x2_ASAP7_75t_R _35085_ (.B(_05468_),
    .C(_05472_),
    .Y(_05474_),
    .A(_05459_));
 INVx2_ASAP7_75t_R _35086_ (.A(net2110),
    .Y(_05475_));
 NOR2x2_ASAP7_75t_R _35087_ (.A(_00578_),
    .B(_05475_),
    .Y(_05476_));
 AND3x2_ASAP7_75t_R _35088_ (.A(_05469_),
    .B(net2110),
    .C(_00578_),
    .Y(_05477_));
 NOR3x2_ASAP7_75t_R _35089_ (.B(_05476_),
    .C(_05477_),
    .Y(_05478_),
    .A(_05474_));
 NAND2x2_ASAP7_75t_R _35090_ (.A(net2112),
    .B(_05478_),
    .Y(_05479_));
 INVx2_ASAP7_75t_R _35091_ (.A(_00578_),
    .Y(_05480_));
 NAND2x2_ASAP7_75t_R _35092_ (.A(net2110),
    .B(_05480_),
    .Y(_05481_));
 INVx2_ASAP7_75t_R _35093_ (.A(net3112),
    .Y(_05482_));
 NAND2x2_ASAP7_75t_R _35094_ (.A(net3122),
    .B(_05482_),
    .Y(_05483_));
 NOR2x2_ASAP7_75t_R _35095_ (.A(_05481_),
    .B(_05483_),
    .Y(_05484_));
 NOR2x2_ASAP7_75t_R _35096_ (.A(net1310),
    .B(net1201),
    .Y(_05485_));
 NAND2x2_ASAP7_75t_R _35097_ (.A(net1034),
    .B(_05485_),
    .Y(_05486_));
 INVx1_ASAP7_75t_R _35098_ (.A(_05486_),
    .Y(_05487_));
 NAND2x1_ASAP7_75t_R _35099_ (.A(_05484_),
    .B(_05487_),
    .Y(_05488_));
 TAPCELL_ASAP7_75t_R PHY_484 ();
 NAND2x2_ASAP7_75t_R _35101_ (.A(net2670),
    .B(_05446_),
    .Y(_05490_));
 TAPCELL_ASAP7_75t_R PHY_483 ();
 NAND2x2_ASAP7_75t_R _35103_ (.A(_05476_),
    .B(_05470_),
    .Y(_05492_));
 AO21x1_ASAP7_75t_R _35104_ (.A1(_05447_),
    .A2(net2548),
    .B(_05492_),
    .Y(_05493_));
 NAND2x1_ASAP7_75t_R _35105_ (.A(_05488_),
    .B(_05493_),
    .Y(_05494_));
 NOR2x2_ASAP7_75t_R _35106_ (.A(_05443_),
    .B(net1205),
    .Y(_05495_));
 CKINVDCx5p33_ASAP7_75t_R _35107_ (.A(_05495_),
    .Y(_05496_));
 NAND2x2_ASAP7_75t_R _35108_ (.A(net2863),
    .B(_05461_),
    .Y(_05497_));
 TAPCELL_ASAP7_75t_R PHY_482 ();
 AO21x1_ASAP7_75t_R _35110_ (.A1(_05496_),
    .A2(net2815),
    .B(_05492_),
    .Y(_05499_));
 CKINVDCx16_ASAP7_75t_R _35111_ (.A(net1201),
    .Y(_05500_));
 NOR2x2_ASAP7_75t_R _35112_ (.A(net1310),
    .B(_05500_),
    .Y(_05501_));
 NAND2x2_ASAP7_75t_R _35113_ (.A(_05501_),
    .B(_05466_),
    .Y(_05502_));
 NAND2x2_ASAP7_75t_R _35114_ (.A(_05485_),
    .B(_05466_),
    .Y(_05503_));
 TAPCELL_ASAP7_75t_R PHY_481 ();
 AO21x1_ASAP7_75t_R _35116_ (.A1(net2153),
    .A2(_05503_),
    .B(_05492_),
    .Y(_05505_));
 NAND2x1_ASAP7_75t_R _35117_ (.A(_05505_),
    .B(_05499_),
    .Y(_05506_));
 NOR2x1_ASAP7_75t_R _35118_ (.A(_05494_),
    .B(_05506_),
    .Y(_05507_));
 NAND2x2_ASAP7_75t_R _35119_ (.A(net3463),
    .B(_05450_),
    .Y(_05508_));
 TAPCELL_ASAP7_75t_R PHY_480 ();
 NOR2x2_ASAP7_75t_R _35121_ (.A(_05432_),
    .B(_05481_),
    .Y(_05510_));
 INVx2_ASAP7_75t_R _35122_ (.A(net3373),
    .Y(_05511_));
 AO21x1_ASAP7_75t_R _35123_ (.A1(net2870),
    .A2(_05496_),
    .B(_05511_),
    .Y(_05512_));
 NAND2x2_ASAP7_75t_R _35124_ (.A(net1311),
    .B(_05500_),
    .Y(_05513_));
 NOR2x2_ASAP7_75t_R _35125_ (.A(_05513_),
    .B(_05440_),
    .Y(_05514_));
 NAND2x2_ASAP7_75t_R _35126_ (.A(net1201),
    .B(_05443_),
    .Y(_05515_));
 NOR2x2_ASAP7_75t_R _35127_ (.A(net3458),
    .B(_05457_),
    .Y(_05516_));
 TAPCELL_ASAP7_75t_R PHY_479 ();
 OAI21x1_ASAP7_75t_R _35129_ (.A1(_05514_),
    .A2(_05516_),
    .B(net3373),
    .Y(_05518_));
 INVx3_ASAP7_75t_R _35130_ (.A(_05485_),
    .Y(_05519_));
 NOR2x2_ASAP7_75t_R _35131_ (.A(_05440_),
    .B(_05519_),
    .Y(_05520_));
 TAPCELL_ASAP7_75t_R PHY_478 ();
 NOR2x2_ASAP7_75t_R _35133_ (.A(net3110),
    .B(_05457_),
    .Y(_05522_));
 OAI21x1_ASAP7_75t_R _35134_ (.A1(net2810),
    .A2(_05522_),
    .B(net3373),
    .Y(_05523_));
 AND3x1_ASAP7_75t_R _35135_ (.A(_05512_),
    .B(_05518_),
    .C(_05523_),
    .Y(_05524_));
 NAND2x1_ASAP7_75t_R _35136_ (.A(_05507_),
    .B(_05524_),
    .Y(_05525_));
 TAPCELL_ASAP7_75t_R PHY_477 ();
 NOR2x2_ASAP7_75t_R _35138_ (.A(_00579_),
    .B(net3112),
    .Y(_05527_));
 NAND2x2_ASAP7_75t_R _35139_ (.A(_05527_),
    .B(_05476_),
    .Y(_05528_));
 TAPCELL_ASAP7_75t_R PHY_476 ();
 NAND2x2_ASAP7_75t_R _35141_ (.A(net1031),
    .B(_05501_),
    .Y(_05530_));
 TAPCELL_ASAP7_75t_R PHY_475 ();
 NAND2x2_ASAP7_75t_R _35143_ (.A(_05455_),
    .B(_05444_),
    .Y(_05532_));
 AO21x1_ASAP7_75t_R _35144_ (.A1(net2036),
    .A2(net1084),
    .B(net2755),
    .Y(_05533_));
 OAI21x1_ASAP7_75t_R _35145_ (.A1(net1124),
    .A2(net2755),
    .B(_05533_),
    .Y(_05534_));
 NAND2x2_ASAP7_75t_R _35146_ (.A(_05444_),
    .B(_05466_),
    .Y(_05535_));
 TAPCELL_ASAP7_75t_R PHY_474 ();
 AO21x1_ASAP7_75t_R _35148_ (.A1(net3462),
    .A2(_05503_),
    .B(net2740),
    .Y(_05537_));
 TAPCELL_ASAP7_75t_R PHY_473 ();
 TAPCELL_ASAP7_75t_R PHY_472 ();
 AOI211x1_ASAP7_75t_R _35151_ (.A1(net2814),
    .A2(net989),
    .B(net2755),
    .C(net1210),
    .Y(_05540_));
 INVx1_ASAP7_75t_R _35152_ (.A(_05540_),
    .Y(_05541_));
 NAND2x1_ASAP7_75t_R _35153_ (.A(_05537_),
    .B(_05541_),
    .Y(_05542_));
 NOR2x1_ASAP7_75t_R _35154_ (.A(_05534_),
    .B(_05542_),
    .Y(_05543_));
 NAND2x2_ASAP7_75t_R _35155_ (.A(net3112),
    .B(_05469_),
    .Y(_05544_));
 NOR2x2_ASAP7_75t_R _35156_ (.A(_05481_),
    .B(_05544_),
    .Y(_05545_));
 TAPCELL_ASAP7_75t_R PHY_471 ();
 NOR2x2_ASAP7_75t_R _35158_ (.A(_00579_),
    .B(_05482_),
    .Y(_05547_));
 NAND2x2_ASAP7_75t_R _35159_ (.A(_05476_),
    .B(_05547_),
    .Y(_05548_));
 TAPCELL_ASAP7_75t_R PHY_470 ();
 NOR2x1_ASAP7_75t_R _35161_ (.A(_05462_),
    .B(_05548_),
    .Y(_05550_));
 NOR2x1_ASAP7_75t_R _35162_ (.A(_05548_),
    .B(net2815),
    .Y(_05551_));
 AOI211x1_ASAP7_75t_R _35163_ (.A1(net2017),
    .A2(_05545_),
    .B(_05550_),
    .C(_05551_),
    .Y(_05552_));
 NOR2x1_ASAP7_75t_R _35164_ (.A(net2036),
    .B(_05548_),
    .Y(_05553_));
 TAPCELL_ASAP7_75t_R PHY_469 ();
 AOI211x1_ASAP7_75t_R _35166_ (.A1(net3110),
    .A2(net989),
    .B(_05548_),
    .C(net2091),
    .Y(_05555_));
 NOR2x1_ASAP7_75t_R _35167_ (.A(_05553_),
    .B(_05555_),
    .Y(_05556_));
 AND2x2_ASAP7_75t_R _35168_ (.A(_05556_),
    .B(_05552_),
    .Y(_05557_));
 NAND2x1_ASAP7_75t_R _35169_ (.A(_05557_),
    .B(_05543_),
    .Y(_05558_));
 NOR2x1_ASAP7_75t_R _35170_ (.A(_05525_),
    .B(_05558_),
    .Y(_05559_));
 NAND2x2_ASAP7_75t_R _35171_ (.A(net2726),
    .B(_05445_),
    .Y(_05560_));
 NOR2x2_ASAP7_75t_R _35172_ (.A(_05515_),
    .B(_05560_),
    .Y(_05561_));
 TAPCELL_ASAP7_75t_R PHY_468 ();
 NAND2x2_ASAP7_75t_R _35174_ (.A(_05527_),
    .B(_05471_),
    .Y(_05563_));
 INVx3_ASAP7_75t_R _35175_ (.A(net2389),
    .Y(_05564_));
 NAND2x1_ASAP7_75t_R _35176_ (.A(net1528),
    .B(_05564_),
    .Y(_05565_));
 NOR2x2_ASAP7_75t_R _35177_ (.A(_05515_),
    .B(net1207),
    .Y(_05566_));
 TAPCELL_ASAP7_75t_R PHY_467 ();
 NOR2x2_ASAP7_75t_R _35179_ (.A(net1202),
    .B(net1212),
    .Y(_05568_));
 OAI21x1_ASAP7_75t_R _35180_ (.A1(_05566_),
    .A2(_05568_),
    .B(_05564_),
    .Y(_05569_));
 NAND2x1_ASAP7_75t_R _35181_ (.A(_05565_),
    .B(_05569_),
    .Y(_05570_));
 TAPCELL_ASAP7_75t_R PHY_466 ();
 NOR2x2_ASAP7_75t_R _35183_ (.A(net2389),
    .B(net3113),
    .Y(_05572_));
 TAPCELL_ASAP7_75t_R PHY_465 ();
 TAPCELL_ASAP7_75t_R PHY_464 ();
 AOI211x1_ASAP7_75t_R _35186_ (.A1(net2814),
    .A2(net989),
    .B(net2389),
    .C(_05457_),
    .Y(_05575_));
 NOR3x1_ASAP7_75t_R _35187_ (.A(_05570_),
    .B(_05572_),
    .C(_05575_),
    .Y(_05576_));
 NOR2x2_ASAP7_75t_R _35188_ (.A(net3116),
    .B(_05544_),
    .Y(_05577_));
 OAI21x1_ASAP7_75t_R _35189_ (.A1(_05441_),
    .A2(_05514_),
    .B(_05577_),
    .Y(_05578_));
 NAND2x2_ASAP7_75t_R _35190_ (.A(net1031),
    .B(_05450_),
    .Y(_05579_));
 NAND2x2_ASAP7_75t_R _35191_ (.A(_05443_),
    .B(net1034),
    .Y(_05580_));
 NAND2x2_ASAP7_75t_R _35192_ (.A(_05547_),
    .B(_05471_),
    .Y(_05581_));
 TAPCELL_ASAP7_75t_R PHY_463 ();
 AO21x1_ASAP7_75t_R _35194_ (.A1(net2833),
    .A2(net3115),
    .B(_05581_),
    .Y(_05583_));
 NAND2x1_ASAP7_75t_R _35195_ (.A(_05578_),
    .B(_05583_),
    .Y(_05584_));
 AO21x1_ASAP7_75t_R _35196_ (.A1(_05535_),
    .A2(net1771),
    .B(_05581_),
    .Y(_05585_));
 AOI211x1_ASAP7_75t_R _35197_ (.A1(net3110),
    .A2(_05500_),
    .B(_05581_),
    .C(net1208),
    .Y(_05586_));
 INVx1_ASAP7_75t_R _35198_ (.A(_05586_),
    .Y(_05587_));
 NAND2x1_ASAP7_75t_R _35199_ (.A(_05585_),
    .B(_05587_),
    .Y(_05588_));
 NOR2x1_ASAP7_75t_R _35200_ (.A(_05584_),
    .B(_05588_),
    .Y(_05589_));
 NAND2x1_ASAP7_75t_R _35201_ (.A(_05576_),
    .B(_05589_),
    .Y(_05590_));
 NAND2x1_ASAP7_75t_R _35202_ (.A(_05463_),
    .B(_05435_),
    .Y(_05591_));
 INVx1_ASAP7_75t_R _35203_ (.A(_05591_),
    .Y(_05592_));
 TAPCELL_ASAP7_75t_R PHY_462 ();
 TAPCELL_ASAP7_75t_R PHY_461 ();
 TAPCELL_ASAP7_75t_R PHY_460 ();
 OAI22x1_ASAP7_75t_R _35207_ (.A1(_05467_),
    .A2(net1000),
    .B1(net1627),
    .B2(_05453_),
    .Y(_05596_));
 NOR2x1_ASAP7_75t_R _35208_ (.A(_05592_),
    .B(_05596_),
    .Y(_05597_));
 NOR2x2_ASAP7_75t_R _35209_ (.A(net2243),
    .B(_05501_),
    .Y(_05598_));
 NOR2x2_ASAP7_75t_R _35210_ (.A(net2090),
    .B(_05472_),
    .Y(_05599_));
 NOR2x2_ASAP7_75t_R _35211_ (.A(net3117),
    .B(_05483_),
    .Y(_05600_));
 NAND2x1_ASAP7_75t_R _35212_ (.A(_05466_),
    .B(_05600_),
    .Y(_05601_));
 NAND2x1_ASAP7_75t_R _35213_ (.A(_05463_),
    .B(_05600_),
    .Y(_05602_));
 OAI21x1_ASAP7_75t_R _35214_ (.A1(_05598_),
    .A2(_05601_),
    .B(_05602_),
    .Y(_05603_));
 AOI21x1_ASAP7_75t_R _35215_ (.A1(_05598_),
    .A2(_05599_),
    .B(_05603_),
    .Y(_05604_));
 NAND2x2_ASAP7_75t_R _35216_ (.A(net3121),
    .B(_05446_),
    .Y(_05605_));
 TAPCELL_ASAP7_75t_R PHY_459 ();
 AO21x1_ASAP7_75t_R _35218_ (.A1(net2191),
    .A2(_05605_),
    .B(_05453_),
    .Y(_05607_));
 AO21x1_ASAP7_75t_R _35219_ (.A1(net2032),
    .A2(net1085),
    .B(_05453_),
    .Y(_05608_));
 AND2x2_ASAP7_75t_R _35220_ (.A(_05607_),
    .B(_05608_),
    .Y(_05609_));
 NAND3x1_ASAP7_75t_R _35221_ (.A(_05597_),
    .B(_05604_),
    .C(_05609_),
    .Y(_05610_));
 NOR2x1_ASAP7_75t_R _35222_ (.A(_05590_),
    .B(_05610_),
    .Y(_05611_));
 NAND2x1_ASAP7_75t_R _35223_ (.A(_05559_),
    .B(_05611_),
    .Y(_05612_));
 NAND2x2_ASAP7_75t_R _35224_ (.A(net2318),
    .B(_05461_),
    .Y(_05613_));
 TAPCELL_ASAP7_75t_R PHY_458 ();
 NOR2x2_ASAP7_75t_R _35226_ (.A(_00578_),
    .B(net2110),
    .Y(_05615_));
 NAND2x2_ASAP7_75t_R _35227_ (.A(_05615_),
    .B(_05470_),
    .Y(_05616_));
 TAPCELL_ASAP7_75t_R PHY_457 ();
 AO21x1_ASAP7_75t_R _35229_ (.A1(net1627),
    .A2(_05613_),
    .B(net2447),
    .Y(_05618_));
 NAND2x2_ASAP7_75t_R _35230_ (.A(net1310),
    .B(_05446_),
    .Y(_05619_));
 TAPCELL_ASAP7_75t_R PHY_456 ();
 AO21x1_ASAP7_75t_R _35232_ (.A1(net2400),
    .A2(_05605_),
    .B(net2447),
    .Y(_05621_));
 TAPCELL_ASAP7_75t_R PHY_455 ();
 AO21x1_ASAP7_75t_R _35234_ (.A1(net2034),
    .A2(net2611),
    .B(net2447),
    .Y(_05623_));
 AND3x1_ASAP7_75t_R _35235_ (.A(_05618_),
    .B(_05621_),
    .C(_05623_),
    .Y(_05624_));
 INVx2_ASAP7_75t_R _35236_ (.A(_05432_),
    .Y(_05625_));
 NAND2x2_ASAP7_75t_R _35237_ (.A(_05615_),
    .B(_05625_),
    .Y(_05626_));
 INVx3_ASAP7_75t_R _35238_ (.A(_05626_),
    .Y(_05627_));
 TAPCELL_ASAP7_75t_R PHY_454 ();
 TAPCELL_ASAP7_75t_R PHY_453 ();
 AOI211x1_ASAP7_75t_R _35241_ (.A1(net2814),
    .A2(net3098),
    .B(_05626_),
    .C(_05457_),
    .Y(_05630_));
 OA21x2_ASAP7_75t_R _35242_ (.A1(net2661),
    .A2(net2810),
    .B(_05627_),
    .Y(_05631_));
 AOI211x1_ASAP7_75t_R _35243_ (.A1(_05566_),
    .A2(_05627_),
    .B(_05630_),
    .C(_05631_),
    .Y(_05632_));
 NAND2x1_ASAP7_75t_R _35244_ (.A(_05624_),
    .B(_05632_),
    .Y(_05633_));
 NAND2x2_ASAP7_75t_R _35245_ (.A(_05527_),
    .B(_05615_),
    .Y(_05634_));
 AO21x1_ASAP7_75t_R _35246_ (.A1(_05462_),
    .A2(_05464_),
    .B(net2461),
    .Y(_05635_));
 NOR2x1_ASAP7_75t_R _35247_ (.A(net2461),
    .B(net3250),
    .Y(_05636_));
 INVx1_ASAP7_75t_R _35248_ (.A(_05636_),
    .Y(_05637_));
 AO21x1_ASAP7_75t_R _35249_ (.A1(net2032),
    .A2(_05440_),
    .B(net2461),
    .Y(_05638_));
 AND3x1_ASAP7_75t_R _35250_ (.A(_05635_),
    .B(_05637_),
    .C(_05638_),
    .Y(_05639_));
 NAND2x2_ASAP7_75t_R _35251_ (.A(_05615_),
    .B(_05547_),
    .Y(_05640_));
 AO21x1_ASAP7_75t_R _35252_ (.A1(net2703),
    .A2(net2870),
    .B(net2618),
    .Y(_05641_));
 NOR2x2_ASAP7_75t_R _35253_ (.A(_05449_),
    .B(net1208),
    .Y(_05642_));
 INVx6_ASAP7_75t_R _35254_ (.A(_05642_),
    .Y(_05643_));
 AO21x1_ASAP7_75t_R _35255_ (.A1(net3350),
    .A2(net2509),
    .B(net2618),
    .Y(_05644_));
 NAND2x1_ASAP7_75t_R _35256_ (.A(_05641_),
    .B(_05644_),
    .Y(_05645_));
 NOR2x2_ASAP7_75t_R _35257_ (.A(net1204),
    .B(_05457_),
    .Y(_05646_));
 INVx3_ASAP7_75t_R _35258_ (.A(_05640_),
    .Y(_05647_));
 NOR2x1_ASAP7_75t_R _35259_ (.A(_05440_),
    .B(_05640_),
    .Y(_05648_));
 AO22x1_ASAP7_75t_R _35260_ (.A1(_05646_),
    .A2(_05647_),
    .B1(_05648_),
    .B2(_05513_),
    .Y(_05649_));
 NOR2x1_ASAP7_75t_R _35261_ (.A(_05645_),
    .B(_05649_),
    .Y(_05650_));
 NAND2x1_ASAP7_75t_R _35262_ (.A(_05639_),
    .B(_05650_),
    .Y(_05651_));
 NOR2x1_ASAP7_75t_R _35263_ (.A(_05633_),
    .B(_05651_),
    .Y(_05652_));
 NOR2x2_ASAP7_75t_R _35264_ (.A(net2110),
    .B(_05480_),
    .Y(_05653_));
 NAND2x2_ASAP7_75t_R _35265_ (.A(_05653_),
    .B(_05470_),
    .Y(_05654_));
 NOR2x2_ASAP7_75t_R _35266_ (.A(_05457_),
    .B(_05654_),
    .Y(_05655_));
 NOR2x2_ASAP7_75t_R _35267_ (.A(net1209),
    .B(_05513_),
    .Y(_05656_));
 INVx2_ASAP7_75t_R _35268_ (.A(_05654_),
    .Y(_05657_));
 OA21x2_ASAP7_75t_R _35269_ (.A1(_05656_),
    .A2(_05566_),
    .B(_05657_),
    .Y(_05658_));
 AO21x1_ASAP7_75t_R _35270_ (.A1(net2814),
    .A2(_05655_),
    .B(_05658_),
    .Y(_05659_));
 NAND2x2_ASAP7_75t_R _35271_ (.A(net3384),
    .B(_05475_),
    .Y(_05660_));
 NOR2x2_ASAP7_75t_R _35272_ (.A(_05432_),
    .B(_05660_),
    .Y(_05661_));
 TAPCELL_ASAP7_75t_R PHY_452 ();
 OA21x2_ASAP7_75t_R _35274_ (.A1(net2809),
    .A2(net2661),
    .B(_05661_),
    .Y(_05663_));
 INVx8_ASAP7_75t_R _35275_ (.A(net2611),
    .Y(_05664_));
 INVx2_ASAP7_75t_R _35276_ (.A(_05580_),
    .Y(_05665_));
 OA21x2_ASAP7_75t_R _35277_ (.A1(_05664_),
    .A2(_05665_),
    .B(_05661_),
    .Y(_05666_));
 NOR2x1_ASAP7_75t_R _35278_ (.A(_05663_),
    .B(_05666_),
    .Y(_05667_));
 TAPCELL_ASAP7_75t_R PHY_451 ();
 NOR2x2_ASAP7_75t_R _35280_ (.A(net1673),
    .B(net2319),
    .Y(_05669_));
 OA21x2_ASAP7_75t_R _35281_ (.A1(_05566_),
    .A2(_05642_),
    .B(_05661_),
    .Y(_05670_));
 AOI21x1_ASAP7_75t_R _35282_ (.A1(_05661_),
    .A2(_05669_),
    .B(_05670_),
    .Y(_05671_));
 NAND2x1_ASAP7_75t_R _35283_ (.A(_05667_),
    .B(_05671_),
    .Y(_05672_));
 NOR2x1_ASAP7_75t_R _35284_ (.A(_05659_),
    .B(_05672_),
    .Y(_05673_));
 NOR2x2_ASAP7_75t_R _35285_ (.A(net3120),
    .B(net1666),
    .Y(_05674_));
 NOR2x2_ASAP7_75t_R _35286_ (.A(_05660_),
    .B(_05544_),
    .Y(_05675_));
 NAND2x2_ASAP7_75t_R _35287_ (.A(net1032),
    .B(net3459),
    .Y(_05676_));
 NAND2x2_ASAP7_75t_R _35288_ (.A(_05653_),
    .B(_05547_),
    .Y(_05677_));
 TAPCELL_ASAP7_75t_R PHY_450 ();
 AO21x1_ASAP7_75t_R _35290_ (.A1(net2698),
    .A2(_05676_),
    .B(_05677_),
    .Y(_05679_));
 INVx1_ASAP7_75t_R _35291_ (.A(_05679_),
    .Y(_05680_));
 AO21x1_ASAP7_75t_R _35292_ (.A1(_05674_),
    .A2(_05675_),
    .B(_05680_),
    .Y(_05681_));
 INVx3_ASAP7_75t_R _35293_ (.A(_05579_),
    .Y(_05682_));
 NAND2x2_ASAP7_75t_R _35294_ (.A(_05527_),
    .B(_05653_),
    .Y(_05683_));
 INVx4_ASAP7_75t_R _35295_ (.A(_05683_),
    .Y(_05684_));
 NAND2x2_ASAP7_75t_R _35296_ (.A(net3109),
    .B(_05461_),
    .Y(_05685_));
 INVx1_ASAP7_75t_R _35297_ (.A(_05685_),
    .Y(_05686_));
 OA21x2_ASAP7_75t_R _35298_ (.A1(_05686_),
    .A2(_05669_),
    .B(_05684_),
    .Y(_05687_));
 AO21x1_ASAP7_75t_R _35299_ (.A1(_05682_),
    .A2(_05684_),
    .B(_05687_),
    .Y(_05688_));
 NOR2x1_ASAP7_75t_R _35300_ (.A(_05681_),
    .B(_05688_),
    .Y(_05689_));
 AND2x2_ASAP7_75t_R _35301_ (.A(_05673_),
    .B(_05689_),
    .Y(_05690_));
 NAND2x2_ASAP7_75t_R _35302_ (.A(_05652_),
    .B(_05690_),
    .Y(_05691_));
 NOR2x2_ASAP7_75t_R _35303_ (.A(_05612_),
    .B(_05691_),
    .Y(_05692_));
 NAND2x2_ASAP7_75t_R _35304_ (.A(_05479_),
    .B(_05692_),
    .Y(_05693_));
 INVx2_ASAP7_75t_R _35305_ (.A(_05693_),
    .Y(_05695_));
 AO21x1_ASAP7_75t_R _35306_ (.A1(_05428_),
    .A2(_05430_),
    .B(_05695_),
    .Y(_05696_));
 INVx1_ASAP7_75t_R _35307_ (.A(_05395_),
    .Y(_05697_));
 NAND2x1_ASAP7_75t_R _35308_ (.A(_05402_),
    .B(_05697_),
    .Y(_05698_));
 INVx1_ASAP7_75t_R _35309_ (.A(_05391_),
    .Y(_05699_));
 NOR2x2_ASAP7_75t_R _35310_ (.A(_05698_),
    .B(_05699_),
    .Y(_05700_));
 INVx1_ASAP7_75t_R _35311_ (.A(_05419_),
    .Y(_05701_));
 NOR2x1_ASAP7_75t_R _35312_ (.A(_05421_),
    .B(_05423_),
    .Y(_05702_));
 NAND2x1_ASAP7_75t_R _35313_ (.A(_05701_),
    .B(_05702_),
    .Y(_05703_));
 NOR2x1_ASAP7_75t_R _35314_ (.A(_05415_),
    .B(_05703_),
    .Y(_05704_));
 NAND2x2_ASAP7_75t_R _35315_ (.A(_05700_),
    .B(_05704_),
    .Y(_05706_));
 INVx1_ASAP7_75t_R _35316_ (.A(_05378_),
    .Y(_05707_));
 NOR2x1_ASAP7_75t_R _35317_ (.A(_05375_),
    .B(_05372_),
    .Y(_05708_));
 NAND2x1_ASAP7_75t_R _35318_ (.A(_05707_),
    .B(_05708_),
    .Y(_05709_));
 INVx1_ASAP7_75t_R _35319_ (.A(_05368_),
    .Y(_05710_));
 NOR2x2_ASAP7_75t_R _35320_ (.A(_05709_),
    .B(_05710_),
    .Y(_05711_));
 INVx1_ASAP7_75t_R _35321_ (.A(_05341_),
    .Y(_05712_));
 NOR2x1_ASAP7_75t_R _35322_ (.A(_05351_),
    .B(_05712_),
    .Y(_05713_));
 NAND2x2_ASAP7_75t_R _35323_ (.A(_05711_),
    .B(_05713_),
    .Y(_05714_));
 NOR2x2_ASAP7_75t_R _35324_ (.A(_05706_),
    .B(_05714_),
    .Y(_05715_));
 NOR3x2_ASAP7_75t_R _35325_ (.B(_05077_),
    .C(_05196_),
    .Y(_05717_),
    .A(_05327_));
 NOR3x2_ASAP7_75t_R _35326_ (.B(_05230_),
    .C(_05195_),
    .Y(_05718_),
    .A(_05148_));
 INVx1_ASAP7_75t_R _35327_ (.A(_05281_),
    .Y(_05719_));
 NOR2x1_ASAP7_75t_R _35328_ (.A(_05288_),
    .B(_05719_),
    .Y(_05720_));
 INVx1_ASAP7_75t_R _35329_ (.A(_05305_),
    .Y(_05721_));
 NAND2x1_ASAP7_75t_R _35330_ (.A(_05311_),
    .B(_05721_),
    .Y(_05722_));
 NOR2x1_ASAP7_75t_R _35331_ (.A(_05297_),
    .B(_05722_),
    .Y(_05723_));
 NAND2x1_ASAP7_75t_R _35332_ (.A(_05720_),
    .B(_05723_),
    .Y(_05724_));
 NOR2x2_ASAP7_75t_R _35333_ (.A(_05269_),
    .B(_05724_),
    .Y(_05725_));
 NAND2x2_ASAP7_75t_R _35334_ (.A(_05718_),
    .B(_05725_),
    .Y(_05726_));
 NOR2x2_ASAP7_75t_R _35335_ (.A(_05717_),
    .B(_05726_),
    .Y(_05728_));
 NAND2x2_ASAP7_75t_R _35336_ (.A(_05715_),
    .B(_05728_),
    .Y(_05729_));
 AOI21x1_ASAP7_75t_R _35337_ (.A1(net3428),
    .A2(_05317_),
    .B(_05715_),
    .Y(_05730_));
 INVx2_ASAP7_75t_R _35338_ (.A(_05730_),
    .Y(_05731_));
 AO21x1_ASAP7_75t_R _35339_ (.A1(_05729_),
    .A2(_05731_),
    .B(_05693_),
    .Y(_05732_));
 TAPCELL_ASAP7_75t_R PHY_449 ();
 INVx3_ASAP7_75t_R _35341_ (.A(_00537_),
    .Y(_05734_));
 NOR2x2_ASAP7_75t_R _35342_ (.A(_00538_),
    .B(_05734_),
    .Y(_05735_));
 TAPCELL_ASAP7_75t_R PHY_448 ();
 NOR2x2_ASAP7_75t_R _35344_ (.A(net1225),
    .B(net1774),
    .Y(_05737_));
 TAPCELL_ASAP7_75t_R PHY_447 ();
 INVx3_ASAP7_75t_R _35346_ (.A(net2338),
    .Y(_05740_));
 NAND2x2_ASAP7_75t_R _35347_ (.A(net2704),
    .B(_05740_),
    .Y(_05741_));
 TAPCELL_ASAP7_75t_R PHY_446 ();
 NOR2x2_ASAP7_75t_R _35349_ (.A(net963),
    .B(_05741_),
    .Y(_05743_));
 INVx1_ASAP7_75t_R _35350_ (.A(_05743_),
    .Y(_05744_));
 INVx3_ASAP7_75t_R _35351_ (.A(_00541_),
    .Y(_05745_));
 NOR2x2_ASAP7_75t_R _35352_ (.A(net2338),
    .B(_05745_),
    .Y(_05746_));
 NAND2x2_ASAP7_75t_R _35353_ (.A(net962),
    .B(_05746_),
    .Y(_05747_));
 NAND2x2_ASAP7_75t_R _35354_ (.A(_00539_),
    .B(_00540_),
    .Y(_05748_));
 NAND2x2_ASAP7_75t_R _35355_ (.A(_00537_),
    .B(_00538_),
    .Y(_05750_));
 NOR2x2_ASAP7_75t_R _35356_ (.A(_05748_),
    .B(_05750_),
    .Y(_05751_));
 CKINVDCx6p67_ASAP7_75t_R _35357_ (.A(_05751_),
    .Y(_05752_));
 AO21x1_ASAP7_75t_R _35358_ (.A1(_05744_),
    .A2(_05747_),
    .B(_05752_),
    .Y(_05753_));
 NAND2x2_ASAP7_75t_R _35359_ (.A(_00541_),
    .B(net2338),
    .Y(_05754_));
 CKINVDCx9p33_ASAP7_75t_R _35360_ (.A(net1774),
    .Y(_05755_));
 TAPCELL_ASAP7_75t_R PHY_445 ();
 NAND2x2_ASAP7_75t_R _35362_ (.A(net1225),
    .B(_05755_),
    .Y(_05757_));
 NOR2x2_ASAP7_75t_R _35363_ (.A(net2569),
    .B(_05757_),
    .Y(_05758_));
 NOR2x2_ASAP7_75t_R _35364_ (.A(net1228),
    .B(_05754_),
    .Y(_05759_));
 OA21x2_ASAP7_75t_R _35365_ (.A1(_05758_),
    .A2(_05759_),
    .B(_05751_),
    .Y(_05761_));
 INVx1_ASAP7_75t_R _35366_ (.A(_05761_),
    .Y(_05762_));
 NAND2x1_ASAP7_75t_R _35367_ (.A(_05753_),
    .B(_05762_),
    .Y(_05763_));
 CKINVDCx16_ASAP7_75t_R _35368_ (.A(net1221),
    .Y(_05764_));
 NOR2x2_ASAP7_75t_R _35369_ (.A(net1774),
    .B(_05764_),
    .Y(_05765_));
 NOR2x2_ASAP7_75t_R _35370_ (.A(_00541_),
    .B(_05740_),
    .Y(_05766_));
 NAND2x2_ASAP7_75t_R _35371_ (.A(_05765_),
    .B(net3475),
    .Y(_05767_));
 TAPCELL_ASAP7_75t_R PHY_444 ();
 TAPCELL_ASAP7_75t_R PHY_443 ();
 AND2x6_ASAP7_75t_R _35374_ (.A(net1223),
    .B(net1778),
    .Y(_05770_));
 NAND2x2_ASAP7_75t_R _35375_ (.A(net1809),
    .B(_05770_),
    .Y(_05772_));
 AO21x1_ASAP7_75t_R _35376_ (.A1(_05767_),
    .A2(_05772_),
    .B(_05752_),
    .Y(_05773_));
 TAPCELL_ASAP7_75t_R PHY_442 ();
 NAND2x2_ASAP7_75t_R _35378_ (.A(net2338),
    .B(_05745_),
    .Y(_05775_));
 NOR2x2_ASAP7_75t_R _35379_ (.A(net1229),
    .B(_05775_),
    .Y(_05776_));
 NAND2x2_ASAP7_75t_R _35380_ (.A(_05751_),
    .B(_05776_),
    .Y(_05777_));
 NOR2x2_ASAP7_75t_R _35381_ (.A(_00541_),
    .B(net2338),
    .Y(_05778_));
 TAPCELL_ASAP7_75t_R PHY_441 ();
 NAND2x2_ASAP7_75t_R _35383_ (.A(net1175),
    .B(_05751_),
    .Y(_05780_));
 NAND3x2_ASAP7_75t_R _35384_ (.B(_05777_),
    .C(_05780_),
    .Y(_05781_),
    .A(_05773_));
 NOR2x2_ASAP7_75t_R _35385_ (.A(_05781_),
    .B(_05763_),
    .Y(_05783_));
 INVx2_ASAP7_75t_R _35386_ (.A(_00539_),
    .Y(_05784_));
 NOR2x2_ASAP7_75t_R _35387_ (.A(net3359),
    .B(_05784_),
    .Y(_05785_));
 INVx3_ASAP7_75t_R _35388_ (.A(_05750_),
    .Y(_05786_));
 NAND2x2_ASAP7_75t_R _35389_ (.A(_05785_),
    .B(_05786_),
    .Y(_05787_));
 TAPCELL_ASAP7_75t_R PHY_440 ();
 INVx4_ASAP7_75t_R _35391_ (.A(_00538_),
    .Y(_05789_));
 OR3x2_ASAP7_75t_R _35392_ (.A(_05734_),
    .B(_05789_),
    .C(_00539_),
    .Y(_05790_));
 NAND3x2_ASAP7_75t_R _35393_ (.B(_05787_),
    .C(_05790_),
    .Y(_05791_),
    .A(_05783_));
 NOR2x1_ASAP7_75t_R _35394_ (.A(_05735_),
    .B(_05791_),
    .Y(_05792_));
 NAND2x2_ASAP7_75t_R _35395_ (.A(_00537_),
    .B(_05792_),
    .Y(_05794_));
 TAPCELL_ASAP7_75t_R PHY_439 ();
 NAND2x2_ASAP7_75t_R _35397_ (.A(net2739),
    .B(net3475),
    .Y(_05796_));
 TAPCELL_ASAP7_75t_R PHY_438 ();
 NOR2x2_ASAP7_75t_R _35399_ (.A(_00537_),
    .B(_00538_),
    .Y(_05798_));
 INVx3_ASAP7_75t_R _35400_ (.A(_05748_),
    .Y(_05799_));
 NAND2x2_ASAP7_75t_R _35401_ (.A(_05798_),
    .B(_05799_),
    .Y(_05800_));
 TAPCELL_ASAP7_75t_R PHY_437 ();
 AO21x1_ASAP7_75t_R _35403_ (.A1(_05767_),
    .A2(net2230),
    .B(_05800_),
    .Y(_05802_));
 NOR2x2_ASAP7_75t_R _35404_ (.A(net1222),
    .B(_05755_),
    .Y(_05803_));
 NAND2x2_ASAP7_75t_R _35405_ (.A(net1174),
    .B(_05803_),
    .Y(_05805_));
 TAPCELL_ASAP7_75t_R PHY_436 ();
 NAND2x2_ASAP7_75t_R _35407_ (.A(net1222),
    .B(net1182),
    .Y(_05807_));
 AO21x1_ASAP7_75t_R _35408_ (.A1(net2288),
    .A2(_05807_),
    .B(_05800_),
    .Y(_05808_));
 TAPCELL_ASAP7_75t_R PHY_435 ();
 NAND2x2_ASAP7_75t_R _35410_ (.A(net1775),
    .B(_05764_),
    .Y(_05810_));
 NOR2x2_ASAP7_75t_R _35411_ (.A(net1444),
    .B(_05810_),
    .Y(_05811_));
 INVx3_ASAP7_75t_R _35412_ (.A(_05800_),
    .Y(_05812_));
 NAND2x1_ASAP7_75t_R _35413_ (.A(_05811_),
    .B(_05812_),
    .Y(_05813_));
 AND3x1_ASAP7_75t_R _35414_ (.A(_05802_),
    .B(_05808_),
    .C(_05813_),
    .Y(_05814_));
 CKINVDCx8_ASAP7_75t_R _35415_ (.A(_05754_),
    .Y(_05816_));
 NAND2x2_ASAP7_75t_R _35416_ (.A(_05803_),
    .B(_05816_),
    .Y(_05817_));
 TAPCELL_ASAP7_75t_R PHY_434 ();
 NAND2x2_ASAP7_75t_R _35418_ (.A(_05746_),
    .B(_05765_),
    .Y(_05819_));
 TAPCELL_ASAP7_75t_R PHY_433 ();
 NAND2x2_ASAP7_75t_R _35420_ (.A(_05785_),
    .B(_05798_),
    .Y(_05821_));
 TAPCELL_ASAP7_75t_R PHY_432 ();
 TAPCELL_ASAP7_75t_R PHY_431 ();
 AO21x1_ASAP7_75t_R _35423_ (.A1(_05817_),
    .A2(_05819_),
    .B(_05821_),
    .Y(_05824_));
 NAND2x2_ASAP7_75t_R _35424_ (.A(_05778_),
    .B(_05765_),
    .Y(_05825_));
 TAPCELL_ASAP7_75t_R PHY_430 ();
 AO21x1_ASAP7_75t_R _35426_ (.A1(net3372),
    .A2(net2288),
    .B(_05821_),
    .Y(_05828_));
 INVx3_ASAP7_75t_R _35427_ (.A(_05821_),
    .Y(_05829_));
 NAND2x1_ASAP7_75t_R _35428_ (.A(net3476),
    .B(_05829_),
    .Y(_05830_));
 AND3x1_ASAP7_75t_R _35429_ (.A(_05824_),
    .B(_05828_),
    .C(_05830_),
    .Y(_05831_));
 NAND2x1_ASAP7_75t_R _35430_ (.A(_05814_),
    .B(_05831_),
    .Y(_05832_));
 NAND2x2_ASAP7_75t_R _35431_ (.A(_05816_),
    .B(_05765_),
    .Y(_05833_));
 TAPCELL_ASAP7_75t_R PHY_429 ();
 INVx6_ASAP7_75t_R _35433_ (.A(_05759_),
    .Y(_05835_));
 TAPCELL_ASAP7_75t_R PHY_428 ();
 NOR2x2_ASAP7_75t_R _35435_ (.A(_00539_),
    .B(net3358),
    .Y(_05838_));
 NAND2x2_ASAP7_75t_R _35436_ (.A(_05838_),
    .B(_05798_),
    .Y(_05839_));
 TAPCELL_ASAP7_75t_R PHY_427 ();
 AO21x1_ASAP7_75t_R _35438_ (.A1(net3467),
    .A2(_05835_),
    .B(_05839_),
    .Y(_05841_));
 TAPCELL_ASAP7_75t_R PHY_426 ();
 AO21x1_ASAP7_75t_R _35440_ (.A1(net980),
    .A2(net2540),
    .B(_05839_),
    .Y(_05843_));
 NAND2x2_ASAP7_75t_R _35441_ (.A(net1774),
    .B(net1222),
    .Y(_05844_));
 NOR2x2_ASAP7_75t_R _35442_ (.A(_05844_),
    .B(net2183),
    .Y(_05845_));
 INVx2_ASAP7_75t_R _35443_ (.A(_05839_),
    .Y(_05846_));
 NAND2x1_ASAP7_75t_R _35444_ (.A(_05845_),
    .B(_05846_),
    .Y(_05847_));
 AND3x1_ASAP7_75t_R _35445_ (.A(_05841_),
    .B(_05843_),
    .C(_05847_),
    .Y(_05849_));
 NAND2x2_ASAP7_75t_R _35446_ (.A(net2489),
    .B(_05770_),
    .Y(_05850_));
 TAPCELL_ASAP7_75t_R PHY_425 ();
 INVx1_ASAP7_75t_R _35448_ (.A(_00540_),
    .Y(_05852_));
 NOR2x2_ASAP7_75t_R _35449_ (.A(_00539_),
    .B(_05852_),
    .Y(_05853_));
 NAND2x2_ASAP7_75t_R _35450_ (.A(_05798_),
    .B(_05853_),
    .Y(_05854_));
 TAPCELL_ASAP7_75t_R PHY_424 ();
 AO21x1_ASAP7_75t_R _35452_ (.A1(_05850_),
    .A2(_05819_),
    .B(_05854_),
    .Y(_05856_));
 NAND2x2_ASAP7_75t_R _35453_ (.A(_05770_),
    .B(_05816_),
    .Y(_05857_));
 TAPCELL_ASAP7_75t_R PHY_423 ();
 NAND2x2_ASAP7_75t_R _35455_ (.A(net2739),
    .B(_05816_),
    .Y(_05860_));
 TAPCELL_ASAP7_75t_R PHY_422 ();
 TAPCELL_ASAP7_75t_R PHY_421 ();
 TAPCELL_ASAP7_75t_R PHY_420 ();
 AO21x1_ASAP7_75t_R _35459_ (.A1(net3357),
    .A2(net2845),
    .B(net2679),
    .Y(_05864_));
 NAND2x1_ASAP7_75t_R _35460_ (.A(_05757_),
    .B(net1810),
    .Y(_05865_));
 NAND2x1_ASAP7_75t_R _35461_ (.A(_05755_),
    .B(net1180),
    .Y(_05866_));
 AO21x1_ASAP7_75t_R _35462_ (.A1(_05865_),
    .A2(_05866_),
    .B(_05854_),
    .Y(_05867_));
 AND3x1_ASAP7_75t_R _35463_ (.A(_05856_),
    .B(_05864_),
    .C(_05867_),
    .Y(_05868_));
 NAND2x1_ASAP7_75t_R _35464_ (.A(_05849_),
    .B(_05868_),
    .Y(_05869_));
 NOR2x2_ASAP7_75t_R _35465_ (.A(_05832_),
    .B(_05869_),
    .Y(_05871_));
 NOR2x2_ASAP7_75t_R _35466_ (.A(_00537_),
    .B(_05789_),
    .Y(_05872_));
 NAND2x2_ASAP7_75t_R _35467_ (.A(_05872_),
    .B(_05838_),
    .Y(_05873_));
 TAPCELL_ASAP7_75t_R PHY_419 ();
 AO21x1_ASAP7_75t_R _35469_ (.A1(_05857_),
    .A2(_05835_),
    .B(_05873_),
    .Y(_05875_));
 NAND2x2_ASAP7_75t_R _35470_ (.A(net1225),
    .B(_05746_),
    .Y(_05876_));
 AO21x1_ASAP7_75t_R _35471_ (.A1(_05876_),
    .A2(net2081),
    .B(_05873_),
    .Y(_05877_));
 INVx3_ASAP7_75t_R _35472_ (.A(_05873_),
    .Y(_05878_));
 NAND2x2_ASAP7_75t_R _35473_ (.A(net1181),
    .B(_05770_),
    .Y(_05879_));
 INVx4_ASAP7_75t_R _35474_ (.A(net2603),
    .Y(_05880_));
 NAND2x1_ASAP7_75t_R _35475_ (.A(_05878_),
    .B(_05880_),
    .Y(_05882_));
 AND3x1_ASAP7_75t_R _35476_ (.A(_05875_),
    .B(_05877_),
    .C(_05882_),
    .Y(_05883_));
 NAND2x2_ASAP7_75t_R _35477_ (.A(_05872_),
    .B(_05853_),
    .Y(_05884_));
 INVx4_ASAP7_75t_R _35478_ (.A(_05884_),
    .Y(_05885_));
 TAPCELL_ASAP7_75t_R PHY_418 ();
 NAND2x2_ASAP7_75t_R _35480_ (.A(net2739),
    .B(_05778_),
    .Y(_05887_));
 AO21x1_ASAP7_75t_R _35481_ (.A1(_05807_),
    .A2(net2736),
    .B(_05884_),
    .Y(_05888_));
 OAI21x1_ASAP7_75t_R _35482_ (.A1(_05884_),
    .A2(net1662),
    .B(_05888_),
    .Y(_05889_));
 AOI21x1_ASAP7_75t_R _35483_ (.A1(_05885_),
    .A2(net3348),
    .B(_05889_),
    .Y(_05890_));
 NAND2x1_ASAP7_75t_R _35484_ (.A(_05883_),
    .B(_05890_),
    .Y(_05891_));
 TAPCELL_ASAP7_75t_R PHY_417 ();
 NAND2x2_ASAP7_75t_R _35486_ (.A(_05799_),
    .B(_05872_),
    .Y(_05894_));
 TAPCELL_ASAP7_75t_R PHY_416 ();
 AOI211x1_ASAP7_75t_R _35488_ (.A1(_05764_),
    .A2(net1776),
    .B(_05894_),
    .C(net2185),
    .Y(_05896_));
 NOR2x2_ASAP7_75t_R _35489_ (.A(net1439),
    .B(_05844_),
    .Y(_05897_));
 INVx5_ASAP7_75t_R _35490_ (.A(_05894_),
    .Y(_05898_));
 NOR2x1_ASAP7_75t_R _35491_ (.A(_05817_),
    .B(_05894_),
    .Y(_05899_));
 AO21x1_ASAP7_75t_R _35492_ (.A1(_05897_),
    .A2(_05898_),
    .B(_05899_),
    .Y(_05900_));
 NOR2x1_ASAP7_75t_R _35493_ (.A(_05896_),
    .B(_05900_),
    .Y(_05901_));
 TAPCELL_ASAP7_75t_R PHY_415 ();
 AO21x1_ASAP7_75t_R _35495_ (.A1(net2876),
    .A2(net2229),
    .B(_05894_),
    .Y(_05904_));
 NAND2x2_ASAP7_75t_R _35496_ (.A(_05764_),
    .B(net1179),
    .Y(_05905_));
 AO21x1_ASAP7_75t_R _35497_ (.A1(net3370),
    .A2(_05905_),
    .B(_05894_),
    .Y(_05906_));
 AND2x2_ASAP7_75t_R _35498_ (.A(_05904_),
    .B(_05906_),
    .Y(_05907_));
 NAND2x2_ASAP7_75t_R _35499_ (.A(_05785_),
    .B(_05872_),
    .Y(_05908_));
 TAPCELL_ASAP7_75t_R PHY_414 ();
 TAPCELL_ASAP7_75t_R PHY_413 ();
 AO21x1_ASAP7_75t_R _35502_ (.A1(_05817_),
    .A2(net3467),
    .B(_05908_),
    .Y(_05911_));
 OA21x2_ASAP7_75t_R _35503_ (.A1(_05908_),
    .A2(_05905_),
    .B(_05911_),
    .Y(_05912_));
 NAND3x1_ASAP7_75t_R _35504_ (.A(_05901_),
    .B(_05907_),
    .C(_05912_),
    .Y(_05913_));
 NOR2x1_ASAP7_75t_R _35505_ (.A(_05891_),
    .B(_05913_),
    .Y(_05915_));
 NAND2x2_ASAP7_75t_R _35506_ (.A(_05871_),
    .B(_05915_),
    .Y(_05916_));
 TAPCELL_ASAP7_75t_R PHY_412 ();
 NAND2x2_ASAP7_75t_R _35508_ (.A(_05764_),
    .B(_05746_),
    .Y(_05918_));
 AO21x1_ASAP7_75t_R _35509_ (.A1(net2271),
    .A2(_05918_),
    .B(_05752_),
    .Y(_05919_));
 OAI21x1_ASAP7_75t_R _35510_ (.A1(_05835_),
    .A2(_05752_),
    .B(_05919_),
    .Y(_05920_));
 NAND2x2_ASAP7_75t_R _35511_ (.A(_05844_),
    .B(net1808),
    .Y(_05921_));
 AO21x1_ASAP7_75t_R _35512_ (.A1(net3370),
    .A2(net2416),
    .B(_05752_),
    .Y(_05922_));
 OAI21x1_ASAP7_75t_R _35513_ (.A1(_05752_),
    .A2(_05921_),
    .B(_05922_),
    .Y(_05923_));
 NOR2x1_ASAP7_75t_R _35514_ (.A(_05920_),
    .B(_05923_),
    .Y(_05924_));
 CKINVDCx9p33_ASAP7_75t_R _35515_ (.A(_05787_),
    .Y(_05926_));
 TAPCELL_ASAP7_75t_R PHY_411 ();
 AND3x1_ASAP7_75t_R _35517_ (.A(_05926_),
    .B(_05764_),
    .C(_05816_),
    .Y(_05928_));
 INVx5_ASAP7_75t_R _35518_ (.A(net962),
    .Y(_05929_));
 NOR2x2_ASAP7_75t_R _35519_ (.A(net2540),
    .B(_05929_),
    .Y(_05930_));
 NOR2x2_ASAP7_75t_R _35520_ (.A(_05844_),
    .B(net2542),
    .Y(_05931_));
 OA21x2_ASAP7_75t_R _35521_ (.A1(_05930_),
    .A2(_05931_),
    .B(_05926_),
    .Y(_05932_));
 AO21x2_ASAP7_75t_R _35522_ (.A1(_05810_),
    .A2(_05757_),
    .B(net2184),
    .Y(_05933_));
 NOR2x1_ASAP7_75t_R _35523_ (.A(_05787_),
    .B(_05933_),
    .Y(_05934_));
 NOR3x1_ASAP7_75t_R _35524_ (.A(_05928_),
    .B(_05932_),
    .C(_05934_),
    .Y(_05935_));
 NAND2x1_ASAP7_75t_R _35525_ (.A(_05924_),
    .B(_05935_),
    .Y(_05937_));
 NAND2x2_ASAP7_75t_R _35526_ (.A(_05853_),
    .B(_05786_),
    .Y(_05938_));
 TAPCELL_ASAP7_75t_R PHY_410 ();
 TAPCELL_ASAP7_75t_R PHY_409 ();
 AO21x1_ASAP7_75t_R _35529_ (.A1(_05879_),
    .A2(_05905_),
    .B(net2520),
    .Y(_05941_));
 OAI21x1_ASAP7_75t_R _35530_ (.A1(net2520),
    .A2(_05921_),
    .B(_05941_),
    .Y(_05942_));
 NAND2x2_ASAP7_75t_R _35531_ (.A(_05803_),
    .B(net2490),
    .Y(_05943_));
 TAPCELL_ASAP7_75t_R PHY_408 ();
 TAPCELL_ASAP7_75t_R PHY_407 ();
 AO21x1_ASAP7_75t_R _35534_ (.A1(net1913),
    .A2(net2271),
    .B(_05938_),
    .Y(_05946_));
 OR3x4_ASAP7_75t_R _35535_ (.A(_05938_),
    .B(net1880),
    .C(_05737_),
    .Y(_05948_));
 NAND2x1_ASAP7_75t_R _35536_ (.A(_05946_),
    .B(_05948_),
    .Y(_05949_));
 NOR2x1_ASAP7_75t_R _35537_ (.A(_05942_),
    .B(_05949_),
    .Y(_05950_));
 NAND2x2_ASAP7_75t_R _35538_ (.A(_05838_),
    .B(_05786_),
    .Y(_05951_));
 TAPCELL_ASAP7_75t_R PHY_406 ();
 INVx2_ASAP7_75t_R _35540_ (.A(net3352),
    .Y(_05953_));
 OAI21x1_ASAP7_75t_R _35541_ (.A1(_05759_),
    .A2(net2518),
    .B(_05953_),
    .Y(_05954_));
 OAI21x1_ASAP7_75t_R _35542_ (.A1(net1913),
    .A2(net3352),
    .B(_05954_),
    .Y(_05955_));
 NOR2x1_ASAP7_75t_R _35543_ (.A(net3352),
    .B(_05772_),
    .Y(_05956_));
 CKINVDCx9p33_ASAP7_75t_R _35544_ (.A(net1174),
    .Y(_05957_));
 TAPCELL_ASAP7_75t_R PHY_405 ();
 AOI211x1_ASAP7_75t_R _35546_ (.A1(_05764_),
    .A2(net1774),
    .B(net3352),
    .C(_05957_),
    .Y(_05960_));
 NOR3x1_ASAP7_75t_R _35547_ (.A(_05955_),
    .B(_05956_),
    .C(_05960_),
    .Y(_05961_));
 NAND2x1_ASAP7_75t_R _35548_ (.A(_05950_),
    .B(_05961_),
    .Y(_05962_));
 NOR2x1_ASAP7_75t_R _35549_ (.A(_05937_),
    .B(_05962_),
    .Y(_05963_));
 NOR2x2_ASAP7_75t_R _35550_ (.A(_05764_),
    .B(net1438),
    .Y(_05964_));
 NAND2x2_ASAP7_75t_R _35551_ (.A(_00537_),
    .B(_05789_),
    .Y(_05965_));
 NOR2x2_ASAP7_75t_R _35552_ (.A(_05748_),
    .B(_05965_),
    .Y(_05966_));
 TAPCELL_ASAP7_75t_R PHY_404 ();
 TAPCELL_ASAP7_75t_R PHY_403 ();
 OA21x2_ASAP7_75t_R _35555_ (.A1(_05845_),
    .A2(_05964_),
    .B(net2636),
    .Y(_05970_));
 NAND2x1_ASAP7_75t_R _35556_ (.A(_05807_),
    .B(net2876),
    .Y(_05971_));
 TAPCELL_ASAP7_75t_R PHY_402 ();
 NAND2x1_ASAP7_75t_R _35558_ (.A(_05796_),
    .B(_05805_),
    .Y(_05973_));
 OA21x2_ASAP7_75t_R _35559_ (.A1(_05971_),
    .A2(_05973_),
    .B(_05966_),
    .Y(_05974_));
 NOR2x1_ASAP7_75t_R _35560_ (.A(_05970_),
    .B(_05974_),
    .Y(_05975_));
 INVx3_ASAP7_75t_R _35561_ (.A(_05887_),
    .Y(_05976_));
 NAND2x2_ASAP7_75t_R _35562_ (.A(_05785_),
    .B(_05735_),
    .Y(_05977_));
 INVx3_ASAP7_75t_R _35563_ (.A(_05977_),
    .Y(_05978_));
 NAND2x1_ASAP7_75t_R _35564_ (.A(_05976_),
    .B(_05978_),
    .Y(_05979_));
 TAPCELL_ASAP7_75t_R PHY_401 ();
 AO21x1_ASAP7_75t_R _35566_ (.A1(net2875),
    .A2(net2229),
    .B(_05977_),
    .Y(_05982_));
 NAND2x1_ASAP7_75t_R _35567_ (.A(_05979_),
    .B(_05982_),
    .Y(_05983_));
 AO21x2_ASAP7_75t_R _35568_ (.A1(_05857_),
    .A2(_05833_),
    .B(_05977_),
    .Y(_05984_));
 NOR2x2_ASAP7_75t_R _35569_ (.A(net1442),
    .B(_05929_),
    .Y(_05985_));
 NAND2x2_ASAP7_75t_R _35570_ (.A(_05985_),
    .B(_05978_),
    .Y(_05986_));
 INVx2_ASAP7_75t_R _35571_ (.A(_05918_),
    .Y(_05987_));
 NAND2x1_ASAP7_75t_R _35572_ (.A(_05987_),
    .B(_05978_),
    .Y(_05988_));
 NAND3x1_ASAP7_75t_R _35573_ (.A(_05984_),
    .B(_05986_),
    .C(_05988_),
    .Y(_05989_));
 NOR2x1_ASAP7_75t_R _35574_ (.A(_05983_),
    .B(_05989_),
    .Y(_05990_));
 NAND2x1_ASAP7_75t_R _35575_ (.A(_05975_),
    .B(_05990_),
    .Y(_05992_));
 NAND2x2_ASAP7_75t_R _35576_ (.A(_05838_),
    .B(_05735_),
    .Y(_05993_));
 TAPCELL_ASAP7_75t_R PHY_400 ();
 TAPCELL_ASAP7_75t_R PHY_399 ();
 TAPCELL_ASAP7_75t_R PHY_398 ();
 AO21x1_ASAP7_75t_R _35580_ (.A1(net3370),
    .A2(net2416),
    .B(_05993_),
    .Y(_05997_));
 OAI21x1_ASAP7_75t_R _35581_ (.A1(net2229),
    .A2(net2525),
    .B(_05997_),
    .Y(_05998_));
 AO21x1_ASAP7_75t_R _35582_ (.A1(net3357),
    .A2(_05833_),
    .B(net2525),
    .Y(_05999_));
 TAPCELL_ASAP7_75t_R PHY_397 ();
 AO21x1_ASAP7_75t_R _35584_ (.A1(_05819_),
    .A2(net2231),
    .B(_05993_),
    .Y(_06001_));
 INVx1_ASAP7_75t_R _35585_ (.A(_05993_),
    .Y(_06003_));
 NAND2x2_ASAP7_75t_R _35586_ (.A(_05985_),
    .B(_06003_),
    .Y(_06004_));
 NAND3x1_ASAP7_75t_R _35587_ (.A(_05999_),
    .B(_06001_),
    .C(_06004_),
    .Y(_06005_));
 NOR2x1_ASAP7_75t_R _35588_ (.A(_05998_),
    .B(_06005_),
    .Y(_06006_));
 NAND2x2_ASAP7_75t_R _35589_ (.A(_05853_),
    .B(_05735_),
    .Y(_06007_));
 TAPCELL_ASAP7_75t_R PHY_396 ();
 AO21x1_ASAP7_75t_R _35591_ (.A1(_05833_),
    .A2(net2485),
    .B(_06007_),
    .Y(_06009_));
 AO21x1_ASAP7_75t_R _35592_ (.A1(net2098),
    .A2(net2231),
    .B(_06007_),
    .Y(_06010_));
 NOR2x1_ASAP7_75t_R _35593_ (.A(_05876_),
    .B(_06007_),
    .Y(_06011_));
 INVx1_ASAP7_75t_R _35594_ (.A(_06011_),
    .Y(_06012_));
 NAND3x1_ASAP7_75t_R _35595_ (.A(_06009_),
    .B(_06010_),
    .C(_06012_),
    .Y(_06014_));
 INVx4_ASAP7_75t_R _35596_ (.A(_05805_),
    .Y(_06015_));
 NAND2x1_ASAP7_75t_R _35597_ (.A(net3360),
    .B(_05784_),
    .Y(_06016_));
 NOR2x2_ASAP7_75t_R _35598_ (.A(_06016_),
    .B(_05965_),
    .Y(_06017_));
 AOI211x1_ASAP7_75t_R _35599_ (.A1(_05764_),
    .A2(net1777),
    .B(_06007_),
    .C(net2543),
    .Y(_06018_));
 AO21x1_ASAP7_75t_R _35600_ (.A1(_06015_),
    .A2(_06017_),
    .B(_06018_),
    .Y(_06019_));
 NOR2x1_ASAP7_75t_R _35601_ (.A(_06019_),
    .B(_06014_),
    .Y(_06020_));
 NAND2x1_ASAP7_75t_R _35602_ (.A(_06020_),
    .B(_06006_),
    .Y(_06021_));
 NOR2x1_ASAP7_75t_R _35603_ (.A(_05992_),
    .B(_06021_),
    .Y(_06022_));
 NAND2x1_ASAP7_75t_R _35604_ (.A(_05963_),
    .B(_06022_),
    .Y(_06023_));
 NOR2x2_ASAP7_75t_R _35605_ (.A(_05916_),
    .B(_06023_),
    .Y(_06025_));
 NAND2x2_ASAP7_75t_R _35606_ (.A(net1978),
    .B(_06025_),
    .Y(_06026_));
 TAPCELL_ASAP7_75t_R PHY_395 ();
 TAPCELL_ASAP7_75t_R PHY_394 ();
 CKINVDCx20_ASAP7_75t_R _35609_ (.A(net1785),
    .Y(_06029_));
 NOR2x2_ASAP7_75t_R _35610_ (.A(net1550),
    .B(_06029_),
    .Y(_06030_));
 TAPCELL_ASAP7_75t_R PHY_393 ();
 TAPCELL_ASAP7_75t_R PHY_392 ();
 INVx2_ASAP7_75t_R _35613_ (.A(_00630_),
    .Y(_06033_));
 NOR2x2_ASAP7_75t_R _35614_ (.A(net1812),
    .B(_06033_),
    .Y(_06034_));
 NAND2x2_ASAP7_75t_R _35615_ (.A(_06030_),
    .B(_06034_),
    .Y(_06036_));
 NOR2x2_ASAP7_75t_R _35616_ (.A(net1812),
    .B(_00630_),
    .Y(_06037_));
 TAPCELL_ASAP7_75t_R PHY_391 ();
 NAND2x2_ASAP7_75t_R _35618_ (.A(_06029_),
    .B(net1093),
    .Y(_06039_));
 INVx3_ASAP7_75t_R _35619_ (.A(net3232),
    .Y(_06040_));
 NOR2x2_ASAP7_75t_R _35620_ (.A(_00626_),
    .B(_06040_),
    .Y(_06041_));
 INVx2_ASAP7_75t_R _35621_ (.A(_00628_),
    .Y(_06042_));
 NOR2x2_ASAP7_75t_R _35622_ (.A(_00627_),
    .B(_06042_),
    .Y(_06043_));
 NAND2x2_ASAP7_75t_R _35623_ (.A(_06041_),
    .B(_06043_),
    .Y(_06044_));
 AO21x1_ASAP7_75t_R _35624_ (.A1(_06036_),
    .A2(_06039_),
    .B(net2786),
    .Y(_06045_));
 NOR2x2_ASAP7_75t_R _35625_ (.A(net1780),
    .B(net1550),
    .Y(_06047_));
 INVx2_ASAP7_75t_R _35626_ (.A(net1812),
    .Y(_06048_));
 NOR2x2_ASAP7_75t_R _35627_ (.A(net2873),
    .B(_06048_),
    .Y(_06049_));
 NAND2x2_ASAP7_75t_R _35628_ (.A(_06047_),
    .B(net2507),
    .Y(_06050_));
 TAPCELL_ASAP7_75t_R PHY_390 ();
 NAND2x2_ASAP7_75t_R _35630_ (.A(net1812),
    .B(net2873),
    .Y(_06052_));
 TAPCELL_ASAP7_75t_R PHY_389 ();
 AO21x1_ASAP7_75t_R _35632_ (.A1(_06050_),
    .A2(_06052_),
    .B(net2786),
    .Y(_06054_));
 AND2x4_ASAP7_75t_R _35633_ (.A(_06045_),
    .B(_06054_),
    .Y(_06055_));
 NOR2x2_ASAP7_75t_R _35634_ (.A(_00627_),
    .B(_00628_),
    .Y(_06056_));
 NAND2x2_ASAP7_75t_R _35635_ (.A(net1782),
    .B(net1550),
    .Y(_06058_));
 AND4x2_ASAP7_75t_R _35636_ (.A(_06041_),
    .B(_06037_),
    .C(_06056_),
    .D(net1663),
    .Y(_06059_));
 TAPCELL_ASAP7_75t_R PHY_388 ();
 CKINVDCx16_ASAP7_75t_R _35638_ (.A(net1550),
    .Y(_06061_));
 TAPCELL_ASAP7_75t_R PHY_387 ();
 NAND2x2_ASAP7_75t_R _35640_ (.A(net2873),
    .B(_06048_),
    .Y(_06063_));
 NAND2x2_ASAP7_75t_R _35641_ (.A(_06041_),
    .B(_06056_),
    .Y(_06064_));
 AOI211x1_ASAP7_75t_R _35642_ (.A1(_06029_),
    .A2(_06061_),
    .B(net1588),
    .C(_06064_),
    .Y(_06065_));
 NOR2x2_ASAP7_75t_R _35643_ (.A(_06059_),
    .B(_06065_),
    .Y(_06066_));
 TAPCELL_ASAP7_75t_R PHY_386 ();
 TAPCELL_ASAP7_75t_R PHY_385 ();
 NAND2x2_ASAP7_75t_R _35646_ (.A(net1276),
    .B(net1297),
    .Y(_06070_));
 AND2x6_ASAP7_75t_R _35647_ (.A(net1814),
    .B(net2873),
    .Y(_06071_));
 NAND2x2_ASAP7_75t_R _35648_ (.A(_06061_),
    .B(_06071_),
    .Y(_06072_));
 TAPCELL_ASAP7_75t_R PHY_384 ();
 TAPCELL_ASAP7_75t_R PHY_383 ();
 AO31x2_ASAP7_75t_R _35651_ (.A1(_06070_),
    .A2(_06050_),
    .A3(_06072_),
    .B(_06064_),
    .Y(_06075_));
 NAND3x2_ASAP7_75t_R _35652_ (.B(_06066_),
    .C(_06075_),
    .Y(_06076_),
    .A(_06055_));
 TAPCELL_ASAP7_75t_R PHY_382 ();
 NAND2x2_ASAP7_75t_R _35654_ (.A(_06030_),
    .B(_06071_),
    .Y(_06078_));
 AND2x6_ASAP7_75t_R _35655_ (.A(_00627_),
    .B(_00628_),
    .Y(_06080_));
 NAND2x2_ASAP7_75t_R _35656_ (.A(_06041_),
    .B(_06080_),
    .Y(_06081_));
 TAPCELL_ASAP7_75t_R PHY_381 ();
 AO21x1_ASAP7_75t_R _35658_ (.A1(_06078_),
    .A2(_06050_),
    .B(_06081_),
    .Y(_06083_));
 NAND2x2_ASAP7_75t_R _35659_ (.A(net1096),
    .B(_06030_),
    .Y(_06084_));
 NAND2x2_ASAP7_75t_R _35660_ (.A(_06037_),
    .B(_06047_),
    .Y(_06085_));
 TAPCELL_ASAP7_75t_R PHY_380 ();
 AO21x1_ASAP7_75t_R _35662_ (.A1(_06084_),
    .A2(_06085_),
    .B(_06081_),
    .Y(_06087_));
 NOR2x2_ASAP7_75t_R _35663_ (.A(net1814),
    .B(net1781),
    .Y(_06088_));
 NAND2x2_ASAP7_75t_R _35664_ (.A(net2874),
    .B(_06088_),
    .Y(_06089_));
 INVx3_ASAP7_75t_R _35665_ (.A(_06089_),
    .Y(_06091_));
 INVx6_ASAP7_75t_R _35666_ (.A(_06081_),
    .Y(_06092_));
 NAND2x2_ASAP7_75t_R _35667_ (.A(_06091_),
    .B(_06092_),
    .Y(_06093_));
 NAND3x2_ASAP7_75t_R _35668_ (.B(_06087_),
    .C(_06093_),
    .Y(_06094_),
    .A(_06083_));
 INVx1_ASAP7_75t_R _35669_ (.A(_06094_),
    .Y(_06095_));
 NAND2x2_ASAP7_75t_R _35670_ (.A(net1782),
    .B(_06061_),
    .Y(_06096_));
 NAND2x2_ASAP7_75t_R _35671_ (.A(net1545),
    .B(_06029_),
    .Y(_06097_));
 NAND2x2_ASAP7_75t_R _35672_ (.A(net1813),
    .B(_06033_),
    .Y(_06098_));
 AO21x2_ASAP7_75t_R _35673_ (.A1(_06096_),
    .A2(net3423),
    .B(_06098_),
    .Y(_06099_));
 NAND2x1_ASAP7_75t_R _35674_ (.A(_06072_),
    .B(_06099_),
    .Y(_06100_));
 INVx1_ASAP7_75t_R _35675_ (.A(_00627_),
    .Y(_06102_));
 NOR2x2_ASAP7_75t_R _35676_ (.A(_00628_),
    .B(_06102_),
    .Y(_06103_));
 NAND2x2_ASAP7_75t_R _35677_ (.A(_06041_),
    .B(_06103_),
    .Y(_06104_));
 INVx4_ASAP7_75t_R _35678_ (.A(_06104_),
    .Y(_06105_));
 NOR2x2_ASAP7_75t_R _35679_ (.A(net1780),
    .B(_06061_),
    .Y(_06106_));
 NAND2x2_ASAP7_75t_R _35680_ (.A(_06106_),
    .B(_06034_),
    .Y(_06107_));
 INVx3_ASAP7_75t_R _35681_ (.A(_06107_),
    .Y(_06108_));
 NOR2x2_ASAP7_75t_R _35682_ (.A(_06096_),
    .B(_06063_),
    .Y(_06109_));
 OA21x2_ASAP7_75t_R _35683_ (.A1(_06108_),
    .A2(_06109_),
    .B(_06105_),
    .Y(_06110_));
 TAPCELL_ASAP7_75t_R PHY_379 ();
 NOR2x1_ASAP7_75t_R _35685_ (.A(_06085_),
    .B(_06104_),
    .Y(_06113_));
 AOI211x1_ASAP7_75t_R _35686_ (.A1(_06100_),
    .A2(_06105_),
    .B(_06110_),
    .C(_06113_),
    .Y(_06114_));
 NAND2x1_ASAP7_75t_R _35687_ (.A(_06095_),
    .B(_06114_),
    .Y(_06115_));
 NOR2x2_ASAP7_75t_R _35688_ (.A(_06076_),
    .B(_06115_),
    .Y(_06116_));
 TAPCELL_ASAP7_75t_R PHY_378 ();
 NAND2x2_ASAP7_75t_R _35690_ (.A(_06047_),
    .B(net1601),
    .Y(_06118_));
 TAPCELL_ASAP7_75t_R PHY_377 ();
 AND2x6_ASAP7_75t_R _35692_ (.A(net3234),
    .B(_00626_),
    .Y(_06120_));
 NAND2x2_ASAP7_75t_R _35693_ (.A(_06056_),
    .B(_06120_),
    .Y(_06121_));
 TAPCELL_ASAP7_75t_R PHY_376 ();
 TAPCELL_ASAP7_75t_R PHY_375 ();
 AO21x1_ASAP7_75t_R _35696_ (.A1(_06107_),
    .A2(net1540),
    .B(_06121_),
    .Y(_06125_));
 NAND2x2_ASAP7_75t_R _35697_ (.A(_06061_),
    .B(net2508),
    .Y(_06126_));
 AO21x1_ASAP7_75t_R _35698_ (.A1(net2530),
    .A2(_06126_),
    .B(_06121_),
    .Y(_06127_));
 AND2x6_ASAP7_75t_R _35699_ (.A(net1781),
    .B(net1545),
    .Y(_06128_));
 NAND2x2_ASAP7_75t_R _35700_ (.A(_06037_),
    .B(_06128_),
    .Y(_06129_));
 TAPCELL_ASAP7_75t_R PHY_374 ();
 NAND2x2_ASAP7_75t_R _35702_ (.A(_06037_),
    .B(_06106_),
    .Y(_06131_));
 TAPCELL_ASAP7_75t_R PHY_373 ();
 AO21x1_ASAP7_75t_R _35704_ (.A1(_06129_),
    .A2(net3434),
    .B(_06121_),
    .Y(_06133_));
 NAND3x1_ASAP7_75t_R _35705_ (.A(_06125_),
    .B(_06127_),
    .C(_06133_),
    .Y(_06135_));
 INVx1_ASAP7_75t_R _35706_ (.A(_06135_),
    .Y(_06136_));
 NAND2x2_ASAP7_75t_R _35707_ (.A(_06029_),
    .B(net2507),
    .Y(_06137_));
 INVx3_ASAP7_75t_R _35708_ (.A(_06137_),
    .Y(_06138_));
 AND2x6_ASAP7_75t_R _35709_ (.A(_06120_),
    .B(_06043_),
    .Y(_06139_));
 TAPCELL_ASAP7_75t_R PHY_372 ();
 INVx11_ASAP7_75t_R _35711_ (.A(net1092),
    .Y(_06141_));
 NOR2x2_ASAP7_75t_R _35712_ (.A(_06096_),
    .B(_06141_),
    .Y(_06142_));
 NOR2x2_ASAP7_75t_R _35713_ (.A(net1591),
    .B(_06128_),
    .Y(_06143_));
 OA21x2_ASAP7_75t_R _35714_ (.A1(_06142_),
    .A2(_06143_),
    .B(_06139_),
    .Y(_06144_));
 NAND2x2_ASAP7_75t_R _35715_ (.A(net2744),
    .B(_06139_),
    .Y(_06146_));
 NOR2x2_ASAP7_75t_R _35716_ (.A(net1759),
    .B(_06146_),
    .Y(_06147_));
 AOI211x1_ASAP7_75t_R _35717_ (.A1(_06138_),
    .A2(_06139_),
    .B(_06144_),
    .C(_06147_),
    .Y(_06148_));
 NAND2x1_ASAP7_75t_R _35718_ (.A(_06136_),
    .B(_06148_),
    .Y(_06149_));
 NAND2x2_ASAP7_75t_R _35719_ (.A(net1782),
    .B(net1093),
    .Y(_06150_));
 NAND2x2_ASAP7_75t_R _35720_ (.A(_06080_),
    .B(_06120_),
    .Y(_06151_));
 AO21x1_ASAP7_75t_R _35721_ (.A1(_06150_),
    .A2(net3434),
    .B(_06151_),
    .Y(_06152_));
 NAND2x2_ASAP7_75t_R _35722_ (.A(net2507),
    .B(_06128_),
    .Y(_06153_));
 AO21x1_ASAP7_75t_R _35723_ (.A1(net1261),
    .A2(_06050_),
    .B(_06151_),
    .Y(_06154_));
 NAND2x1_ASAP7_75t_R _35724_ (.A(_06152_),
    .B(_06154_),
    .Y(_06155_));
 INVx1_ASAP7_75t_R _35725_ (.A(_06155_),
    .Y(_06157_));
 NAND2x2_ASAP7_75t_R _35726_ (.A(_06103_),
    .B(_06120_),
    .Y(_06158_));
 CKINVDCx8_ASAP7_75t_R _35727_ (.A(net3472),
    .Y(_06159_));
 TAPCELL_ASAP7_75t_R PHY_371 ();
 NAND2x2_ASAP7_75t_R _35729_ (.A(net1599),
    .B(_06159_),
    .Y(_06161_));
 TAPCELL_ASAP7_75t_R PHY_370 ();
 AO21x1_ASAP7_75t_R _35731_ (.A1(_06150_),
    .A2(_06085_),
    .B(net2344),
    .Y(_06163_));
 NAND2x2_ASAP7_75t_R _35732_ (.A(_06161_),
    .B(_06163_),
    .Y(_06164_));
 AO21x2_ASAP7_75t_R _35733_ (.A1(net1261),
    .A2(_06050_),
    .B(net2344),
    .Y(_06165_));
 AOI211x1_ASAP7_75t_R _35734_ (.A1(_06029_),
    .A2(_06061_),
    .B(net2344),
    .C(net1603),
    .Y(_06166_));
 INVx1_ASAP7_75t_R _35735_ (.A(_06166_),
    .Y(_06168_));
 NAND2x2_ASAP7_75t_R _35736_ (.A(_06165_),
    .B(_06168_),
    .Y(_06169_));
 NOR2x1_ASAP7_75t_R _35737_ (.A(_06164_),
    .B(_06169_),
    .Y(_06170_));
 NAND2x1_ASAP7_75t_R _35738_ (.A(_06157_),
    .B(_06170_),
    .Y(_06171_));
 NOR2x1_ASAP7_75t_R _35739_ (.A(_06149_),
    .B(_06171_),
    .Y(_06172_));
 NAND2x1_ASAP7_75t_R _35740_ (.A(_06116_),
    .B(_06172_),
    .Y(_06173_));
 INVx3_ASAP7_75t_R _35741_ (.A(_00626_),
    .Y(_06174_));
 NOR2x2_ASAP7_75t_R _35742_ (.A(net3232),
    .B(_06174_),
    .Y(_06175_));
 NAND2x2_ASAP7_75t_R _35743_ (.A(_06175_),
    .B(_06103_),
    .Y(_06176_));
 AO21x1_ASAP7_75t_R _35744_ (.A1(_06129_),
    .A2(_06085_),
    .B(_06176_),
    .Y(_06177_));
 AO21x2_ASAP7_75t_R _35745_ (.A1(_06036_),
    .A2(_06107_),
    .B(_06176_),
    .Y(_06179_));
 NAND2x1_ASAP7_75t_R _35746_ (.A(_06177_),
    .B(_06179_),
    .Y(_06180_));
 NAND2x2_ASAP7_75t_R _35747_ (.A(net2507),
    .B(_06106_),
    .Y(_06181_));
 NAND2x2_ASAP7_75t_R _35748_ (.A(_06047_),
    .B(_06071_),
    .Y(_06182_));
 AO21x1_ASAP7_75t_R _35749_ (.A1(_06181_),
    .A2(_06182_),
    .B(_06176_),
    .Y(_06183_));
 TAPCELL_ASAP7_75t_R PHY_369 ();
 AO21x1_ASAP7_75t_R _35751_ (.A1(_06078_),
    .A2(_06050_),
    .B(_06176_),
    .Y(_06185_));
 NAND2x1_ASAP7_75t_R _35752_ (.A(_06183_),
    .B(_06185_),
    .Y(_06186_));
 NOR2x1_ASAP7_75t_R _35753_ (.A(_06180_),
    .B(_06186_),
    .Y(_06187_));
 NOR2x2_ASAP7_75t_R _35754_ (.A(_06058_),
    .B(_06052_),
    .Y(_06188_));
 CKINVDCx6p67_ASAP7_75t_R _35755_ (.A(_06188_),
    .Y(_06190_));
 NAND2x2_ASAP7_75t_R _35756_ (.A(_06175_),
    .B(_06080_),
    .Y(_06191_));
 AO21x1_ASAP7_75t_R _35757_ (.A1(_06190_),
    .A2(_06182_),
    .B(_06191_),
    .Y(_06192_));
 NOR2x2_ASAP7_75t_R _35758_ (.A(_06096_),
    .B(_06098_),
    .Y(_06193_));
 INVx4_ASAP7_75t_R _35759_ (.A(_06191_),
    .Y(_06194_));
 NAND2x1_ASAP7_75t_R _35760_ (.A(_06193_),
    .B(_06194_),
    .Y(_06195_));
 NAND2x2_ASAP7_75t_R _35761_ (.A(net1782),
    .B(net1598),
    .Y(_06196_));
 INVx2_ASAP7_75t_R _35762_ (.A(_06196_),
    .Y(_06197_));
 NAND2x1_ASAP7_75t_R _35763_ (.A(_06197_),
    .B(_06194_),
    .Y(_06198_));
 AND3x1_ASAP7_75t_R _35764_ (.A(_06192_),
    .B(_06195_),
    .C(_06198_),
    .Y(_06199_));
 NAND2x1_ASAP7_75t_R _35765_ (.A(_06187_),
    .B(_06199_),
    .Y(_06201_));
 TAPCELL_ASAP7_75t_R PHY_368 ();
 NAND2x2_ASAP7_75t_R _35767_ (.A(_06043_),
    .B(_06175_),
    .Y(_06203_));
 TAPCELL_ASAP7_75t_R PHY_367 ();
 AO21x1_ASAP7_75t_R _35769_ (.A1(_06107_),
    .A2(_06196_),
    .B(_06203_),
    .Y(_06205_));
 AO21x1_ASAP7_75t_R _35770_ (.A1(_06131_),
    .A2(_06150_),
    .B(_06203_),
    .Y(_06206_));
 INVx5_ASAP7_75t_R _35771_ (.A(_06203_),
    .Y(_06207_));
 NAND2x1_ASAP7_75t_R _35772_ (.A(net2856),
    .B(_06207_),
    .Y(_06208_));
 AND3x1_ASAP7_75t_R _35773_ (.A(_06205_),
    .B(_06206_),
    .C(_06208_),
    .Y(_06209_));
 NAND2x2_ASAP7_75t_R _35774_ (.A(_06056_),
    .B(_06175_),
    .Y(_06210_));
 INVx3_ASAP7_75t_R _35775_ (.A(_06210_),
    .Y(_06212_));
 NOR2x2_ASAP7_75t_R _35776_ (.A(_06097_),
    .B(_06141_),
    .Y(_06213_));
 NOR2x1_ASAP7_75t_R _35777_ (.A(_06091_),
    .B(_06213_),
    .Y(_06214_));
 INVx1_ASAP7_75t_R _35778_ (.A(_06214_),
    .Y(_06215_));
 TAPCELL_ASAP7_75t_R PHY_366 ();
 TAPCELL_ASAP7_75t_R PHY_365 ();
 AOI211x1_ASAP7_75t_R _35781_ (.A1(_06029_),
    .A2(net1548),
    .B(_06210_),
    .C(_06098_),
    .Y(_06218_));
 NAND2x2_ASAP7_75t_R _35782_ (.A(net1784),
    .B(net3429),
    .Y(_06219_));
 NOR2x1_ASAP7_75t_R _35783_ (.A(_06210_),
    .B(_06219_),
    .Y(_06220_));
 AOI211x1_ASAP7_75t_R _35784_ (.A1(_06212_),
    .A2(_06215_),
    .B(_06218_),
    .C(_06220_),
    .Y(_06221_));
 NAND2x1_ASAP7_75t_R _35785_ (.A(_06209_),
    .B(_06221_),
    .Y(_06223_));
 NOR2x1_ASAP7_75t_R _35786_ (.A(_06201_),
    .B(_06223_),
    .Y(_06224_));
 TAPCELL_ASAP7_75t_R PHY_364 ();
 NAND2x2_ASAP7_75t_R _35788_ (.A(_06106_),
    .B(_06071_),
    .Y(_06226_));
 TAPCELL_ASAP7_75t_R PHY_363 ();
 NOR2x2_ASAP7_75t_R _35790_ (.A(net3232),
    .B(_00626_),
    .Y(_06228_));
 NAND2x2_ASAP7_75t_R _35791_ (.A(_06228_),
    .B(_06103_),
    .Y(_06229_));
 TAPCELL_ASAP7_75t_R PHY_362 ();
 AO21x1_ASAP7_75t_R _35793_ (.A1(_06181_),
    .A2(_06226_),
    .B(_06229_),
    .Y(_06231_));
 TAPCELL_ASAP7_75t_R PHY_361 ();
 AO21x1_ASAP7_75t_R _35795_ (.A1(_06150_),
    .A2(_06085_),
    .B(_06229_),
    .Y(_06234_));
 NOR2x1_ASAP7_75t_R _35796_ (.A(_06229_),
    .B(_06118_),
    .Y(_06235_));
 INVx1_ASAP7_75t_R _35797_ (.A(_06235_),
    .Y(_06236_));
 NAND3x1_ASAP7_75t_R _35798_ (.A(_06231_),
    .B(_06234_),
    .C(_06236_),
    .Y(_06237_));
 TAPCELL_ASAP7_75t_R PHY_360 ();
 NAND2x2_ASAP7_75t_R _35800_ (.A(_06058_),
    .B(net1296),
    .Y(_06239_));
 NAND2x2_ASAP7_75t_R _35801_ (.A(_06228_),
    .B(_06080_),
    .Y(_06240_));
 TAPCELL_ASAP7_75t_R PHY_359 ();
 AO21x1_ASAP7_75t_R _35803_ (.A1(_06190_),
    .A2(_06239_),
    .B(_06240_),
    .Y(_06242_));
 AO21x1_ASAP7_75t_R _35804_ (.A1(_06084_),
    .A2(_06039_),
    .B(_06240_),
    .Y(_06243_));
 INVx3_ASAP7_75t_R _35805_ (.A(_06240_),
    .Y(_06245_));
 NAND2x2_ASAP7_75t_R _35806_ (.A(_06197_),
    .B(_06245_),
    .Y(_06246_));
 NAND3x1_ASAP7_75t_R _35807_ (.A(_06242_),
    .B(_06243_),
    .C(_06246_),
    .Y(_06247_));
 NOR2x1_ASAP7_75t_R _35808_ (.A(_06237_),
    .B(_06247_),
    .Y(_06248_));
 INVx1_ASAP7_75t_R _35809_ (.A(_06248_),
    .Y(_06249_));
 NAND2x2_ASAP7_75t_R _35810_ (.A(_06056_),
    .B(_06228_),
    .Y(_06250_));
 INVx6_ASAP7_75t_R _35811_ (.A(_06250_),
    .Y(_06251_));
 NAND2x1_ASAP7_75t_R _35812_ (.A(_06109_),
    .B(_06251_),
    .Y(_06252_));
 AO21x1_ASAP7_75t_R _35813_ (.A1(_06129_),
    .A2(_06131_),
    .B(_06250_),
    .Y(_06253_));
 NAND2x1_ASAP7_75t_R _35814_ (.A(_06252_),
    .B(_06253_),
    .Y(_06254_));
 NOR2x2_ASAP7_75t_R _35815_ (.A(net1603),
    .B(_06096_),
    .Y(_06256_));
 TAPCELL_ASAP7_75t_R PHY_358 ();
 OAI21x1_ASAP7_75t_R _35817_ (.A1(net2856),
    .A2(_06256_),
    .B(_06251_),
    .Y(_06258_));
 NOR2x2_ASAP7_75t_R _35818_ (.A(net1603),
    .B(net3424),
    .Y(_06259_));
 NAND2x1_ASAP7_75t_R _35819_ (.A(_06259_),
    .B(_06251_),
    .Y(_06260_));
 NOR2x2_ASAP7_75t_R _35820_ (.A(_06029_),
    .B(_06098_),
    .Y(_06261_));
 NAND2x1_ASAP7_75t_R _35821_ (.A(_06261_),
    .B(_06251_),
    .Y(_06262_));
 NAND3x1_ASAP7_75t_R _35822_ (.A(_06258_),
    .B(_06260_),
    .C(_06262_),
    .Y(_06263_));
 NOR2x1_ASAP7_75t_R _35823_ (.A(_06254_),
    .B(_06263_),
    .Y(_06264_));
 TAPCELL_ASAP7_75t_R PHY_357 ();
 TAPCELL_ASAP7_75t_R PHY_356 ();
 NAND2x2_ASAP7_75t_R _35826_ (.A(_06228_),
    .B(_06043_),
    .Y(_06268_));
 AOI211x1_ASAP7_75t_R _35827_ (.A1(net1276),
    .A2(_06061_),
    .B(net1592),
    .C(_06268_),
    .Y(_06269_));
 INVx2_ASAP7_75t_R _35828_ (.A(_06085_),
    .Y(_06270_));
 TAPCELL_ASAP7_75t_R PHY_355 ();
 NOR2x1_ASAP7_75t_R _35830_ (.A(net1665),
    .B(_06141_),
    .Y(_06272_));
 INVx3_ASAP7_75t_R _35831_ (.A(_06268_),
    .Y(_06273_));
 OA21x2_ASAP7_75t_R _35832_ (.A1(_06270_),
    .A2(_06272_),
    .B(_06273_),
    .Y(_06274_));
 NOR2x1_ASAP7_75t_R _35833_ (.A(_06269_),
    .B(_06274_),
    .Y(_06275_));
 AO21x1_ASAP7_75t_R _35834_ (.A1(_06226_),
    .A2(_06219_),
    .B(_06268_),
    .Y(_06276_));
 NAND2x2_ASAP7_75t_R _35835_ (.A(_06030_),
    .B(net2507),
    .Y(_06278_));
 AO21x1_ASAP7_75t_R _35836_ (.A1(net1215),
    .A2(net1628),
    .B(_06268_),
    .Y(_06279_));
 AND2x2_ASAP7_75t_R _35837_ (.A(_06276_),
    .B(_06279_),
    .Y(_06280_));
 NAND2x1_ASAP7_75t_R _35838_ (.A(_06275_),
    .B(_06280_),
    .Y(_06281_));
 INVx1_ASAP7_75t_R _35839_ (.A(_06281_),
    .Y(_06282_));
 NAND2x1_ASAP7_75t_R _35840_ (.A(_06264_),
    .B(_06282_),
    .Y(_06283_));
 NOR2x2_ASAP7_75t_R _35841_ (.A(_06249_),
    .B(_06283_),
    .Y(_06284_));
 NAND2x2_ASAP7_75t_R _35842_ (.A(_06224_),
    .B(_06284_),
    .Y(_06285_));
 NOR2x2_ASAP7_75t_R _35843_ (.A(_06173_),
    .B(_06285_),
    .Y(_06286_));
 XOR2x1_ASAP7_75t_R _35844_ (.A(_06026_),
    .Y(_06287_),
    .B(_06286_));
 AOI21x1_ASAP7_75t_R _35845_ (.A1(_05696_),
    .A2(_05732_),
    .B(_06287_),
    .Y(_06289_));
 NOR2x2_ASAP7_75t_R _35846_ (.A(net3368),
    .B(_05693_),
    .Y(_06290_));
 AND2x4_ASAP7_75t_R _35847_ (.A(_05693_),
    .B(net3368),
    .Y(_06291_));
 OAI21x1_ASAP7_75t_R _35848_ (.A1(_06290_),
    .A2(_06291_),
    .B(_05715_),
    .Y(_06292_));
 INVx1_ASAP7_75t_R _35849_ (.A(_05728_),
    .Y(_06293_));
 NOR2x2_ASAP7_75t_R _35850_ (.A(_06293_),
    .B(_05693_),
    .Y(_06294_));
 NOR2x1_ASAP7_75t_R _35851_ (.A(net3368),
    .B(_05695_),
    .Y(_06295_));
 OAI21x1_ASAP7_75t_R _35852_ (.A1(_06294_),
    .A2(_06295_),
    .B(_05427_),
    .Y(_06296_));
 INVx1_ASAP7_75t_R _35853_ (.A(_06287_),
    .Y(_06297_));
 AOI21x1_ASAP7_75t_R _35854_ (.A1(_06292_),
    .A2(_06296_),
    .B(_06297_),
    .Y(_06298_));
 OAI21x1_ASAP7_75t_R _35855_ (.A1(_06289_),
    .A2(_06298_),
    .B(net394),
    .Y(_06300_));
 NAND2x1_ASAP7_75t_R _35856_ (.A(_05052_),
    .B(_06300_),
    .Y(_06301_));
 XOR2x1_ASAP7_75t_R _35857_ (.A(_06301_),
    .Y(_00105_),
    .B(_08779_));
 AND2x2_ASAP7_75t_R _35858_ (.A(net388),
    .B(_00850_),
    .Y(_06302_));
 TAPCELL_ASAP7_75t_R PHY_354 ();
 AO21x1_ASAP7_75t_R _35860_ (.A1(_05206_),
    .A2(net3102),
    .B(_05306_),
    .Y(_06304_));
 TAPCELL_ASAP7_75t_R PHY_353 ();
 AO21x1_ASAP7_75t_R _35862_ (.A1(net2126),
    .A2(net1091),
    .B(_05306_),
    .Y(_06306_));
 TAPCELL_ASAP7_75t_R PHY_352 ();
 TAPCELL_ASAP7_75t_R PHY_351 ();
 AO21x1_ASAP7_75t_R _35865_ (.A1(net1835),
    .A2(net1946),
    .B(_05306_),
    .Y(_06310_));
 AND3x1_ASAP7_75t_R _35866_ (.A(_06304_),
    .B(_06306_),
    .C(_06310_),
    .Y(_06311_));
 AOI211x1_ASAP7_75t_R _35867_ (.A1(net3436),
    .A2(_05068_),
    .B(_05153_),
    .C(_05177_),
    .Y(_06312_));
 INVx1_ASAP7_75t_R _35868_ (.A(_06312_),
    .Y(_06313_));
 AO21x1_ASAP7_75t_R _35869_ (.A1(net1835),
    .A2(_05345_),
    .B(_05153_),
    .Y(_06314_));
 AND3x1_ASAP7_75t_R _35870_ (.A(_06313_),
    .B(_05167_),
    .C(_06314_),
    .Y(_06315_));
 NAND2x1_ASAP7_75t_R _35871_ (.A(_06311_),
    .B(_06315_),
    .Y(_06316_));
 TAPCELL_ASAP7_75t_R PHY_350 ();
 AOI211x1_ASAP7_75t_R _35873_ (.A1(net3436),
    .A2(net1147),
    .B(_05215_),
    .C(_05090_),
    .Y(_06318_));
 AOI211x1_ASAP7_75t_R _35874_ (.A1(_05173_),
    .A2(_05420_),
    .B(_06318_),
    .C(_05291_),
    .Y(_06319_));
 NOR2x2_ASAP7_75t_R _35875_ (.A(net3097),
    .B(_05177_),
    .Y(_06321_));
 NAND2x1_ASAP7_75t_R _35876_ (.A(_05217_),
    .B(_05162_),
    .Y(_06322_));
 INVx1_ASAP7_75t_R _35877_ (.A(_06322_),
    .Y(_06323_));
 OAI21x1_ASAP7_75t_R _35878_ (.A1(_06321_),
    .A2(_06323_),
    .B(_05247_),
    .Y(_06324_));
 OA21x2_ASAP7_75t_R _35879_ (.A1(_05215_),
    .A2(_05122_),
    .B(_05234_),
    .Y(_06325_));
 NAND3x1_ASAP7_75t_R _35880_ (.A(_06319_),
    .B(_06324_),
    .C(_06325_),
    .Y(_06326_));
 NOR2x1_ASAP7_75t_R _35881_ (.A(_06316_),
    .B(_06326_),
    .Y(_06327_));
 NOR2x2_ASAP7_75t_R _35882_ (.A(net1522),
    .B(net3455),
    .Y(_06328_));
 OA21x2_ASAP7_75t_R _35883_ (.A1(_05173_),
    .A2(_05151_),
    .B(_05175_),
    .Y(_06329_));
 AOI211x1_ASAP7_75t_R _35884_ (.A1(net1304),
    .A2(_06328_),
    .B(_06329_),
    .C(_05272_),
    .Y(_06330_));
 TAPCELL_ASAP7_75t_R PHY_349 ();
 OR3x1_ASAP7_75t_R _35886_ (.A(_05086_),
    .B(_05345_),
    .C(_05184_),
    .Y(_06333_));
 AO21x1_ASAP7_75t_R _35887_ (.A1(net2126),
    .A2(_05233_),
    .B(_05086_),
    .Y(_06334_));
 TAPCELL_ASAP7_75t_R PHY_348 ();
 TAPCELL_ASAP7_75t_R PHY_347 ();
 AO21x1_ASAP7_75t_R _35890_ (.A1(net1822),
    .A2(net3096),
    .B(_05086_),
    .Y(_06337_));
 AND3x1_ASAP7_75t_R _35891_ (.A(_06333_),
    .B(_06334_),
    .C(_06337_),
    .Y(_06338_));
 NAND2x1_ASAP7_75t_R _35892_ (.A(_06330_),
    .B(_06338_),
    .Y(_06339_));
 TAPCELL_ASAP7_75t_R PHY_346 ();
 AO21x1_ASAP7_75t_R _35894_ (.A1(net1822),
    .A2(_05211_),
    .B(net3108),
    .Y(_06341_));
 TAPCELL_ASAP7_75t_R PHY_345 ();
 TAPCELL_ASAP7_75t_R PHY_344 ();
 AO21x1_ASAP7_75t_R _35897_ (.A1(_05185_),
    .A2(net2645),
    .B(net3108),
    .Y(_06345_));
 INVx4_ASAP7_75t_R _35898_ (.A(net3096),
    .Y(_06346_));
 NAND2x2_ASAP7_75t_R _35899_ (.A(_06346_),
    .B(_05171_),
    .Y(_06347_));
 AND3x2_ASAP7_75t_R _35900_ (.A(_06341_),
    .B(_06345_),
    .C(_06347_),
    .Y(_06348_));
 NAND2x1_ASAP7_75t_R _35901_ (.A(net2225),
    .B(_05108_),
    .Y(_06349_));
 TAPCELL_ASAP7_75t_R PHY_343 ();
 AO21x1_ASAP7_75t_R _35903_ (.A1(net1403),
    .A2(net1945),
    .B(_05107_),
    .Y(_06351_));
 NAND2x1_ASAP7_75t_R _35904_ (.A(_06349_),
    .B(_06351_),
    .Y(_06352_));
 TAPCELL_ASAP7_75t_R PHY_342 ();
 AO21x1_ASAP7_75t_R _35906_ (.A1(net3446),
    .A2(net3105),
    .B(_05107_),
    .Y(_06355_));
 AO21x1_ASAP7_75t_R _35907_ (.A1(net3449),
    .A2(_05271_),
    .B(_05107_),
    .Y(_06356_));
 NAND2x1_ASAP7_75t_R _35908_ (.A(_06355_),
    .B(_06356_),
    .Y(_06357_));
 NOR2x2_ASAP7_75t_R _35909_ (.A(_06352_),
    .B(_06357_),
    .Y(_06358_));
 TAPCELL_ASAP7_75t_R PHY_341 ();
 AO21x1_ASAP7_75t_R _35911_ (.A1(_05206_),
    .A2(net1237),
    .B(net2493),
    .Y(_06360_));
 NAND3x2_ASAP7_75t_R _35912_ (.B(_06358_),
    .C(_06360_),
    .Y(_06361_),
    .A(_06348_));
 NOR2x2_ASAP7_75t_R _35913_ (.A(_06339_),
    .B(_06361_),
    .Y(_06362_));
 NAND2x2_ASAP7_75t_R _35914_ (.A(_06327_),
    .B(_06362_),
    .Y(_06363_));
 AO21x1_ASAP7_75t_R _35915_ (.A1(net1822),
    .A2(net1877),
    .B(_05208_),
    .Y(_06365_));
 OAI21x1_ASAP7_75t_R _35916_ (.A1(net964),
    .A2(_05208_),
    .B(_06365_),
    .Y(_06366_));
 TAPCELL_ASAP7_75t_R PHY_340 ();
 OAI21x1_ASAP7_75t_R _35918_ (.A1(_05208_),
    .A2(net2146),
    .B(_05263_),
    .Y(_06368_));
 TAPCELL_ASAP7_75t_R PHY_339 ();
 AO21x1_ASAP7_75t_R _35920_ (.A1(_05360_),
    .A2(_05345_),
    .B(_05198_),
    .Y(_06370_));
 TAPCELL_ASAP7_75t_R PHY_338 ();
 AO21x1_ASAP7_75t_R _35922_ (.A1(net3440),
    .A2(net2149),
    .B(_05198_),
    .Y(_06372_));
 NAND2x1_ASAP7_75t_R _35923_ (.A(_06370_),
    .B(_06372_),
    .Y(_06373_));
 OR3x1_ASAP7_75t_R _35924_ (.A(_06366_),
    .B(_06368_),
    .C(_06373_),
    .Y(_06374_));
 AO21x1_ASAP7_75t_R _35925_ (.A1(net3101),
    .A2(_05143_),
    .B(_05256_),
    .Y(_06376_));
 TAPCELL_ASAP7_75t_R PHY_337 ();
 AO21x1_ASAP7_75t_R _35927_ (.A1(_05360_),
    .A2(net1793),
    .B(_05256_),
    .Y(_06378_));
 NOR2x1_ASAP7_75t_R _35928_ (.A(net1768),
    .B(_05256_),
    .Y(_06379_));
 INVx1_ASAP7_75t_R _35929_ (.A(_06379_),
    .Y(_06380_));
 NAND3x1_ASAP7_75t_R _35930_ (.A(_06376_),
    .B(_06378_),
    .C(_06380_),
    .Y(_06381_));
 TAPCELL_ASAP7_75t_R PHY_336 ();
 AO31x2_ASAP7_75t_R _35932_ (.A1(_05206_),
    .A2(net1091),
    .A3(net2146),
    .B(_05240_),
    .Y(_06383_));
 AO21x1_ASAP7_75t_R _35933_ (.A1(net3426),
    .A2(net1793),
    .B(_05240_),
    .Y(_06384_));
 AO21x1_ASAP7_75t_R _35934_ (.A1(net992),
    .A2(net1944),
    .B(_05240_),
    .Y(_06385_));
 NAND3x1_ASAP7_75t_R _35935_ (.A(_06383_),
    .B(_06384_),
    .C(_06385_),
    .Y(_06387_));
 OR2x2_ASAP7_75t_R _35936_ (.A(_06381_),
    .B(_06387_),
    .Y(_06388_));
 NOR2x1_ASAP7_75t_R _35937_ (.A(_06374_),
    .B(_06388_),
    .Y(_06389_));
 TAPCELL_ASAP7_75t_R PHY_335 ();
 TAPCELL_ASAP7_75t_R PHY_334 ();
 AO21x1_ASAP7_75t_R _35940_ (.A1(net1766),
    .A2(net2149),
    .B(_05138_),
    .Y(_06392_));
 AO21x1_ASAP7_75t_R _35941_ (.A1(net1944),
    .A2(net2644),
    .B(_05138_),
    .Y(_06393_));
 INVx1_ASAP7_75t_R _35942_ (.A(_05138_),
    .Y(_06394_));
 NAND2x1_ASAP7_75t_R _35943_ (.A(_06394_),
    .B(_05096_),
    .Y(_06395_));
 AND3x1_ASAP7_75t_R _35944_ (.A(_06392_),
    .B(_06393_),
    .C(_06395_),
    .Y(_06396_));
 AO21x1_ASAP7_75t_R _35945_ (.A1(net1877),
    .A2(_05360_),
    .B(_05118_),
    .Y(_06398_));
 AO21x1_ASAP7_75t_R _35946_ (.A1(_05185_),
    .A2(net2643),
    .B(_05118_),
    .Y(_06399_));
 NAND2x1_ASAP7_75t_R _35947_ (.A(_05191_),
    .B(_05201_),
    .Y(_06400_));
 AND3x1_ASAP7_75t_R _35948_ (.A(_06398_),
    .B(_06399_),
    .C(_06400_),
    .Y(_06401_));
 NAND2x2_ASAP7_75t_R _35949_ (.A(_06396_),
    .B(_06401_),
    .Y(_06402_));
 AOI211x1_ASAP7_75t_R _35950_ (.A1(net1324),
    .A2(net1153),
    .B(net3410),
    .C(net2274),
    .Y(_06403_));
 OA21x2_ASAP7_75t_R _35951_ (.A1(_05203_),
    .A2(_05218_),
    .B(_05127_),
    .Y(_06404_));
 NOR2x1_ASAP7_75t_R _35952_ (.A(_06403_),
    .B(_06404_),
    .Y(_06405_));
 AO21x1_ASAP7_75t_R _35953_ (.A1(net3454),
    .A2(net964),
    .B(net3410),
    .Y(_06406_));
 OA21x2_ASAP7_75t_R _35954_ (.A1(_05128_),
    .A2(net3445),
    .B(_06406_),
    .Y(_06407_));
 NAND2x2_ASAP7_75t_R _35955_ (.A(_06405_),
    .B(_06407_),
    .Y(_06409_));
 TAPCELL_ASAP7_75t_R PHY_333 ();
 AO31x2_ASAP7_75t_R _35957_ (.A1(_05259_),
    .A2(net2027),
    .A3(net3454),
    .B(_05062_),
    .Y(_06411_));
 AO21x1_ASAP7_75t_R _35958_ (.A1(_05206_),
    .A2(net1140),
    .B(_05062_),
    .Y(_06412_));
 TAPCELL_ASAP7_75t_R PHY_332 ();
 AO21x1_ASAP7_75t_R _35960_ (.A1(net1768),
    .A2(net1237),
    .B(_05062_),
    .Y(_06414_));
 NAND3x2_ASAP7_75t_R _35961_ (.B(_06412_),
    .C(_06414_),
    .Y(_06415_),
    .A(_06411_));
 NOR3x2_ASAP7_75t_R _35962_ (.B(_06409_),
    .C(_06415_),
    .Y(_06416_),
    .A(_06402_));
 NAND2x2_ASAP7_75t_R _35963_ (.A(_06389_),
    .B(_06416_),
    .Y(_06417_));
 NOR2x1_ASAP7_75t_R _35964_ (.A(_06363_),
    .B(_06417_),
    .Y(_06418_));
 NAND2x2_ASAP7_75t_R _35965_ (.A(_05329_),
    .B(_06418_),
    .Y(_06420_));
 AOI21x1_ASAP7_75t_R _35966_ (.A1(_05430_),
    .A2(_05428_),
    .B(net3435),
    .Y(_06421_));
 NOR3x2_ASAP7_75t_R _35967_ (.B(net3437),
    .C(_06417_),
    .Y(_06422_),
    .A(net3353));
 AOI21x1_ASAP7_75t_R _35968_ (.A1(_05731_),
    .A2(_05729_),
    .B(_06422_),
    .Y(_06423_));
 NOR2x1_ASAP7_75t_R _35969_ (.A(_06421_),
    .B(_06423_),
    .Y(_06424_));
 NOR3x2_ASAP7_75t_R _35970_ (.B(_05734_),
    .C(_05789_),
    .Y(_06425_),
    .A(_05791_));
 NAND2x2_ASAP7_75t_R _35971_ (.A(_05755_),
    .B(_05816_),
    .Y(_06426_));
 NAND2x2_ASAP7_75t_R _35972_ (.A(_05844_),
    .B(net2489),
    .Y(_06427_));
 AO21x1_ASAP7_75t_R _35973_ (.A1(_06426_),
    .A2(_06427_),
    .B(_05821_),
    .Y(_06428_));
 NAND2x2_ASAP7_75t_R _35974_ (.A(_05803_),
    .B(_05766_),
    .Y(_06429_));
 TAPCELL_ASAP7_75t_R PHY_331 ();
 TAPCELL_ASAP7_75t_R PHY_330 ();
 TAPCELL_ASAP7_75t_R PHY_329 ();
 AO31x2_ASAP7_75t_R _35978_ (.A1(net1037),
    .A2(net2423),
    .A3(net2737),
    .B(_05821_),
    .Y(_06434_));
 NAND2x1_ASAP7_75t_R _35979_ (.A(_06428_),
    .B(_06434_),
    .Y(_06435_));
 NOR2x2_ASAP7_75t_R _35980_ (.A(net1775),
    .B(net2183),
    .Y(_06436_));
 NOR2x1_ASAP7_75t_R _35981_ (.A(_05897_),
    .B(_06436_),
    .Y(_06437_));
 AO21x1_ASAP7_75t_R _35982_ (.A1(_06437_),
    .A2(net2485),
    .B(_05800_),
    .Y(_06438_));
 NOR2x1_ASAP7_75t_R _35983_ (.A(net2230),
    .B(_05800_),
    .Y(_06439_));
 AOI211x1_ASAP7_75t_R _35984_ (.A1(net1224),
    .A2(_05755_),
    .B(_05800_),
    .C(_05957_),
    .Y(_06440_));
 NOR2x1_ASAP7_75t_R _35985_ (.A(_06439_),
    .B(_06440_),
    .Y(_06442_));
 NAND2x1_ASAP7_75t_R _35986_ (.A(_06438_),
    .B(_06442_),
    .Y(_06443_));
 NOR2x1_ASAP7_75t_R _35987_ (.A(_06435_),
    .B(_06443_),
    .Y(_06444_));
 AOI21x1_ASAP7_75t_R _35988_ (.A1(_05905_),
    .A2(net1560),
    .B(_05839_),
    .Y(_06445_));
 NOR2x1_ASAP7_75t_R _35989_ (.A(_05839_),
    .B(net2098),
    .Y(_06446_));
 NOR2x2_ASAP7_75t_R _35990_ (.A(_05839_),
    .B(_05876_),
    .Y(_06447_));
 OR3x1_ASAP7_75t_R _35991_ (.A(_06445_),
    .B(_06446_),
    .C(_06447_),
    .Y(_06448_));
 NAND2x2_ASAP7_75t_R _35992_ (.A(net1222),
    .B(net3474),
    .Y(_06449_));
 TAPCELL_ASAP7_75t_R PHY_328 ();
 AOI21x1_ASAP7_75t_R _35994_ (.A1(_06449_),
    .A2(net1807),
    .B(_05854_),
    .Y(_06451_));
 AO21x1_ASAP7_75t_R _35995_ (.A1(_05929_),
    .A2(_05844_),
    .B(_05957_),
    .Y(_06453_));
 NOR2x1_ASAP7_75t_R _35996_ (.A(_05854_),
    .B(_06453_),
    .Y(_06454_));
 NOR2x1_ASAP7_75t_R _35997_ (.A(_06451_),
    .B(_06454_),
    .Y(_06455_));
 OAI21x1_ASAP7_75t_R _35998_ (.A1(net1913),
    .A2(net2679),
    .B(_06455_),
    .Y(_06456_));
 NOR2x1_ASAP7_75t_R _35999_ (.A(_06448_),
    .B(_06456_),
    .Y(_06457_));
 NAND2x2_ASAP7_75t_R _36000_ (.A(_06444_),
    .B(_06457_),
    .Y(_06458_));
 NOR2x1_ASAP7_75t_R _36001_ (.A(net2185),
    .B(_05894_),
    .Y(_06459_));
 AO21x2_ASAP7_75t_R _36002_ (.A1(_06459_),
    .A2(_05810_),
    .B(_05899_),
    .Y(_06460_));
 NAND2x2_ASAP7_75t_R _36003_ (.A(_05976_),
    .B(_05898_),
    .Y(_06461_));
 AO21x1_ASAP7_75t_R _36004_ (.A1(net1662),
    .A2(net1037),
    .B(_05894_),
    .Y(_06462_));
 NAND2x2_ASAP7_75t_R _36005_ (.A(_06461_),
    .B(_06462_),
    .Y(_06464_));
 AO21x1_ASAP7_75t_R _36006_ (.A1(net1786),
    .A2(_05957_),
    .B(_05908_),
    .Y(_06465_));
 AO21x1_ASAP7_75t_R _36007_ (.A1(_05817_),
    .A2(_05876_),
    .B(_05908_),
    .Y(_06466_));
 NAND2x2_ASAP7_75t_R _36008_ (.A(_06465_),
    .B(_06466_),
    .Y(_06467_));
 NOR3x2_ASAP7_75t_R _36009_ (.B(_06464_),
    .C(_06467_),
    .Y(_06468_),
    .A(_06460_));
 AO21x1_ASAP7_75t_R _36010_ (.A1(net1118),
    .A2(net980),
    .B(_05873_),
    .Y(_06469_));
 AO21x1_ASAP7_75t_R _36011_ (.A1(net2876),
    .A2(net2229),
    .B(_05873_),
    .Y(_06470_));
 NAND2x1_ASAP7_75t_R _36012_ (.A(_06469_),
    .B(_06470_),
    .Y(_06471_));
 NOR2x2_ASAP7_75t_R _36013_ (.A(_05810_),
    .B(net2184),
    .Y(_06472_));
 NAND2x1_ASAP7_75t_R _36014_ (.A(_06472_),
    .B(_05878_),
    .Y(_06473_));
 TAPCELL_ASAP7_75t_R PHY_327 ();
 AO21x1_ASAP7_75t_R _36016_ (.A1(_05857_),
    .A2(_05817_),
    .B(_05873_),
    .Y(_06476_));
 NAND2x1_ASAP7_75t_R _36017_ (.A(_06473_),
    .B(_06476_),
    .Y(_06477_));
 NOR2x1_ASAP7_75t_R _36018_ (.A(_06477_),
    .B(_06471_),
    .Y(_06478_));
 AO21x1_ASAP7_75t_R _36019_ (.A1(net3467),
    .A2(_05835_),
    .B(_05884_),
    .Y(_06479_));
 AO21x1_ASAP7_75t_R _36020_ (.A1(net1786),
    .A2(net1560),
    .B(_05884_),
    .Y(_06480_));
 INVx4_ASAP7_75t_R _36021_ (.A(_05819_),
    .Y(_06481_));
 NAND2x1_ASAP7_75t_R _36022_ (.A(_06481_),
    .B(_05885_),
    .Y(_06482_));
 AND3x1_ASAP7_75t_R _36023_ (.A(_06479_),
    .B(_06480_),
    .C(_06482_),
    .Y(_06483_));
 NAND2x2_ASAP7_75t_R _36024_ (.A(_06478_),
    .B(_06483_),
    .Y(_06484_));
 INVx2_ASAP7_75t_R _36025_ (.A(_06484_),
    .Y(_06486_));
 NAND2x1_ASAP7_75t_R _36026_ (.A(_06468_),
    .B(_06486_),
    .Y(_06487_));
 NOR2x1_ASAP7_75t_R _36027_ (.A(_06458_),
    .B(_06487_),
    .Y(_06488_));
 OAI21x1_ASAP7_75t_R _36028_ (.A1(_05759_),
    .A2(_05743_),
    .B(_05751_),
    .Y(_06489_));
 NAND2x2_ASAP7_75t_R _36029_ (.A(_05764_),
    .B(net3475),
    .Y(_06490_));
 AO21x1_ASAP7_75t_R _36030_ (.A1(_06490_),
    .A2(_05957_),
    .B(_05752_),
    .Y(_06491_));
 NAND2x2_ASAP7_75t_R _36031_ (.A(_06489_),
    .B(_06491_),
    .Y(_06492_));
 NAND2x1_ASAP7_75t_R _36032_ (.A(_06015_),
    .B(_05926_),
    .Y(_06493_));
 NOR2x2_ASAP7_75t_R _36033_ (.A(_05810_),
    .B(net2540),
    .Y(_06494_));
 OAI21x1_ASAP7_75t_R _36034_ (.A1(_06494_),
    .A2(_05930_),
    .B(_05926_),
    .Y(_06495_));
 NAND2x2_ASAP7_75t_R _36035_ (.A(_06493_),
    .B(_06495_),
    .Y(_06497_));
 NAND2x1_ASAP7_75t_R _36036_ (.A(_05964_),
    .B(_05926_),
    .Y(_06498_));
 OAI21x1_ASAP7_75t_R _36037_ (.A1(_05845_),
    .A2(_06472_),
    .B(_05926_),
    .Y(_06499_));
 NAND2x2_ASAP7_75t_R _36038_ (.A(_06498_),
    .B(_06499_),
    .Y(_06500_));
 NOR3x2_ASAP7_75t_R _36039_ (.B(_06497_),
    .C(_06500_),
    .Y(_06501_),
    .A(_06492_));
 NAND2x2_ASAP7_75t_R _36040_ (.A(_06436_),
    .B(_05953_),
    .Y(_06502_));
 NAND2x2_ASAP7_75t_R _36041_ (.A(_06502_),
    .B(_05954_),
    .Y(_06503_));
 AOI211x1_ASAP7_75t_R _36042_ (.A1(_05764_),
    .A2(net1774),
    .B(net3352),
    .C(_05775_),
    .Y(_06504_));
 AOI211x1_ASAP7_75t_R _36043_ (.A1(_05764_),
    .A2(_05755_),
    .B(net3352),
    .C(_05957_),
    .Y(_06505_));
 NOR3x2_ASAP7_75t_R _36044_ (.B(_06504_),
    .C(_06505_),
    .Y(_06506_),
    .A(_06503_));
 AO21x1_ASAP7_75t_R _36045_ (.A1(_05817_),
    .A2(_05860_),
    .B(_05938_),
    .Y(_06508_));
 INVx2_ASAP7_75t_R _36046_ (.A(_05938_),
    .Y(_06509_));
 NAND2x2_ASAP7_75t_R _36047_ (.A(net2359),
    .B(_06509_),
    .Y(_06510_));
 NAND2x1_ASAP7_75t_R _36048_ (.A(_05897_),
    .B(_06509_),
    .Y(_06511_));
 AND3x2_ASAP7_75t_R _36049_ (.A(_06508_),
    .B(_06510_),
    .C(_06511_),
    .Y(_06512_));
 NAND3x1_ASAP7_75t_R _36050_ (.A(_06501_),
    .B(_06506_),
    .C(_06512_),
    .Y(_06513_));
 AO21x1_ASAP7_75t_R _36051_ (.A1(net2422),
    .A2(_05887_),
    .B(_05977_),
    .Y(_06514_));
 INVx2_ASAP7_75t_R _36052_ (.A(_06449_),
    .Y(_06515_));
 OAI21x1_ASAP7_75t_R _36053_ (.A1(_06494_),
    .A2(_06515_),
    .B(_05978_),
    .Y(_06516_));
 NOR2x2_ASAP7_75t_R _36054_ (.A(net2183),
    .B(_05929_),
    .Y(_06517_));
 OAI21x1_ASAP7_75t_R _36055_ (.A1(_05897_),
    .A2(net2404),
    .B(_05978_),
    .Y(_06519_));
 NAND3x2_ASAP7_75t_R _36056_ (.B(_06516_),
    .C(_06519_),
    .Y(_06520_),
    .A(_06514_));
 INVx3_ASAP7_75t_R _36057_ (.A(net3370),
    .Y(_06521_));
 OAI21x1_ASAP7_75t_R _36058_ (.A1(_06521_),
    .A2(_06015_),
    .B(_05966_),
    .Y(_06522_));
 NOR2x2_ASAP7_75t_R _36059_ (.A(_05757_),
    .B(net2540),
    .Y(_06523_));
 OAI21x1_ASAP7_75t_R _36060_ (.A1(_05776_),
    .A2(_06523_),
    .B(_05966_),
    .Y(_06524_));
 NAND2x2_ASAP7_75t_R _36061_ (.A(net2636),
    .B(_05931_),
    .Y(_06525_));
 NAND3x2_ASAP7_75t_R _36062_ (.B(_06524_),
    .C(_06525_),
    .Y(_06526_),
    .A(_06522_));
 NAND2x2_ASAP7_75t_R _36063_ (.A(net2636),
    .B(net2360),
    .Y(_06527_));
 NAND2x2_ASAP7_75t_R _36064_ (.A(_05985_),
    .B(_05966_),
    .Y(_06528_));
 NAND2x2_ASAP7_75t_R _36065_ (.A(_05966_),
    .B(net2519),
    .Y(_06530_));
 NAND3x2_ASAP7_75t_R _36066_ (.B(_06528_),
    .C(_06530_),
    .Y(_06531_),
    .A(_06527_));
 NOR3x1_ASAP7_75t_R _36067_ (.A(_06520_),
    .B(_06526_),
    .C(_06531_),
    .Y(_06532_));
 NAND2x1_ASAP7_75t_R _36068_ (.A(_06017_),
    .B(_06015_),
    .Y(_06533_));
 AO21x1_ASAP7_75t_R _36069_ (.A1(net1037),
    .A2(net2229),
    .B(_06007_),
    .Y(_06534_));
 NAND2x1_ASAP7_75t_R _36070_ (.A(_06533_),
    .B(_06534_),
    .Y(_06535_));
 AO21x2_ASAP7_75t_R _36071_ (.A1(_05833_),
    .A2(_05835_),
    .B(_06007_),
    .Y(_06536_));
 AO21x1_ASAP7_75t_R _36072_ (.A1(net1913),
    .A2(_05850_),
    .B(_06007_),
    .Y(_06537_));
 NAND2x1_ASAP7_75t_R _36073_ (.A(_06536_),
    .B(_06537_),
    .Y(_06538_));
 NOR2x1_ASAP7_75t_R _36074_ (.A(_06535_),
    .B(_06538_),
    .Y(_06539_));
 NOR2x1_ASAP7_75t_R _36075_ (.A(_05957_),
    .B(_05993_),
    .Y(_06541_));
 NAND2x1_ASAP7_75t_R _36076_ (.A(_05844_),
    .B(_06541_),
    .Y(_06542_));
 AO21x1_ASAP7_75t_R _36077_ (.A1(_05850_),
    .A2(_06426_),
    .B(_05993_),
    .Y(_06543_));
 AO21x1_ASAP7_75t_R _36078_ (.A1(net1662),
    .A2(net1807),
    .B(_05993_),
    .Y(_06544_));
 AND3x1_ASAP7_75t_R _36079_ (.A(_06542_),
    .B(_06543_),
    .C(_06544_),
    .Y(_06545_));
 NAND2x1_ASAP7_75t_R _36080_ (.A(_06539_),
    .B(_06545_),
    .Y(_06546_));
 INVx1_ASAP7_75t_R _36081_ (.A(_06546_),
    .Y(_06547_));
 NAND2x1_ASAP7_75t_R _36082_ (.A(_06532_),
    .B(_06547_),
    .Y(_06548_));
 NOR2x1_ASAP7_75t_R _36083_ (.A(_06513_),
    .B(_06548_),
    .Y(_06549_));
 NAND2x1_ASAP7_75t_R _36084_ (.A(_06488_),
    .B(_06549_),
    .Y(_06550_));
 NOR2x2_ASAP7_75t_R _36085_ (.A(_06425_),
    .B(_06550_),
    .Y(_06552_));
 AO21x1_ASAP7_75t_R _36086_ (.A1(net2033),
    .A2(net2611),
    .B(_05683_),
    .Y(_06553_));
 TAPCELL_ASAP7_75t_R PHY_326 ();
 AO21x1_ASAP7_75t_R _36088_ (.A1(net2698),
    .A2(net2548),
    .B(_05683_),
    .Y(_06555_));
 NAND2x1_ASAP7_75t_R _36089_ (.A(_06553_),
    .B(_06555_),
    .Y(_06556_));
 NAND2x1_ASAP7_75t_R _36090_ (.A(net3450),
    .B(_05684_),
    .Y(_06557_));
 AO21x1_ASAP7_75t_R _36091_ (.A1(net3356),
    .A2(_05613_),
    .B(_05683_),
    .Y(_06558_));
 NAND2x1_ASAP7_75t_R _36092_ (.A(_06557_),
    .B(_06558_),
    .Y(_06559_));
 NOR2x1_ASAP7_75t_R _36093_ (.A(_06556_),
    .B(_06559_),
    .Y(_06560_));
 AO21x1_ASAP7_75t_R _36094_ (.A1(_05462_),
    .A2(_05464_),
    .B(_05677_),
    .Y(_06561_));
 AO21x1_ASAP7_75t_R _36095_ (.A1(net2548),
    .A2(net2115),
    .B(_05677_),
    .Y(_06563_));
 NOR2x1_ASAP7_75t_R _36096_ (.A(_05677_),
    .B(net2703),
    .Y(_06564_));
 INVx1_ASAP7_75t_R _36097_ (.A(_06564_),
    .Y(_06565_));
 AND3x1_ASAP7_75t_R _36098_ (.A(_06561_),
    .B(_06563_),
    .C(_06565_),
    .Y(_06566_));
 NAND2x1_ASAP7_75t_R _36099_ (.A(_06560_),
    .B(_06566_),
    .Y(_06567_));
 NAND2x2_ASAP7_75t_R _36100_ (.A(net1312),
    .B(net2016),
    .Y(_06568_));
 TAPCELL_ASAP7_75t_R PHY_325 ();
 AO21x1_ASAP7_75t_R _36102_ (.A1(_05613_),
    .A2(_06568_),
    .B(_05654_),
    .Y(_06570_));
 AO21x1_ASAP7_75t_R _36103_ (.A1(net2115),
    .A2(_05457_),
    .B(_05654_),
    .Y(_06571_));
 AND2x2_ASAP7_75t_R _36104_ (.A(_06570_),
    .B(_06571_),
    .Y(_06572_));
 NAND2x2_ASAP7_75t_R _36105_ (.A(_05446_),
    .B(_05501_),
    .Y(_06574_));
 TAPCELL_ASAP7_75t_R PHY_324 ();
 NAND2x2_ASAP7_75t_R _36107_ (.A(_05653_),
    .B(_05625_),
    .Y(_06576_));
 TAPCELL_ASAP7_75t_R PHY_323 ();
 AO21x1_ASAP7_75t_R _36109_ (.A1(net2698),
    .A2(net2003),
    .B(_06576_),
    .Y(_06578_));
 TAPCELL_ASAP7_75t_R PHY_322 ();
 NOR2x1_ASAP7_75t_R _36111_ (.A(net2477),
    .B(_06576_),
    .Y(_06580_));
 INVx1_ASAP7_75t_R _36112_ (.A(_06580_),
    .Y(_06581_));
 OAI21x1_ASAP7_75t_R _36113_ (.A1(_05566_),
    .A2(_05669_),
    .B(_05661_),
    .Y(_06582_));
 AND3x1_ASAP7_75t_R _36114_ (.A(_06578_),
    .B(_06581_),
    .C(_06582_),
    .Y(_06583_));
 NAND2x1_ASAP7_75t_R _36115_ (.A(_06572_),
    .B(_06583_),
    .Y(_06585_));
 NOR2x1_ASAP7_75t_R _36116_ (.A(_06567_),
    .B(_06585_),
    .Y(_06586_));
 TAPCELL_ASAP7_75t_R PHY_321 ();
 AOI21x1_ASAP7_75t_R _36118_ (.A1(_05619_),
    .A2(net2003),
    .B(net2618),
    .Y(_06588_));
 OAI21x1_ASAP7_75t_R _36119_ (.A1(net2865),
    .A2(_05450_),
    .B(net1035),
    .Y(_06589_));
 NOR2x2_ASAP7_75t_R _36120_ (.A(_05640_),
    .B(_06589_),
    .Y(_06590_));
 AOI211x1_ASAP7_75t_R _36121_ (.A1(_05647_),
    .A2(net1528),
    .B(_06588_),
    .C(_06590_),
    .Y(_06591_));
 NOR2x2_ASAP7_75t_R _36122_ (.A(net3121),
    .B(net1666),
    .Y(_06592_));
 INVx3_ASAP7_75t_R _36123_ (.A(_05634_),
    .Y(_06593_));
 OA21x2_ASAP7_75t_R _36124_ (.A1(net1528),
    .A2(_06592_),
    .B(_06593_),
    .Y(_06594_));
 TAPCELL_ASAP7_75t_R PHY_320 ();
 NOR2x2_ASAP7_75t_R _36126_ (.A(net2461),
    .B(net3461),
    .Y(_06597_));
 AOI21x1_ASAP7_75t_R _36127_ (.A1(net2477),
    .A2(net2033),
    .B(net2461),
    .Y(_06598_));
 NOR3x2_ASAP7_75t_R _36128_ (.B(_06597_),
    .C(_06598_),
    .Y(_06599_),
    .A(_06594_));
 NAND2x2_ASAP7_75t_R _36129_ (.A(_06591_),
    .B(_06599_),
    .Y(_06600_));
 NOR2x1_ASAP7_75t_R _36130_ (.A(net2548),
    .B(_05626_),
    .Y(_06601_));
 OA21x2_ASAP7_75t_R _36131_ (.A1(_05682_),
    .A2(_05665_),
    .B(_05627_),
    .Y(_06602_));
 NOR2x1_ASAP7_75t_R _36132_ (.A(_06601_),
    .B(_06602_),
    .Y(_06603_));
 TAPCELL_ASAP7_75t_R PHY_319 ();
 AO21x1_ASAP7_75t_R _36134_ (.A1(net3356),
    .A2(net2816),
    .B(net2411),
    .Y(_06605_));
 TAPCELL_ASAP7_75t_R PHY_318 ();
 AO21x1_ASAP7_75t_R _36136_ (.A1(net2703),
    .A2(net2659),
    .B(net2411),
    .Y(_06608_));
 AND2x2_ASAP7_75t_R _36137_ (.A(_06605_),
    .B(_06608_),
    .Y(_06609_));
 NAND2x2_ASAP7_75t_R _36138_ (.A(_06603_),
    .B(_06609_),
    .Y(_06610_));
 TAPCELL_ASAP7_75t_R PHY_317 ();
 AO31x2_ASAP7_75t_R _36140_ (.A1(net2220),
    .A2(net2478),
    .A3(net1083),
    .B(net2447),
    .Y(_06612_));
 CKINVDCx8_ASAP7_75t_R _36141_ (.A(_05616_),
    .Y(_06613_));
 TAPCELL_ASAP7_75t_R PHY_316 ();
 AOI211x1_ASAP7_75t_R _36143_ (.A1(net1000),
    .A2(net989),
    .B(_05616_),
    .C(net1671),
    .Y(_06615_));
 AOI21x1_ASAP7_75t_R _36144_ (.A1(_06613_),
    .A2(_05568_),
    .B(_06615_),
    .Y(_06616_));
 NAND2x2_ASAP7_75t_R _36145_ (.A(_06612_),
    .B(_06616_),
    .Y(_06618_));
 NOR3x2_ASAP7_75t_R _36146_ (.B(_06610_),
    .C(_06618_),
    .Y(_06619_),
    .A(_06600_));
 NAND2x2_ASAP7_75t_R _36147_ (.A(_06586_),
    .B(_06619_),
    .Y(_06620_));
 AND3x2_ASAP7_75t_R _36148_ (.A(_05545_),
    .B(_05449_),
    .C(_05461_),
    .Y(_06621_));
 OA21x2_ASAP7_75t_R _36149_ (.A1(_05516_),
    .A2(_05441_),
    .B(_05545_),
    .Y(_06622_));
 OA21x2_ASAP7_75t_R _36150_ (.A1(net1528),
    .A2(_05674_),
    .B(_05545_),
    .Y(_06623_));
 NOR3x1_ASAP7_75t_R _36151_ (.A(_06621_),
    .B(_06622_),
    .C(_06623_),
    .Y(_06624_));
 TAPCELL_ASAP7_75t_R PHY_315 ();
 INVx1_ASAP7_75t_R _36153_ (.A(_06574_),
    .Y(_06626_));
 INVx5_ASAP7_75t_R _36154_ (.A(net3118),
    .Y(_06627_));
 TAPCELL_ASAP7_75t_R PHY_314 ();
 OA21x2_ASAP7_75t_R _36156_ (.A1(_06626_),
    .A2(_05514_),
    .B(_06627_),
    .Y(_06630_));
 AOI211x1_ASAP7_75t_R _36157_ (.A1(net1315),
    .A2(net1202),
    .B(_05528_),
    .C(_05457_),
    .Y(_06631_));
 OA21x2_ASAP7_75t_R _36158_ (.A1(_05674_),
    .A2(_05568_),
    .B(_06627_),
    .Y(_06632_));
 NOR3x1_ASAP7_75t_R _36159_ (.A(_06630_),
    .B(_06631_),
    .C(_06632_),
    .Y(_06633_));
 NAND2x1_ASAP7_75t_R _36160_ (.A(_06624_),
    .B(_06633_),
    .Y(_06634_));
 TAPCELL_ASAP7_75t_R PHY_313 ();
 AOI211x1_ASAP7_75t_R _36162_ (.A1(net2814),
    .A2(net3098),
    .B(_05492_),
    .C(net2091),
    .Y(_06636_));
 NOR2x2_ASAP7_75t_R _36163_ (.A(net1666),
    .B(_05519_),
    .Y(_06637_));
 OA21x2_ASAP7_75t_R _36164_ (.A1(_06637_),
    .A2(_05642_),
    .B(_05484_),
    .Y(_06638_));
 NOR2x1_ASAP7_75t_R _36165_ (.A(_05492_),
    .B(_06589_),
    .Y(_06640_));
 NOR3x1_ASAP7_75t_R _36166_ (.A(_06636_),
    .B(_06638_),
    .C(_06640_),
    .Y(_06641_));
 AO21x1_ASAP7_75t_R _36167_ (.A1(_05462_),
    .A2(net2815),
    .B(_05511_),
    .Y(_06642_));
 OA21x2_ASAP7_75t_R _36168_ (.A1(_05561_),
    .A2(_06592_),
    .B(net3373),
    .Y(_06643_));
 INVx1_ASAP7_75t_R _36169_ (.A(_06643_),
    .Y(_06644_));
 NAND2x1_ASAP7_75t_R _36170_ (.A(_06642_),
    .B(_06644_),
    .Y(_06645_));
 OAI21x1_ASAP7_75t_R _36171_ (.A1(_05516_),
    .A2(_05664_),
    .B(net3373),
    .Y(_06646_));
 NOR2x2_ASAP7_75t_R _36172_ (.A(_05500_),
    .B(net2092),
    .Y(_06647_));
 OAI21x1_ASAP7_75t_R _36173_ (.A1(_06647_),
    .A2(_05514_),
    .B(net3373),
    .Y(_06648_));
 NAND2x1_ASAP7_75t_R _36174_ (.A(net3373),
    .B(_05520_),
    .Y(_06649_));
 NAND3x1_ASAP7_75t_R _36175_ (.A(_06646_),
    .B(_06648_),
    .C(_06649_),
    .Y(_06651_));
 NOR2x1_ASAP7_75t_R _36176_ (.A(_06645_),
    .B(_06651_),
    .Y(_06652_));
 NAND2x1_ASAP7_75t_R _36177_ (.A(_06641_),
    .B(_06652_),
    .Y(_06653_));
 NOR2x1_ASAP7_75t_R _36178_ (.A(_06634_),
    .B(_06653_),
    .Y(_06654_));
 TAPCELL_ASAP7_75t_R PHY_312 ();
 AO21x1_ASAP7_75t_R _36180_ (.A1(net3249),
    .A2(net2836),
    .B(_05472_),
    .Y(_06656_));
 AO21x1_ASAP7_75t_R _36181_ (.A1(_05605_),
    .A2(net2035),
    .B(_05472_),
    .Y(_06657_));
 NAND2x1_ASAP7_75t_R _36182_ (.A(_05495_),
    .B(_05600_),
    .Y(_06658_));
 AND3x1_ASAP7_75t_R _36183_ (.A(_06656_),
    .B(_06657_),
    .C(_06658_),
    .Y(_06659_));
 OAI21x1_ASAP7_75t_R _36184_ (.A1(net2863),
    .A2(_05467_),
    .B(_05591_),
    .Y(_06660_));
 AOI211x1_ASAP7_75t_R _36185_ (.A1(_05435_),
    .A2(_05441_),
    .B(_06660_),
    .C(_05458_),
    .Y(_06662_));
 NAND2x1_ASAP7_75t_R _36186_ (.A(_06659_),
    .B(_06662_),
    .Y(_06663_));
 AOI211x1_ASAP7_75t_R _36187_ (.A1(net1000),
    .A2(net3111),
    .B(_05581_),
    .C(net1208),
    .Y(_06664_));
 INVx1_ASAP7_75t_R _36188_ (.A(_06664_),
    .Y(_06665_));
 AO21x2_ASAP7_75t_R _36189_ (.A1(net2835),
    .A2(_06568_),
    .B(_05581_),
    .Y(_06666_));
 AND2x2_ASAP7_75t_R _36190_ (.A(_06665_),
    .B(_06666_),
    .Y(_06667_));
 AO21x1_ASAP7_75t_R _36191_ (.A1(_05535_),
    .A2(_05503_),
    .B(net2389),
    .Y(_06668_));
 AND2x2_ASAP7_75t_R _36192_ (.A(_06668_),
    .B(_05569_),
    .Y(_06669_));
 AOI211x1_ASAP7_75t_R _36193_ (.A1(net2814),
    .A2(net3111),
    .B(net2389),
    .C(_05457_),
    .Y(_06670_));
 INVx2_ASAP7_75t_R _36194_ (.A(_05619_),
    .Y(_06671_));
 OA21x2_ASAP7_75t_R _36195_ (.A1(_06671_),
    .A2(_05520_),
    .B(_05564_),
    .Y(_06673_));
 NOR2x1_ASAP7_75t_R _36196_ (.A(_06670_),
    .B(_06673_),
    .Y(_06674_));
 NAND3x1_ASAP7_75t_R _36197_ (.A(_06667_),
    .B(_06669_),
    .C(_06674_),
    .Y(_06675_));
 NOR2x1_ASAP7_75t_R _36198_ (.A(_06663_),
    .B(_06675_),
    .Y(_06676_));
 NAND2x2_ASAP7_75t_R _36199_ (.A(_06654_),
    .B(_06676_),
    .Y(_06677_));
 NOR2x2_ASAP7_75t_R _36200_ (.A(_06620_),
    .B(_06677_),
    .Y(_06678_));
 NAND2x2_ASAP7_75t_R _36201_ (.A(_05479_),
    .B(_06678_),
    .Y(_06679_));
 NOR2x1_ASAP7_75t_R _36202_ (.A(_06552_),
    .B(_06679_),
    .Y(_06680_));
 AOI211x1_ASAP7_75t_R _36203_ (.A1(_05478_),
    .A2(net2113),
    .B(_06620_),
    .C(_06677_),
    .Y(_06681_));
 INVx1_ASAP7_75t_R _36204_ (.A(_06501_),
    .Y(_06682_));
 NAND2x1_ASAP7_75t_R _36205_ (.A(_06512_),
    .B(_06506_),
    .Y(_06684_));
 NOR2x1_ASAP7_75t_R _36206_ (.A(_06682_),
    .B(_06684_),
    .Y(_06685_));
 INVx1_ASAP7_75t_R _36207_ (.A(_06520_),
    .Y(_06686_));
 NOR2x1_ASAP7_75t_R _36208_ (.A(_06531_),
    .B(_06526_),
    .Y(_06687_));
 NAND2x1_ASAP7_75t_R _36209_ (.A(_06686_),
    .B(_06687_),
    .Y(_06688_));
 NOR2x1_ASAP7_75t_R _36210_ (.A(_06546_),
    .B(_06688_),
    .Y(_06689_));
 NAND2x1_ASAP7_75t_R _36211_ (.A(_06685_),
    .B(_06689_),
    .Y(_06690_));
 INVx1_ASAP7_75t_R _36212_ (.A(_06468_),
    .Y(_06691_));
 NOR2x1_ASAP7_75t_R _36213_ (.A(_06484_),
    .B(_06691_),
    .Y(_06692_));
 INVx1_ASAP7_75t_R _36214_ (.A(_06458_),
    .Y(_06693_));
 NAND2x1_ASAP7_75t_R _36215_ (.A(_06692_),
    .B(_06693_),
    .Y(_06695_));
 NOR2x1_ASAP7_75t_R _36216_ (.A(_06695_),
    .B(_06690_),
    .Y(_06696_));
 NAND2x2_ASAP7_75t_R _36217_ (.A(_05794_),
    .B(_06696_),
    .Y(_06697_));
 NOR2x1_ASAP7_75t_R _36218_ (.A(net1927),
    .B(_06697_),
    .Y(_06698_));
 INVx1_ASAP7_75t_R _36219_ (.A(_06055_),
    .Y(_06699_));
 NAND2x1_ASAP7_75t_R _36220_ (.A(_06075_),
    .B(_06066_),
    .Y(_06700_));
 NOR2x1_ASAP7_75t_R _36221_ (.A(_06700_),
    .B(_06699_),
    .Y(_06701_));
 TAPCELL_ASAP7_75t_R PHY_311 ();
 AO21x1_ASAP7_75t_R _36223_ (.A1(_06099_),
    .A2(_06072_),
    .B(_06104_),
    .Y(_06703_));
 NOR2x1_ASAP7_75t_R _36224_ (.A(_06113_),
    .B(_06110_),
    .Y(_06704_));
 NAND2x1_ASAP7_75t_R _36225_ (.A(_06703_),
    .B(_06704_),
    .Y(_06706_));
 NOR2x1_ASAP7_75t_R _36226_ (.A(_06094_),
    .B(_06706_),
    .Y(_06707_));
 NAND2x2_ASAP7_75t_R _36227_ (.A(_06701_),
    .B(_06707_),
    .Y(_06708_));
 NOR3x1_ASAP7_75t_R _36228_ (.A(_06169_),
    .B(_06155_),
    .C(_06164_),
    .Y(_06709_));
 NAND2x2_ASAP7_75t_R _36229_ (.A(_06043_),
    .B(_06120_),
    .Y(_06710_));
 OR3x2_ASAP7_75t_R _36230_ (.A(_06710_),
    .B(net1603),
    .C(net1758),
    .Y(_06711_));
 INVx1_ASAP7_75t_R _36231_ (.A(_06144_),
    .Y(_06712_));
 NAND2x1_ASAP7_75t_R _36232_ (.A(_06138_),
    .B(_06139_),
    .Y(_06713_));
 NAND3x1_ASAP7_75t_R _36233_ (.A(_06711_),
    .B(_06712_),
    .C(_06713_),
    .Y(_06714_));
 NOR2x1_ASAP7_75t_R _36234_ (.A(_06135_),
    .B(_06714_),
    .Y(_06715_));
 NAND2x1_ASAP7_75t_R _36235_ (.A(_06709_),
    .B(_06715_),
    .Y(_06717_));
 NOR2x1_ASAP7_75t_R _36236_ (.A(_06717_),
    .B(_06708_),
    .Y(_06718_));
 INVx1_ASAP7_75t_R _36237_ (.A(_06254_),
    .Y(_06719_));
 INVx1_ASAP7_75t_R _36238_ (.A(_06263_),
    .Y(_06720_));
 NAND2x1_ASAP7_75t_R _36239_ (.A(_06719_),
    .B(_06720_),
    .Y(_06721_));
 NOR2x1_ASAP7_75t_R _36240_ (.A(_06281_),
    .B(_06721_),
    .Y(_06722_));
 NAND2x1_ASAP7_75t_R _36241_ (.A(_06248_),
    .B(_06722_),
    .Y(_06723_));
 INVx1_ASAP7_75t_R _36242_ (.A(_06201_),
    .Y(_06724_));
 INVx1_ASAP7_75t_R _36243_ (.A(_06223_),
    .Y(_06725_));
 NAND2x1_ASAP7_75t_R _36244_ (.A(_06724_),
    .B(_06725_),
    .Y(_06726_));
 NOR2x1_ASAP7_75t_R _36245_ (.A(_06723_),
    .B(_06726_),
    .Y(_06728_));
 NAND2x2_ASAP7_75t_R _36246_ (.A(_06718_),
    .B(_06728_),
    .Y(_06729_));
 TAPCELL_ASAP7_75t_R PHY_310 ();
 AOI21x1_ASAP7_75t_R _36248_ (.A1(net2764),
    .A2(net2399),
    .B(net1217),
    .Y(_06731_));
 NAND2x2_ASAP7_75t_R _36249_ (.A(net3422),
    .B(net1295),
    .Y(_06732_));
 AOI21x1_ASAP7_75t_R _36250_ (.A1(_06732_),
    .A2(_06226_),
    .B(_06191_),
    .Y(_06733_));
 TAPCELL_ASAP7_75t_R PHY_309 ();
 NOR2x1_ASAP7_75t_R _36252_ (.A(net2764),
    .B(_06078_),
    .Y(_06735_));
 AOI211x1_ASAP7_75t_R _36253_ (.A1(_06731_),
    .A2(_06042_),
    .B(_06733_),
    .C(_06735_),
    .Y(_06736_));
 TAPCELL_ASAP7_75t_R PHY_308 ();
 NOR2x2_ASAP7_75t_R _36255_ (.A(net1783),
    .B(net1604),
    .Y(_06739_));
 OR3x1_ASAP7_75t_R _36256_ (.A(net2482),
    .B(_06143_),
    .C(_06739_),
    .Y(_06740_));
 NOR2x2_ASAP7_75t_R _36257_ (.A(net1758),
    .B(_06128_),
    .Y(_06741_));
 NOR2x1_ASAP7_75t_R _36258_ (.A(_06741_),
    .B(_06161_),
    .Y(_06742_));
 AOI21x1_ASAP7_75t_R _36259_ (.A1(_06251_),
    .A2(_06740_),
    .B(_06742_),
    .Y(_06743_));
 NAND2x1_ASAP7_75t_R _36260_ (.A(_06736_),
    .B(_06743_),
    .Y(_06744_));
 NOR2x1_ASAP7_75t_R _36261_ (.A(_06278_),
    .B(net2344),
    .Y(_06745_));
 AOI21x1_ASAP7_75t_R _36262_ (.A1(_06240_),
    .A2(net2399),
    .B(net1540),
    .Y(_06746_));
 NOR2x1_ASAP7_75t_R _36263_ (.A(_06745_),
    .B(_06746_),
    .Y(_06747_));
 INVx1_ASAP7_75t_R _36264_ (.A(_06747_),
    .Y(_06748_));
 NAND2x2_ASAP7_75t_R _36265_ (.A(net1096),
    .B(_06097_),
    .Y(_06750_));
 AO21x2_ASAP7_75t_R _36266_ (.A1(_06036_),
    .A2(_06750_),
    .B(_06203_),
    .Y(_06751_));
 TAPCELL_ASAP7_75t_R PHY_307 ();
 TAPCELL_ASAP7_75t_R PHY_306 ();
 AO21x1_ASAP7_75t_R _36269_ (.A1(net2764),
    .A2(_06250_),
    .B(net1262),
    .Y(_06754_));
 NAND2x1_ASAP7_75t_R _36270_ (.A(_06751_),
    .B(_06754_),
    .Y(_06755_));
 NOR2x1_ASAP7_75t_R _36271_ (.A(_06748_),
    .B(_06755_),
    .Y(_06756_));
 NOR2x1_ASAP7_75t_R _36272_ (.A(_06141_),
    .B(_06268_),
    .Y(_06757_));
 TAPCELL_ASAP7_75t_R PHY_305 ();
 TAPCELL_ASAP7_75t_R PHY_304 ();
 TAPCELL_ASAP7_75t_R PHY_303 ();
 NOR2x1_ASAP7_75t_R _36276_ (.A(net2639),
    .B(_06240_),
    .Y(_06762_));
 AO21x1_ASAP7_75t_R _36277_ (.A1(_06757_),
    .A2(_06061_),
    .B(_06762_),
    .Y(_06763_));
 INVx2_ASAP7_75t_R _36278_ (.A(_06121_),
    .Y(_06764_));
 NOR2x2_ASAP7_75t_R _36279_ (.A(_06058_),
    .B(_06063_),
    .Y(_06765_));
 TAPCELL_ASAP7_75t_R PHY_302 ();
 TAPCELL_ASAP7_75t_R PHY_301 ();
 AOI21x1_ASAP7_75t_R _36282_ (.A1(net1541),
    .A2(_06036_),
    .B(_06191_),
    .Y(_06768_));
 AOI21x1_ASAP7_75t_R _36283_ (.A1(_06764_),
    .A2(net3431),
    .B(_06768_),
    .Y(_06769_));
 INVx1_ASAP7_75t_R _36284_ (.A(_06769_),
    .Y(_06770_));
 NOR2x1_ASAP7_75t_R _36285_ (.A(_06763_),
    .B(_06770_),
    .Y(_06772_));
 NAND2x1_ASAP7_75t_R _36286_ (.A(_06756_),
    .B(_06772_),
    .Y(_06773_));
 NOR2x1_ASAP7_75t_R _36287_ (.A(_06744_),
    .B(_06773_),
    .Y(_06774_));
 INVx4_ASAP7_75t_R _36288_ (.A(_06229_),
    .Y(_06775_));
 AO22x1_ASAP7_75t_R _36289_ (.A1(_06251_),
    .A2(net3431),
    .B1(_06775_),
    .B2(net2084),
    .Y(_06776_));
 NAND2x1_ASAP7_75t_R _36290_ (.A(_06037_),
    .B(_06139_),
    .Y(_06777_));
 AO21x1_ASAP7_75t_R _36291_ (.A1(net2639),
    .A2(_06085_),
    .B(_06176_),
    .Y(_06778_));
 OAI21x1_ASAP7_75t_R _36292_ (.A1(net1664),
    .A2(_06777_),
    .B(_06778_),
    .Y(_06779_));
 NOR2x1_ASAP7_75t_R _36293_ (.A(_06776_),
    .B(_06779_),
    .Y(_06780_));
 INVx5_ASAP7_75t_R _36294_ (.A(_06176_),
    .Y(_06781_));
 AND2x6_ASAP7_75t_R _36295_ (.A(_06080_),
    .B(_06120_),
    .Y(_06783_));
 AO22x1_ASAP7_75t_R _36296_ (.A1(_06781_),
    .A2(_06256_),
    .B1(_06783_),
    .B2(_06739_),
    .Y(_06784_));
 NAND2x1_ASAP7_75t_R _36297_ (.A(net2744),
    .B(_06273_),
    .Y(_06785_));
 TAPCELL_ASAP7_75t_R PHY_300 ();
 TAPCELL_ASAP7_75t_R PHY_299 ();
 AO21x1_ASAP7_75t_R _36300_ (.A1(net3328),
    .A2(net3231),
    .B(_06240_),
    .Y(_06788_));
 OAI21x1_ASAP7_75t_R _36301_ (.A1(_06741_),
    .A2(_06785_),
    .B(_06788_),
    .Y(_06789_));
 NOR2x1_ASAP7_75t_R _36302_ (.A(_06784_),
    .B(_06789_),
    .Y(_06790_));
 NAND2x1_ASAP7_75t_R _36303_ (.A(_06780_),
    .B(_06790_),
    .Y(_06791_));
 AO21x1_ASAP7_75t_R _36304_ (.A1(_06036_),
    .A2(_06226_),
    .B(_06240_),
    .Y(_06792_));
 NAND2x2_ASAP7_75t_R _36305_ (.A(_06029_),
    .B(_06071_),
    .Y(_06794_));
 AO21x1_ASAP7_75t_R _36306_ (.A1(net2530),
    .A2(_06794_),
    .B(_06121_),
    .Y(_06795_));
 AO21x1_ASAP7_75t_R _36307_ (.A1(net3434),
    .A2(_06085_),
    .B(_06710_),
    .Y(_06796_));
 NAND3x1_ASAP7_75t_R _36308_ (.A(_06792_),
    .B(_06795_),
    .C(_06796_),
    .Y(_06797_));
 TAPCELL_ASAP7_75t_R PHY_298 ();
 NOR2x2_ASAP7_75t_R _36310_ (.A(_06098_),
    .B(net3421),
    .Y(_06799_));
 AOI22x1_ASAP7_75t_R _36311_ (.A1(_06783_),
    .A2(net2813),
    .B1(_06139_),
    .B2(_06799_),
    .Y(_06800_));
 NOR2x2_ASAP7_75t_R _36312_ (.A(_06029_),
    .B(_06052_),
    .Y(_06801_));
 NAND3x2_ASAP7_75t_R _36313_ (.B(net1549),
    .C(_06801_),
    .Y(_06802_),
    .A(_06092_));
 AO21x1_ASAP7_75t_R _36314_ (.A1(_06129_),
    .A2(net3231),
    .B(_06121_),
    .Y(_06803_));
 NAND3x1_ASAP7_75t_R _36315_ (.A(_06800_),
    .B(_06802_),
    .C(_06803_),
    .Y(_06805_));
 NOR2x1_ASAP7_75t_R _36316_ (.A(_06797_),
    .B(_06805_),
    .Y(_06806_));
 INVx1_ASAP7_75t_R _36317_ (.A(_06806_),
    .Y(_06807_));
 NOR2x1_ASAP7_75t_R _36318_ (.A(_06791_),
    .B(_06807_),
    .Y(_06808_));
 NAND2x1_ASAP7_75t_R _36319_ (.A(_06774_),
    .B(_06808_),
    .Y(_06809_));
 OA21x2_ASAP7_75t_R _36320_ (.A1(_06193_),
    .A2(net2084),
    .B(_06783_),
    .Y(_06810_));
 AOI211x1_ASAP7_75t_R _36321_ (.A1(net1276),
    .A2(net1546),
    .B(_06191_),
    .C(_06141_),
    .Y(_06811_));
 TAPCELL_ASAP7_75t_R PHY_297 ();
 AOI21x1_ASAP7_75t_R _36323_ (.A1(_06118_),
    .A2(_06196_),
    .B(net2786),
    .Y(_06813_));
 OR3x2_ASAP7_75t_R _36324_ (.A(_06810_),
    .B(_06811_),
    .C(_06813_),
    .Y(_06814_));
 INVx5_ASAP7_75t_R _36325_ (.A(_06064_),
    .Y(_06816_));
 INVx4_ASAP7_75t_R _36326_ (.A(_06118_),
    .Y(_06817_));
 OA21x2_ASAP7_75t_R _36327_ (.A1(_06142_),
    .A2(_06213_),
    .B(_06816_),
    .Y(_06818_));
 AOI21x1_ASAP7_75t_R _36328_ (.A1(_06816_),
    .A2(_06817_),
    .B(_06818_),
    .Y(_06819_));
 INVx1_ASAP7_75t_R _36329_ (.A(_06143_),
    .Y(_06820_));
 TAPCELL_ASAP7_75t_R PHY_296 ();
 OAI22x1_ASAP7_75t_R _36331_ (.A1(_06820_),
    .A2(_06710_),
    .B1(net3235),
    .B2(_06732_),
    .Y(_06822_));
 NOR2x1_ASAP7_75t_R _36332_ (.A(_06822_),
    .B(_06147_),
    .Y(_06823_));
 NAND2x2_ASAP7_75t_R _36333_ (.A(_06819_),
    .B(_06823_),
    .Y(_06824_));
 NOR2x1_ASAP7_75t_R _36334_ (.A(_06210_),
    .B(net3328),
    .Y(_06825_));
 AOI21x1_ASAP7_75t_R _36335_ (.A1(net3473),
    .A2(_06159_),
    .B(_06825_),
    .Y(_06827_));
 NOR2x2_ASAP7_75t_R _36336_ (.A(net1552),
    .B(net1588),
    .Y(_06828_));
 OAI21x1_ASAP7_75t_R _36337_ (.A1(_06142_),
    .A2(_06828_),
    .B(_06092_),
    .Y(_06829_));
 AOI21x1_ASAP7_75t_R _36338_ (.A1(_06131_),
    .A2(_06129_),
    .B(_06081_),
    .Y(_06830_));
 INVx1_ASAP7_75t_R _36339_ (.A(_06830_),
    .Y(_06831_));
 NAND2x2_ASAP7_75t_R _36340_ (.A(_06829_),
    .B(_06831_),
    .Y(_06832_));
 INVx1_ASAP7_75t_R _36341_ (.A(_06832_),
    .Y(_06833_));
 NAND2x2_ASAP7_75t_R _36342_ (.A(_06827_),
    .B(_06833_),
    .Y(_06834_));
 NOR3x1_ASAP7_75t_R _36343_ (.A(_06814_),
    .B(_06824_),
    .C(_06834_),
    .Y(_06835_));
 AOI22x1_ASAP7_75t_R _36344_ (.A1(_06159_),
    .A2(_06739_),
    .B1(_06783_),
    .B2(_06143_),
    .Y(_06836_));
 AOI22x1_ASAP7_75t_R _36345_ (.A1(_06783_),
    .A2(_06138_),
    .B1(_06251_),
    .B2(_06256_),
    .Y(_06838_));
 NAND2x1_ASAP7_75t_R _36346_ (.A(_06836_),
    .B(_06838_),
    .Y(_06839_));
 INVx1_ASAP7_75t_R _36347_ (.A(_06839_),
    .Y(_06840_));
 NAND2x2_ASAP7_75t_R _36348_ (.A(net3423),
    .B(net3429),
    .Y(_06841_));
 AO21x1_ASAP7_75t_R _36349_ (.A1(_06841_),
    .A2(_06137_),
    .B(_06104_),
    .Y(_06842_));
 AO21x1_ASAP7_75t_R _36350_ (.A1(_06278_),
    .A2(net3433),
    .B(net2412),
    .Y(_06843_));
 NAND2x2_ASAP7_75t_R _36351_ (.A(_06842_),
    .B(_06843_),
    .Y(_06844_));
 NOR2x1_ASAP7_75t_R _36352_ (.A(net3433),
    .B(_06030_),
    .Y(_06845_));
 OAI21x1_ASAP7_75t_R _36353_ (.A1(_06261_),
    .A2(_06845_),
    .B(_06273_),
    .Y(_06846_));
 NAND2x2_ASAP7_75t_R _36354_ (.A(net2855),
    .B(_06194_),
    .Y(_06847_));
 NAND2x2_ASAP7_75t_R _36355_ (.A(_06259_),
    .B(_06775_),
    .Y(_06849_));
 NAND3x2_ASAP7_75t_R _36356_ (.B(_06847_),
    .C(_06849_),
    .Y(_06850_),
    .A(_06846_));
 NOR2x1_ASAP7_75t_R _36357_ (.A(_06844_),
    .B(_06850_),
    .Y(_06851_));
 NAND2x1_ASAP7_75t_R _36358_ (.A(_06840_),
    .B(_06851_),
    .Y(_06852_));
 NAND2x2_ASAP7_75t_R _36359_ (.A(net1545),
    .B(net1295),
    .Y(_06853_));
 AO21x1_ASAP7_75t_R _36360_ (.A1(_06853_),
    .A2(_06126_),
    .B(net2786),
    .Y(_06854_));
 AO21x1_ASAP7_75t_R _36361_ (.A1(_06190_),
    .A2(net2530),
    .B(_06064_),
    .Y(_06855_));
 NAND2x1_ASAP7_75t_R _36362_ (.A(_06854_),
    .B(_06855_),
    .Y(_06856_));
 NOR2x1_ASAP7_75t_R _36363_ (.A(net2530),
    .B(_06044_),
    .Y(_06857_));
 NOR2x1_ASAP7_75t_R _36364_ (.A(_06121_),
    .B(_06181_),
    .Y(_06858_));
 AOI211x1_ASAP7_75t_R _36365_ (.A1(_06193_),
    .A2(_06139_),
    .B(_06857_),
    .C(_06858_),
    .Y(_06860_));
 INVx1_ASAP7_75t_R _36366_ (.A(_06860_),
    .Y(_06861_));
 NOR2x1_ASAP7_75t_R _36367_ (.A(_06856_),
    .B(_06861_),
    .Y(_06862_));
 NAND2x2_ASAP7_75t_R _36368_ (.A(_06096_),
    .B(net2744),
    .Y(_06863_));
 OAI22x1_ASAP7_75t_R _36369_ (.A1(_06863_),
    .A2(_06210_),
    .B1(_06084_),
    .B2(net2412),
    .Y(_06864_));
 OAI22x1_ASAP7_75t_R _36370_ (.A1(_06104_),
    .A2(_06036_),
    .B1(_06064_),
    .B2(_06126_),
    .Y(_06865_));
 NOR2x1_ASAP7_75t_R _36371_ (.A(_06864_),
    .B(_06865_),
    .Y(_06866_));
 OAI22x1_ASAP7_75t_R _36372_ (.A1(_06176_),
    .A2(_06226_),
    .B1(net2787),
    .B2(net3434),
    .Y(_06867_));
 OAI22x1_ASAP7_75t_R _36373_ (.A1(net1261),
    .A2(_06203_),
    .B1(net1217),
    .B2(_06121_),
    .Y(_06868_));
 NOR2x1_ASAP7_75t_R _36374_ (.A(_06867_),
    .B(_06868_),
    .Y(_06869_));
 NAND2x1_ASAP7_75t_R _36375_ (.A(_06866_),
    .B(_06869_),
    .Y(_06871_));
 INVx1_ASAP7_75t_R _36376_ (.A(_06871_),
    .Y(_06872_));
 NAND2x1_ASAP7_75t_R _36377_ (.A(_06862_),
    .B(_06872_),
    .Y(_06873_));
 NOR2x1_ASAP7_75t_R _36378_ (.A(_06852_),
    .B(_06873_),
    .Y(_06874_));
 NAND2x1_ASAP7_75t_R _36379_ (.A(_06835_),
    .B(_06874_),
    .Y(_06875_));
 NOR2x2_ASAP7_75t_R _36380_ (.A(_06809_),
    .B(_06875_),
    .Y(_06876_));
 NAND2x1_ASAP7_75t_R _36381_ (.A(_06729_),
    .B(_06876_),
    .Y(_06877_));
 AO21x2_ASAP7_75t_R _36382_ (.A1(_06131_),
    .A2(_06750_),
    .B(_06151_),
    .Y(_06878_));
 OAI21x1_ASAP7_75t_R _36383_ (.A1(_06765_),
    .A2(_06109_),
    .B(_06783_),
    .Y(_06879_));
 NAND2x2_ASAP7_75t_R _36384_ (.A(_06091_),
    .B(_06783_),
    .Y(_06880_));
 NAND3x2_ASAP7_75t_R _36385_ (.B(_06879_),
    .C(_06880_),
    .Y(_06882_),
    .A(_06878_));
 AO21x2_ASAP7_75t_R _36386_ (.A1(_06153_),
    .A2(_06278_),
    .B(_06151_),
    .Y(_06883_));
 AO21x2_ASAP7_75t_R _36387_ (.A1(_06072_),
    .A2(_06794_),
    .B(_06151_),
    .Y(_06884_));
 NAND2x2_ASAP7_75t_R _36388_ (.A(_06138_),
    .B(_06783_),
    .Y(_06885_));
 NAND3x2_ASAP7_75t_R _36389_ (.B(_06884_),
    .C(_06885_),
    .Y(_06886_),
    .A(_06883_));
 NOR2x2_ASAP7_75t_R _36390_ (.A(_06882_),
    .B(_06886_),
    .Y(_06887_));
 OR3x2_ASAP7_75t_R _36391_ (.A(_06040_),
    .B(_06174_),
    .C(_00627_),
    .Y(_06888_));
 NAND3x2_ASAP7_75t_R _36392_ (.B(net2343),
    .C(_06888_),
    .Y(_06889_),
    .A(_06887_));
 NOR3x2_ASAP7_75t_R _36393_ (.B(_06040_),
    .C(_06174_),
    .Y(_06890_),
    .A(net3441));
 INVx1_ASAP7_75t_R _36394_ (.A(_06744_),
    .Y(_06891_));
 NAND3x1_ASAP7_75t_R _36395_ (.A(_06747_),
    .B(_06751_),
    .C(_06754_),
    .Y(_06893_));
 INVx1_ASAP7_75t_R _36396_ (.A(_06763_),
    .Y(_06894_));
 NAND2x1_ASAP7_75t_R _36397_ (.A(_06769_),
    .B(_06894_),
    .Y(_06895_));
 NOR2x1_ASAP7_75t_R _36398_ (.A(_06893_),
    .B(_06895_),
    .Y(_06896_));
 NAND2x1_ASAP7_75t_R _36399_ (.A(_06891_),
    .B(_06896_),
    .Y(_06897_));
 INVx1_ASAP7_75t_R _36400_ (.A(_06791_),
    .Y(_06898_));
 NAND2x1_ASAP7_75t_R _36401_ (.A(_06806_),
    .B(_06898_),
    .Y(_06899_));
 NOR2x1_ASAP7_75t_R _36402_ (.A(_06897_),
    .B(_06899_),
    .Y(_06900_));
 NOR3x1_ASAP7_75t_R _36403_ (.A(_06839_),
    .B(_06850_),
    .C(_06844_),
    .Y(_06901_));
 INVx1_ASAP7_75t_R _36404_ (.A(_06856_),
    .Y(_06902_));
 NAND2x1_ASAP7_75t_R _36405_ (.A(_06860_),
    .B(_06902_),
    .Y(_06904_));
 NOR2x1_ASAP7_75t_R _36406_ (.A(_06871_),
    .B(_06904_),
    .Y(_06905_));
 NAND2x1_ASAP7_75t_R _36407_ (.A(_06901_),
    .B(_06905_),
    .Y(_06906_));
 INVx1_ASAP7_75t_R _36408_ (.A(_06814_),
    .Y(_06907_));
 NOR2x1_ASAP7_75t_R _36409_ (.A(_06834_),
    .B(_06824_),
    .Y(_06908_));
 NAND2x1_ASAP7_75t_R _36410_ (.A(_06907_),
    .B(_06908_),
    .Y(_06909_));
 NOR2x1_ASAP7_75t_R _36411_ (.A(_06906_),
    .B(_06909_),
    .Y(_06910_));
 NAND2x2_ASAP7_75t_R _36412_ (.A(_06900_),
    .B(_06910_),
    .Y(_06911_));
 OAI21x1_ASAP7_75t_R _36413_ (.A1(_06890_),
    .A2(_06911_),
    .B(_06286_),
    .Y(_06912_));
 NAND2x2_ASAP7_75t_R _36414_ (.A(_06877_),
    .B(_06912_),
    .Y(_06913_));
 OAI21x1_ASAP7_75t_R _36415_ (.A1(_06680_),
    .A2(_06698_),
    .B(_06913_),
    .Y(_06915_));
 NOR2x1_ASAP7_75t_R _36416_ (.A(_06697_),
    .B(_06679_),
    .Y(_06916_));
 NOR2x1_ASAP7_75t_R _36417_ (.A(_06552_),
    .B(net1928),
    .Y(_06917_));
 NOR2x1_ASAP7_75t_R _36418_ (.A(_06911_),
    .B(_06286_),
    .Y(_06918_));
 NOR2x1_ASAP7_75t_R _36419_ (.A(_06041_),
    .B(_06889_),
    .Y(_06919_));
 NAND2x2_ASAP7_75t_R _36420_ (.A(net3233),
    .B(_06919_),
    .Y(_06920_));
 AOI21x1_ASAP7_75t_R _36421_ (.A1(_06920_),
    .A2(_06876_),
    .B(_06729_),
    .Y(_06921_));
 NOR2x1_ASAP7_75t_R _36422_ (.A(_06918_),
    .B(_06921_),
    .Y(_06922_));
 OAI21x1_ASAP7_75t_R _36423_ (.A1(_06916_),
    .A2(_06917_),
    .B(_06922_),
    .Y(_06923_));
 NAND2x1_ASAP7_75t_R _36424_ (.A(_06915_),
    .B(_06923_),
    .Y(_06924_));
 NAND2x1_ASAP7_75t_R _36425_ (.A(_06424_),
    .B(_06924_),
    .Y(_06926_));
 NOR2x1_ASAP7_75t_R _36426_ (.A(_06424_),
    .B(_06924_),
    .Y(_06927_));
 INVx1_ASAP7_75t_R _36427_ (.A(_06927_),
    .Y(_06928_));
 AOI21x1_ASAP7_75t_R _36428_ (.A1(_06926_),
    .A2(_06928_),
    .B(net388),
    .Y(_06929_));
 INVx1_ASAP7_75t_R _36429_ (.A(_00499_),
    .Y(_06930_));
 OAI21x1_ASAP7_75t_R _36430_ (.A1(_06302_),
    .A2(_06929_),
    .B(_06930_),
    .Y(_06931_));
 NOR3x1_ASAP7_75t_R _36431_ (.A(_05726_),
    .B(net3114),
    .C(net3354),
    .Y(_06932_));
 OAI21x1_ASAP7_75t_R _36432_ (.A1(_05730_),
    .A2(_06932_),
    .B(net3419),
    .Y(_06933_));
 NOR3x1_ASAP7_75t_R _36433_ (.A(_05726_),
    .B(_05715_),
    .C(net3354),
    .Y(_06934_));
 OAI21x1_ASAP7_75t_R _36434_ (.A1(_05429_),
    .A2(_06934_),
    .B(_06422_),
    .Y(_06935_));
 NAND2x1_ASAP7_75t_R _36435_ (.A(_06933_),
    .B(_06935_),
    .Y(_06937_));
 AOI21x1_ASAP7_75t_R _36436_ (.A1(_06915_),
    .A2(_06923_),
    .B(_06937_),
    .Y(_06938_));
 OAI21x1_ASAP7_75t_R _36437_ (.A1(_06927_),
    .A2(_06938_),
    .B(net394),
    .Y(_06939_));
 INVx1_ASAP7_75t_R _36438_ (.A(_06302_),
    .Y(_06940_));
 NAND3x2_ASAP7_75t_R _36439_ (.B(_00499_),
    .C(_06940_),
    .Y(_06941_),
    .A(_06939_));
 NAND2x2_ASAP7_75t_R _36440_ (.A(_06931_),
    .B(_06941_),
    .Y(_00106_));
 NOR2x1_ASAP7_75t_R _36441_ (.A(net394),
    .B(_00849_),
    .Y(_06942_));
 AO21x1_ASAP7_75t_R _36442_ (.A1(net1877),
    .A2(_05360_),
    .B(net3095),
    .Y(_06943_));
 AO21x1_ASAP7_75t_R _36443_ (.A1(_05185_),
    .A2(net990),
    .B(net3095),
    .Y(_06944_));
 AND2x2_ASAP7_75t_R _36444_ (.A(_06943_),
    .B(_06944_),
    .Y(_06945_));
 AO21x1_ASAP7_75t_R _36445_ (.A1(net1764),
    .A2(net2149),
    .B(net3095),
    .Y(_06947_));
 AND2x2_ASAP7_75t_R _36446_ (.A(_05254_),
    .B(_06947_),
    .Y(_06948_));
 NAND2x1_ASAP7_75t_R _36447_ (.A(_06945_),
    .B(_06948_),
    .Y(_06949_));
 AO21x1_ASAP7_75t_R _36448_ (.A1(net992),
    .A2(net990),
    .B(_05256_),
    .Y(_06950_));
 OA21x2_ASAP7_75t_R _36449_ (.A1(_05256_),
    .A2(net1878),
    .B(_06950_),
    .Y(_06951_));
 OA211x2_ASAP7_75t_R _36450_ (.A1(net3436),
    .A2(net3442),
    .B(_05181_),
    .C(net2171),
    .Y(_06952_));
 INVx1_ASAP7_75t_R _36451_ (.A(_06952_),
    .Y(_06953_));
 NAND2x1_ASAP7_75t_R _36452_ (.A(_06953_),
    .B(_06951_),
    .Y(_06954_));
 NOR2x1_ASAP7_75t_R _36453_ (.A(_06949_),
    .B(_06954_),
    .Y(_06955_));
 NOR2x2_ASAP7_75t_R _36454_ (.A(net1521),
    .B(net3100),
    .Y(_06956_));
 OA21x2_ASAP7_75t_R _36455_ (.A1(net2171),
    .A2(_06956_),
    .B(_05332_),
    .Y(_06958_));
 NAND2x1_ASAP7_75t_R _36456_ (.A(_05059_),
    .B(_05332_),
    .Y(_06959_));
 NAND2x2_ASAP7_75t_R _36457_ (.A(_05151_),
    .B(_05332_),
    .Y(_06960_));
 NAND3x1_ASAP7_75t_R _36458_ (.A(_05331_),
    .B(_06959_),
    .C(_06960_),
    .Y(_06961_));
 NOR2x1_ASAP7_75t_R _36459_ (.A(_06958_),
    .B(_06961_),
    .Y(_06962_));
 AO21x1_ASAP7_75t_R _36460_ (.A1(_05360_),
    .A2(net1793),
    .B(_05198_),
    .Y(_06963_));
 NAND2x1_ASAP7_75t_R _36461_ (.A(_05059_),
    .B(_05199_),
    .Y(_06964_));
 NAND2x1_ASAP7_75t_R _36462_ (.A(_05142_),
    .B(_05199_),
    .Y(_06965_));
 AND3x1_ASAP7_75t_R _36463_ (.A(_06963_),
    .B(_06964_),
    .C(_06965_),
    .Y(_06966_));
 AND2x2_ASAP7_75t_R _36464_ (.A(_06962_),
    .B(_06966_),
    .Y(_06967_));
 NAND2x1_ASAP7_75t_R _36465_ (.A(_06967_),
    .B(_06955_),
    .Y(_06969_));
 AO21x1_ASAP7_75t_R _36466_ (.A1(net2417),
    .A2(net2643),
    .B(_05138_),
    .Y(_06970_));
 OAI21x1_ASAP7_75t_R _36467_ (.A1(net1838),
    .A2(_05138_),
    .B(_06970_),
    .Y(_06971_));
 AO21x1_ASAP7_75t_R _36468_ (.A1(_05206_),
    .A2(_05165_),
    .B(_05138_),
    .Y(_06972_));
 OAI21x1_ASAP7_75t_R _36469_ (.A1(net2150),
    .A2(_05138_),
    .B(_06972_),
    .Y(_06973_));
 NOR2x1_ASAP7_75t_R _36470_ (.A(_06971_),
    .B(_06973_),
    .Y(_06974_));
 AO21x1_ASAP7_75t_R _36471_ (.A1(net1765),
    .A2(net1894),
    .B(net3444),
    .Y(_06975_));
 AO21x1_ASAP7_75t_R _36472_ (.A1(net1822),
    .A2(net1877),
    .B(net3444),
    .Y(_06976_));
 AND3x1_ASAP7_75t_R _36473_ (.A(_05374_),
    .B(_06975_),
    .C(_06976_),
    .Y(_06977_));
 AND2x2_ASAP7_75t_R _36474_ (.A(_06974_),
    .B(_06977_),
    .Y(_06978_));
 AO31x2_ASAP7_75t_R _36475_ (.A1(net2150),
    .A2(net1237),
    .A3(net1091),
    .B(_05062_),
    .Y(_06980_));
 AO21x1_ASAP7_75t_R _36476_ (.A1(net2146),
    .A2(net1140),
    .B(_05062_),
    .Y(_06981_));
 NAND2x1_ASAP7_75t_R _36477_ (.A(_05065_),
    .B(net3456),
    .Y(_06982_));
 AOI21x1_ASAP7_75t_R _36478_ (.A1(net1836),
    .A2(_06982_),
    .B(_05062_),
    .Y(_06983_));
 INVx1_ASAP7_75t_R _36479_ (.A(_06983_),
    .Y(_06984_));
 NAND3x1_ASAP7_75t_R _36480_ (.A(_06980_),
    .B(_06981_),
    .C(_06984_),
    .Y(_06985_));
 NAND2x2_ASAP7_75t_R _36481_ (.A(_05191_),
    .B(_05127_),
    .Y(_06986_));
 NAND2x1_ASAP7_75t_R _36482_ (.A(_05239_),
    .B(_05127_),
    .Y(_06987_));
 NAND2x1_ASAP7_75t_R _36483_ (.A(_06986_),
    .B(_06987_),
    .Y(_06988_));
 NAND2x2_ASAP7_75t_R _36484_ (.A(_05218_),
    .B(_05127_),
    .Y(_06989_));
 AO21x2_ASAP7_75t_R _36485_ (.A1(_05163_),
    .A2(_05165_),
    .B(_05126_),
    .Y(_06991_));
 NAND2x1_ASAP7_75t_R _36486_ (.A(_06989_),
    .B(_06991_),
    .Y(_06992_));
 NOR2x1_ASAP7_75t_R _36487_ (.A(_06988_),
    .B(_06992_),
    .Y(_06993_));
 AO21x1_ASAP7_75t_R _36488_ (.A1(net3427),
    .A2(net1877),
    .B(_05126_),
    .Y(_06994_));
 NAND2x1_ASAP7_75t_R _36489_ (.A(_05422_),
    .B(_05127_),
    .Y(_06995_));
 AO21x1_ASAP7_75t_R _36490_ (.A1(net1945),
    .A2(net2643),
    .B(_05126_),
    .Y(_06996_));
 AND3x1_ASAP7_75t_R _36491_ (.A(_06994_),
    .B(_06995_),
    .C(_06996_),
    .Y(_06997_));
 NAND2x1_ASAP7_75t_R _36492_ (.A(_06993_),
    .B(_06997_),
    .Y(_06998_));
 NOR2x1_ASAP7_75t_R _36493_ (.A(_06985_),
    .B(_06998_),
    .Y(_06999_));
 NAND2x2_ASAP7_75t_R _36494_ (.A(_06978_),
    .B(_06999_),
    .Y(_07000_));
 NOR2x1_ASAP7_75t_R _36495_ (.A(_06969_),
    .B(_07000_),
    .Y(_07002_));
 TAPCELL_ASAP7_75t_R PHY_295 ();
 OA21x2_ASAP7_75t_R _36497_ (.A1(net3446),
    .A2(net2529),
    .B(_05274_),
    .Y(_07004_));
 AO21x1_ASAP7_75t_R _36498_ (.A1(_05211_),
    .A2(net2027),
    .B(net3455),
    .Y(_07005_));
 AO21x1_ASAP7_75t_R _36499_ (.A1(net1403),
    .A2(net1947),
    .B(net2529),
    .Y(_07006_));
 AND2x2_ASAP7_75t_R _36500_ (.A(_07005_),
    .B(_07006_),
    .Y(_07007_));
 AND2x2_ASAP7_75t_R _36501_ (.A(_07004_),
    .B(_07007_),
    .Y(_07008_));
 AO21x1_ASAP7_75t_R _36502_ (.A1(net3369),
    .A2(net2146),
    .B(net2621),
    .Y(_07009_));
 AO21x1_ASAP7_75t_R _36503_ (.A1(net990),
    .A2(net964),
    .B(net2621),
    .Y(_07010_));
 NAND2x2_ASAP7_75t_R _36504_ (.A(_06346_),
    .B(_05108_),
    .Y(_07011_));
 NAND3x2_ASAP7_75t_R _36505_ (.B(_07010_),
    .C(_07011_),
    .Y(_07013_),
    .A(_07009_));
 AO21x1_ASAP7_75t_R _36506_ (.A1(net1867),
    .A2(net1140),
    .B(net2493),
    .Y(_07014_));
 AO21x1_ASAP7_75t_R _36507_ (.A1(net992),
    .A2(net964),
    .B(net2493),
    .Y(_07015_));
 NAND3x2_ASAP7_75t_R _36508_ (.B(_07015_),
    .C(_06347_),
    .Y(_07016_),
    .A(_07014_));
 NOR2x2_ASAP7_75t_R _36509_ (.A(_07013_),
    .B(_07016_),
    .Y(_07017_));
 AO21x1_ASAP7_75t_R _36510_ (.A1(net1140),
    .A2(_05122_),
    .B(net3104),
    .Y(_07018_));
 AO21x1_ASAP7_75t_R _36511_ (.A1(_05360_),
    .A2(net992),
    .B(net3104),
    .Y(_07019_));
 AND2x2_ASAP7_75t_R _36512_ (.A(_07018_),
    .B(_07019_),
    .Y(_07020_));
 NAND3x2_ASAP7_75t_R _36513_ (.B(_07017_),
    .C(_07020_),
    .Y(_07021_),
    .A(_07008_));
 AO31x2_ASAP7_75t_R _36514_ (.A1(net964),
    .A2(net2138),
    .A3(net992),
    .B(_05215_),
    .Y(_07022_));
 AO21x1_ASAP7_75t_R _36515_ (.A1(_05206_),
    .A2(net3101),
    .B(_05215_),
    .Y(_07024_));
 AO21x1_ASAP7_75t_R _36516_ (.A1(net1867),
    .A2(net1764),
    .B(_05215_),
    .Y(_07025_));
 NAND3x1_ASAP7_75t_R _36517_ (.A(_07022_),
    .B(_07024_),
    .C(_07025_),
    .Y(_07026_));
 AO21x1_ASAP7_75t_R _36518_ (.A1(net3096),
    .A2(_05360_),
    .B(_05186_),
    .Y(_07027_));
 OA21x2_ASAP7_75t_R _36519_ (.A1(net964),
    .A2(_05186_),
    .B(_07027_),
    .Y(_07028_));
 NOR2x1_ASAP7_75t_R _36520_ (.A(_05177_),
    .B(_05186_),
    .Y(_07029_));
 OA31x2_ASAP7_75t_R _36521_ (.A1(_05205_),
    .A2(_05203_),
    .A3(_05218_),
    .B1(_05247_),
    .Y(_07030_));
 NOR2x1_ASAP7_75t_R _36522_ (.A(_07029_),
    .B(_07030_),
    .Y(_07031_));
 NAND2x1_ASAP7_75t_R _36523_ (.A(_07028_),
    .B(_07031_),
    .Y(_07032_));
 NOR2x1_ASAP7_75t_R _36524_ (.A(_07026_),
    .B(_07032_),
    .Y(_07033_));
 NAND2x1_ASAP7_75t_R _36525_ (.A(_06346_),
    .B(_05154_),
    .Y(_07035_));
 OAI21x1_ASAP7_75t_R _36526_ (.A1(net2784),
    .A2(_05319_),
    .B(_07035_),
    .Y(_07036_));
 AO21x1_ASAP7_75t_R _36527_ (.A1(_05163_),
    .A2(net3102),
    .B(_05153_),
    .Y(_07037_));
 NAND2x1_ASAP7_75t_R _36528_ (.A(_05168_),
    .B(_07037_),
    .Y(_07038_));
 OR2x2_ASAP7_75t_R _36529_ (.A(_07036_),
    .B(_07038_),
    .Y(_07039_));
 AO21x1_ASAP7_75t_R _36530_ (.A1(net1091),
    .A2(net1140),
    .B(_05306_),
    .Y(_07040_));
 NOR2x1_ASAP7_75t_R _36531_ (.A(_05058_),
    .B(_05306_),
    .Y(_07041_));
 OA211x2_ASAP7_75t_R _36532_ (.A1(net1321),
    .A2(net3442),
    .B(_05100_),
    .C(net2224),
    .Y(_07042_));
 NOR2x1_ASAP7_75t_R _36533_ (.A(_07041_),
    .B(_07042_),
    .Y(_07043_));
 NAND2x1_ASAP7_75t_R _36534_ (.A(_07040_),
    .B(_07043_),
    .Y(_07044_));
 NOR2x1_ASAP7_75t_R _36535_ (.A(_07039_),
    .B(_07044_),
    .Y(_07046_));
 NAND2x1_ASAP7_75t_R _36536_ (.A(_07033_),
    .B(_07046_),
    .Y(_07047_));
 NOR2x2_ASAP7_75t_R _36537_ (.A(_07021_),
    .B(_07047_),
    .Y(_07048_));
 NAND2x2_ASAP7_75t_R _36538_ (.A(_07002_),
    .B(_07048_),
    .Y(_07049_));
 INVx2_ASAP7_75t_R _36539_ (.A(_07049_),
    .Y(_07050_));
 AO21x1_ASAP7_75t_R _36540_ (.A1(net1902),
    .A2(net2815),
    .B(_05492_),
    .Y(_07051_));
 TAPCELL_ASAP7_75t_R PHY_294 ();
 AO21x1_ASAP7_75t_R _36542_ (.A1(net1084),
    .A2(_05486_),
    .B(_05492_),
    .Y(_07053_));
 NOR2x1_ASAP7_75t_R _36543_ (.A(_05492_),
    .B(net2003),
    .Y(_07054_));
 INVx1_ASAP7_75t_R _36544_ (.A(_07054_),
    .Y(_07055_));
 AND3x1_ASAP7_75t_R _36545_ (.A(_07051_),
    .B(_07053_),
    .C(_07055_),
    .Y(_07057_));
 AO21x1_ASAP7_75t_R _36546_ (.A1(net1902),
    .A2(_05613_),
    .B(_05511_),
    .Y(_07058_));
 AO21x1_ASAP7_75t_R _36547_ (.A1(_06574_),
    .A2(_05580_),
    .B(_05511_),
    .Y(_07059_));
 AND2x2_ASAP7_75t_R _36548_ (.A(_07058_),
    .B(_07059_),
    .Y(_07060_));
 AND2x2_ASAP7_75t_R _36549_ (.A(_07057_),
    .B(_07060_),
    .Y(_07061_));
 AO21x1_ASAP7_75t_R _36550_ (.A1(net2400),
    .A2(net2610),
    .B(net2755),
    .Y(_07062_));
 NOR2x1_ASAP7_75t_R _36551_ (.A(_05528_),
    .B(net2815),
    .Y(_07063_));
 INVx1_ASAP7_75t_R _36552_ (.A(_07063_),
    .Y(_07064_));
 NAND3x1_ASAP7_75t_R _36553_ (.A(_05537_),
    .B(_07062_),
    .C(_07064_),
    .Y(_07065_));
 NOR2x2_ASAP7_75t_R _36554_ (.A(_05513_),
    .B(net1666),
    .Y(_07066_));
 OA21x2_ASAP7_75t_R _36555_ (.A1(_06637_),
    .A2(_07066_),
    .B(_05545_),
    .Y(_07068_));
 NOR2x1_ASAP7_75t_R _36556_ (.A(_05550_),
    .B(_07068_),
    .Y(_07069_));
 AO21x1_ASAP7_75t_R _36557_ (.A1(net2663),
    .A2(net1124),
    .B(_05548_),
    .Y(_07070_));
 AO21x1_ASAP7_75t_R _36558_ (.A1(net2032),
    .A2(net2610),
    .B(_05548_),
    .Y(_07071_));
 NAND3x1_ASAP7_75t_R _36559_ (.A(_07069_),
    .B(_07070_),
    .C(_07071_),
    .Y(_07072_));
 NOR2x1_ASAP7_75t_R _36560_ (.A(_07065_),
    .B(_07072_),
    .Y(_07073_));
 NAND2x2_ASAP7_75t_R _36561_ (.A(_07061_),
    .B(_07073_),
    .Y(_07074_));
 INVx2_ASAP7_75t_R _36562_ (.A(_07074_),
    .Y(_07075_));
 AO21x1_ASAP7_75t_R _36563_ (.A1(net3349),
    .A2(_05613_),
    .B(_05453_),
    .Y(_07076_));
 OAI21x1_ASAP7_75t_R _36564_ (.A1(net1000),
    .A2(_05467_),
    .B(_07076_),
    .Y(_07077_));
 AO22x1_ASAP7_75t_R _36565_ (.A1(_05435_),
    .A2(_06626_),
    .B1(_05458_),
    .B2(_05515_),
    .Y(_07079_));
 NOR2x1_ASAP7_75t_R _36566_ (.A(_07077_),
    .B(_07079_),
    .Y(_07080_));
 AO21x1_ASAP7_75t_R _36567_ (.A1(net2191),
    .A2(net3113),
    .B(_05472_),
    .Y(_07081_));
 AO21x1_ASAP7_75t_R _36568_ (.A1(net2153),
    .A2(net2815),
    .B(_05472_),
    .Y(_07082_));
 AO21x1_ASAP7_75t_R _36569_ (.A1(net2833),
    .A2(net1084),
    .B(_05472_),
    .Y(_07083_));
 NAND2x1_ASAP7_75t_R _36570_ (.A(_05600_),
    .B(net2809),
    .Y(_07084_));
 AND4x1_ASAP7_75t_R _36571_ (.A(_07081_),
    .B(_07082_),
    .C(_07083_),
    .D(_07084_),
    .Y(_07085_));
 NAND2x2_ASAP7_75t_R _36572_ (.A(_07080_),
    .B(_07085_),
    .Y(_07086_));
 AO21x1_ASAP7_75t_R _36573_ (.A1(_05643_),
    .A2(_05462_),
    .B(net2390),
    .Y(_07087_));
 AO21x1_ASAP7_75t_R _36574_ (.A1(net1627),
    .A2(net1771),
    .B(net2390),
    .Y(_07088_));
 AO21x1_ASAP7_75t_R _36575_ (.A1(net1085),
    .A2(_05486_),
    .B(net2390),
    .Y(_07090_));
 INVx1_ASAP7_75t_R _36576_ (.A(_05572_),
    .Y(_07091_));
 AND4x2_ASAP7_75t_R _36577_ (.A(_07087_),
    .B(_07088_),
    .C(_07090_),
    .D(_07091_),
    .Y(_07092_));
 NAND2x1_ASAP7_75t_R _36578_ (.A(_05577_),
    .B(_06637_),
    .Y(_07093_));
 NAND2x1_ASAP7_75t_R _36579_ (.A(_07093_),
    .B(_06666_),
    .Y(_07094_));
 OA211x2_ASAP7_75t_R _36580_ (.A1(net1000),
    .A2(net3098),
    .B(_05577_),
    .C(_05461_),
    .Y(_07095_));
 NOR2x2_ASAP7_75t_R _36581_ (.A(_07094_),
    .B(_07095_),
    .Y(_07096_));
 AO21x1_ASAP7_75t_R _36582_ (.A1(net1083),
    .A2(net2400),
    .B(_05581_),
    .Y(_07097_));
 OA21x2_ASAP7_75t_R _36583_ (.A1(_05486_),
    .A2(_05581_),
    .B(_07097_),
    .Y(_07098_));
 NAND3x2_ASAP7_75t_R _36584_ (.B(_07096_),
    .C(_07098_),
    .Y(_07099_),
    .A(_07092_));
 NOR2x1_ASAP7_75t_R _36585_ (.A(_07086_),
    .B(_07099_),
    .Y(_07101_));
 NAND2x2_ASAP7_75t_R _36586_ (.A(_07075_),
    .B(_07101_),
    .Y(_07102_));
 AO21x1_ASAP7_75t_R _36587_ (.A1(net1083),
    .A2(net2115),
    .B(_05683_),
    .Y(_07103_));
 AO21x1_ASAP7_75t_R _36588_ (.A1(net2567),
    .A2(net2032),
    .B(_05683_),
    .Y(_07104_));
 AND2x2_ASAP7_75t_R _36589_ (.A(_07103_),
    .B(_07104_),
    .Y(_07105_));
 AO21x1_ASAP7_75t_R _36590_ (.A1(net1627),
    .A2(net2870),
    .B(_05683_),
    .Y(_07106_));
 NAND2x1_ASAP7_75t_R _36591_ (.A(_05684_),
    .B(_05686_),
    .Y(_07107_));
 AND3x1_ASAP7_75t_R _36592_ (.A(_07106_),
    .B(_07107_),
    .C(_06557_),
    .Y(_07108_));
 NAND2x2_ASAP7_75t_R _36593_ (.A(_07105_),
    .B(_07108_),
    .Y(_07109_));
 NOR2x1_ASAP7_75t_R _36594_ (.A(net1206),
    .B(_06576_),
    .Y(_07110_));
 AO21x2_ASAP7_75t_R _36595_ (.A1(_05445_),
    .A2(net3121),
    .B(net2726),
    .Y(_07112_));
 NOR2x1_ASAP7_75t_R _36596_ (.A(_07112_),
    .B(_06576_),
    .Y(_07113_));
 AOI221x1_ASAP7_75t_R _36597_ (.A1(_05661_),
    .A2(net3463),
    .B1(net3460),
    .B2(_07110_),
    .C(_07113_),
    .Y(_07114_));
 AO21x1_ASAP7_75t_R _36598_ (.A1(net2400),
    .A2(net3461),
    .B(_05654_),
    .Y(_07115_));
 NAND2x1_ASAP7_75t_R _36599_ (.A(_05463_),
    .B(_05657_),
    .Y(_07116_));
 NAND2x1_ASAP7_75t_R _36600_ (.A(_05522_),
    .B(_05657_),
    .Y(_07117_));
 AND3x1_ASAP7_75t_R _36601_ (.A(_07115_),
    .B(_07116_),
    .C(_07117_),
    .Y(_07118_));
 NAND2x2_ASAP7_75t_R _36602_ (.A(_07114_),
    .B(_07118_),
    .Y(_07119_));
 AO21x1_ASAP7_75t_R _36603_ (.A1(net2032),
    .A2(net2611),
    .B(_05677_),
    .Y(_07120_));
 OA21x2_ASAP7_75t_R _36604_ (.A1(_05677_),
    .A2(net1083),
    .B(_07120_),
    .Y(_07121_));
 OA211x2_ASAP7_75t_R _36605_ (.A1(net2814),
    .A2(net3098),
    .B(_05675_),
    .C(net3463),
    .Y(_07123_));
 INVx1_ASAP7_75t_R _36606_ (.A(_07123_),
    .Y(_07124_));
 NAND2x2_ASAP7_75t_R _36607_ (.A(_07121_),
    .B(_07124_),
    .Y(_07125_));
 NOR3x2_ASAP7_75t_R _36608_ (.B(_07119_),
    .C(_07125_),
    .Y(_07126_),
    .A(_07109_));
 AO21x1_ASAP7_75t_R _36609_ (.A1(net2220),
    .A2(net3115),
    .B(net2447),
    .Y(_07127_));
 AO21x1_ASAP7_75t_R _36610_ (.A1(net2191),
    .A2(net1083),
    .B(net2447),
    .Y(_07128_));
 NAND2x1_ASAP7_75t_R _36611_ (.A(_07127_),
    .B(_07128_),
    .Y(_07129_));
 AO21x1_ASAP7_75t_R _36612_ (.A1(net1773),
    .A2(net1267),
    .B(net2447),
    .Y(_07130_));
 NAND2x2_ASAP7_75t_R _36613_ (.A(net2702),
    .B(_06613_),
    .Y(_07131_));
 NAND2x2_ASAP7_75t_R _36614_ (.A(_05463_),
    .B(_06613_),
    .Y(_07132_));
 NAND3x1_ASAP7_75t_R _36615_ (.A(_07130_),
    .B(_07131_),
    .C(_07132_),
    .Y(_07134_));
 NOR2x1_ASAP7_75t_R _36616_ (.A(_07129_),
    .B(_07134_),
    .Y(_07135_));
 OR3x1_ASAP7_75t_R _36617_ (.A(_05626_),
    .B(_05450_),
    .C(_07112_),
    .Y(_07136_));
 AO21x1_ASAP7_75t_R _36618_ (.A1(_05613_),
    .A2(net2816),
    .B(net2411),
    .Y(_07137_));
 AO21x1_ASAP7_75t_R _36619_ (.A1(net2870),
    .A2(net1773),
    .B(net2411),
    .Y(_07138_));
 AND3x1_ASAP7_75t_R _36620_ (.A(_07137_),
    .B(_07138_),
    .C(_06608_),
    .Y(_07139_));
 AND3x2_ASAP7_75t_R _36621_ (.A(_07135_),
    .B(_07136_),
    .C(_07139_),
    .Y(_07140_));
 AO21x1_ASAP7_75t_R _36622_ (.A1(net2191),
    .A2(net1083),
    .B(net2617),
    .Y(_07141_));
 AO21x1_ASAP7_75t_R _36623_ (.A1(net1772),
    .A2(net1267),
    .B(net2617),
    .Y(_07142_));
 NOR2x1_ASAP7_75t_R _36624_ (.A(_05676_),
    .B(net2617),
    .Y(_07143_));
 INVx1_ASAP7_75t_R _36625_ (.A(_07143_),
    .Y(_07145_));
 AND3x1_ASAP7_75t_R _36626_ (.A(_07141_),
    .B(_07142_),
    .C(_07145_),
    .Y(_07146_));
 INVx1_ASAP7_75t_R _36627_ (.A(_07146_),
    .Y(_07147_));
 AO21x1_ASAP7_75t_R _36628_ (.A1(net1083),
    .A2(net1124),
    .B(net2461),
    .Y(_07148_));
 AO21x1_ASAP7_75t_R _36629_ (.A1(net2611),
    .A2(net2477),
    .B(net2461),
    .Y(_07149_));
 AND2x2_ASAP7_75t_R _36630_ (.A(_07148_),
    .B(_07149_),
    .Y(_07150_));
 NAND2x2_ASAP7_75t_R _36631_ (.A(_06592_),
    .B(_06593_),
    .Y(_07151_));
 NOR2x2_ASAP7_75t_R _36632_ (.A(net1208),
    .B(_05519_),
    .Y(_07152_));
 OA21x2_ASAP7_75t_R _36633_ (.A1(_07152_),
    .A2(net2834),
    .B(_06593_),
    .Y(_07153_));
 INVx1_ASAP7_75t_R _36634_ (.A(_07153_),
    .Y(_07154_));
 NAND3x2_ASAP7_75t_R _36635_ (.B(_07151_),
    .C(_07154_),
    .Y(_07156_),
    .A(_07150_));
 NOR2x2_ASAP7_75t_R _36636_ (.A(_07147_),
    .B(_07156_),
    .Y(_07157_));
 NAND3x2_ASAP7_75t_R _36637_ (.B(_07140_),
    .C(_07157_),
    .Y(_07158_),
    .A(_07126_));
 NOR2x2_ASAP7_75t_R _36638_ (.A(_07102_),
    .B(_07158_),
    .Y(_07159_));
 NAND2x2_ASAP7_75t_R _36639_ (.A(_07159_),
    .B(_07050_),
    .Y(_07160_));
 NOR3x2_ASAP7_75t_R _36640_ (.B(_07099_),
    .C(_07086_),
    .Y(_07161_),
    .A(_07074_));
 INVx1_ASAP7_75t_R _36641_ (.A(_07126_),
    .Y(_07162_));
 NAND2x1_ASAP7_75t_R _36642_ (.A(_07157_),
    .B(_07140_),
    .Y(_07163_));
 NOR2x1_ASAP7_75t_R _36643_ (.A(_07163_),
    .B(_07162_),
    .Y(_07164_));
 NAND2x2_ASAP7_75t_R _36644_ (.A(_07161_),
    .B(_07164_),
    .Y(_07165_));
 NAND2x2_ASAP7_75t_R _36645_ (.A(net3165),
    .B(_07165_),
    .Y(_07167_));
 INVx2_ASAP7_75t_R _36646_ (.A(_06436_),
    .Y(_07168_));
 AO21x1_ASAP7_75t_R _36647_ (.A1(_05918_),
    .A2(_07168_),
    .B(_05884_),
    .Y(_07169_));
 NAND2x1_ASAP7_75t_R _36648_ (.A(_06494_),
    .B(_05885_),
    .Y(_07170_));
 AO21x1_ASAP7_75t_R _36649_ (.A1(net1118),
    .A2(net3375),
    .B(_05884_),
    .Y(_07171_));
 AND3x1_ASAP7_75t_R _36650_ (.A(_07169_),
    .B(_07170_),
    .C(_07171_),
    .Y(_07172_));
 AO21x1_ASAP7_75t_R _36651_ (.A1(net2603),
    .A2(net980),
    .B(_05873_),
    .Y(_07173_));
 AO21x1_ASAP7_75t_R _36652_ (.A1(net1037),
    .A2(net1787),
    .B(_05873_),
    .Y(_07174_));
 NAND2x1_ASAP7_75t_R _36653_ (.A(_07173_),
    .B(_07174_),
    .Y(_07175_));
 INVx1_ASAP7_75t_R _36654_ (.A(_05875_),
    .Y(_07176_));
 NOR2x1_ASAP7_75t_R _36655_ (.A(_05764_),
    .B(net2185),
    .Y(_07178_));
 OA21x2_ASAP7_75t_R _36656_ (.A1(_06472_),
    .A2(_07178_),
    .B(_05878_),
    .Y(_07179_));
 NOR3x1_ASAP7_75t_R _36657_ (.A(_07175_),
    .B(_07176_),
    .C(_07179_),
    .Y(_07180_));
 NAND2x1_ASAP7_75t_R _36658_ (.A(_07172_),
    .B(_07180_),
    .Y(_07181_));
 AO21x1_ASAP7_75t_R _36659_ (.A1(net2423),
    .A2(net1118),
    .B(_05908_),
    .Y(_07182_));
 AO21x1_ASAP7_75t_R _36660_ (.A1(net1786),
    .A2(net1560),
    .B(_05908_),
    .Y(_07183_));
 INVx1_ASAP7_75t_R _36661_ (.A(_05908_),
    .Y(_07184_));
 NAND2x1_ASAP7_75t_R _36662_ (.A(_05759_),
    .B(_07184_),
    .Y(_07185_));
 AND3x1_ASAP7_75t_R _36663_ (.A(_07182_),
    .B(_07183_),
    .C(_07185_),
    .Y(_07186_));
 NAND2x1_ASAP7_75t_R _36664_ (.A(_05810_),
    .B(_05816_),
    .Y(_07187_));
 AO21x1_ASAP7_75t_R _36665_ (.A1(_07187_),
    .A2(net2186),
    .B(_05894_),
    .Y(_07189_));
 AO21x1_ASAP7_75t_R _36666_ (.A1(net2422),
    .A2(net3370),
    .B(_05894_),
    .Y(_07190_));
 NAND2x1_ASAP7_75t_R _36667_ (.A(_06515_),
    .B(_05898_),
    .Y(_07191_));
 NAND2x2_ASAP7_75t_R _36668_ (.A(_05776_),
    .B(_05898_),
    .Y(_07192_));
 AND4x1_ASAP7_75t_R _36669_ (.A(_07189_),
    .B(_07190_),
    .C(_07191_),
    .D(_07192_),
    .Y(_07193_));
 NAND2x1_ASAP7_75t_R _36670_ (.A(_07186_),
    .B(_07193_),
    .Y(_07194_));
 NOR2x1_ASAP7_75t_R _36671_ (.A(_07181_),
    .B(_07194_),
    .Y(_07195_));
 AO21x1_ASAP7_75t_R _36672_ (.A1(net1662),
    .A2(net1037),
    .B(_05821_),
    .Y(_07196_));
 AO21x1_ASAP7_75t_R _36673_ (.A1(net2423),
    .A2(_05905_),
    .B(_05821_),
    .Y(_07197_));
 AND2x2_ASAP7_75t_R _36674_ (.A(_07196_),
    .B(_07197_),
    .Y(_07198_));
 AO21x1_ASAP7_75t_R _36675_ (.A1(_05817_),
    .A2(net2845),
    .B(_05821_),
    .Y(_07200_));
 NAND2x1_ASAP7_75t_R _36676_ (.A(_05758_),
    .B(_05829_),
    .Y(_07201_));
 NAND2x1_ASAP7_75t_R _36677_ (.A(_05987_),
    .B(_05829_),
    .Y(_07202_));
 AND3x1_ASAP7_75t_R _36678_ (.A(_07200_),
    .B(_07201_),
    .C(_07202_),
    .Y(_07203_));
 NAND2x2_ASAP7_75t_R _36679_ (.A(_07198_),
    .B(_07203_),
    .Y(_07204_));
 INVx2_ASAP7_75t_R _36680_ (.A(_05854_),
    .Y(_07205_));
 OA21x2_ASAP7_75t_R _36681_ (.A1(_06523_),
    .A2(_06494_),
    .B(_07205_),
    .Y(_07206_));
 NAND2x2_ASAP7_75t_R _36682_ (.A(net1176),
    .B(_05810_),
    .Y(_07207_));
 NOR2x2_ASAP7_75t_R _36683_ (.A(_07207_),
    .B(net2679),
    .Y(_07208_));
 NOR2x2_ASAP7_75t_R _36684_ (.A(_05854_),
    .B(_05918_),
    .Y(_07209_));
 NOR3x2_ASAP7_75t_R _36685_ (.B(_07208_),
    .C(_07209_),
    .Y(_07211_),
    .A(_07206_));
 OA21x2_ASAP7_75t_R _36686_ (.A1(_05985_),
    .A2(_05897_),
    .B(_05846_),
    .Y(_07212_));
 INVx1_ASAP7_75t_R _36687_ (.A(_05866_),
    .Y(_07213_));
 OA21x2_ASAP7_75t_R _36688_ (.A1(_07213_),
    .A2(_05776_),
    .B(_05846_),
    .Y(_07214_));
 NOR3x2_ASAP7_75t_R _36689_ (.B(_07214_),
    .C(_06447_),
    .Y(_07215_),
    .A(_07212_));
 NAND2x2_ASAP7_75t_R _36690_ (.A(_07211_),
    .B(_07215_),
    .Y(_07216_));
 AO21x1_ASAP7_75t_R _36691_ (.A1(_05850_),
    .A2(_06427_),
    .B(_05800_),
    .Y(_07217_));
 AO21x1_ASAP7_75t_R _36692_ (.A1(_05817_),
    .A2(net2485),
    .B(_05800_),
    .Y(_07218_));
 NAND2x1_ASAP7_75t_R _36693_ (.A(_05745_),
    .B(_05765_),
    .Y(_07219_));
 AO21x2_ASAP7_75t_R _36694_ (.A1(_06490_),
    .A2(_07219_),
    .B(_05800_),
    .Y(_07220_));
 NAND3x2_ASAP7_75t_R _36695_ (.B(_07218_),
    .C(_07220_),
    .Y(_07222_),
    .A(_07217_));
 NOR3x2_ASAP7_75t_R _36696_ (.B(_07216_),
    .C(_07222_),
    .Y(_07223_),
    .A(_07204_));
 NAND2x1_ASAP7_75t_R _36697_ (.A(_07195_),
    .B(_07223_),
    .Y(_07224_));
 AO21x1_ASAP7_75t_R _36698_ (.A1(net1037),
    .A2(_06449_),
    .B(_05938_),
    .Y(_07225_));
 OAI21x1_ASAP7_75t_R _36699_ (.A1(_05938_),
    .A2(_05887_),
    .B(_07225_),
    .Y(_07226_));
 OA211x2_ASAP7_75t_R _36700_ (.A1(_05740_),
    .A2(_05810_),
    .B(_06509_),
    .C(_00541_),
    .Y(_07227_));
 NOR2x1_ASAP7_75t_R _36701_ (.A(_07226_),
    .B(_07227_),
    .Y(_07228_));
 INVx4_ASAP7_75t_R _36702_ (.A(_05964_),
    .Y(_07229_));
 AO31x2_ASAP7_75t_R _36703_ (.A1(_07229_),
    .A2(net2098),
    .A3(_05819_),
    .B(net3352),
    .Y(_07230_));
 INVx1_ASAP7_75t_R _36704_ (.A(_05956_),
    .Y(_07231_));
 AO21x1_ASAP7_75t_R _36705_ (.A1(_05825_),
    .A2(net3355),
    .B(net3352),
    .Y(_07233_));
 AND3x1_ASAP7_75t_R _36706_ (.A(_07230_),
    .B(_07231_),
    .C(_07233_),
    .Y(_07234_));
 NAND2x1_ASAP7_75t_R _36707_ (.A(_07228_),
    .B(_07234_),
    .Y(_07235_));
 AO21x1_ASAP7_75t_R _36708_ (.A1(_05817_),
    .A2(_05833_),
    .B(_05752_),
    .Y(_07236_));
 AO21x1_ASAP7_75t_R _36709_ (.A1(net1807),
    .A2(_07207_),
    .B(_05752_),
    .Y(_07237_));
 NAND2x1_ASAP7_75t_R _36710_ (.A(_05751_),
    .B(_05987_),
    .Y(_07238_));
 AND3x1_ASAP7_75t_R _36711_ (.A(_07236_),
    .B(_07237_),
    .C(_07238_),
    .Y(_07239_));
 TAPCELL_ASAP7_75t_R PHY_293 ();
 AO21x1_ASAP7_75t_R _36713_ (.A1(net1662),
    .A2(net1804),
    .B(_05787_),
    .Y(_07241_));
 AO21x1_ASAP7_75t_R _36714_ (.A1(net2098),
    .A2(net2846),
    .B(_05787_),
    .Y(_07242_));
 NOR2x1_ASAP7_75t_R _36715_ (.A(_05807_),
    .B(_05787_),
    .Y(_07244_));
 INVx1_ASAP7_75t_R _36716_ (.A(_07244_),
    .Y(_07245_));
 NAND2x1_ASAP7_75t_R _36717_ (.A(_05930_),
    .B(_05926_),
    .Y(_07246_));
 AND4x1_ASAP7_75t_R _36718_ (.A(_07241_),
    .B(_07242_),
    .C(_07245_),
    .D(_07246_),
    .Y(_07247_));
 NAND2x1_ASAP7_75t_R _36719_ (.A(_07239_),
    .B(_07247_),
    .Y(_07248_));
 NOR2x1_ASAP7_75t_R _36720_ (.A(_07235_),
    .B(_07248_),
    .Y(_07249_));
 AO21x1_ASAP7_75t_R _36721_ (.A1(net1787),
    .A2(net3370),
    .B(_05993_),
    .Y(_07250_));
 AND3x1_ASAP7_75t_R _36722_ (.A(_06001_),
    .B(_07250_),
    .C(_06004_),
    .Y(_07251_));
 AO21x1_ASAP7_75t_R _36723_ (.A1(_05819_),
    .A2(net2231),
    .B(_06007_),
    .Y(_07252_));
 AO21x1_ASAP7_75t_R _36724_ (.A1(net1804),
    .A2(net1560),
    .B(_06007_),
    .Y(_07253_));
 AO21x1_ASAP7_75t_R _36725_ (.A1(net3370),
    .A2(net2416),
    .B(_06007_),
    .Y(_07255_));
 NAND2x1_ASAP7_75t_R _36726_ (.A(net2517),
    .B(_06017_),
    .Y(_07256_));
 AND4x1_ASAP7_75t_R _36727_ (.A(_07252_),
    .B(_07253_),
    .C(_07255_),
    .D(_07256_),
    .Y(_07257_));
 NAND2x1_ASAP7_75t_R _36728_ (.A(_07251_),
    .B(_07257_),
    .Y(_07258_));
 OA21x2_ASAP7_75t_R _36729_ (.A1(_06015_),
    .A2(_05976_),
    .B(net2636),
    .Y(_07259_));
 NAND2x2_ASAP7_75t_R _36730_ (.A(_05811_),
    .B(_05966_),
    .Y(_07260_));
 NAND2x2_ASAP7_75t_R _36731_ (.A(_05966_),
    .B(_06481_),
    .Y(_07261_));
 NAND2x1_ASAP7_75t_R _36732_ (.A(_07260_),
    .B(_07261_),
    .Y(_07262_));
 AOI211x1_ASAP7_75t_R _36733_ (.A1(net2636),
    .A2(_06494_),
    .B(_07259_),
    .C(_07262_),
    .Y(_07263_));
 AO21x1_ASAP7_75t_R _36734_ (.A1(net2271),
    .A2(net2485),
    .B(_05977_),
    .Y(_07264_));
 AO21x1_ASAP7_75t_R _36735_ (.A1(net1118),
    .A2(_05887_),
    .B(_05977_),
    .Y(_07266_));
 OA211x2_ASAP7_75t_R _36736_ (.A1(net1037),
    .A2(_05977_),
    .B(_07264_),
    .C(_07266_),
    .Y(_07267_));
 NAND2x1_ASAP7_75t_R _36737_ (.A(_07263_),
    .B(_07267_),
    .Y(_07268_));
 NOR2x1_ASAP7_75t_R _36738_ (.A(_07258_),
    .B(_07268_),
    .Y(_07269_));
 NAND2x1_ASAP7_75t_R _36739_ (.A(_07249_),
    .B(_07269_),
    .Y(_07270_));
 NOR2x2_ASAP7_75t_R _36740_ (.A(_07224_),
    .B(_07270_),
    .Y(_07271_));
 INVx2_ASAP7_75t_R _36741_ (.A(_07271_),
    .Y(_07272_));
 AOI21x1_ASAP7_75t_R _36742_ (.A1(_07160_),
    .A2(_07167_),
    .B(_07272_),
    .Y(_07273_));
 NAND2x2_ASAP7_75t_R _36743_ (.A(_07159_),
    .B(_07049_),
    .Y(_07274_));
 NAND2x2_ASAP7_75t_R _36744_ (.A(_07050_),
    .B(_07165_),
    .Y(_07275_));
 AOI21x1_ASAP7_75t_R _36745_ (.A1(_07274_),
    .A2(_07275_),
    .B(_07271_),
    .Y(_07277_));
 NAND2x1_ASAP7_75t_R _36746_ (.A(_06817_),
    .B(_06245_),
    .Y(_07278_));
 AO21x1_ASAP7_75t_R _36747_ (.A1(_06129_),
    .A2(_06039_),
    .B(_06240_),
    .Y(_07279_));
 NAND2x1_ASAP7_75t_R _36748_ (.A(_07278_),
    .B(_07279_),
    .Y(_07280_));
 AO21x1_ASAP7_75t_R _36749_ (.A1(net1215),
    .A2(_06050_),
    .B(_06240_),
    .Y(_07281_));
 TAPCELL_ASAP7_75t_R PHY_292 ();
 AO21x1_ASAP7_75t_R _36751_ (.A1(_06190_),
    .A2(net2590),
    .B(_06240_),
    .Y(_07283_));
 NAND2x1_ASAP7_75t_R _36752_ (.A(_07281_),
    .B(_07283_),
    .Y(_07284_));
 NOR2x1_ASAP7_75t_R _36753_ (.A(_07280_),
    .B(_07284_),
    .Y(_07285_));
 AO21x1_ASAP7_75t_R _36754_ (.A1(_06078_),
    .A2(net2590),
    .B(_06229_),
    .Y(_07286_));
 AO21x1_ASAP7_75t_R _36755_ (.A1(net1215),
    .A2(net1628),
    .B(_06229_),
    .Y(_07288_));
 NAND2x1_ASAP7_75t_R _36756_ (.A(_07286_),
    .B(_07288_),
    .Y(_07289_));
 AO21x1_ASAP7_75t_R _36757_ (.A1(_06129_),
    .A2(_06085_),
    .B(_06229_),
    .Y(_07290_));
 OAI21x1_ASAP7_75t_R _36758_ (.A1(net2412),
    .A2(net3330),
    .B(_07290_),
    .Y(_07291_));
 NOR2x1_ASAP7_75t_R _36759_ (.A(_07289_),
    .B(_07291_),
    .Y(_07292_));
 NAND2x1_ASAP7_75t_R _36760_ (.A(_07285_),
    .B(_07292_),
    .Y(_07293_));
 OA21x2_ASAP7_75t_R _36761_ (.A1(_06108_),
    .A2(_06197_),
    .B(_06273_),
    .Y(_07294_));
 NOR2x1_ASAP7_75t_R _36762_ (.A(_06274_),
    .B(_07294_),
    .Y(_07295_));
 OA21x2_ASAP7_75t_R _36763_ (.A1(_06799_),
    .A2(_06261_),
    .B(_06251_),
    .Y(_07296_));
 INVx2_ASAP7_75t_R _36764_ (.A(_06039_),
    .Y(_07297_));
 OA21x2_ASAP7_75t_R _36765_ (.A1(_06817_),
    .A2(_07297_),
    .B(_06251_),
    .Y(_07299_));
 NOR2x1_ASAP7_75t_R _36766_ (.A(_07296_),
    .B(_07299_),
    .Y(_07300_));
 TAPCELL_ASAP7_75t_R PHY_291 ();
 NOR2x1_ASAP7_75t_R _36768_ (.A(_06268_),
    .B(_06181_),
    .Y(_07302_));
 INVx1_ASAP7_75t_R _36769_ (.A(_07302_),
    .Y(_07303_));
 NAND3x1_ASAP7_75t_R _36770_ (.A(_07295_),
    .B(_07300_),
    .C(_07303_),
    .Y(_07304_));
 NOR2x1_ASAP7_75t_R _36771_ (.A(_07293_),
    .B(_07304_),
    .Y(_07305_));
 AO21x1_ASAP7_75t_R _36772_ (.A1(_06096_),
    .A2(net3425),
    .B(_06063_),
    .Y(_07306_));
 AO21x1_ASAP7_75t_R _36773_ (.A1(_07306_),
    .A2(net1217),
    .B(_06191_),
    .Y(_07307_));
 INVx1_ASAP7_75t_R _36774_ (.A(_06733_),
    .Y(_07308_));
 AND2x2_ASAP7_75t_R _36775_ (.A(_07307_),
    .B(_07308_),
    .Y(_07310_));
 TAPCELL_ASAP7_75t_R PHY_290 ();
 AO21x2_ASAP7_75t_R _36777_ (.A1(net2242),
    .A2(net1214),
    .B(_06176_),
    .Y(_07312_));
 AO21x1_ASAP7_75t_R _36778_ (.A1(_06196_),
    .A2(net3329),
    .B(_06176_),
    .Y(_07313_));
 NAND2x1_ASAP7_75t_R _36779_ (.A(_06259_),
    .B(_06781_),
    .Y(_07314_));
 AND3x1_ASAP7_75t_R _36780_ (.A(_07312_),
    .B(_07313_),
    .C(_07314_),
    .Y(_07315_));
 NAND2x1_ASAP7_75t_R _36781_ (.A(_07310_),
    .B(_07315_),
    .Y(_07316_));
 NAND2x1_ASAP7_75t_R _36782_ (.A(net1547),
    .B(net2744),
    .Y(_07317_));
 AO21x1_ASAP7_75t_R _36783_ (.A1(_06181_),
    .A2(_07317_),
    .B(net3235),
    .Y(_07318_));
 AO21x1_ASAP7_75t_R _36784_ (.A1(_06036_),
    .A2(net1540),
    .B(net3235),
    .Y(_07319_));
 AO21x1_ASAP7_75t_R _36785_ (.A1(net3231),
    .A2(net2639),
    .B(net3235),
    .Y(_07321_));
 AND3x1_ASAP7_75t_R _36786_ (.A(_07318_),
    .B(_07319_),
    .C(_07321_),
    .Y(_07322_));
 AND3x2_ASAP7_75t_R _36787_ (.A(_06207_),
    .B(_06097_),
    .C(net1598),
    .Y(_07323_));
 OA21x2_ASAP7_75t_R _36788_ (.A1(_06256_),
    .A2(_06739_),
    .B(_06207_),
    .Y(_07324_));
 NOR2x1_ASAP7_75t_R _36789_ (.A(net1214),
    .B(_06203_),
    .Y(_07325_));
 NOR3x1_ASAP7_75t_R _36790_ (.A(_07323_),
    .B(_07324_),
    .C(_07325_),
    .Y(_07326_));
 NAND2x1_ASAP7_75t_R _36791_ (.A(_07322_),
    .B(_07326_),
    .Y(_07327_));
 NOR2x1_ASAP7_75t_R _36792_ (.A(_07316_),
    .B(_07327_),
    .Y(_07328_));
 NAND2x1_ASAP7_75t_R _36793_ (.A(_07305_),
    .B(_07328_),
    .Y(_07329_));
 OA21x2_ASAP7_75t_R _36794_ (.A1(_06121_),
    .A2(_06126_),
    .B(_06795_),
    .Y(_07330_));
 NOR2x2_ASAP7_75t_R _36795_ (.A(_06047_),
    .B(_06098_),
    .Y(_07332_));
 NAND2x2_ASAP7_75t_R _36796_ (.A(_07332_),
    .B(_06139_),
    .Y(_07333_));
 OA21x2_ASAP7_75t_R _36797_ (.A1(_06146_),
    .A2(_06030_),
    .B(_07333_),
    .Y(_07334_));
 AOI211x1_ASAP7_75t_R _36798_ (.A1(_06029_),
    .A2(net1545),
    .B(_06121_),
    .C(net3433),
    .Y(_07335_));
 AOI211x1_ASAP7_75t_R _36799_ (.A1(_06029_),
    .A2(_06061_),
    .B(_06121_),
    .C(_06141_),
    .Y(_07336_));
 NOR2x1_ASAP7_75t_R _36800_ (.A(_07335_),
    .B(_07336_),
    .Y(_07337_));
 NAND3x1_ASAP7_75t_R _36801_ (.A(_07330_),
    .B(_07334_),
    .C(_07337_),
    .Y(_07338_));
 AO21x1_ASAP7_75t_R _36802_ (.A1(_06190_),
    .A2(_06078_),
    .B(_06158_),
    .Y(_07339_));
 AO21x1_ASAP7_75t_R _36803_ (.A1(net2480),
    .A2(_06181_),
    .B(_06158_),
    .Y(_07340_));
 TAPCELL_ASAP7_75t_R PHY_289 ();
 AO21x1_ASAP7_75t_R _36805_ (.A1(net2639),
    .A2(net3331),
    .B(_06158_),
    .Y(_07343_));
 AND3x1_ASAP7_75t_R _36806_ (.A(_07339_),
    .B(_07340_),
    .C(_07343_),
    .Y(_07344_));
 INVx2_ASAP7_75t_R _36807_ (.A(_07332_),
    .Y(_07345_));
 TAPCELL_ASAP7_75t_R PHY_288 ();
 AO21x1_ASAP7_75t_R _36809_ (.A1(_07345_),
    .A2(_06794_),
    .B(_06151_),
    .Y(_07347_));
 AND3x1_ASAP7_75t_R _36810_ (.A(_07347_),
    .B(_06878_),
    .C(_06880_),
    .Y(_07348_));
 NAND2x1_ASAP7_75t_R _36811_ (.A(_07344_),
    .B(_07348_),
    .Y(_07349_));
 NOR2x1_ASAP7_75t_R _36812_ (.A(_07338_),
    .B(_07349_),
    .Y(_07350_));
 NOR2x2_ASAP7_75t_R _36813_ (.A(_06052_),
    .B(net2786),
    .Y(_07351_));
 NOR2x2_ASAP7_75t_R _36814_ (.A(_06853_),
    .B(net2786),
    .Y(_07352_));
 AOI21x1_ASAP7_75t_R _36815_ (.A1(net1663),
    .A2(_07351_),
    .B(_07352_),
    .Y(_07354_));
 AO21x1_ASAP7_75t_R _36816_ (.A1(net2639),
    .A2(_06089_),
    .B(net2786),
    .Y(_07355_));
 AND2x2_ASAP7_75t_R _36817_ (.A(_07354_),
    .B(_07355_),
    .Y(_07356_));
 INVx1_ASAP7_75t_R _36818_ (.A(_06059_),
    .Y(_07357_));
 AO21x1_ASAP7_75t_R _36819_ (.A1(net2480),
    .A2(_06072_),
    .B(_06064_),
    .Y(_07358_));
 AO21x1_ASAP7_75t_R _36820_ (.A1(_06036_),
    .A2(net3330),
    .B(_06064_),
    .Y(_07359_));
 AND3x1_ASAP7_75t_R _36821_ (.A(_07357_),
    .B(_07358_),
    .C(_07359_),
    .Y(_07360_));
 NAND2x1_ASAP7_75t_R _36822_ (.A(_07356_),
    .B(_07360_),
    .Y(_07361_));
 NAND2x1_ASAP7_75t_R _36823_ (.A(net1602),
    .B(_06092_),
    .Y(_07362_));
 AO21x1_ASAP7_75t_R _36824_ (.A1(_06084_),
    .A2(_06131_),
    .B(_06081_),
    .Y(_07363_));
 NAND2x1_ASAP7_75t_R _36825_ (.A(_07362_),
    .B(_07363_),
    .Y(_07365_));
 NAND2x1_ASAP7_75t_R _36826_ (.A(_07332_),
    .B(_06092_),
    .Y(_07366_));
 AO21x1_ASAP7_75t_R _36827_ (.A1(_06078_),
    .A2(net2590),
    .B(_06081_),
    .Y(_07367_));
 NAND2x1_ASAP7_75t_R _36828_ (.A(_07366_),
    .B(_07367_),
    .Y(_07368_));
 NOR2x1_ASAP7_75t_R _36829_ (.A(_07365_),
    .B(_07368_),
    .Y(_07369_));
 AOI211x1_ASAP7_75t_R _36830_ (.A1(_06029_),
    .A2(_06061_),
    .B(net1589),
    .C(_06104_),
    .Y(_07370_));
 INVx1_ASAP7_75t_R _36831_ (.A(_07370_),
    .Y(_07371_));
 TAPCELL_ASAP7_75t_R PHY_287 ();
 AO21x1_ASAP7_75t_R _36833_ (.A1(_06190_),
    .A2(_06050_),
    .B(_06104_),
    .Y(_07373_));
 AO21x1_ASAP7_75t_R _36834_ (.A1(net3328),
    .A2(_06085_),
    .B(_06104_),
    .Y(_07374_));
 AND3x1_ASAP7_75t_R _36835_ (.A(_07371_),
    .B(_07373_),
    .C(_07374_),
    .Y(_07376_));
 NAND2x1_ASAP7_75t_R _36836_ (.A(_07369_),
    .B(_07376_),
    .Y(_07377_));
 NOR2x1_ASAP7_75t_R _36837_ (.A(_07361_),
    .B(_07377_),
    .Y(_07378_));
 NAND2x1_ASAP7_75t_R _36838_ (.A(_07350_),
    .B(_07378_),
    .Y(_07379_));
 NOR2x1_ASAP7_75t_R _36839_ (.A(_07329_),
    .B(_07379_),
    .Y(_07380_));
 NAND2x2_ASAP7_75t_R _36840_ (.A(_06920_),
    .B(_07380_),
    .Y(_07381_));
 XOR2x1_ASAP7_75t_R _36841_ (.A(net3435),
    .Y(_07382_),
    .B(_07381_));
 OAI21x1_ASAP7_75t_R _36842_ (.A1(_07273_),
    .A2(_07277_),
    .B(_07382_),
    .Y(_07383_));
 AOI21x1_ASAP7_75t_R _36843_ (.A1(_07274_),
    .A2(_07275_),
    .B(_07272_),
    .Y(_07384_));
 AOI21x1_ASAP7_75t_R _36844_ (.A1(_07160_),
    .A2(_07167_),
    .B(_07271_),
    .Y(_07385_));
 INVx1_ASAP7_75t_R _36845_ (.A(_07382_),
    .Y(_07387_));
 OAI21x1_ASAP7_75t_R _36846_ (.A1(_07384_),
    .A2(_07385_),
    .B(_07387_),
    .Y(_07388_));
 AOI21x1_ASAP7_75t_R _36847_ (.A1(_07383_),
    .A2(_07388_),
    .B(net388),
    .Y(_07389_));
 NOR2x2_ASAP7_75t_R _36848_ (.A(_06942_),
    .B(_07389_),
    .Y(_07390_));
 XOR2x1_ASAP7_75t_R _36849_ (.A(_07390_),
    .Y(_00107_),
    .B(_00385_));
 NOR2x2_ASAP7_75t_R _36850_ (.A(net394),
    .B(_00848_),
    .Y(_07391_));
 OR3x1_ASAP7_75t_R _36851_ (.A(_06191_),
    .B(net2756),
    .C(_06259_),
    .Y(_07392_));
 INVx2_ASAP7_75t_R _36852_ (.A(_06150_),
    .Y(_07393_));
 NAND2x1_ASAP7_75t_R _36853_ (.A(_07393_),
    .B(_06781_),
    .Y(_07394_));
 NAND2x1_ASAP7_75t_R _36854_ (.A(_06739_),
    .B(_06781_),
    .Y(_07395_));
 AO21x1_ASAP7_75t_R _36855_ (.A1(_06196_),
    .A2(net1540),
    .B(_06176_),
    .Y(_07397_));
 AND4x1_ASAP7_75t_R _36856_ (.A(_07392_),
    .B(_07394_),
    .C(_07395_),
    .D(_07397_),
    .Y(_07398_));
 AO21x1_ASAP7_75t_R _36857_ (.A1(_06107_),
    .A2(_06196_),
    .B(_06210_),
    .Y(_07399_));
 AO21x1_ASAP7_75t_R _36858_ (.A1(_06129_),
    .A2(_06131_),
    .B(_06210_),
    .Y(_07400_));
 AND2x2_ASAP7_75t_R _36859_ (.A(_07399_),
    .B(_07400_),
    .Y(_07401_));
 INVx1_ASAP7_75t_R _36860_ (.A(_06863_),
    .Y(_07402_));
 AOI211x1_ASAP7_75t_R _36861_ (.A1(_06029_),
    .A2(_06061_),
    .B(_06210_),
    .C(_06098_),
    .Y(_07403_));
 AOI21x1_ASAP7_75t_R _36862_ (.A1(_06212_),
    .A2(_07402_),
    .B(_07403_),
    .Y(_07404_));
 NAND2x1_ASAP7_75t_R _36863_ (.A(_07401_),
    .B(_07404_),
    .Y(_07405_));
 OA21x2_ASAP7_75t_R _36864_ (.A1(net3327),
    .A2(net2482),
    .B(_06207_),
    .Y(_07406_));
 NOR2x1_ASAP7_75t_R _36865_ (.A(_06203_),
    .B(net3330),
    .Y(_07408_));
 NOR2x1_ASAP7_75t_R _36866_ (.A(_06239_),
    .B(_06203_),
    .Y(_07409_));
 OR3x1_ASAP7_75t_R _36867_ (.A(_07406_),
    .B(_07408_),
    .C(_07409_),
    .Y(_07410_));
 NOR2x1_ASAP7_75t_R _36868_ (.A(_07405_),
    .B(_07410_),
    .Y(_07411_));
 NAND2x1_ASAP7_75t_R _36869_ (.A(_07398_),
    .B(_07411_),
    .Y(_07412_));
 AO21x1_ASAP7_75t_R _36870_ (.A1(_06190_),
    .A2(net2590),
    .B(_06250_),
    .Y(_07413_));
 AND2x2_ASAP7_75t_R _36871_ (.A(_07413_),
    .B(_06262_),
    .Y(_07414_));
 AO21x1_ASAP7_75t_R _36872_ (.A1(_06084_),
    .A2(_06085_),
    .B(_06250_),
    .Y(_07415_));
 OA21x2_ASAP7_75t_R _36873_ (.A1(_06250_),
    .A2(_06089_),
    .B(_07415_),
    .Y(_07416_));
 NAND2x1_ASAP7_75t_R _36874_ (.A(_07414_),
    .B(_07416_),
    .Y(_07417_));
 INVx1_ASAP7_75t_R _36875_ (.A(_06750_),
    .Y(_07419_));
 NAND2x1_ASAP7_75t_R _36876_ (.A(_07419_),
    .B(_06273_),
    .Y(_07420_));
 AO21x1_ASAP7_75t_R _36877_ (.A1(_06036_),
    .A2(_06107_),
    .B(_06268_),
    .Y(_07421_));
 NAND2x1_ASAP7_75t_R _36878_ (.A(_07420_),
    .B(_07421_),
    .Y(_07422_));
 AO21x1_ASAP7_75t_R _36879_ (.A1(_06273_),
    .A2(_06138_),
    .B(_07422_),
    .Y(_07423_));
 NOR2x1_ASAP7_75t_R _36880_ (.A(_07417_),
    .B(_07423_),
    .Y(_07424_));
 AO21x1_ASAP7_75t_R _36881_ (.A1(net1260),
    .A2(_06239_),
    .B(_06240_),
    .Y(_07425_));
 AO21x1_ASAP7_75t_R _36882_ (.A1(_06226_),
    .A2(net2614),
    .B(_06240_),
    .Y(_07426_));
 AND2x2_ASAP7_75t_R _36883_ (.A(_07425_),
    .B(_07426_),
    .Y(_07427_));
 AO21x1_ASAP7_75t_R _36884_ (.A1(_06084_),
    .A2(_06089_),
    .B(_06240_),
    .Y(_07428_));
 OA21x2_ASAP7_75t_R _36885_ (.A1(_06240_),
    .A2(_06036_),
    .B(_07428_),
    .Y(_07430_));
 NAND2x1_ASAP7_75t_R _36886_ (.A(_07427_),
    .B(_07430_),
    .Y(_07431_));
 AO21x1_ASAP7_75t_R _36887_ (.A1(_06036_),
    .A2(_06107_),
    .B(_06229_),
    .Y(_07432_));
 AO21x1_ASAP7_75t_R _36888_ (.A1(_06129_),
    .A2(_06039_),
    .B(_06229_),
    .Y(_07433_));
 AND2x2_ASAP7_75t_R _36889_ (.A(_07432_),
    .B(_07433_),
    .Y(_07434_));
 AO21x1_ASAP7_75t_R _36890_ (.A1(_06226_),
    .A2(net2614),
    .B(_06229_),
    .Y(_07435_));
 NOR2x2_ASAP7_75t_R _36891_ (.A(_06229_),
    .B(net1628),
    .Y(_07436_));
 INVx1_ASAP7_75t_R _36892_ (.A(_07436_),
    .Y(_07437_));
 NAND2x1_ASAP7_75t_R _36893_ (.A(_06256_),
    .B(_06775_),
    .Y(_07438_));
 AND3x1_ASAP7_75t_R _36894_ (.A(_07435_),
    .B(_07437_),
    .C(_07438_),
    .Y(_07439_));
 NAND2x1_ASAP7_75t_R _36895_ (.A(_07434_),
    .B(_07439_),
    .Y(_07441_));
 NOR2x1_ASAP7_75t_R _36896_ (.A(_07431_),
    .B(_07441_),
    .Y(_07442_));
 NAND2x2_ASAP7_75t_R _36897_ (.A(_07424_),
    .B(_07442_),
    .Y(_07443_));
 NOR2x2_ASAP7_75t_R _36898_ (.A(_07412_),
    .B(_07443_),
    .Y(_07444_));
 AO21x1_ASAP7_75t_R _36899_ (.A1(net1215),
    .A2(net2590),
    .B(net2399),
    .Y(_07445_));
 AO21x1_ASAP7_75t_R _36900_ (.A1(_06084_),
    .A2(net1217),
    .B(net2399),
    .Y(_07446_));
 NAND2x1_ASAP7_75t_R _36901_ (.A(_06108_),
    .B(_06105_),
    .Y(_07447_));
 NAND3x1_ASAP7_75t_R _36902_ (.A(_07445_),
    .B(_07446_),
    .C(_07447_),
    .Y(_07448_));
 OA21x2_ASAP7_75t_R _36903_ (.A1(_06270_),
    .A2(_06213_),
    .B(_06092_),
    .Y(_07449_));
 AO21x1_ASAP7_75t_R _36904_ (.A1(_06092_),
    .A2(_06108_),
    .B(_07449_),
    .Y(_07450_));
 OA21x2_ASAP7_75t_R _36905_ (.A1(_06193_),
    .A2(_06259_),
    .B(_06092_),
    .Y(_07452_));
 NOR3x1_ASAP7_75t_R _36906_ (.A(_07448_),
    .B(_07450_),
    .C(_07452_),
    .Y(_07453_));
 INVx1_ASAP7_75t_R _36907_ (.A(_06126_),
    .Y(_07454_));
 INVx4_ASAP7_75t_R _36908_ (.A(net2786),
    .Y(_07455_));
 OA21x2_ASAP7_75t_R _36909_ (.A1(_07454_),
    .A2(_06256_),
    .B(_07455_),
    .Y(_07456_));
 OA21x2_ASAP7_75t_R _36910_ (.A1(_06817_),
    .A2(net3432),
    .B(_07455_),
    .Y(_07457_));
 OA21x2_ASAP7_75t_R _36911_ (.A1(net3327),
    .A2(net2482),
    .B(_07455_),
    .Y(_07458_));
 OR3x1_ASAP7_75t_R _36912_ (.A(_07456_),
    .B(_07457_),
    .C(_07458_),
    .Y(_07459_));
 AO21x1_ASAP7_75t_R _36913_ (.A1(net1215),
    .A2(_06050_),
    .B(_06064_),
    .Y(_07460_));
 INVx5_ASAP7_75t_R _36914_ (.A(net2614),
    .Y(_07461_));
 NAND2x1_ASAP7_75t_R _36915_ (.A(_06816_),
    .B(_07461_),
    .Y(_07463_));
 AND2x2_ASAP7_75t_R _36916_ (.A(_07460_),
    .B(_07463_),
    .Y(_07464_));
 NAND2x1_ASAP7_75t_R _36917_ (.A(_06142_),
    .B(_06816_),
    .Y(_07465_));
 OA21x2_ASAP7_75t_R _36918_ (.A1(_06109_),
    .A2(net3432),
    .B(_06816_),
    .Y(_07466_));
 INVx1_ASAP7_75t_R _36919_ (.A(_07466_),
    .Y(_07467_));
 NAND3x1_ASAP7_75t_R _36920_ (.A(_07464_),
    .B(_07465_),
    .C(_07467_),
    .Y(_07468_));
 NOR2x1_ASAP7_75t_R _36921_ (.A(_07459_),
    .B(_07468_),
    .Y(_07469_));
 NAND2x1_ASAP7_75t_R _36922_ (.A(_07453_),
    .B(_07469_),
    .Y(_07470_));
 AO21x1_ASAP7_75t_R _36923_ (.A1(_06078_),
    .A2(_06226_),
    .B(_06151_),
    .Y(_07471_));
 AO21x2_ASAP7_75t_R _36924_ (.A1(_06107_),
    .A2(_06750_),
    .B(_06151_),
    .Y(_07472_));
 NAND3x2_ASAP7_75t_R _36925_ (.B(_07472_),
    .C(_06885_),
    .Y(_07474_),
    .A(_07471_));
 NAND2x2_ASAP7_75t_R _36926_ (.A(_06034_),
    .B(_06128_),
    .Y(_07475_));
 AO21x1_ASAP7_75t_R _36927_ (.A1(_06036_),
    .A2(_07475_),
    .B(net2346),
    .Y(_07476_));
 NAND2x1_ASAP7_75t_R _36928_ (.A(_07393_),
    .B(_06159_),
    .Y(_07477_));
 NAND2x1_ASAP7_75t_R _36929_ (.A(_06817_),
    .B(_06159_),
    .Y(_07478_));
 NAND3x1_ASAP7_75t_R _36930_ (.A(_07476_),
    .B(_07477_),
    .C(_07478_),
    .Y(_07479_));
 NOR2x1_ASAP7_75t_R _36931_ (.A(_06182_),
    .B(net2346),
    .Y(_07480_));
 AO21x1_ASAP7_75t_R _36932_ (.A1(_06799_),
    .A2(_06159_),
    .B(_07480_),
    .Y(_07481_));
 NOR3x1_ASAP7_75t_R _36933_ (.A(_07474_),
    .B(_07479_),
    .C(_07481_),
    .Y(_07482_));
 AOI21x1_ASAP7_75t_R _36934_ (.A1(_06219_),
    .A2(_06099_),
    .B(_06121_),
    .Y(_07483_));
 OA21x2_ASAP7_75t_R _36935_ (.A1(net3327),
    .A2(_06270_),
    .B(_06764_),
    .Y(_07485_));
 NOR2x1_ASAP7_75t_R _36936_ (.A(_06121_),
    .B(_07475_),
    .Y(_07486_));
 OR3x1_ASAP7_75t_R _36937_ (.A(_07483_),
    .B(_07485_),
    .C(_07486_),
    .Y(_07487_));
 AO21x1_ASAP7_75t_R _36938_ (.A1(_07345_),
    .A2(_06050_),
    .B(_06710_),
    .Y(_07488_));
 OA21x2_ASAP7_75t_R _36939_ (.A1(_06710_),
    .A2(_06841_),
    .B(_07488_),
    .Y(_07489_));
 AO21x1_ASAP7_75t_R _36940_ (.A1(_07475_),
    .A2(_06036_),
    .B(_06710_),
    .Y(_07490_));
 NAND2x1_ASAP7_75t_R _36941_ (.A(_06139_),
    .B(_06108_),
    .Y(_07491_));
 NAND2x1_ASAP7_75t_R _36942_ (.A(_06270_),
    .B(_06139_),
    .Y(_07492_));
 AND3x1_ASAP7_75t_R _36943_ (.A(_07490_),
    .B(_07491_),
    .C(_07492_),
    .Y(_07493_));
 NAND2x1_ASAP7_75t_R _36944_ (.A(_07489_),
    .B(_07493_),
    .Y(_07494_));
 NOR2x1_ASAP7_75t_R _36945_ (.A(_07487_),
    .B(_07494_),
    .Y(_07496_));
 NAND2x1_ASAP7_75t_R _36946_ (.A(_07482_),
    .B(_07496_),
    .Y(_07497_));
 NOR2x2_ASAP7_75t_R _36947_ (.A(_07470_),
    .B(_07497_),
    .Y(_07498_));
 NAND2x2_ASAP7_75t_R _36948_ (.A(_07444_),
    .B(_07498_),
    .Y(_07499_));
 XOR2x2_ASAP7_75t_R _36949_ (.A(_07499_),
    .B(_06729_),
    .Y(_07500_));
 AO21x2_ASAP7_75t_R _36950_ (.A1(_05929_),
    .A2(_05844_),
    .B(net2184),
    .Y(_07501_));
 AO21x1_ASAP7_75t_R _36951_ (.A1(_07501_),
    .A2(net2423),
    .B(net3352),
    .Y(_07502_));
 NAND2x1_ASAP7_75t_R _36952_ (.A(net2518),
    .B(_06509_),
    .Y(_07503_));
 NOR2x1_ASAP7_75t_R _36953_ (.A(net3371),
    .B(_05938_),
    .Y(_07504_));
 INVx1_ASAP7_75t_R _36954_ (.A(_07504_),
    .Y(_07505_));
 AO21x1_ASAP7_75t_R _36955_ (.A1(net2271),
    .A2(_05747_),
    .B(_05938_),
    .Y(_07507_));
 AND4x1_ASAP7_75t_R _36956_ (.A(_07502_),
    .B(_07503_),
    .C(_07505_),
    .D(_07507_),
    .Y(_07508_));
 AO31x2_ASAP7_75t_R _36957_ (.A1(net1560),
    .A2(net2423),
    .A3(net3375),
    .B(_05752_),
    .Y(_07509_));
 AO21x1_ASAP7_75t_R _36958_ (.A1(net1913),
    .A2(net2271),
    .B(_05752_),
    .Y(_07510_));
 AO21x1_ASAP7_75t_R _36959_ (.A1(_05833_),
    .A2(net2485),
    .B(_05752_),
    .Y(_07511_));
 NAND3x1_ASAP7_75t_R _36960_ (.A(_07509_),
    .B(_07510_),
    .C(_07511_),
    .Y(_07512_));
 AOI21x1_ASAP7_75t_R _36961_ (.A1(_05926_),
    .A2(_05880_),
    .B(_05932_),
    .Y(_07513_));
 AND3x1_ASAP7_75t_R _36962_ (.A(_05926_),
    .B(_05816_),
    .C(_05757_),
    .Y(_07514_));
 AOI21x1_ASAP7_75t_R _36963_ (.A1(_05926_),
    .A2(_07178_),
    .B(_07514_),
    .Y(_07515_));
 NAND2x1_ASAP7_75t_R _36964_ (.A(_07513_),
    .B(_07515_),
    .Y(_07516_));
 NOR2x1_ASAP7_75t_R _36965_ (.A(_07512_),
    .B(_07516_),
    .Y(_07518_));
 NAND2x1_ASAP7_75t_R _36966_ (.A(_07508_),
    .B(_07518_),
    .Y(_07519_));
 OA21x2_ASAP7_75t_R _36967_ (.A1(_05880_),
    .A2(_06015_),
    .B(net2636),
    .Y(_07520_));
 AO21x1_ASAP7_75t_R _36968_ (.A1(net2636),
    .A2(_06523_),
    .B(_07520_),
    .Y(_07521_));
 INVx1_ASAP7_75t_R _36969_ (.A(_05966_),
    .Y(_07522_));
 AO21x1_ASAP7_75t_R _36970_ (.A1(net2743),
    .A2(_05835_),
    .B(_07522_),
    .Y(_07523_));
 NAND2x1_ASAP7_75t_R _36971_ (.A(_06527_),
    .B(_07523_),
    .Y(_07524_));
 AO21x1_ASAP7_75t_R _36972_ (.A1(_07168_),
    .A2(net2485),
    .B(_05977_),
    .Y(_07525_));
 OAI21x1_ASAP7_75t_R _36973_ (.A1(net2706),
    .A2(_05977_),
    .B(_07525_),
    .Y(_07526_));
 NOR3x1_ASAP7_75t_R _36974_ (.A(_07521_),
    .B(_07524_),
    .C(_07526_),
    .Y(_07527_));
 AO21x1_ASAP7_75t_R _36975_ (.A1(net1913),
    .A2(net2271),
    .B(net2525),
    .Y(_07529_));
 AND2x2_ASAP7_75t_R _36976_ (.A(_07529_),
    .B(_06004_),
    .Y(_07530_));
 AO21x1_ASAP7_75t_R _36977_ (.A1(net1804),
    .A2(net1037),
    .B(net2525),
    .Y(_07531_));
 OA21x2_ASAP7_75t_R _36978_ (.A1(net1118),
    .A2(net2525),
    .B(_07531_),
    .Y(_07532_));
 NAND2x1_ASAP7_75t_R _36979_ (.A(_07530_),
    .B(_07532_),
    .Y(_07533_));
 AO21x1_ASAP7_75t_R _36980_ (.A1(net2875),
    .A2(net2229),
    .B(_06007_),
    .Y(_07534_));
 AO21x1_ASAP7_75t_R _36981_ (.A1(net1118),
    .A2(_05905_),
    .B(_06007_),
    .Y(_07535_));
 AND2x2_ASAP7_75t_R _36982_ (.A(_07534_),
    .B(_07535_),
    .Y(_07536_));
 NAND2x1_ASAP7_75t_R _36983_ (.A(_06017_),
    .B(_06481_),
    .Y(_07537_));
 NAND3x1_ASAP7_75t_R _36984_ (.A(_07536_),
    .B(_07537_),
    .C(_06536_),
    .Y(_07538_));
 NOR2x1_ASAP7_75t_R _36985_ (.A(_07533_),
    .B(_07538_),
    .Y(_07540_));
 NAND2x1_ASAP7_75t_R _36986_ (.A(_07527_),
    .B(_07540_),
    .Y(_07541_));
 NOR2x1_ASAP7_75t_R _36987_ (.A(_07519_),
    .B(_07541_),
    .Y(_07542_));
 AO21x1_ASAP7_75t_R _36988_ (.A1(_05850_),
    .A2(_07187_),
    .B(_05894_),
    .Y(_07543_));
 AO21x1_ASAP7_75t_R _36989_ (.A1(net1118),
    .A2(net980),
    .B(_05894_),
    .Y(_07544_));
 NAND3x1_ASAP7_75t_R _36990_ (.A(_07543_),
    .B(_07544_),
    .C(_07192_),
    .Y(_07545_));
 AO21x1_ASAP7_75t_R _36991_ (.A1(_07168_),
    .A2(_05835_),
    .B(_05908_),
    .Y(_07546_));
 NAND2x1_ASAP7_75t_R _36992_ (.A(net1177),
    .B(_07184_),
    .Y(_07547_));
 AO21x2_ASAP7_75t_R _36993_ (.A1(net2876),
    .A2(net3466),
    .B(_05908_),
    .Y(_07548_));
 NAND3x1_ASAP7_75t_R _36994_ (.A(_07546_),
    .B(_07547_),
    .C(_07548_),
    .Y(_07549_));
 NOR2x1_ASAP7_75t_R _36995_ (.A(_07545_),
    .B(_07549_),
    .Y(_07551_));
 AO21x1_ASAP7_75t_R _36996_ (.A1(net1037),
    .A2(net2738),
    .B(_05884_),
    .Y(_07552_));
 AO21x1_ASAP7_75t_R _36997_ (.A1(_07501_),
    .A2(_05835_),
    .B(_05884_),
    .Y(_07553_));
 NAND2x1_ASAP7_75t_R _36998_ (.A(_07552_),
    .B(_07553_),
    .Y(_07554_));
 AO21x1_ASAP7_75t_R _36999_ (.A1(net1806),
    .A2(net1560),
    .B(_05873_),
    .Y(_07555_));
 AO21x1_ASAP7_75t_R _37000_ (.A1(net1118),
    .A2(_05905_),
    .B(_05873_),
    .Y(_07556_));
 AND2x2_ASAP7_75t_R _37001_ (.A(_07555_),
    .B(_07556_),
    .Y(_07557_));
 AO21x1_ASAP7_75t_R _37002_ (.A1(net3470),
    .A2(net2845),
    .B(_05873_),
    .Y(_07558_));
 AO21x1_ASAP7_75t_R _37003_ (.A1(net2098),
    .A2(net2082),
    .B(_05873_),
    .Y(_07559_));
 NAND2x1_ASAP7_75t_R _37004_ (.A(_05845_),
    .B(_05878_),
    .Y(_07560_));
 AND3x1_ASAP7_75t_R _37005_ (.A(_07558_),
    .B(_07559_),
    .C(_07560_),
    .Y(_07562_));
 NAND2x1_ASAP7_75t_R _37006_ (.A(_07557_),
    .B(_07562_),
    .Y(_07563_));
 NOR2x1_ASAP7_75t_R _37007_ (.A(_07554_),
    .B(_07563_),
    .Y(_07564_));
 NAND2x1_ASAP7_75t_R _37008_ (.A(_07551_),
    .B(_07564_),
    .Y(_07565_));
 AO21x1_ASAP7_75t_R _37009_ (.A1(_05850_),
    .A2(net2081),
    .B(net3351),
    .Y(_07566_));
 AO21x1_ASAP7_75t_R _37010_ (.A1(net1560),
    .A2(_05905_),
    .B(net3351),
    .Y(_07567_));
 NAND3x1_ASAP7_75t_R _37011_ (.A(_07566_),
    .B(_07567_),
    .C(_07201_),
    .Y(_07568_));
 NOR2x2_ASAP7_75t_R _37012_ (.A(net1694),
    .B(_05800_),
    .Y(_07569_));
 AOI211x1_ASAP7_75t_R _37013_ (.A1(net1183),
    .A2(_05812_),
    .B(_06439_),
    .C(_07569_),
    .Y(_07570_));
 NAND2x1_ASAP7_75t_R _37014_ (.A(net3348),
    .B(_05812_),
    .Y(_07571_));
 AO21x1_ASAP7_75t_R _37015_ (.A1(_07229_),
    .A2(net2485),
    .B(_05800_),
    .Y(_07573_));
 NAND3x1_ASAP7_75t_R _37016_ (.A(_07570_),
    .B(_07571_),
    .C(_07573_),
    .Y(_07574_));
 NOR2x1_ASAP7_75t_R _37017_ (.A(_07568_),
    .B(_07574_),
    .Y(_07575_));
 AO21x1_ASAP7_75t_R _37018_ (.A1(net2743),
    .A2(_05835_),
    .B(_05839_),
    .Y(_07576_));
 AO21x1_ASAP7_75t_R _37019_ (.A1(_05850_),
    .A2(net2081),
    .B(_05839_),
    .Y(_07577_));
 AO21x1_ASAP7_75t_R _37020_ (.A1(_05921_),
    .A2(net3375),
    .B(_05839_),
    .Y(_07578_));
 NAND3x1_ASAP7_75t_R _37021_ (.A(_07576_),
    .B(_07577_),
    .C(_07578_),
    .Y(_07579_));
 AO21x1_ASAP7_75t_R _37022_ (.A1(net1695),
    .A2(net1560),
    .B(_05854_),
    .Y(_07580_));
 AO21x1_ASAP7_75t_R _37023_ (.A1(net2288),
    .A2(net2737),
    .B(_05854_),
    .Y(_07581_));
 NAND2x1_ASAP7_75t_R _37024_ (.A(_07205_),
    .B(_05880_),
    .Y(_07582_));
 AND3x1_ASAP7_75t_R _37025_ (.A(_07580_),
    .B(_07581_),
    .C(_07582_),
    .Y(_07584_));
 AO21x1_ASAP7_75t_R _37026_ (.A1(_05817_),
    .A2(net3467),
    .B(_05854_),
    .Y(_07585_));
 NOR2x1_ASAP7_75t_R _37027_ (.A(_05854_),
    .B(net2098),
    .Y(_07586_));
 INVx1_ASAP7_75t_R _37028_ (.A(_07586_),
    .Y(_07587_));
 AND3x1_ASAP7_75t_R _37029_ (.A(_05856_),
    .B(_07585_),
    .C(_07587_),
    .Y(_07588_));
 NAND2x1_ASAP7_75t_R _37030_ (.A(_07584_),
    .B(_07588_),
    .Y(_07589_));
 NOR2x1_ASAP7_75t_R _37031_ (.A(_07579_),
    .B(_07589_),
    .Y(_07590_));
 NAND2x1_ASAP7_75t_R _37032_ (.A(_07575_),
    .B(_07590_),
    .Y(_07591_));
 NOR2x2_ASAP7_75t_R _37033_ (.A(_07565_),
    .B(_07591_),
    .Y(_07592_));
 NAND2x2_ASAP7_75t_R _37034_ (.A(_07592_),
    .B(_07542_),
    .Y(_07593_));
 XOR2x1_ASAP7_75t_R _37035_ (.A(_07500_),
    .Y(_07595_),
    .B(_07593_));
 XOR2x2_ASAP7_75t_R _37036_ (.A(net3165),
    .B(_05715_),
    .Y(_07596_));
 AO21x1_ASAP7_75t_R _37037_ (.A1(net2146),
    .A2(net1140),
    .B(net2621),
    .Y(_07597_));
 NAND2x1_ASAP7_75t_R _37038_ (.A(_05205_),
    .B(_05108_),
    .Y(_07598_));
 NAND3x1_ASAP7_75t_R _37039_ (.A(_06356_),
    .B(_07597_),
    .C(_07598_),
    .Y(_07599_));
 NOR2x2_ASAP7_75t_R _37040_ (.A(net3105),
    .B(net3107),
    .Y(_07600_));
 NOR2x1_ASAP7_75t_R _37041_ (.A(net2469),
    .B(net2493),
    .Y(_07601_));
 NOR2x1_ASAP7_75t_R _37042_ (.A(_05122_),
    .B(net2493),
    .Y(_07602_));
 OR3x1_ASAP7_75t_R _37043_ (.A(_07600_),
    .B(_07601_),
    .C(_07602_),
    .Y(_07603_));
 INVx1_ASAP7_75t_R _37044_ (.A(net3426),
    .Y(_07604_));
 OA21x2_ASAP7_75t_R _37045_ (.A1(_07604_),
    .A2(_05113_),
    .B(_05108_),
    .Y(_07606_));
 NOR3x1_ASAP7_75t_R _37046_ (.A(_07599_),
    .B(_07603_),
    .C(_07606_),
    .Y(_07607_));
 AO21x1_ASAP7_75t_R _37047_ (.A1(net1867),
    .A2(net1091),
    .B(_05086_),
    .Y(_07608_));
 NAND2x1_ASAP7_75t_R _37048_ (.A(net1149),
    .B(net2225),
    .Y(_07609_));
 AO21x1_ASAP7_75t_R _37049_ (.A1(_07609_),
    .A2(net992),
    .B(_05086_),
    .Y(_07610_));
 NAND2x1_ASAP7_75t_R _37050_ (.A(_05203_),
    .B(_05087_),
    .Y(_07611_));
 NAND3x1_ASAP7_75t_R _37051_ (.A(_07608_),
    .B(_07610_),
    .C(_07611_),
    .Y(_07612_));
 AOI22x1_ASAP7_75t_R _37052_ (.A1(_06328_),
    .A2(net1304),
    .B1(_05308_),
    .B2(_05175_),
    .Y(_07613_));
 NAND2x2_ASAP7_75t_R _37053_ (.A(_05110_),
    .B(_05175_),
    .Y(_07614_));
 AO21x1_ASAP7_75t_R _37054_ (.A1(net992),
    .A2(_05259_),
    .B(net2529),
    .Y(_07615_));
 NAND3x1_ASAP7_75t_R _37055_ (.A(_07613_),
    .B(_07614_),
    .C(_07615_),
    .Y(_07617_));
 NOR2x1_ASAP7_75t_R _37056_ (.A(_07612_),
    .B(_07617_),
    .Y(_07618_));
 NAND2x1_ASAP7_75t_R _37057_ (.A(_07607_),
    .B(_07618_),
    .Y(_07619_));
 AO31x2_ASAP7_75t_R _37058_ (.A1(net1794),
    .A2(net3453),
    .A3(net990),
    .B(_05153_),
    .Y(_07620_));
 NOR2x1_ASAP7_75t_R _37059_ (.A(_05233_),
    .B(_05153_),
    .Y(_07621_));
 INVx1_ASAP7_75t_R _37060_ (.A(_07621_),
    .Y(_07622_));
 AO21x1_ASAP7_75t_R _37061_ (.A1(net1867),
    .A2(net1091),
    .B(_05153_),
    .Y(_07623_));
 NAND3x1_ASAP7_75t_R _37062_ (.A(_07620_),
    .B(_07622_),
    .C(_07623_),
    .Y(_07624_));
 OA21x2_ASAP7_75t_R _37063_ (.A1(_06323_),
    .A2(_05238_),
    .B(_05100_),
    .Y(_07625_));
 NOR2x1_ASAP7_75t_R _37064_ (.A(net3451),
    .B(_05306_),
    .Y(_07626_));
 INVx1_ASAP7_75t_R _37065_ (.A(_05101_),
    .Y(_07628_));
 OR3x1_ASAP7_75t_R _37066_ (.A(_07625_),
    .B(_07626_),
    .C(_07628_),
    .Y(_07629_));
 NOR2x1_ASAP7_75t_R _37067_ (.A(_07624_),
    .B(_07629_),
    .Y(_07630_));
 OA21x2_ASAP7_75t_R _37068_ (.A1(_05178_),
    .A2(net2161),
    .B(_05420_),
    .Y(_07631_));
 AO21x1_ASAP7_75t_R _37069_ (.A1(_05422_),
    .A2(_05420_),
    .B(_07631_),
    .Y(_07632_));
 INVx1_ASAP7_75t_R _37070_ (.A(_05309_),
    .Y(_07633_));
 NOR2x1_ASAP7_75t_R _37071_ (.A(net1894),
    .B(_05186_),
    .Y(_07634_));
 NOR2x1_ASAP7_75t_R _37072_ (.A(_05186_),
    .B(net3102),
    .Y(_07635_));
 OR3x1_ASAP7_75t_R _37073_ (.A(_07633_),
    .B(_07634_),
    .C(_07635_),
    .Y(_07636_));
 AOI211x1_ASAP7_75t_R _37074_ (.A1(_05106_),
    .A2(_05247_),
    .B(_07632_),
    .C(_07636_),
    .Y(_07637_));
 NAND2x1_ASAP7_75t_R _37075_ (.A(_07630_),
    .B(_07637_),
    .Y(_07639_));
 NOR2x1_ASAP7_75t_R _37076_ (.A(_07619_),
    .B(_07639_),
    .Y(_07640_));
 OA21x2_ASAP7_75t_R _37077_ (.A1(_05200_),
    .A2(_05218_),
    .B(_05201_),
    .Y(_07641_));
 NAND2x1_ASAP7_75t_R _37078_ (.A(_06400_),
    .B(_05121_),
    .Y(_07642_));
 NOR2x1_ASAP7_75t_R _37079_ (.A(_07641_),
    .B(_07642_),
    .Y(_07643_));
 AOI211x1_ASAP7_75t_R _37080_ (.A1(net1324),
    .A2(net3442),
    .B(_05118_),
    .C(_05345_),
    .Y(_07644_));
 NAND2x1_ASAP7_75t_R _37081_ (.A(_05096_),
    .B(_05201_),
    .Y(_07645_));
 INVx1_ASAP7_75t_R _37082_ (.A(_05360_),
    .Y(_07646_));
 NAND2x1_ASAP7_75t_R _37083_ (.A(_07646_),
    .B(_05201_),
    .Y(_07647_));
 NAND2x1_ASAP7_75t_R _37084_ (.A(_07645_),
    .B(_07647_),
    .Y(_07648_));
 NOR2x1_ASAP7_75t_R _37085_ (.A(_07644_),
    .B(_07648_),
    .Y(_07650_));
 NAND2x1_ASAP7_75t_R _37086_ (.A(_07643_),
    .B(_07650_),
    .Y(_07651_));
 AO21x1_ASAP7_75t_R _37087_ (.A1(_05206_),
    .A2(_05143_),
    .B(_05138_),
    .Y(_07652_));
 AO21x1_ASAP7_75t_R _37088_ (.A1(net1921),
    .A2(net1237),
    .B(_05138_),
    .Y(_07653_));
 AND2x2_ASAP7_75t_R _37089_ (.A(_07652_),
    .B(_07653_),
    .Y(_07654_));
 AO21x1_ASAP7_75t_R _37090_ (.A1(net1822),
    .A2(net1836),
    .B(_05138_),
    .Y(_07655_));
 OA21x2_ASAP7_75t_R _37091_ (.A1(net990),
    .A2(_05138_),
    .B(_07655_),
    .Y(_07656_));
 NAND2x1_ASAP7_75t_R _37092_ (.A(_07654_),
    .B(_07656_),
    .Y(_07657_));
 NOR2x1_ASAP7_75t_R _37093_ (.A(_07651_),
    .B(_07657_),
    .Y(_07658_));
 AO21x1_ASAP7_75t_R _37094_ (.A1(_05360_),
    .A2(net2027),
    .B(_05062_),
    .Y(_07659_));
 OA21x2_ASAP7_75t_R _37095_ (.A1(_05345_),
    .A2(_05062_),
    .B(_07659_),
    .Y(_07661_));
 AO21x1_ASAP7_75t_R _37096_ (.A1(_05265_),
    .A2(_05165_),
    .B(_05062_),
    .Y(_07662_));
 OA21x2_ASAP7_75t_R _37097_ (.A1(net1921),
    .A2(_05062_),
    .B(_07662_),
    .Y(_07663_));
 NAND2x1_ASAP7_75t_R _37098_ (.A(_07661_),
    .B(_07663_),
    .Y(_07664_));
 INVx2_ASAP7_75t_R _37099_ (.A(_06996_),
    .Y(_07665_));
 NOR2x1_ASAP7_75t_R _37100_ (.A(_05356_),
    .B(_07665_),
    .Y(_07666_));
 AO21x1_ASAP7_75t_R _37101_ (.A1(net1921),
    .A2(net1237),
    .B(net3412),
    .Y(_07667_));
 NAND3x1_ASAP7_75t_R _37102_ (.A(_07666_),
    .B(_06989_),
    .C(_07667_),
    .Y(_07668_));
 NOR2x1_ASAP7_75t_R _37103_ (.A(_07664_),
    .B(_07668_),
    .Y(_07669_));
 NAND2x2_ASAP7_75t_R _37104_ (.A(_07658_),
    .B(_07669_),
    .Y(_07670_));
 AO21x1_ASAP7_75t_R _37105_ (.A1(_05143_),
    .A2(_05122_),
    .B(_05198_),
    .Y(_07672_));
 NAND2x1_ASAP7_75t_R _37106_ (.A(net1485),
    .B(_05199_),
    .Y(_07673_));
 NAND3x1_ASAP7_75t_R _37107_ (.A(_05338_),
    .B(_07672_),
    .C(_07673_),
    .Y(_07674_));
 OA21x2_ASAP7_75t_R _37108_ (.A1(_05178_),
    .A2(_06956_),
    .B(_05332_),
    .Y(_07675_));
 AO21x1_ASAP7_75t_R _37109_ (.A1(net992),
    .A2(net990),
    .B(_05208_),
    .Y(_07676_));
 NAND2x1_ASAP7_75t_R _37110_ (.A(_06960_),
    .B(_07676_),
    .Y(_07677_));
 NOR3x1_ASAP7_75t_R _37111_ (.A(_07674_),
    .B(_07675_),
    .C(_07677_),
    .Y(_07678_));
 AO21x1_ASAP7_75t_R _37112_ (.A1(net1921),
    .A2(net1894),
    .B(_05256_),
    .Y(_07679_));
 INVx1_ASAP7_75t_R _37113_ (.A(_07679_),
    .Y(_07680_));
 NOR2x1_ASAP7_75t_R _37114_ (.A(_05143_),
    .B(_05256_),
    .Y(_07681_));
 AOI21x1_ASAP7_75t_R _37115_ (.A1(net964),
    .A2(net1879),
    .B(_05256_),
    .Y(_07683_));
 OR3x1_ASAP7_75t_R _37116_ (.A(_07680_),
    .B(_07681_),
    .C(_07683_),
    .Y(_07684_));
 AO21x1_ASAP7_75t_R _37117_ (.A1(net2139),
    .A2(net1793),
    .B(net3095),
    .Y(_07685_));
 AO21x1_ASAP7_75t_R _37118_ (.A1(net992),
    .A2(_05259_),
    .B(net3095),
    .Y(_07686_));
 AND2x2_ASAP7_75t_R _37119_ (.A(_07685_),
    .B(_07686_),
    .Y(_07687_));
 AO21x1_ASAP7_75t_R _37120_ (.A1(net1766),
    .A2(net1237),
    .B(_05240_),
    .Y(_07688_));
 AO21x1_ASAP7_75t_R _37121_ (.A1(net3101),
    .A2(net2314),
    .B(_05240_),
    .Y(_07689_));
 NAND2x1_ASAP7_75t_R _37122_ (.A(_05178_),
    .B(_05241_),
    .Y(_07690_));
 AND3x1_ASAP7_75t_R _37123_ (.A(_07688_),
    .B(_07689_),
    .C(_07690_),
    .Y(_07691_));
 NAND2x1_ASAP7_75t_R _37124_ (.A(_07687_),
    .B(_07691_),
    .Y(_07692_));
 NOR2x1_ASAP7_75t_R _37125_ (.A(_07684_),
    .B(_07692_),
    .Y(_07694_));
 NAND2x1_ASAP7_75t_R _37126_ (.A(_07678_),
    .B(_07694_),
    .Y(_07695_));
 NOR2x2_ASAP7_75t_R _37127_ (.A(_07670_),
    .B(_07695_),
    .Y(_07696_));
 NAND2x2_ASAP7_75t_R _37128_ (.A(_07640_),
    .B(_07696_),
    .Y(_07697_));
 AO21x1_ASAP7_75t_R _37129_ (.A1(net1627),
    .A2(net1267),
    .B(_05581_),
    .Y(_07698_));
 NAND2x1_ASAP7_75t_R _37130_ (.A(_05656_),
    .B(_05577_),
    .Y(_07699_));
 NAND2x2_ASAP7_75t_R _37131_ (.A(_05577_),
    .B(_05664_),
    .Y(_07700_));
 AND3x1_ASAP7_75t_R _37132_ (.A(_07698_),
    .B(_07699_),
    .C(_07700_),
    .Y(_07701_));
 AO21x1_ASAP7_75t_R _37133_ (.A1(net2658),
    .A2(net1267),
    .B(net2389),
    .Y(_07702_));
 OA21x2_ASAP7_75t_R _37134_ (.A1(net2568),
    .A2(net2389),
    .B(_07702_),
    .Y(_07703_));
 AND2x2_ASAP7_75t_R _37135_ (.A(_07701_),
    .B(_07703_),
    .Y(_07705_));
 AO21x1_ASAP7_75t_R _37136_ (.A1(net2663),
    .A2(net1124),
    .B(_05472_),
    .Y(_07706_));
 AO21x1_ASAP7_75t_R _37137_ (.A1(_05685_),
    .A2(_06568_),
    .B(_05472_),
    .Y(_07707_));
 NAND2x2_ASAP7_75t_R _37138_ (.A(_05600_),
    .B(_05682_),
    .Y(_07708_));
 NAND3x2_ASAP7_75t_R _37139_ (.B(_07707_),
    .C(_07708_),
    .Y(_07709_),
    .A(_07706_));
 AO21x1_ASAP7_75t_R _37140_ (.A1(net3349),
    .A2(net2509),
    .B(_05453_),
    .Y(_07710_));
 AO21x1_ASAP7_75t_R _37141_ (.A1(net1627),
    .A2(net2153),
    .B(_05453_),
    .Y(_07711_));
 NAND2x2_ASAP7_75t_R _37142_ (.A(_07710_),
    .B(_07711_),
    .Y(_07712_));
 AO21x1_ASAP7_75t_R _37143_ (.A1(net2568),
    .A2(net2032),
    .B(_05453_),
    .Y(_07713_));
 OAI21x1_ASAP7_75t_R _37144_ (.A1(net1124),
    .A2(_05453_),
    .B(_07713_),
    .Y(_07714_));
 NOR3x2_ASAP7_75t_R _37145_ (.B(_07712_),
    .C(_07714_),
    .Y(_07716_),
    .A(_07709_));
 NAND2x2_ASAP7_75t_R _37146_ (.A(_07705_),
    .B(_07716_),
    .Y(_07717_));
 AO21x2_ASAP7_75t_R _37147_ (.A1(net1627),
    .A2(net2659),
    .B(_05492_),
    .Y(_07718_));
 NAND2x2_ASAP7_75t_R _37148_ (.A(_05484_),
    .B(_07152_),
    .Y(_07719_));
 NAND2x2_ASAP7_75t_R _37149_ (.A(_05439_),
    .B(_05484_),
    .Y(_07720_));
 NAND3x2_ASAP7_75t_R _37150_ (.B(_07719_),
    .C(_07720_),
    .Y(_07721_),
    .A(_07718_));
 OA21x2_ASAP7_75t_R _37151_ (.A1(net2834),
    .A2(_05463_),
    .B(net3373),
    .Y(_07722_));
 NOR2x2_ASAP7_75t_R _37152_ (.A(_07722_),
    .B(_06643_),
    .Y(_07723_));
 AO21x1_ASAP7_75t_R _37153_ (.A1(net2220),
    .A2(net2032),
    .B(_05511_),
    .Y(_07724_));
 NAND2x2_ASAP7_75t_R _37154_ (.A(net3164),
    .B(net2511),
    .Y(_07725_));
 NAND3x2_ASAP7_75t_R _37155_ (.B(_07724_),
    .C(_07725_),
    .Y(_07727_),
    .A(_07723_));
 NOR2x2_ASAP7_75t_R _37156_ (.A(_07721_),
    .B(_07727_),
    .Y(_07728_));
 AO21x1_ASAP7_75t_R _37157_ (.A1(net3462),
    .A2(net2836),
    .B(net2755),
    .Y(_07729_));
 OAI21x1_ASAP7_75t_R _37158_ (.A1(_06647_),
    .A2(net3106),
    .B(_06627_),
    .Y(_07730_));
 AND3x1_ASAP7_75t_R _37159_ (.A(_07729_),
    .B(_07064_),
    .C(_07730_),
    .Y(_07731_));
 AO21x1_ASAP7_75t_R _37160_ (.A1(net1084),
    .A2(_05580_),
    .B(_05548_),
    .Y(_07732_));
 OA21x2_ASAP7_75t_R _37161_ (.A1(_05520_),
    .A2(_05514_),
    .B(_05545_),
    .Y(_07733_));
 INVx1_ASAP7_75t_R _37162_ (.A(_07733_),
    .Y(_07734_));
 NAND2x1_ASAP7_75t_R _37163_ (.A(_07732_),
    .B(_07734_),
    .Y(_07735_));
 NAND2x1_ASAP7_75t_R _37164_ (.A(_07066_),
    .B(_05545_),
    .Y(_07736_));
 INVx1_ASAP7_75t_R _37165_ (.A(_06621_),
    .Y(_07738_));
 NAND2x1_ASAP7_75t_R _37166_ (.A(_07736_),
    .B(_07738_),
    .Y(_07739_));
 NOR2x1_ASAP7_75t_R _37167_ (.A(_07735_),
    .B(_07739_),
    .Y(_07740_));
 NAND2x2_ASAP7_75t_R _37168_ (.A(_07731_),
    .B(_07740_),
    .Y(_07741_));
 INVx1_ASAP7_75t_R _37169_ (.A(_07741_),
    .Y(_07742_));
 NAND2x2_ASAP7_75t_R _37170_ (.A(_07728_),
    .B(_07742_),
    .Y(_07743_));
 NOR2x2_ASAP7_75t_R _37171_ (.A(_07717_),
    .B(_07743_),
    .Y(_07744_));
 AO21x1_ASAP7_75t_R _37172_ (.A1(net2658),
    .A2(net1267),
    .B(_05616_),
    .Y(_07745_));
 AO21x1_ASAP7_75t_R _37173_ (.A1(net1124),
    .A2(net3115),
    .B(net2447),
    .Y(_07746_));
 NAND3x1_ASAP7_75t_R _37174_ (.A(_07745_),
    .B(_07746_),
    .C(_07131_),
    .Y(_07747_));
 NOR2x2_ASAP7_75t_R _37175_ (.A(net2116),
    .B(_05626_),
    .Y(_07749_));
 AOI211x1_ASAP7_75t_R _37176_ (.A1(net1033),
    .A2(_05627_),
    .B(_07749_),
    .C(_06601_),
    .Y(_07750_));
 NAND2x1_ASAP7_75t_R _37177_ (.A(_05674_),
    .B(_05627_),
    .Y(_07751_));
 AO21x1_ASAP7_75t_R _37178_ (.A1(_05496_),
    .A2(net2509),
    .B(_05626_),
    .Y(_07752_));
 NAND3x1_ASAP7_75t_R _37179_ (.A(_07750_),
    .B(_07751_),
    .C(_07752_),
    .Y(_07753_));
 NOR2x1_ASAP7_75t_R _37180_ (.A(_07747_),
    .B(_07753_),
    .Y(_07754_));
 AO21x1_ASAP7_75t_R _37181_ (.A1(net2220),
    .A2(_05580_),
    .B(net2616),
    .Y(_07755_));
 AO21x1_ASAP7_75t_R _37182_ (.A1(net2400),
    .A2(net1124),
    .B(net2616),
    .Y(_07756_));
 AND2x2_ASAP7_75t_R _37183_ (.A(_07755_),
    .B(_07756_),
    .Y(_07757_));
 AOI211x1_ASAP7_75t_R _37184_ (.A1(net2814),
    .A2(net3098),
    .B(net2616),
    .C(net1668),
    .Y(_07758_));
 INVx1_ASAP7_75t_R _37185_ (.A(_05598_),
    .Y(_07760_));
 AND3x1_ASAP7_75t_R _37186_ (.A(_07760_),
    .B(_05461_),
    .C(_05647_),
    .Y(_07761_));
 NOR2x1_ASAP7_75t_R _37187_ (.A(_07758_),
    .B(_07761_),
    .Y(_07762_));
 NAND2x1_ASAP7_75t_R _37188_ (.A(_07757_),
    .B(_07762_),
    .Y(_07763_));
 AOI211x1_ASAP7_75t_R _37189_ (.A1(net1000),
    .A2(net989),
    .B(_05634_),
    .C(_05440_),
    .Y(_07764_));
 AOI21x1_ASAP7_75t_R _37190_ (.A1(_05516_),
    .A2(_06593_),
    .B(_07764_),
    .Y(_07765_));
 AO21x1_ASAP7_75t_R _37191_ (.A1(net3350),
    .A2(_05464_),
    .B(net2462),
    .Y(_07766_));
 AO21x1_ASAP7_75t_R _37192_ (.A1(net2658),
    .A2(net1267),
    .B(net2462),
    .Y(_07767_));
 NAND3x1_ASAP7_75t_R _37193_ (.A(_07765_),
    .B(_07766_),
    .C(_07767_),
    .Y(_07768_));
 NOR2x1_ASAP7_75t_R _37194_ (.A(_07763_),
    .B(_07768_),
    .Y(_07769_));
 NAND2x2_ASAP7_75t_R _37195_ (.A(_07754_),
    .B(_07769_),
    .Y(_07771_));
 AOI21x1_ASAP7_75t_R _37196_ (.A1(net2698),
    .A2(_06574_),
    .B(_05654_),
    .Y(_07772_));
 NOR2x1_ASAP7_75t_R _37197_ (.A(_05655_),
    .B(_07772_),
    .Y(_07773_));
 AO21x1_ASAP7_75t_R _37198_ (.A1(net1627),
    .A2(net1267),
    .B(_05654_),
    .Y(_07774_));
 OA21x2_ASAP7_75t_R _37199_ (.A1(_05464_),
    .A2(_05654_),
    .B(_07774_),
    .Y(_07775_));
 NAND2x1_ASAP7_75t_R _37200_ (.A(_07773_),
    .B(_07775_),
    .Y(_07776_));
 NAND2x1_ASAP7_75t_R _37201_ (.A(_05461_),
    .B(_05661_),
    .Y(_07777_));
 NAND2x1_ASAP7_75t_R _37202_ (.A(_05674_),
    .B(_05661_),
    .Y(_07778_));
 OAI21x1_ASAP7_75t_R _37203_ (.A1(net2320),
    .A2(_07777_),
    .B(_07778_),
    .Y(_07779_));
 OA21x2_ASAP7_75t_R _37204_ (.A1(_05664_),
    .A2(_05516_),
    .B(_05661_),
    .Y(_07780_));
 NOR2x2_ASAP7_75t_R _37205_ (.A(_05605_),
    .B(_06576_),
    .Y(_07782_));
 NOR3x1_ASAP7_75t_R _37206_ (.A(_07779_),
    .B(_07780_),
    .C(_07782_),
    .Y(_07783_));
 INVx1_ASAP7_75t_R _37207_ (.A(_07783_),
    .Y(_07784_));
 NOR2x1_ASAP7_75t_R _37208_ (.A(_07776_),
    .B(_07784_),
    .Y(_07785_));
 AO21x1_ASAP7_75t_R _37209_ (.A1(net2003),
    .A2(net2477),
    .B(_05677_),
    .Y(_07786_));
 INVx1_ASAP7_75t_R _37210_ (.A(_07786_),
    .Y(_07787_));
 AO21x1_ASAP7_75t_R _37211_ (.A1(net3250),
    .A2(_05503_),
    .B(_05677_),
    .Y(_07788_));
 OAI21x1_ASAP7_75t_R _37212_ (.A1(_05464_),
    .A2(_05677_),
    .B(_07788_),
    .Y(_07789_));
 NOR2x1_ASAP7_75t_R _37213_ (.A(_07787_),
    .B(_07789_),
    .Y(_07790_));
 INVx1_ASAP7_75t_R _37214_ (.A(_07790_),
    .Y(_07791_));
 AOI211x1_ASAP7_75t_R _37215_ (.A1(net1000),
    .A2(net3111),
    .B(_05683_),
    .C(net1674),
    .Y(_07793_));
 INVx1_ASAP7_75t_R _37216_ (.A(_07793_),
    .Y(_07794_));
 AO21x1_ASAP7_75t_R _37217_ (.A1(net3349),
    .A2(net2509),
    .B(_05683_),
    .Y(_07795_));
 AND2x2_ASAP7_75t_R _37218_ (.A(_07794_),
    .B(_07795_),
    .Y(_07796_));
 AO21x1_ASAP7_75t_R _37219_ (.A1(net2401),
    .A2(net3461),
    .B(_05683_),
    .Y(_07797_));
 AO21x1_ASAP7_75t_R _37220_ (.A1(net2033),
    .A2(net2477),
    .B(_05683_),
    .Y(_07798_));
 NAND2x2_ASAP7_75t_R _37221_ (.A(net3106),
    .B(_05684_),
    .Y(_07799_));
 AND3x2_ASAP7_75t_R _37222_ (.A(_07797_),
    .B(_07798_),
    .C(_07799_),
    .Y(_07800_));
 NAND2x1_ASAP7_75t_R _37223_ (.A(_07796_),
    .B(_07800_),
    .Y(_07801_));
 NOR2x1_ASAP7_75t_R _37224_ (.A(_07791_),
    .B(_07801_),
    .Y(_07802_));
 NAND2x1_ASAP7_75t_R _37225_ (.A(_07785_),
    .B(_07802_),
    .Y(_07804_));
 NOR2x2_ASAP7_75t_R _37226_ (.A(_07771_),
    .B(_07804_),
    .Y(_07805_));
 NAND2x2_ASAP7_75t_R _37227_ (.A(_07744_),
    .B(_07805_),
    .Y(_07806_));
 XOR2x2_ASAP7_75t_R _37228_ (.A(_07697_),
    .B(_07806_),
    .Y(_07807_));
 XOR2x1_ASAP7_75t_R _37229_ (.A(_07596_),
    .Y(_07808_),
    .B(_07807_));
 NOR2x1_ASAP7_75t_R _37230_ (.A(_07595_),
    .B(_07808_),
    .Y(_07809_));
 INVx1_ASAP7_75t_R _37231_ (.A(_07593_),
    .Y(_07810_));
 XOR2x1_ASAP7_75t_R _37232_ (.A(_07500_),
    .Y(_07811_),
    .B(_07810_));
 XOR2x2_ASAP7_75t_R _37233_ (.A(net3165),
    .B(_05427_),
    .Y(_07812_));
 XOR2x1_ASAP7_75t_R _37234_ (.A(_07812_),
    .Y(_07813_),
    .B(_07807_));
 NOR2x1_ASAP7_75t_R _37235_ (.A(_07811_),
    .B(_07813_),
    .Y(_07815_));
 OAI21x1_ASAP7_75t_R _37236_ (.A1(_07809_),
    .A2(_07815_),
    .B(net394),
    .Y(_07816_));
 INVx1_ASAP7_75t_R _37237_ (.A(_07816_),
    .Y(_07817_));
 OAI21x1_ASAP7_75t_R _37238_ (.A1(_07391_),
    .A2(_07817_),
    .B(_00386_),
    .Y(_07818_));
 INVx1_ASAP7_75t_R _37239_ (.A(_07391_),
    .Y(_07819_));
 NAND3x1_ASAP7_75t_R _37240_ (.A(_07816_),
    .B(_17145_),
    .C(_07819_),
    .Y(_07820_));
 NAND2x1_ASAP7_75t_R _37241_ (.A(_07820_),
    .B(_07818_),
    .Y(_00108_));
 AND2x2_ASAP7_75t_R _37242_ (.A(net388),
    .B(_00847_),
    .Y(_07821_));
 NOR2x1_ASAP7_75t_R _37243_ (.A(net1215),
    .B(net2786),
    .Y(_07822_));
 AOI21x1_ASAP7_75t_R _37244_ (.A1(_06058_),
    .A2(_07351_),
    .B(_07822_),
    .Y(_07823_));
 NAND2x2_ASAP7_75t_R _37245_ (.A(_06828_),
    .B(_07455_),
    .Y(_07825_));
 AO21x1_ASAP7_75t_R _37246_ (.A1(net3231),
    .A2(_06039_),
    .B(net2786),
    .Y(_07826_));
 NAND3x1_ASAP7_75t_R _37247_ (.A(_07823_),
    .B(_07825_),
    .C(_07826_),
    .Y(_07827_));
 AO21x1_ASAP7_75t_R _37248_ (.A1(net1215),
    .A2(_06181_),
    .B(_06064_),
    .Y(_07828_));
 AND2x2_ASAP7_75t_R _37249_ (.A(_07828_),
    .B(_07463_),
    .Y(_07829_));
 AO21x1_ASAP7_75t_R _37250_ (.A1(_07475_),
    .A2(net3330),
    .B(_06064_),
    .Y(_07830_));
 AND2x2_ASAP7_75t_R _37251_ (.A(_07830_),
    .B(_07465_),
    .Y(_07831_));
 NAND2x1_ASAP7_75t_R _37252_ (.A(_07829_),
    .B(_07831_),
    .Y(_07832_));
 NOR2x1_ASAP7_75t_R _37253_ (.A(_07827_),
    .B(_07832_),
    .Y(_07833_));
 AO21x1_ASAP7_75t_R _37254_ (.A1(_06092_),
    .A2(_06109_),
    .B(_06830_),
    .Y(_07834_));
 AOI211x1_ASAP7_75t_R _37255_ (.A1(net1276),
    .A2(_06061_),
    .B(_06052_),
    .C(_06081_),
    .Y(_07836_));
 INVx1_ASAP7_75t_R _37256_ (.A(_07836_),
    .Y(_07837_));
 NAND2x1_ASAP7_75t_R _37257_ (.A(_07366_),
    .B(_07837_),
    .Y(_07838_));
 NOR2x1_ASAP7_75t_R _37258_ (.A(_07834_),
    .B(_07838_),
    .Y(_07839_));
 AO21x1_ASAP7_75t_R _37259_ (.A1(net1215),
    .A2(net2234),
    .B(_06104_),
    .Y(_07840_));
 AO21x1_ASAP7_75t_R _37260_ (.A1(_06029_),
    .A2(_00630_),
    .B(net1812),
    .Y(_07841_));
 AO21x1_ASAP7_75t_R _37261_ (.A1(_06089_),
    .A2(_07841_),
    .B(_06104_),
    .Y(_07842_));
 NAND2x2_ASAP7_75t_R _37262_ (.A(_07461_),
    .B(_06105_),
    .Y(_07843_));
 AND3x1_ASAP7_75t_R _37263_ (.A(_07840_),
    .B(_07842_),
    .C(_07843_),
    .Y(_07844_));
 AND2x2_ASAP7_75t_R _37264_ (.A(_07839_),
    .B(_07844_),
    .Y(_07845_));
 NAND2x1_ASAP7_75t_R _37265_ (.A(_07833_),
    .B(_07845_),
    .Y(_07847_));
 AO21x1_ASAP7_75t_R _37266_ (.A1(_06278_),
    .A2(net2234),
    .B(_06710_),
    .Y(_07848_));
 NAND2x1_ASAP7_75t_R _37267_ (.A(_06256_),
    .B(_06139_),
    .Y(_07849_));
 NAND2x1_ASAP7_75t_R _37268_ (.A(net2813),
    .B(_06139_),
    .Y(_07850_));
 AND3x1_ASAP7_75t_R _37269_ (.A(_07848_),
    .B(_07849_),
    .C(_07850_),
    .Y(_07851_));
 AO21x1_ASAP7_75t_R _37270_ (.A1(net2480),
    .A2(_06050_),
    .B(_06121_),
    .Y(_07852_));
 OA21x2_ASAP7_75t_R _37271_ (.A1(_06121_),
    .A2(net3328),
    .B(_07852_),
    .Y(_07853_));
 AND2x2_ASAP7_75t_R _37272_ (.A(_07851_),
    .B(_07853_),
    .Y(_07854_));
 AO21x1_ASAP7_75t_R _37273_ (.A1(net3328),
    .A2(net2639),
    .B(_06151_),
    .Y(_07855_));
 OA21x2_ASAP7_75t_R _37274_ (.A1(net1541),
    .A2(_06151_),
    .B(_07855_),
    .Y(_07856_));
 AO21x1_ASAP7_75t_R _37275_ (.A1(_06278_),
    .A2(_06181_),
    .B(_06151_),
    .Y(_07858_));
 OA21x2_ASAP7_75t_R _37276_ (.A1(_06072_),
    .A2(_06151_),
    .B(_07858_),
    .Y(_07859_));
 NAND2x1_ASAP7_75t_R _37277_ (.A(_07856_),
    .B(_07859_),
    .Y(_07860_));
 NOR2x1_ASAP7_75t_R _37278_ (.A(_06129_),
    .B(net2344),
    .Y(_07861_));
 OA21x2_ASAP7_75t_R _37279_ (.A1(_07402_),
    .A2(_06261_),
    .B(_06159_),
    .Y(_07862_));
 OR3x1_ASAP7_75t_R _37280_ (.A(_06742_),
    .B(_07861_),
    .C(_07862_),
    .Y(_07863_));
 NOR2x1_ASAP7_75t_R _37281_ (.A(_07860_),
    .B(_07863_),
    .Y(_07864_));
 NAND2x2_ASAP7_75t_R _37282_ (.A(_07854_),
    .B(_07864_),
    .Y(_07865_));
 NOR2x2_ASAP7_75t_R _37283_ (.A(_07847_),
    .B(_07865_),
    .Y(_07866_));
 AO21x1_ASAP7_75t_R _37284_ (.A1(_07306_),
    .A2(net3329),
    .B(_06176_),
    .Y(_07867_));
 AO21x1_ASAP7_75t_R _37285_ (.A1(net1214),
    .A2(net2234),
    .B(_06176_),
    .Y(_07869_));
 NAND3x1_ASAP7_75t_R _37286_ (.A(_07867_),
    .B(_07395_),
    .C(_07869_),
    .Y(_07870_));
 OA21x2_ASAP7_75t_R _37287_ (.A1(net3327),
    .A2(net2482),
    .B(_06194_),
    .Y(_07871_));
 AOI21x1_ASAP7_75t_R _37288_ (.A1(_06841_),
    .A2(net2242),
    .B(_06191_),
    .Y(_07872_));
 NOR2x1_ASAP7_75t_R _37289_ (.A(_06089_),
    .B(_06191_),
    .Y(_07873_));
 OR3x1_ASAP7_75t_R _37290_ (.A(_07871_),
    .B(_07872_),
    .C(_07873_),
    .Y(_07874_));
 NOR2x1_ASAP7_75t_R _37291_ (.A(_07870_),
    .B(_07874_),
    .Y(_07875_));
 AO21x1_ASAP7_75t_R _37292_ (.A1(net2242),
    .A2(net2234),
    .B(_06203_),
    .Y(_07876_));
 AO21x1_ASAP7_75t_R _37293_ (.A1(net3330),
    .A2(net1217),
    .B(_06203_),
    .Y(_07877_));
 NAND2x1_ASAP7_75t_R _37294_ (.A(_06739_),
    .B(_06207_),
    .Y(_07878_));
 NAND3x1_ASAP7_75t_R _37295_ (.A(_07876_),
    .B(_07877_),
    .C(_07878_),
    .Y(_07880_));
 AOI211x1_ASAP7_75t_R _37296_ (.A1(net1276),
    .A2(net1548),
    .B(net3235),
    .C(net3329),
    .Y(_07881_));
 OA21x2_ASAP7_75t_R _37297_ (.A1(_06817_),
    .A2(net3432),
    .B(_06212_),
    .Y(_07882_));
 NOR2x1_ASAP7_75t_R _37298_ (.A(_07881_),
    .B(_07882_),
    .Y(_07883_));
 AOI211x1_ASAP7_75t_R _37299_ (.A1(net1276),
    .A2(_06061_),
    .B(net3235),
    .C(_06098_),
    .Y(_07884_));
 NOR2x1_ASAP7_75t_R _37300_ (.A(net3235),
    .B(net2590),
    .Y(_07885_));
 AOI211x1_ASAP7_75t_R _37301_ (.A1(_06256_),
    .A2(_06212_),
    .B(_07884_),
    .C(_07885_),
    .Y(_07886_));
 NAND2x1_ASAP7_75t_R _37302_ (.A(_07883_),
    .B(_07886_),
    .Y(_07887_));
 NOR2x1_ASAP7_75t_R _37303_ (.A(_07880_),
    .B(_07887_),
    .Y(_07888_));
 NAND2x1_ASAP7_75t_R _37304_ (.A(_07875_),
    .B(_07888_),
    .Y(_07889_));
 AO21x1_ASAP7_75t_R _37305_ (.A1(_06214_),
    .A2(_06036_),
    .B(_06250_),
    .Y(_07891_));
 AO21x1_ASAP7_75t_R _37306_ (.A1(net2480),
    .A2(net2234),
    .B(_06250_),
    .Y(_07892_));
 AO21x1_ASAP7_75t_R _37307_ (.A1(_06190_),
    .A2(_06794_),
    .B(_06250_),
    .Y(_07893_));
 NAND3x1_ASAP7_75t_R _37308_ (.A(_07891_),
    .B(_07892_),
    .C(_07893_),
    .Y(_07894_));
 AO21x1_ASAP7_75t_R _37309_ (.A1(_06196_),
    .A2(_06118_),
    .B(_06268_),
    .Y(_07895_));
 AO21x1_ASAP7_75t_R _37310_ (.A1(net3328),
    .A2(net3230),
    .B(_06268_),
    .Y(_07896_));
 AND2x2_ASAP7_75t_R _37311_ (.A(_07896_),
    .B(_07895_),
    .Y(_07897_));
 AO21x1_ASAP7_75t_R _37312_ (.A1(_06078_),
    .A2(_06226_),
    .B(_06268_),
    .Y(_07898_));
 AO21x1_ASAP7_75t_R _37313_ (.A1(_06181_),
    .A2(_06070_),
    .B(_06268_),
    .Y(_07899_));
 NAND3x1_ASAP7_75t_R _37314_ (.A(_07897_),
    .B(_07898_),
    .C(_07899_),
    .Y(_07900_));
 NOR2x1_ASAP7_75t_R _37315_ (.A(_07894_),
    .B(_07900_),
    .Y(_07902_));
 NAND2x1_ASAP7_75t_R _37316_ (.A(_06246_),
    .B(_07278_),
    .Y(_07903_));
 AO21x1_ASAP7_75t_R _37317_ (.A1(net1095),
    .A2(_06245_),
    .B(_07903_),
    .Y(_07904_));
 AO21x1_ASAP7_75t_R _37318_ (.A1(_06190_),
    .A2(_06078_),
    .B(_06240_),
    .Y(_07905_));
 NAND2x1_ASAP7_75t_R _37319_ (.A(_07461_),
    .B(_06245_),
    .Y(_07906_));
 INVx1_ASAP7_75t_R _37320_ (.A(_06153_),
    .Y(_07907_));
 NAND2x1_ASAP7_75t_R _37321_ (.A(_06245_),
    .B(_07907_),
    .Y(_07908_));
 NAND3x1_ASAP7_75t_R _37322_ (.A(_07905_),
    .B(_07906_),
    .C(_07908_),
    .Y(_07909_));
 AO21x1_ASAP7_75t_R _37323_ (.A1(net1260),
    .A2(net2234),
    .B(net2412),
    .Y(_07910_));
 AO21x1_ASAP7_75t_R _37324_ (.A1(_06118_),
    .A2(_06039_),
    .B(net2412),
    .Y(_07911_));
 NAND3x1_ASAP7_75t_R _37325_ (.A(_07910_),
    .B(_07911_),
    .C(_07438_),
    .Y(_07913_));
 NOR3x1_ASAP7_75t_R _37326_ (.A(_07904_),
    .B(_07909_),
    .C(_07913_),
    .Y(_07914_));
 NAND2x1_ASAP7_75t_R _37327_ (.A(_07914_),
    .B(_07902_),
    .Y(_07915_));
 NOR2x1_ASAP7_75t_R _37328_ (.A(_07889_),
    .B(_07915_),
    .Y(_07916_));
 NAND2x2_ASAP7_75t_R _37329_ (.A(_07866_),
    .B(_07916_),
    .Y(_07917_));
 XOR2x2_ASAP7_75t_R _37330_ (.A(_07917_),
    .B(_06729_),
    .Y(_07918_));
 NAND2x2_ASAP7_75t_R _37331_ (.A(net1204),
    .B(net1036),
    .Y(_07919_));
 AO21x1_ASAP7_75t_R _37332_ (.A1(net2191),
    .A2(_07919_),
    .B(_05472_),
    .Y(_07920_));
 AO21x1_ASAP7_75t_R _37333_ (.A1(_06568_),
    .A2(net1267),
    .B(_05472_),
    .Y(_07921_));
 NAND2x1_ASAP7_75t_R _37334_ (.A(_05600_),
    .B(_07152_),
    .Y(_07922_));
 AND3x1_ASAP7_75t_R _37335_ (.A(_07920_),
    .B(_07921_),
    .C(_07922_),
    .Y(_07924_));
 OA21x2_ASAP7_75t_R _37336_ (.A1(_05453_),
    .A2(net2658),
    .B(_05465_),
    .Y(_07925_));
 NOR2x1_ASAP7_75t_R _37337_ (.A(net3113),
    .B(_05453_),
    .Y(_07926_));
 AO21x1_ASAP7_75t_R _37338_ (.A1(_05458_),
    .A2(_05515_),
    .B(_07926_),
    .Y(_07927_));
 INVx1_ASAP7_75t_R _37339_ (.A(_07927_),
    .Y(_07928_));
 NAND3x1_ASAP7_75t_R _37340_ (.A(_07924_),
    .B(_07925_),
    .C(_07928_),
    .Y(_07929_));
 AO21x1_ASAP7_75t_R _37341_ (.A1(net1627),
    .A2(net2658),
    .B(net2389),
    .Y(_07930_));
 AO21x1_ASAP7_75t_R _37342_ (.A1(net2191),
    .A2(net3115),
    .B(net2389),
    .Y(_07931_));
 NAND2x1_ASAP7_75t_R _37343_ (.A(_06637_),
    .B(_05564_),
    .Y(_07932_));
 AND3x1_ASAP7_75t_R _37344_ (.A(_07930_),
    .B(_07931_),
    .C(_07932_),
    .Y(_07933_));
 AND2x2_ASAP7_75t_R _37345_ (.A(_05587_),
    .B(_06666_),
    .Y(_07935_));
 AO21x1_ASAP7_75t_R _37346_ (.A1(net2663),
    .A2(net1124),
    .B(_05581_),
    .Y(_07936_));
 NAND2x1_ASAP7_75t_R _37347_ (.A(_05455_),
    .B(_05577_),
    .Y(_07937_));
 AND2x2_ASAP7_75t_R _37348_ (.A(_07936_),
    .B(_07937_),
    .Y(_07938_));
 NAND3x1_ASAP7_75t_R _37349_ (.A(_07933_),
    .B(_07935_),
    .C(_07938_),
    .Y(_07939_));
 NOR2x1_ASAP7_75t_R _37350_ (.A(_07929_),
    .B(_07939_),
    .Y(_07940_));
 NAND2x1_ASAP7_75t_R _37351_ (.A(_05545_),
    .B(_05561_),
    .Y(_07941_));
 AO21x1_ASAP7_75t_R _37352_ (.A1(net3350),
    .A2(net2509),
    .B(_05548_),
    .Y(_07942_));
 NAND2x1_ASAP7_75t_R _37353_ (.A(_07941_),
    .B(_07942_),
    .Y(_07943_));
 AOI211x1_ASAP7_75t_R _37354_ (.A1(net2814),
    .A2(net3111),
    .B(_05548_),
    .C(_05457_),
    .Y(_07944_));
 NOR3x1_ASAP7_75t_R _37355_ (.A(_07943_),
    .B(_07733_),
    .C(_07944_),
    .Y(_07946_));
 AO21x1_ASAP7_75t_R _37356_ (.A1(_06574_),
    .A2(_05619_),
    .B(_05528_),
    .Y(_07947_));
 AO21x1_ASAP7_75t_R _37357_ (.A1(net2833),
    .A2(net2610),
    .B(_05528_),
    .Y(_07948_));
 AO21x1_ASAP7_75t_R _37358_ (.A1(net2032),
    .A2(_05486_),
    .B(_05528_),
    .Y(_07949_));
 NAND3x1_ASAP7_75t_R _37359_ (.A(_07947_),
    .B(_07948_),
    .C(_07949_),
    .Y(_07950_));
 AO21x1_ASAP7_75t_R _37360_ (.A1(net3462),
    .A2(net2870),
    .B(net2755),
    .Y(_07951_));
 AO21x2_ASAP7_75t_R _37361_ (.A1(net2153),
    .A2(_05503_),
    .B(net3118),
    .Y(_07952_));
 NAND2x1_ASAP7_75t_R _37362_ (.A(net2834),
    .B(_06627_),
    .Y(_07953_));
 NAND3x1_ASAP7_75t_R _37363_ (.A(_07951_),
    .B(_07952_),
    .C(_07953_),
    .Y(_07954_));
 NOR2x1_ASAP7_75t_R _37364_ (.A(_07950_),
    .B(_07954_),
    .Y(_07955_));
 NAND2x1_ASAP7_75t_R _37365_ (.A(_07955_),
    .B(_07946_),
    .Y(_07957_));
 OA21x2_ASAP7_75t_R _37366_ (.A1(net1528),
    .A2(_05674_),
    .B(net3374),
    .Y(_07958_));
 NAND2x1_ASAP7_75t_R _37367_ (.A(_06649_),
    .B(_06648_),
    .Y(_07959_));
 AOI211x1_ASAP7_75t_R _37368_ (.A1(net3374),
    .A2(_07152_),
    .B(_07958_),
    .C(_07959_),
    .Y(_07960_));
 AO21x1_ASAP7_75t_R _37369_ (.A1(_05605_),
    .A2(net2036),
    .B(_05492_),
    .Y(_07961_));
 NAND2x1_ASAP7_75t_R _37370_ (.A(_05495_),
    .B(_05484_),
    .Y(_07962_));
 NAND2x1_ASAP7_75t_R _37371_ (.A(_07066_),
    .B(_05484_),
    .Y(_07963_));
 AND4x1_ASAP7_75t_R _37372_ (.A(_05505_),
    .B(_07961_),
    .C(_07962_),
    .D(_07963_),
    .Y(_07964_));
 NAND2x1_ASAP7_75t_R _37373_ (.A(_07960_),
    .B(_07964_),
    .Y(_07965_));
 NOR2x1_ASAP7_75t_R _37374_ (.A(_07957_),
    .B(_07965_),
    .Y(_07966_));
 NAND2x1_ASAP7_75t_R _37375_ (.A(_07940_),
    .B(_07966_),
    .Y(_07968_));
 NOR2x1_ASAP7_75t_R _37376_ (.A(net2411),
    .B(_05496_),
    .Y(_07969_));
 INVx1_ASAP7_75t_R _37377_ (.A(_07969_),
    .Y(_07970_));
 AND3x1_ASAP7_75t_R _37378_ (.A(_07136_),
    .B(_07970_),
    .C(_07138_),
    .Y(_07971_));
 OAI21x1_ASAP7_75t_R _37379_ (.A1(_05642_),
    .A2(_05656_),
    .B(_06613_),
    .Y(_07972_));
 NAND2x2_ASAP7_75t_R _37380_ (.A(_05561_),
    .B(_06613_),
    .Y(_07973_));
 NAND2x1_ASAP7_75t_R _37381_ (.A(_05566_),
    .B(_06613_),
    .Y(_07974_));
 NAND3x1_ASAP7_75t_R _37382_ (.A(_07972_),
    .B(_07973_),
    .C(_07974_),
    .Y(_07975_));
 OA21x2_ASAP7_75t_R _37383_ (.A1(net2661),
    .A2(_05441_),
    .B(_06613_),
    .Y(_07976_));
 AO21x1_ASAP7_75t_R _37384_ (.A1(_05665_),
    .A2(_06613_),
    .B(_07976_),
    .Y(_07977_));
 NOR2x1_ASAP7_75t_R _37385_ (.A(_07975_),
    .B(_07977_),
    .Y(_07979_));
 NAND2x1_ASAP7_75t_R _37386_ (.A(_07971_),
    .B(_07979_),
    .Y(_07980_));
 AO21x1_ASAP7_75t_R _37387_ (.A1(_05613_),
    .A2(net2816),
    .B(net2618),
    .Y(_07981_));
 AO21x1_ASAP7_75t_R _37388_ (.A1(net1903),
    .A2(net1267),
    .B(net2618),
    .Y(_07982_));
 NAND2x1_ASAP7_75t_R _37389_ (.A(_05656_),
    .B(_05647_),
    .Y(_07983_));
 AND3x2_ASAP7_75t_R _37390_ (.A(_07981_),
    .B(_07982_),
    .C(_07983_),
    .Y(_07984_));
 AO21x1_ASAP7_75t_R _37391_ (.A1(net2191),
    .A2(_05457_),
    .B(net2461),
    .Y(_07985_));
 AND2x2_ASAP7_75t_R _37392_ (.A(_07985_),
    .B(_05637_),
    .Y(_07986_));
 OAI21x1_ASAP7_75t_R _37393_ (.A1(_06671_),
    .A2(_05646_),
    .B(_05647_),
    .Y(_07987_));
 NAND3x2_ASAP7_75t_R _37394_ (.B(_07986_),
    .C(_07987_),
    .Y(_07988_),
    .A(_07984_));
 NOR2x2_ASAP7_75t_R _37395_ (.A(_07980_),
    .B(_07988_),
    .Y(_07990_));
 AO21x1_ASAP7_75t_R _37396_ (.A1(net1772),
    .A2(net2509),
    .B(_05654_),
    .Y(_07991_));
 AO21x1_ASAP7_75t_R _37397_ (.A1(_05605_),
    .A2(_05676_),
    .B(_05654_),
    .Y(_07992_));
 AND2x2_ASAP7_75t_R _37398_ (.A(_07991_),
    .B(_07992_),
    .Y(_07993_));
 NOR2x1_ASAP7_75t_R _37399_ (.A(_07782_),
    .B(_05666_),
    .Y(_07994_));
 NAND3x1_ASAP7_75t_R _37400_ (.A(_07993_),
    .B(_07994_),
    .C(_06582_),
    .Y(_07995_));
 AO21x1_ASAP7_75t_R _37401_ (.A1(net1627),
    .A2(_05613_),
    .B(_05683_),
    .Y(_07996_));
 AO21x1_ASAP7_75t_R _37402_ (.A1(net2191),
    .A2(net1083),
    .B(_05683_),
    .Y(_07997_));
 AND3x1_ASAP7_75t_R _37403_ (.A(_07996_),
    .B(_07997_),
    .C(_07799_),
    .Y(_07998_));
 AO21x1_ASAP7_75t_R _37404_ (.A1(net3349),
    .A2(_05613_),
    .B(_05677_),
    .Y(_07999_));
 OA211x2_ASAP7_75t_R _37405_ (.A1(net1267),
    .A2(_05677_),
    .B(_07999_),
    .C(_05679_),
    .Y(_08001_));
 NAND2x1_ASAP7_75t_R _37406_ (.A(_07998_),
    .B(_08001_),
    .Y(_08002_));
 NOR2x1_ASAP7_75t_R _37407_ (.A(_07995_),
    .B(_08002_),
    .Y(_08003_));
 NAND2x2_ASAP7_75t_R _37408_ (.A(_07990_),
    .B(_08003_),
    .Y(_08004_));
 NOR2x2_ASAP7_75t_R _37409_ (.A(_07968_),
    .B(_08004_),
    .Y(_08005_));
 AO21x1_ASAP7_75t_R _37410_ (.A1(_05807_),
    .A2(_05905_),
    .B(_05938_),
    .Y(_08006_));
 AO21x1_ASAP7_75t_R _37411_ (.A1(_05772_),
    .A2(_05796_),
    .B(net2521),
    .Y(_08007_));
 NAND2x1_ASAP7_75t_R _37412_ (.A(_08006_),
    .B(_08007_),
    .Y(_08008_));
 NAND2x1_ASAP7_75t_R _37413_ (.A(_06510_),
    .B(_05948_),
    .Y(_08009_));
 NOR2x1_ASAP7_75t_R _37414_ (.A(_08008_),
    .B(_08009_),
    .Y(_08010_));
 AO21x1_ASAP7_75t_R _37415_ (.A1(net980),
    .A2(net3355),
    .B(net3352),
    .Y(_08012_));
 OAI21x1_ASAP7_75t_R _37416_ (.A1(net1662),
    .A2(net3352),
    .B(_08012_),
    .Y(_08013_));
 OA211x2_ASAP7_75t_R _37417_ (.A1(net1225),
    .A2(_05755_),
    .B(_05953_),
    .C(net2490),
    .Y(_08014_));
 NOR2x1_ASAP7_75t_R _37418_ (.A(_08013_),
    .B(_08014_),
    .Y(_08015_));
 NAND2x1_ASAP7_75t_R _37419_ (.A(_08010_),
    .B(_08015_),
    .Y(_08016_));
 OAI22x1_ASAP7_75t_R _37420_ (.A1(_05780_),
    .A2(net2761),
    .B1(_05772_),
    .B2(_05752_),
    .Y(_08017_));
 AOI211x1_ASAP7_75t_R _37421_ (.A1(net3348),
    .A2(_05751_),
    .B(_08017_),
    .C(_05761_),
    .Y(_08018_));
 AO21x1_ASAP7_75t_R _37422_ (.A1(_05747_),
    .A2(_05876_),
    .B(_05787_),
    .Y(_08019_));
 AO21x1_ASAP7_75t_R _37423_ (.A1(net2423),
    .A2(net3375),
    .B(_05787_),
    .Y(_08020_));
 NAND2x2_ASAP7_75t_R _37424_ (.A(_05985_),
    .B(_05926_),
    .Y(_08021_));
 NAND2x1_ASAP7_75t_R _37425_ (.A(_06523_),
    .B(_05926_),
    .Y(_08023_));
 AND4x1_ASAP7_75t_R _37426_ (.A(_08019_),
    .B(_08020_),
    .C(_08021_),
    .D(_08023_),
    .Y(_08024_));
 NAND2x1_ASAP7_75t_R _37427_ (.A(_08018_),
    .B(_08024_),
    .Y(_08025_));
 NOR2x2_ASAP7_75t_R _37428_ (.A(_08016_),
    .B(_08025_),
    .Y(_08026_));
 AO21x1_ASAP7_75t_R _37429_ (.A1(net2271),
    .A2(_05918_),
    .B(_05977_),
    .Y(_08027_));
 AO21x1_ASAP7_75t_R _37430_ (.A1(_06490_),
    .A2(net3375),
    .B(_05977_),
    .Y(_08028_));
 AND3x1_ASAP7_75t_R _37431_ (.A(_05984_),
    .B(_08027_),
    .C(_08028_),
    .Y(_08029_));
 AND2x2_ASAP7_75t_R _37432_ (.A(_06524_),
    .B(_06525_),
    .Y(_08030_));
 AO21x1_ASAP7_75t_R _37433_ (.A1(_05850_),
    .A2(net1913),
    .B(_07522_),
    .Y(_08031_));
 AND2x2_ASAP7_75t_R _37434_ (.A(_06528_),
    .B(_08031_),
    .Y(_08032_));
 NAND3x1_ASAP7_75t_R _37435_ (.A(_08029_),
    .B(_08030_),
    .C(_08032_),
    .Y(_08034_));
 AO21x1_ASAP7_75t_R _37436_ (.A1(_05876_),
    .A2(_05918_),
    .B(net2525),
    .Y(_08035_));
 OAI21x1_ASAP7_75t_R _37437_ (.A1(net2743),
    .A2(net2525),
    .B(_08035_),
    .Y(_08036_));
 AO21x1_ASAP7_75t_R _37438_ (.A1(net3471),
    .A2(_06449_),
    .B(_05993_),
    .Y(_08037_));
 OAI21x1_ASAP7_75t_R _37439_ (.A1(_05957_),
    .A2(net2525),
    .B(_08037_),
    .Y(_08038_));
 NOR2x1_ASAP7_75t_R _37440_ (.A(_08036_),
    .B(_08038_),
    .Y(_08039_));
 AO21x1_ASAP7_75t_R _37441_ (.A1(net2422),
    .A2(net1118),
    .B(_06007_),
    .Y(_08040_));
 AND3x1_ASAP7_75t_R _37442_ (.A(_07534_),
    .B(_08040_),
    .C(_06533_),
    .Y(_08041_));
 NOR2x1_ASAP7_75t_R _37443_ (.A(net2098),
    .B(_06007_),
    .Y(_08042_));
 NOR2x2_ASAP7_75t_R _37444_ (.A(net2485),
    .B(_06007_),
    .Y(_08043_));
 AOI211x1_ASAP7_75t_R _37445_ (.A1(_05897_),
    .A2(_06017_),
    .B(_08042_),
    .C(_08043_),
    .Y(_08045_));
 NAND3x1_ASAP7_75t_R _37446_ (.A(_08039_),
    .B(_08041_),
    .C(_08045_),
    .Y(_08046_));
 NOR2x1_ASAP7_75t_R _37447_ (.A(_08046_),
    .B(_08034_),
    .Y(_08047_));
 NAND2x2_ASAP7_75t_R _37448_ (.A(_08026_),
    .B(_08047_),
    .Y(_08048_));
 AO21x1_ASAP7_75t_R _37449_ (.A1(_06490_),
    .A2(_07207_),
    .B(_05908_),
    .Y(_08049_));
 AO21x1_ASAP7_75t_R _37450_ (.A1(net1913),
    .A2(net2485),
    .B(_05908_),
    .Y(_08050_));
 NAND2x1_ASAP7_75t_R _37451_ (.A(_08049_),
    .B(_08050_),
    .Y(_08051_));
 NAND2x1_ASAP7_75t_R _37452_ (.A(_07192_),
    .B(_05906_),
    .Y(_08052_));
 OR3x1_ASAP7_75t_R _37453_ (.A(_06460_),
    .B(_08051_),
    .C(_08052_),
    .Y(_08053_));
 AO21x1_ASAP7_75t_R _37454_ (.A1(net1662),
    .A2(net1037),
    .B(_05873_),
    .Y(_08054_));
 AO21x1_ASAP7_75t_R _37455_ (.A1(_05817_),
    .A2(net2271),
    .B(_05873_),
    .Y(_08056_));
 NAND2x1_ASAP7_75t_R _37456_ (.A(_06521_),
    .B(_05878_),
    .Y(_08057_));
 AND3x1_ASAP7_75t_R _37457_ (.A(_08054_),
    .B(_08056_),
    .C(_08057_),
    .Y(_08058_));
 OA21x2_ASAP7_75t_R _37458_ (.A1(_05811_),
    .A2(net2517),
    .B(_05885_),
    .Y(_08059_));
 AO21x1_ASAP7_75t_R _37459_ (.A1(net2403),
    .A2(_05885_),
    .B(_08059_),
    .Y(_08060_));
 NOR2x1_ASAP7_75t_R _37460_ (.A(_05889_),
    .B(_08060_),
    .Y(_08061_));
 NAND2x1_ASAP7_75t_R _37461_ (.A(_08058_),
    .B(_08061_),
    .Y(_08062_));
 NOR2x1_ASAP7_75t_R _37462_ (.A(_08053_),
    .B(_08062_),
    .Y(_08063_));
 AO21x1_ASAP7_75t_R _37463_ (.A1(_05850_),
    .A2(net1913),
    .B(_05800_),
    .Y(_08064_));
 NAND2x1_ASAP7_75t_R _37464_ (.A(_05964_),
    .B(_05812_),
    .Y(_08065_));
 NAND3x1_ASAP7_75t_R _37465_ (.A(_08064_),
    .B(_07220_),
    .C(_08065_),
    .Y(_08067_));
 AO21x1_ASAP7_75t_R _37466_ (.A1(net2743),
    .A2(net3467),
    .B(net3351),
    .Y(_08068_));
 NAND2x1_ASAP7_75t_R _37467_ (.A(_06472_),
    .B(_05829_),
    .Y(_08069_));
 NAND2x1_ASAP7_75t_R _37468_ (.A(_05811_),
    .B(_05829_),
    .Y(_08070_));
 NAND3x1_ASAP7_75t_R _37469_ (.A(_08068_),
    .B(_08069_),
    .C(_08070_),
    .Y(_08071_));
 AO21x1_ASAP7_75t_R _37470_ (.A1(net1662),
    .A2(_06490_),
    .B(net3351),
    .Y(_08072_));
 OAI21x1_ASAP7_75t_R _37471_ (.A1(net3351),
    .A2(_05905_),
    .B(_08072_),
    .Y(_08073_));
 NOR3x1_ASAP7_75t_R _37472_ (.A(_08067_),
    .B(_08071_),
    .C(_08073_),
    .Y(_08074_));
 AOI211x1_ASAP7_75t_R _37473_ (.A1(net1227),
    .A2(net1775),
    .B(net2679),
    .C(net1443),
    .Y(_08075_));
 OA21x2_ASAP7_75t_R _37474_ (.A1(_06481_),
    .A2(net2403),
    .B(_07205_),
    .Y(_08076_));
 NOR2x1_ASAP7_75t_R _37475_ (.A(_08075_),
    .B(_08076_),
    .Y(_08078_));
 AO21x1_ASAP7_75t_R _37476_ (.A1(net1662),
    .A2(_05957_),
    .B(_05839_),
    .Y(_08079_));
 AND2x2_ASAP7_75t_R _37477_ (.A(_08079_),
    .B(_05847_),
    .Y(_08080_));
 AO21x1_ASAP7_75t_R _37478_ (.A1(net1787),
    .A2(_05866_),
    .B(net2679),
    .Y(_08081_));
 NAND3x1_ASAP7_75t_R _37479_ (.A(_08078_),
    .B(_08080_),
    .C(_08081_),
    .Y(_08082_));
 INVx1_ASAP7_75t_R _37480_ (.A(_08082_),
    .Y(_08083_));
 AND2x4_ASAP7_75t_R _37481_ (.A(_08074_),
    .B(_08083_),
    .Y(_08084_));
 NAND2x2_ASAP7_75t_R _37482_ (.A(_08063_),
    .B(_08084_),
    .Y(_08085_));
 NOR2x2_ASAP7_75t_R _37483_ (.A(_08048_),
    .B(_08085_),
    .Y(_08086_));
 XOR2x2_ASAP7_75t_R _37484_ (.A(_08005_),
    .B(_08086_),
    .Y(_08087_));
 XNOR2x2_ASAP7_75t_R _37485_ (.A(_07918_),
    .B(_08087_),
    .Y(_08089_));
 XOR2x2_ASAP7_75t_R _37486_ (.A(_07697_),
    .B(_05427_),
    .Y(_08090_));
 AO21x1_ASAP7_75t_R _37487_ (.A1(net2146),
    .A2(net3101),
    .B(_05256_),
    .Y(_08091_));
 NAND2x1_ASAP7_75t_R _37488_ (.A(_05181_),
    .B(net2094),
    .Y(_08092_));
 AND3x1_ASAP7_75t_R _37489_ (.A(_08091_),
    .B(_05258_),
    .C(_08092_),
    .Y(_08093_));
 AO21x1_ASAP7_75t_R _37490_ (.A1(net1867),
    .A2(net2146),
    .B(net3095),
    .Y(_08094_));
 AO21x1_ASAP7_75t_R _37491_ (.A1(net3426),
    .A2(net1877),
    .B(net3095),
    .Y(_08095_));
 NAND2x1_ASAP7_75t_R _37492_ (.A(_05106_),
    .B(_05241_),
    .Y(_08096_));
 AND3x1_ASAP7_75t_R _37493_ (.A(_08094_),
    .B(_08095_),
    .C(_08096_),
    .Y(_08097_));
 NAND2x1_ASAP7_75t_R _37494_ (.A(_08093_),
    .B(_08097_),
    .Y(_08098_));
 AO21x1_ASAP7_75t_R _37495_ (.A1(net1091),
    .A2(net1140),
    .B(_05198_),
    .Y(_08100_));
 AO21x1_ASAP7_75t_R _37496_ (.A1(net1877),
    .A2(net1793),
    .B(_05198_),
    .Y(_08101_));
 AO21x1_ASAP7_75t_R _37497_ (.A1(net964),
    .A2(_05058_),
    .B(_05198_),
    .Y(_08102_));
 AND3x1_ASAP7_75t_R _37498_ (.A(_08100_),
    .B(_08101_),
    .C(_08102_),
    .Y(_08103_));
 NAND2x1_ASAP7_75t_R _37499_ (.A(_06960_),
    .B(_05261_),
    .Y(_08104_));
 NOR2x1_ASAP7_75t_R _37500_ (.A(_08104_),
    .B(_06368_),
    .Y(_08105_));
 NAND2x1_ASAP7_75t_R _37501_ (.A(_08103_),
    .B(_08105_),
    .Y(_08106_));
 NOR2x1_ASAP7_75t_R _37502_ (.A(_08098_),
    .B(_08106_),
    .Y(_08107_));
 AO21x1_ASAP7_75t_R _37503_ (.A1(net1922),
    .A2(net1765),
    .B(_05062_),
    .Y(_08108_));
 NAND2x1_ASAP7_75t_R _37504_ (.A(_05264_),
    .B(_05063_),
    .Y(_08109_));
 AND3x2_ASAP7_75t_R _37505_ (.A(_08108_),
    .B(_08109_),
    .C(_06984_),
    .Y(_08111_));
 AOI211x1_ASAP7_75t_R _37506_ (.A1(net1324),
    .A2(net1153),
    .B(net3412),
    .C(_05090_),
    .Y(_08112_));
 NOR2x2_ASAP7_75t_R _37507_ (.A(_08112_),
    .B(_07665_),
    .Y(_08113_));
 AO21x1_ASAP7_75t_R _37508_ (.A1(net2146),
    .A2(_05265_),
    .B(_05126_),
    .Y(_08114_));
 AND2x2_ASAP7_75t_R _37509_ (.A(_08114_),
    .B(_06986_),
    .Y(_08115_));
 NAND3x2_ASAP7_75t_R _37510_ (.B(_08113_),
    .C(_08115_),
    .Y(_08116_),
    .A(_08111_));
 NAND2x1_ASAP7_75t_R _37511_ (.A(_07647_),
    .B(_05134_),
    .Y(_08117_));
 OA21x2_ASAP7_75t_R _37512_ (.A1(_05308_),
    .A2(net2161),
    .B(_05201_),
    .Y(_08118_));
 AO21x1_ASAP7_75t_R _37513_ (.A1(_05217_),
    .A2(net2783),
    .B(net2468),
    .Y(_08119_));
 AOI21x1_ASAP7_75t_R _37514_ (.A1(net2126),
    .A2(_08119_),
    .B(_05138_),
    .Y(_08120_));
 AOI211x1_ASAP7_75t_R _37515_ (.A1(net1323),
    .A2(net1152),
    .B(net1526),
    .C(_05118_),
    .Y(_08122_));
 OR4x2_ASAP7_75t_R _37516_ (.A(_08117_),
    .B(_08118_),
    .C(_08120_),
    .D(_08122_),
    .Y(_08123_));
 NOR2x2_ASAP7_75t_R _37517_ (.A(_08116_),
    .B(_08123_),
    .Y(_08124_));
 NAND2x2_ASAP7_75t_R _37518_ (.A(_08107_),
    .B(_08124_),
    .Y(_08125_));
 NAND2x1_ASAP7_75t_R _37519_ (.A(_05092_),
    .B(_05154_),
    .Y(_08126_));
 OAI21x1_ASAP7_75t_R _37520_ (.A1(net2784),
    .A2(_05319_),
    .B(_08126_),
    .Y(_08127_));
 INVx1_ASAP7_75t_R _37521_ (.A(_05321_),
    .Y(_08128_));
 AOI211x1_ASAP7_75t_R _37522_ (.A1(_05178_),
    .A2(_05154_),
    .B(_08127_),
    .C(_08128_),
    .Y(_08129_));
 AO21x1_ASAP7_75t_R _37523_ (.A1(net2149),
    .A2(net1237),
    .B(_05306_),
    .Y(_08130_));
 AO21x1_ASAP7_75t_R _37524_ (.A1(net3453),
    .A2(net990),
    .B(_05306_),
    .Y(_08131_));
 NOR2x2_ASAP7_75t_R _37525_ (.A(net2315),
    .B(_05306_),
    .Y(_08133_));
 INVx1_ASAP7_75t_R _37526_ (.A(_08133_),
    .Y(_08134_));
 NOR2x1_ASAP7_75t_R _37527_ (.A(net1822),
    .B(_05306_),
    .Y(_08135_));
 INVx1_ASAP7_75t_R _37528_ (.A(_08135_),
    .Y(_08136_));
 AND4x1_ASAP7_75t_R _37529_ (.A(_08130_),
    .B(_08131_),
    .C(_08134_),
    .D(_08136_),
    .Y(_08137_));
 NAND2x1_ASAP7_75t_R _37530_ (.A(_08129_),
    .B(_08137_),
    .Y(_08138_));
 AO21x1_ASAP7_75t_R _37531_ (.A1(net2126),
    .A2(net1867),
    .B(_05215_),
    .Y(_08139_));
 AO21x1_ASAP7_75t_R _37532_ (.A1(net3426),
    .A2(_05259_),
    .B(_05215_),
    .Y(_08140_));
 NAND2x1_ASAP7_75t_R _37533_ (.A(net2094),
    .B(_05420_),
    .Y(_08141_));
 AND3x1_ASAP7_75t_R _37534_ (.A(_08139_),
    .B(_08140_),
    .C(_08141_),
    .Y(_08142_));
 OA21x2_ASAP7_75t_R _37535_ (.A1(_05096_),
    .A2(_05092_),
    .B(_05247_),
    .Y(_08144_));
 AO21x1_ASAP7_75t_R _37536_ (.A1(_05247_),
    .A2(_06321_),
    .B(_05245_),
    .Y(_08145_));
 AOI211x1_ASAP7_75t_R _37537_ (.A1(net1489),
    .A2(_05247_),
    .B(_08144_),
    .C(_08145_),
    .Y(_08146_));
 NAND2x1_ASAP7_75t_R _37538_ (.A(_08142_),
    .B(_08146_),
    .Y(_08147_));
 NOR2x1_ASAP7_75t_R _37539_ (.A(_08138_),
    .B(_08147_),
    .Y(_08148_));
 NAND2x1_ASAP7_75t_R _37540_ (.A(_05308_),
    .B(_05171_),
    .Y(_08149_));
 NAND2x1_ASAP7_75t_R _37541_ (.A(_05264_),
    .B(_05171_),
    .Y(_08150_));
 AND3x2_ASAP7_75t_R _37542_ (.A(_05081_),
    .B(_08149_),
    .C(_08150_),
    .Y(_08151_));
 AO21x1_ASAP7_75t_R _37543_ (.A1(net1140),
    .A2(_05271_),
    .B(net2621),
    .Y(_08152_));
 AND2x2_ASAP7_75t_R _37544_ (.A(_08152_),
    .B(_06349_),
    .Y(_08153_));
 AO21x1_ASAP7_75t_R _37545_ (.A1(net1837),
    .A2(net990),
    .B(net2493),
    .Y(_08155_));
 NAND3x2_ASAP7_75t_R _37546_ (.B(_08153_),
    .C(_08155_),
    .Y(_08156_),
    .A(_08151_));
 AO21x1_ASAP7_75t_R _37547_ (.A1(net990),
    .A2(_05058_),
    .B(net2529),
    .Y(_08157_));
 NAND2x1_ASAP7_75t_R _37548_ (.A(_07614_),
    .B(_08157_),
    .Y(_08158_));
 AO21x1_ASAP7_75t_R _37549_ (.A1(_05206_),
    .A2(net1140),
    .B(net2529),
    .Y(_08159_));
 OAI21x1_ASAP7_75t_R _37550_ (.A1(net1091),
    .A2(net2529),
    .B(_08159_),
    .Y(_08160_));
 NOR2x2_ASAP7_75t_R _37551_ (.A(_08158_),
    .B(_08160_),
    .Y(_08161_));
 OA21x2_ASAP7_75t_R _37552_ (.A1(_05239_),
    .A2(_05191_),
    .B(_05087_),
    .Y(_08162_));
 AOI211x1_ASAP7_75t_R _37553_ (.A1(_05238_),
    .A2(_05087_),
    .B(_08162_),
    .C(_05207_),
    .Y(_08163_));
 AND2x2_ASAP7_75t_R _37554_ (.A(_05387_),
    .B(_05389_),
    .Y(_08164_));
 NAND3x2_ASAP7_75t_R _37555_ (.B(_08163_),
    .C(_08164_),
    .Y(_08166_),
    .A(_08161_));
 NOR2x2_ASAP7_75t_R _37556_ (.A(_08156_),
    .B(_08166_),
    .Y(_08167_));
 NAND2x2_ASAP7_75t_R _37557_ (.A(_08148_),
    .B(_08167_),
    .Y(_08168_));
 NOR2x2_ASAP7_75t_R _37558_ (.A(_08125_),
    .B(_08168_),
    .Y(_08169_));
 INVx1_ASAP7_75t_R _37559_ (.A(_08169_),
    .Y(_08170_));
 XOR2x2_ASAP7_75t_R _37560_ (.A(_08090_),
    .B(_08170_),
    .Y(_08171_));
 INVx2_ASAP7_75t_R _37561_ (.A(_08171_),
    .Y(_08172_));
 NAND2x1_ASAP7_75t_R _37562_ (.A(_08172_),
    .B(_08089_),
    .Y(_08173_));
 INVx2_ASAP7_75t_R _37563_ (.A(_08089_),
    .Y(_08174_));
 NAND2x1_ASAP7_75t_R _37564_ (.A(_08171_),
    .B(_08174_),
    .Y(_08175_));
 AOI21x1_ASAP7_75t_R _37565_ (.A1(_08173_),
    .A2(_08175_),
    .B(net388),
    .Y(_08177_));
 INVx1_ASAP7_75t_R _37566_ (.A(_00387_),
    .Y(_08178_));
 OAI21x1_ASAP7_75t_R _37567_ (.A1(_07821_),
    .A2(_08177_),
    .B(_08178_),
    .Y(_08179_));
 NOR2x1_ASAP7_75t_R _37568_ (.A(_00528_),
    .B(_00847_),
    .Y(_08180_));
 NAND2x1_ASAP7_75t_R _37569_ (.A(_08171_),
    .B(_08089_),
    .Y(_08181_));
 NAND2x1_ASAP7_75t_R _37570_ (.A(_08172_),
    .B(_08174_),
    .Y(_08182_));
 AOI21x1_ASAP7_75t_R _37571_ (.A1(_08181_),
    .A2(_08182_),
    .B(net388),
    .Y(_08183_));
 OAI21x1_ASAP7_75t_R _37572_ (.A1(_08180_),
    .A2(_08183_),
    .B(_00387_),
    .Y(_08184_));
 NAND2x1_ASAP7_75t_R _37573_ (.A(_08184_),
    .B(_08179_),
    .Y(_00109_));
 NOR2x1_ASAP7_75t_R _37574_ (.A(_00528_),
    .B(_00846_),
    .Y(_08185_));
 OAI21x1_ASAP7_75t_R _37575_ (.A1(net2786),
    .A2(_06150_),
    .B(_06252_),
    .Y(_08187_));
 AO22x1_ASAP7_75t_R _37576_ (.A1(net1094),
    .A2(_06251_),
    .B1(_06816_),
    .B2(net2507),
    .Y(_08188_));
 NOR2x1_ASAP7_75t_R _37577_ (.A(_08187_),
    .B(_08188_),
    .Y(_08189_));
 OAI21x1_ASAP7_75t_R _37578_ (.A1(net2399),
    .A2(net1628),
    .B(_07333_),
    .Y(_08190_));
 AO22x2_ASAP7_75t_R _37579_ (.A1(_06816_),
    .A2(_06188_),
    .B1(_06775_),
    .B2(_07297_),
    .Y(_08191_));
 NOR2x1_ASAP7_75t_R _37580_ (.A(_08190_),
    .B(_08191_),
    .Y(_08192_));
 NAND2x1_ASAP7_75t_R _37581_ (.A(_08189_),
    .B(_08192_),
    .Y(_08193_));
 AO22x1_ASAP7_75t_R _37582_ (.A1(_07907_),
    .A2(_06251_),
    .B1(_06245_),
    .B2(_06801_),
    .Y(_08194_));
 INVx1_ASAP7_75t_R _37583_ (.A(_06047_),
    .Y(_08195_));
 NOR2x1_ASAP7_75t_R _37584_ (.A(_06098_),
    .B(_08195_),
    .Y(_08196_));
 AO22x1_ASAP7_75t_R _37585_ (.A1(_06207_),
    .A2(_08196_),
    .B1(_06105_),
    .B2(_06213_),
    .Y(_08198_));
 NOR2x1_ASAP7_75t_R _37586_ (.A(_08194_),
    .B(_08198_),
    .Y(_08199_));
 NOR2x1_ASAP7_75t_R _37587_ (.A(_06084_),
    .B(_06210_),
    .Y(_08200_));
 NOR2x1_ASAP7_75t_R _37588_ (.A(_06182_),
    .B(_06081_),
    .Y(_08201_));
 NOR2x1_ASAP7_75t_R _37589_ (.A(_08200_),
    .B(_08201_),
    .Y(_08202_));
 NAND2x1_ASAP7_75t_R _37590_ (.A(_06193_),
    .B(_06105_),
    .Y(_08203_));
 AND3x1_ASAP7_75t_R _37591_ (.A(_08202_),
    .B(_08203_),
    .C(_07825_),
    .Y(_08204_));
 NAND2x1_ASAP7_75t_R _37592_ (.A(_08199_),
    .B(_08204_),
    .Y(_08205_));
 NOR2x2_ASAP7_75t_R _37593_ (.A(_08205_),
    .B(_08193_),
    .Y(_08206_));
 INVx1_ASAP7_75t_R _37594_ (.A(_06811_),
    .Y(_08207_));
 INVx1_ASAP7_75t_R _37595_ (.A(_07351_),
    .Y(_08209_));
 NAND2x2_ASAP7_75t_R _37596_ (.A(net1598),
    .B(_06139_),
    .Y(_08210_));
 AO21x1_ASAP7_75t_R _37597_ (.A1(_08209_),
    .A2(_08210_),
    .B(_06741_),
    .Y(_08211_));
 NAND2x1_ASAP7_75t_R _37598_ (.A(_08207_),
    .B(_08211_),
    .Y(_08212_));
 AO21x1_ASAP7_75t_R _37599_ (.A1(net2764),
    .A2(_06240_),
    .B(_06853_),
    .Y(_08213_));
 NAND2x1_ASAP7_75t_R _37600_ (.A(_07419_),
    .B(_06781_),
    .Y(_08214_));
 AND2x2_ASAP7_75t_R _37601_ (.A(_08213_),
    .B(_08214_),
    .Y(_08215_));
 NOR2x1_ASAP7_75t_R _37602_ (.A(_06219_),
    .B(_06104_),
    .Y(_08216_));
 AO21x1_ASAP7_75t_R _37603_ (.A1(_06193_),
    .A2(_06212_),
    .B(_08216_),
    .Y(_08217_));
 AO22x1_ASAP7_75t_R _37604_ (.A1(_06273_),
    .A2(_07454_),
    .B1(_06212_),
    .B2(_06259_),
    .Y(_08218_));
 NOR2x1_ASAP7_75t_R _37605_ (.A(_08217_),
    .B(_08218_),
    .Y(_08220_));
 NAND2x1_ASAP7_75t_R _37606_ (.A(_08215_),
    .B(_08220_),
    .Y(_08221_));
 NOR2x2_ASAP7_75t_R _37607_ (.A(_08212_),
    .B(_08221_),
    .Y(_08222_));
 AO21x1_ASAP7_75t_R _37608_ (.A1(_06107_),
    .A2(_07841_),
    .B(_06064_),
    .Y(_08223_));
 OA21x2_ASAP7_75t_R _37609_ (.A1(_06151_),
    .A2(_06750_),
    .B(_08223_),
    .Y(_08224_));
 NOR2x1_ASAP7_75t_R _37610_ (.A(_06268_),
    .B(_06196_),
    .Y(_08225_));
 AOI221x1_ASAP7_75t_R _37611_ (.A1(_06781_),
    .A2(_06091_),
    .B1(_06765_),
    .B2(_06783_),
    .C(_08225_),
    .Y(_08226_));
 NAND2x1_ASAP7_75t_R _37612_ (.A(_08224_),
    .B(_08226_),
    .Y(_08227_));
 NAND2x1_ASAP7_75t_R _37613_ (.A(net2084),
    .B(_06159_),
    .Y(_08228_));
 AND2x2_ASAP7_75t_R _37614_ (.A(_06884_),
    .B(_08228_),
    .Y(_08229_));
 AND3x1_ASAP7_75t_R _37615_ (.A(_07852_),
    .B(_06777_),
    .C(_07362_),
    .Y(_08231_));
 NAND2x2_ASAP7_75t_R _37616_ (.A(_08229_),
    .B(_08231_),
    .Y(_08232_));
 NOR2x2_ASAP7_75t_R _37617_ (.A(_08227_),
    .B(_08232_),
    .Y(_08233_));
 NAND3x2_ASAP7_75t_R _37618_ (.B(_08222_),
    .C(_08233_),
    .Y(_08234_),
    .A(_08206_));
 OA21x2_ASAP7_75t_R _37619_ (.A1(net1261),
    .A2(_06151_),
    .B(_06711_),
    .Y(_08235_));
 NAND2x1_ASAP7_75t_R _37620_ (.A(_07308_),
    .B(_06751_),
    .Y(_08236_));
 AO21x1_ASAP7_75t_R _37621_ (.A1(_06061_),
    .A2(_06757_),
    .B(_06745_),
    .Y(_08237_));
 NOR2x1_ASAP7_75t_R _37622_ (.A(_08236_),
    .B(_08237_),
    .Y(_08238_));
 OA21x2_ASAP7_75t_R _37623_ (.A1(net1276),
    .A2(_06785_),
    .B(_06183_),
    .Y(_08239_));
 AND3x2_ASAP7_75t_R _37624_ (.A(_08235_),
    .B(_08238_),
    .C(_08239_),
    .Y(_08240_));
 AOI22x1_ASAP7_75t_R _37625_ (.A1(_06159_),
    .A2(_07461_),
    .B1(_07455_),
    .B2(net2482),
    .Y(_08242_));
 NAND2x2_ASAP7_75t_R _37626_ (.A(_08242_),
    .B(_07430_),
    .Y(_08243_));
 OR3x2_ASAP7_75t_R _37627_ (.A(net2412),
    .B(_06096_),
    .C(_06063_),
    .Y(_08244_));
 AO21x1_ASAP7_75t_R _37628_ (.A1(_06078_),
    .A2(_06226_),
    .B(_06203_),
    .Y(_08245_));
 NAND2x2_ASAP7_75t_R _37629_ (.A(_06029_),
    .B(_07352_),
    .Y(_08246_));
 NAND3x2_ASAP7_75t_R _37630_ (.B(_08245_),
    .C(_08246_),
    .Y(_08247_),
    .A(_08244_));
 NAND2x2_ASAP7_75t_R _37631_ (.A(net1548),
    .B(_07436_),
    .Y(_08248_));
 NAND3x2_ASAP7_75t_R _37632_ (.B(_06165_),
    .C(_06849_),
    .Y(_08249_),
    .A(_08248_));
 NOR3x2_ASAP7_75t_R _37633_ (.B(_08247_),
    .C(_08249_),
    .Y(_08250_),
    .A(_08243_));
 INVx1_ASAP7_75t_R _37634_ (.A(_07861_),
    .Y(_08251_));
 OA21x2_ASAP7_75t_R _37635_ (.A1(_06268_),
    .A2(_06078_),
    .B(_08251_),
    .Y(_08253_));
 NAND2x2_ASAP7_75t_R _37636_ (.A(net3430),
    .B(_06159_),
    .Y(_08254_));
 AO21x1_ASAP7_75t_R _37637_ (.A1(_06036_),
    .A2(net3330),
    .B(_06210_),
    .Y(_08255_));
 NAND3x2_ASAP7_75t_R _37638_ (.B(_08254_),
    .C(_08255_),
    .Y(_08256_),
    .A(_08253_));
 AO21x1_ASAP7_75t_R _37639_ (.A1(_06191_),
    .A2(net2399),
    .B(net3331),
    .Y(_08257_));
 AO21x1_ASAP7_75t_R _37640_ (.A1(net3434),
    .A2(net1217),
    .B(_06121_),
    .Y(_08258_));
 AND2x2_ASAP7_75t_R _37641_ (.A(_08257_),
    .B(_08258_),
    .Y(_08259_));
 AO21x1_ASAP7_75t_R _37642_ (.A1(net1214),
    .A2(_06036_),
    .B(_06121_),
    .Y(_08260_));
 AO21x1_ASAP7_75t_R _37643_ (.A1(_06219_),
    .A2(net3331),
    .B(net2412),
    .Y(_08261_));
 NAND3x2_ASAP7_75t_R _37644_ (.B(_08260_),
    .C(_08261_),
    .Y(_08262_),
    .A(_08259_));
 NOR2x2_ASAP7_75t_R _37645_ (.A(_08256_),
    .B(_08262_),
    .Y(_08264_));
 NAND3x2_ASAP7_75t_R _37646_ (.B(_08250_),
    .C(_08264_),
    .Y(_08265_),
    .A(_08240_));
 NOR2x2_ASAP7_75t_R _37647_ (.A(_08234_),
    .B(_08265_),
    .Y(_08266_));
 NAND2x2_ASAP7_75t_R _37648_ (.A(_08169_),
    .B(_08266_),
    .Y(_08267_));
 OAI22x1_ASAP7_75t_R _37649_ (.A1(_08265_),
    .A2(_08234_),
    .B1(_08125_),
    .B2(_08168_),
    .Y(_08268_));
 OAI21x1_ASAP7_75t_R _37650_ (.A1(_05873_),
    .A2(net2083),
    .B(_05875_),
    .Y(_08269_));
 AOI211x1_ASAP7_75t_R _37651_ (.A1(net1227),
    .A2(_05755_),
    .B(net2541),
    .C(_05873_),
    .Y(_08270_));
 AOI211x1_ASAP7_75t_R _37652_ (.A1(_05764_),
    .A2(_05755_),
    .B(_05957_),
    .C(_05873_),
    .Y(_08271_));
 NOR3x2_ASAP7_75t_R _37653_ (.B(_08270_),
    .C(_08271_),
    .Y(_08272_),
    .A(_08269_));
 AO21x1_ASAP7_75t_R _37654_ (.A1(net3357),
    .A2(_05876_),
    .B(_05908_),
    .Y(_08273_));
 NAND2x1_ASAP7_75t_R _37655_ (.A(_08273_),
    .B(_07548_),
    .Y(_08275_));
 AO21x1_ASAP7_75t_R _37656_ (.A1(net1662),
    .A2(_06490_),
    .B(_05894_),
    .Y(_08276_));
 AO21x1_ASAP7_75t_R _37657_ (.A1(net2604),
    .A2(net2736),
    .B(_05894_),
    .Y(_08277_));
 NAND2x2_ASAP7_75t_R _37658_ (.A(net2483),
    .B(_05898_),
    .Y(_08278_));
 NAND3x2_ASAP7_75t_R _37659_ (.B(_08277_),
    .C(_08278_),
    .Y(_08279_),
    .A(_08276_));
 NOR2x2_ASAP7_75t_R _37660_ (.A(_08275_),
    .B(_08279_),
    .Y(_08280_));
 AO21x1_ASAP7_75t_R _37661_ (.A1(_05817_),
    .A2(_07229_),
    .B(_05884_),
    .Y(_08281_));
 AO21x1_ASAP7_75t_R _37662_ (.A1(_06490_),
    .A2(_05905_),
    .B(_05884_),
    .Y(_08282_));
 NAND2x1_ASAP7_75t_R _37663_ (.A(_06472_),
    .B(_05885_),
    .Y(_08283_));
 AND3x2_ASAP7_75t_R _37664_ (.A(_08281_),
    .B(_08282_),
    .C(_08283_),
    .Y(_08284_));
 NAND3x2_ASAP7_75t_R _37665_ (.B(_08280_),
    .C(_08284_),
    .Y(_08286_),
    .A(_08272_));
 AO21x1_ASAP7_75t_R _37666_ (.A1(net1806),
    .A2(net1807),
    .B(_05800_),
    .Y(_08287_));
 OAI21x1_ASAP7_75t_R _37667_ (.A1(net1118),
    .A2(_05800_),
    .B(_08287_),
    .Y(_08288_));
 AO21x1_ASAP7_75t_R _37668_ (.A1(net1787),
    .A2(net1560),
    .B(net3351),
    .Y(_08289_));
 AO21x1_ASAP7_75t_R _37669_ (.A1(net2098),
    .A2(net1441),
    .B(net3351),
    .Y(_08290_));
 NAND2x2_ASAP7_75t_R _37670_ (.A(_08289_),
    .B(_08290_),
    .Y(_08291_));
 AOI21x1_ASAP7_75t_R _37671_ (.A1(net1443),
    .A2(_05933_),
    .B(_05800_),
    .Y(_08292_));
 NOR3x2_ASAP7_75t_R _37672_ (.B(_08291_),
    .C(_08292_),
    .Y(_08293_),
    .A(_08288_));
 AO21x1_ASAP7_75t_R _37673_ (.A1(_05876_),
    .A2(net2081),
    .B(_05839_),
    .Y(_08294_));
 OA21x2_ASAP7_75t_R _37674_ (.A1(net3469),
    .A2(_05839_),
    .B(_08294_),
    .Y(_08295_));
 AO21x1_ASAP7_75t_R _37675_ (.A1(net2603),
    .A2(_05805_),
    .B(_05839_),
    .Y(_08297_));
 OA21x2_ASAP7_75t_R _37676_ (.A1(net1037),
    .A2(_05839_),
    .B(_08297_),
    .Y(_08298_));
 AND2x2_ASAP7_75t_R _37677_ (.A(_08295_),
    .B(_08298_),
    .Y(_08299_));
 NOR2x1_ASAP7_75t_R _37678_ (.A(_05854_),
    .B(_07229_),
    .Y(_08300_));
 AO21x1_ASAP7_75t_R _37679_ (.A1(net3348),
    .A2(_07205_),
    .B(_08300_),
    .Y(_08301_));
 AOI21x1_ASAP7_75t_R _37680_ (.A1(_05973_),
    .A2(_07205_),
    .B(_08301_),
    .Y(_08302_));
 NAND3x2_ASAP7_75t_R _37681_ (.B(_08299_),
    .C(_08302_),
    .Y(_08303_),
    .A(_08293_));
 NOR2x2_ASAP7_75t_R _37682_ (.A(_08303_),
    .B(_08286_),
    .Y(_08304_));
 NAND2x2_ASAP7_75t_R _37683_ (.A(_06517_),
    .B(_05966_),
    .Y(_08305_));
 NAND3x2_ASAP7_75t_R _37684_ (.B(_07260_),
    .C(_08305_),
    .Y(_08306_),
    .A(_07261_));
 AO21x1_ASAP7_75t_R _37685_ (.A1(net1804),
    .A2(_06490_),
    .B(_05977_),
    .Y(_08308_));
 AO21x1_ASAP7_75t_R _37686_ (.A1(_05744_),
    .A2(net2846),
    .B(_05977_),
    .Y(_08309_));
 NAND2x2_ASAP7_75t_R _37687_ (.A(_08308_),
    .B(_08309_),
    .Y(_08310_));
 NOR3x2_ASAP7_75t_R _37688_ (.B(_08310_),
    .C(_05974_),
    .Y(_08311_),
    .A(_08306_));
 INVx1_ASAP7_75t_R _37689_ (.A(_08042_),
    .Y(_08312_));
 NAND2x1_ASAP7_75t_R _37690_ (.A(_06017_),
    .B(_07213_),
    .Y(_08313_));
 AND4x2_ASAP7_75t_R _37691_ (.A(_06536_),
    .B(_07534_),
    .C(_08312_),
    .D(_08313_),
    .Y(_08314_));
 AO21x1_ASAP7_75t_R _37692_ (.A1(_05833_),
    .A2(_05918_),
    .B(_05993_),
    .Y(_08315_));
 AO21x1_ASAP7_75t_R _37693_ (.A1(net1787),
    .A2(net1560),
    .B(_05993_),
    .Y(_08316_));
 AND3x2_ASAP7_75t_R _37694_ (.A(_08315_),
    .B(_05997_),
    .C(_08316_),
    .Y(_08317_));
 NAND3x2_ASAP7_75t_R _37695_ (.B(_08314_),
    .C(_08317_),
    .Y(_08319_),
    .A(_08311_));
 OR3x1_ASAP7_75t_R _37696_ (.A(_05938_),
    .B(net1880),
    .C(net2761),
    .Y(_08320_));
 NAND2x2_ASAP7_75t_R _37697_ (.A(_06510_),
    .B(_08320_),
    .Y(_08321_));
 AO21x1_ASAP7_75t_R _37698_ (.A1(_05879_),
    .A2(net3375),
    .B(net2521),
    .Y(_08322_));
 OAI21x1_ASAP7_75t_R _37699_ (.A1(_05775_),
    .A2(net2521),
    .B(_08322_),
    .Y(_08323_));
 AO21x1_ASAP7_75t_R _37700_ (.A1(net1560),
    .A2(_05957_),
    .B(net3352),
    .Y(_08324_));
 OAI21x1_ASAP7_75t_R _37701_ (.A1(_05817_),
    .A2(net3352),
    .B(_08324_),
    .Y(_08325_));
 NOR3x2_ASAP7_75t_R _37702_ (.B(_08323_),
    .C(_08325_),
    .Y(_08326_),
    .A(_08321_));
 OAI21x1_ASAP7_75t_R _37703_ (.A1(net1804),
    .A2(_05787_),
    .B(_06495_),
    .Y(_08327_));
 AO21x2_ASAP7_75t_R _37704_ (.A1(_05850_),
    .A2(_05747_),
    .B(_05787_),
    .Y(_08328_));
 NAND2x2_ASAP7_75t_R _37705_ (.A(_08021_),
    .B(_08328_),
    .Y(_08330_));
 OA21x2_ASAP7_75t_R _37706_ (.A1(_06521_),
    .A2(_06015_),
    .B(_05926_),
    .Y(_08331_));
 NOR3x2_ASAP7_75t_R _37707_ (.B(_08330_),
    .C(_08331_),
    .Y(_08332_),
    .A(_08327_));
 AOI221x1_ASAP7_75t_R _37708_ (.A1(net1229),
    .A2(_05755_),
    .B1(_05775_),
    .B2(_05957_),
    .C(_05752_),
    .Y(_08333_));
 AOI211x1_ASAP7_75t_R _37709_ (.A1(_05743_),
    .A2(_05751_),
    .B(_08333_),
    .C(_05761_),
    .Y(_08334_));
 NAND3x2_ASAP7_75t_R _37710_ (.B(_08332_),
    .C(_08334_),
    .Y(_08335_),
    .A(_08326_));
 NOR2x2_ASAP7_75t_R _37711_ (.A(_08319_),
    .B(_08335_),
    .Y(_08336_));
 NAND2x2_ASAP7_75t_R _37712_ (.A(_08304_),
    .B(_08336_),
    .Y(_08337_));
 NOR2x2_ASAP7_75t_R _37713_ (.A(_06425_),
    .B(_08337_),
    .Y(_08338_));
 NAND3x2_ASAP7_75t_R _37714_ (.B(_08268_),
    .C(net2774),
    .Y(_08339_),
    .A(_08267_));
 AO21x1_ASAP7_75t_R _37715_ (.A1(_08267_),
    .A2(_08268_),
    .B(net2774),
    .Y(_08341_));
 AO21x1_ASAP7_75t_R _37716_ (.A1(net2003),
    .A2(net2663),
    .B(net2410),
    .Y(_08342_));
 OAI21x1_ASAP7_75t_R _37717_ (.A1(net1086),
    .A2(net2410),
    .B(_08342_),
    .Y(_08343_));
 AO21x1_ASAP7_75t_R _37718_ (.A1(net1902),
    .A2(net2153),
    .B(net2410),
    .Y(_08344_));
 OAI21x1_ASAP7_75t_R _37719_ (.A1(net1211),
    .A2(net2410),
    .B(_08344_),
    .Y(_08345_));
 NOR2x1_ASAP7_75t_R _37720_ (.A(_08343_),
    .B(_08345_),
    .Y(_08346_));
 NOR2x2_ASAP7_75t_R _37721_ (.A(net2548),
    .B(_05616_),
    .Y(_08347_));
 AO21x1_ASAP7_75t_R _37722_ (.A1(_06671_),
    .A2(_06613_),
    .B(_08347_),
    .Y(_08348_));
 NAND3x1_ASAP7_75t_R _37723_ (.A(_07972_),
    .B(_07973_),
    .C(_07132_),
    .Y(_08349_));
 NOR2x1_ASAP7_75t_R _37724_ (.A(_08348_),
    .B(_08349_),
    .Y(_08350_));
 NAND2x2_ASAP7_75t_R _37725_ (.A(_08346_),
    .B(_08350_),
    .Y(_08352_));
 AO21x1_ASAP7_75t_R _37726_ (.A1(_06568_),
    .A2(_05503_),
    .B(_05634_),
    .Y(_08353_));
 OAI21x1_ASAP7_75t_R _37727_ (.A1(_05634_),
    .A2(net3349),
    .B(_08353_),
    .Y(_08354_));
 AO21x1_ASAP7_75t_R _37728_ (.A1(net2032),
    .A2(net3461),
    .B(_05640_),
    .Y(_08355_));
 AO21x1_ASAP7_75t_R _37729_ (.A1(net2658),
    .A2(_05496_),
    .B(_05640_),
    .Y(_08356_));
 NAND2x1_ASAP7_75t_R _37730_ (.A(_08355_),
    .B(_08356_),
    .Y(_08357_));
 AOI21x1_ASAP7_75t_R _37731_ (.A1(_07919_),
    .A2(net1083),
    .B(_05634_),
    .Y(_08358_));
 OR3x1_ASAP7_75t_R _37732_ (.A(_08354_),
    .B(_08357_),
    .C(_08358_),
    .Y(_08359_));
 NOR2x2_ASAP7_75t_R _37733_ (.A(_08352_),
    .B(_08359_),
    .Y(_08360_));
 OA21x2_ASAP7_75t_R _37734_ (.A1(_06592_),
    .A2(net2834),
    .B(_05657_),
    .Y(_08361_));
 NOR2x1_ASAP7_75t_R _37735_ (.A(_07772_),
    .B(_08361_),
    .Y(_08363_));
 AO21x1_ASAP7_75t_R _37736_ (.A1(net2191),
    .A2(_05605_),
    .B(_06576_),
    .Y(_08364_));
 AO21x1_ASAP7_75t_R _37737_ (.A1(net2567),
    .A2(net2477),
    .B(_06576_),
    .Y(_08365_));
 NAND2x1_ASAP7_75t_R _37738_ (.A(_05661_),
    .B(_07152_),
    .Y(_08366_));
 AND3x1_ASAP7_75t_R _37739_ (.A(_08364_),
    .B(_08365_),
    .C(_08366_),
    .Y(_08367_));
 NAND2x1_ASAP7_75t_R _37740_ (.A(_08363_),
    .B(_08367_),
    .Y(_08368_));
 AOI211x1_ASAP7_75t_R _37741_ (.A1(net2814),
    .A2(net3098),
    .B(_05677_),
    .C(net1205),
    .Y(_08369_));
 AND3x1_ASAP7_75t_R _37742_ (.A(_05675_),
    .B(_05439_),
    .C(net2814),
    .Y(_08370_));
 AOI211x1_ASAP7_75t_R _37743_ (.A1(_05675_),
    .A2(net1528),
    .B(_08369_),
    .C(_08370_),
    .Y(_08371_));
 AOI211x1_ASAP7_75t_R _37744_ (.A1(net1000),
    .A2(net3098),
    .B(_05683_),
    .C(_05440_),
    .Y(_08372_));
 INVx1_ASAP7_75t_R _37745_ (.A(_08372_),
    .Y(_08374_));
 AO21x1_ASAP7_75t_R _37746_ (.A1(_05685_),
    .A2(_05503_),
    .B(_05683_),
    .Y(_08375_));
 OAI21x1_ASAP7_75t_R _37747_ (.A1(_05516_),
    .A2(_05522_),
    .B(_05684_),
    .Y(_08376_));
 AND3x1_ASAP7_75t_R _37748_ (.A(_08374_),
    .B(_08375_),
    .C(_08376_),
    .Y(_08377_));
 NAND2x1_ASAP7_75t_R _37749_ (.A(_08371_),
    .B(_08377_),
    .Y(_08378_));
 NOR2x1_ASAP7_75t_R _37750_ (.A(_08368_),
    .B(_08378_),
    .Y(_08379_));
 NAND2x2_ASAP7_75t_R _37751_ (.A(_08360_),
    .B(_08379_),
    .Y(_08380_));
 OA211x2_ASAP7_75t_R _37752_ (.A1(net2712),
    .A2(net989),
    .B(_05577_),
    .C(_05439_),
    .Y(_08381_));
 AO21x1_ASAP7_75t_R _37753_ (.A1(_05496_),
    .A2(net2509),
    .B(_05581_),
    .Y(_08382_));
 NAND2x1_ASAP7_75t_R _37754_ (.A(_08382_),
    .B(_06666_),
    .Y(_08383_));
 AO21x1_ASAP7_75t_R _37755_ (.A1(_05490_),
    .A2(_05457_),
    .B(net2389),
    .Y(_08385_));
 OAI21x1_ASAP7_75t_R _37756_ (.A1(net2389),
    .A2(_05613_),
    .B(_08385_),
    .Y(_08386_));
 OR3x1_ASAP7_75t_R _37757_ (.A(_08381_),
    .B(_08383_),
    .C(_08386_),
    .Y(_08387_));
 AOI221x1_ASAP7_75t_R _37758_ (.A1(net1000),
    .A2(net3098),
    .B1(_05440_),
    .B2(_05457_),
    .C(_05453_),
    .Y(_08388_));
 OAI21x1_ASAP7_75t_R _37759_ (.A1(net2864),
    .A2(_05467_),
    .B(_05465_),
    .Y(_08389_));
 NOR2x1_ASAP7_75t_R _37760_ (.A(_08388_),
    .B(_08389_),
    .Y(_08390_));
 AO21x1_ASAP7_75t_R _37761_ (.A1(net2657),
    .A2(_05605_),
    .B(_05472_),
    .Y(_08391_));
 AO21x1_ASAP7_75t_R _37762_ (.A1(net2032),
    .A2(net2610),
    .B(_05472_),
    .Y(_08392_));
 AND2x2_ASAP7_75t_R _37763_ (.A(_08391_),
    .B(_08392_),
    .Y(_08393_));
 OA21x2_ASAP7_75t_R _37764_ (.A1(_05601_),
    .A2(_07760_),
    .B(_07922_),
    .Y(_08394_));
 AND2x2_ASAP7_75t_R _37765_ (.A(_08393_),
    .B(_08394_),
    .Y(_08396_));
 NAND2x1_ASAP7_75t_R _37766_ (.A(_08390_),
    .B(_08396_),
    .Y(_08397_));
 NOR2x1_ASAP7_75t_R _37767_ (.A(_08387_),
    .B(_08397_),
    .Y(_08398_));
 OA21x2_ASAP7_75t_R _37768_ (.A1(_06637_),
    .A2(_07066_),
    .B(net3373),
    .Y(_08399_));
 NAND2x1_ASAP7_75t_R _37769_ (.A(_05518_),
    .B(_05523_),
    .Y(_08400_));
 AOI211x1_ASAP7_75t_R _37770_ (.A1(net3373),
    .A2(_05566_),
    .B(_08399_),
    .C(_08400_),
    .Y(_08401_));
 AOI211x1_ASAP7_75t_R _37771_ (.A1(net2814),
    .A2(net3098),
    .B(_05492_),
    .C(net1669),
    .Y(_08402_));
 INVx1_ASAP7_75t_R _37772_ (.A(_08402_),
    .Y(_08403_));
 AO21x1_ASAP7_75t_R _37773_ (.A1(net2663),
    .A2(_05605_),
    .B(_05492_),
    .Y(_08404_));
 AND3x1_ASAP7_75t_R _37774_ (.A(_08403_),
    .B(_07719_),
    .C(_08404_),
    .Y(_08405_));
 NAND2x1_ASAP7_75t_R _37775_ (.A(_08401_),
    .B(_08405_),
    .Y(_08407_));
 NAND2x1_ASAP7_75t_R _37776_ (.A(_05656_),
    .B(_06627_),
    .Y(_08408_));
 NAND2x2_ASAP7_75t_R _37777_ (.A(_08408_),
    .B(_07952_),
    .Y(_08409_));
 OA21x2_ASAP7_75t_R _37778_ (.A1(net3106),
    .A2(_05516_),
    .B(_06627_),
    .Y(_08410_));
 OA21x2_ASAP7_75t_R _37779_ (.A1(_06671_),
    .A2(_05520_),
    .B(_06627_),
    .Y(_08411_));
 NOR3x2_ASAP7_75t_R _37780_ (.B(_08410_),
    .C(_08411_),
    .Y(_08412_),
    .A(_08409_));
 NAND2x1_ASAP7_75t_R _37781_ (.A(_07941_),
    .B(_07738_),
    .Y(_08413_));
 AO21x1_ASAP7_75t_R _37782_ (.A1(_05646_),
    .A2(_05545_),
    .B(_07733_),
    .Y(_08414_));
 NOR2x1_ASAP7_75t_R _37783_ (.A(_08413_),
    .B(_08414_),
    .Y(_08415_));
 NAND2x2_ASAP7_75t_R _37784_ (.A(_08412_),
    .B(_08415_),
    .Y(_08416_));
 NOR2x2_ASAP7_75t_R _37785_ (.A(_08407_),
    .B(_08416_),
    .Y(_08418_));
 NAND2x2_ASAP7_75t_R _37786_ (.A(_08398_),
    .B(_08418_),
    .Y(_08419_));
 AOI211x1_ASAP7_75t_R _37787_ (.A1(_05478_),
    .A2(net2111),
    .B(_08380_),
    .C(_08419_),
    .Y(_08420_));
 AO21x1_ASAP7_75t_R _37788_ (.A1(net2137),
    .A2(net1836),
    .B(_05240_),
    .Y(_08421_));
 AO21x1_ASAP7_75t_R _37789_ (.A1(net1944),
    .A2(_05058_),
    .B(_05240_),
    .Y(_08422_));
 NAND2x1_ASAP7_75t_R _37790_ (.A(net2161),
    .B(_05241_),
    .Y(_08423_));
 AND4x2_ASAP7_75t_R _37791_ (.A(_05254_),
    .B(_08421_),
    .C(_08422_),
    .D(_08423_),
    .Y(_08424_));
 AO21x1_ASAP7_75t_R _37792_ (.A1(_05206_),
    .A2(net2149),
    .B(_05198_),
    .Y(_08425_));
 NAND2x1_ASAP7_75t_R _37793_ (.A(_08425_),
    .B(_05338_),
    .Y(_08426_));
 AO21x1_ASAP7_75t_R _37794_ (.A1(net2056),
    .A2(net1836),
    .B(_05208_),
    .Y(_08427_));
 AO21x1_ASAP7_75t_R _37795_ (.A1(_05185_),
    .A2(net2643),
    .B(_05208_),
    .Y(_08429_));
 NAND2x2_ASAP7_75t_R _37796_ (.A(_05203_),
    .B(_05332_),
    .Y(_08430_));
 NAND3x2_ASAP7_75t_R _37797_ (.B(_08429_),
    .C(_08430_),
    .Y(_08431_),
    .A(_08427_));
 NOR2x2_ASAP7_75t_R _37798_ (.A(_08426_),
    .B(_08431_),
    .Y(_08432_));
 OA21x2_ASAP7_75t_R _37799_ (.A1(_05200_),
    .A2(_05264_),
    .B(_05181_),
    .Y(_08433_));
 AND3x1_ASAP7_75t_R _37800_ (.A(_05181_),
    .B(_05065_),
    .C(net3436),
    .Y(_08434_));
 AOI211x1_ASAP7_75t_R _37801_ (.A1(_05181_),
    .A2(net3409),
    .B(_08433_),
    .C(_08434_),
    .Y(_08435_));
 NAND3x2_ASAP7_75t_R _37802_ (.B(_08432_),
    .C(_08435_),
    .Y(_08436_),
    .A(_08424_));
 AO21x1_ASAP7_75t_R _37803_ (.A1(net3369),
    .A2(net1091),
    .B(_05062_),
    .Y(_08437_));
 AO21x1_ASAP7_75t_R _37804_ (.A1(_05211_),
    .A2(net1877),
    .B(_05062_),
    .Y(_08438_));
 NAND2x1_ASAP7_75t_R _37805_ (.A(_05106_),
    .B(_05063_),
    .Y(_08440_));
 NAND2x1_ASAP7_75t_R _37806_ (.A(_05162_),
    .B(_05063_),
    .Y(_08441_));
 AND4x2_ASAP7_75t_R _37807_ (.A(_08437_),
    .B(_08438_),
    .C(_08440_),
    .D(_08441_),
    .Y(_08442_));
 AO21x1_ASAP7_75t_R _37808_ (.A1(net2027),
    .A2(net1945),
    .B(net3444),
    .Y(_08443_));
 AO21x1_ASAP7_75t_R _37809_ (.A1(net1922),
    .A2(_05265_),
    .B(net3444),
    .Y(_08444_));
 NAND2x1_ASAP7_75t_R _37810_ (.A(_08443_),
    .B(_08444_),
    .Y(_08445_));
 AO21x1_ASAP7_75t_R _37811_ (.A1(net1877),
    .A2(_05112_),
    .B(_05138_),
    .Y(_08446_));
 AO21x1_ASAP7_75t_R _37812_ (.A1(_05119_),
    .A2(net1894),
    .B(_05138_),
    .Y(_08447_));
 INVx1_ASAP7_75t_R _37813_ (.A(_05226_),
    .Y(_08448_));
 NAND3x2_ASAP7_75t_R _37814_ (.B(_08447_),
    .C(_08448_),
    .Y(_08449_),
    .A(_08446_));
 NOR2x2_ASAP7_75t_R _37815_ (.A(_08445_),
    .B(_08449_),
    .Y(_08451_));
 OA211x2_ASAP7_75t_R _37816_ (.A1(net1323),
    .A2(net3442),
    .B(_05127_),
    .C(net2223),
    .Y(_08452_));
 NAND2x2_ASAP7_75t_R _37817_ (.A(_05264_),
    .B(_05127_),
    .Y(_08453_));
 NAND3x2_ASAP7_75t_R _37818_ (.B(_06986_),
    .C(_08453_),
    .Y(_08454_),
    .A(_06991_));
 NOR2x2_ASAP7_75t_R _37819_ (.A(_08452_),
    .B(_08454_),
    .Y(_08455_));
 NAND3x2_ASAP7_75t_R _37820_ (.B(_08451_),
    .C(_08455_),
    .Y(_08456_),
    .A(_08442_));
 NOR2x2_ASAP7_75t_R _37821_ (.A(_08436_),
    .B(_08456_),
    .Y(_08457_));
 AO21x1_ASAP7_75t_R _37822_ (.A1(net1403),
    .A2(net2645),
    .B(net3455),
    .Y(_08458_));
 NAND2x1_ASAP7_75t_R _37823_ (.A(_07614_),
    .B(_08458_),
    .Y(_08459_));
 NOR2x1_ASAP7_75t_R _37824_ (.A(net1767),
    .B(net3455),
    .Y(_08460_));
 AO21x1_ASAP7_75t_R _37825_ (.A1(_06328_),
    .A2(_05089_),
    .B(_08460_),
    .Y(_08462_));
 NOR2x1_ASAP7_75t_R _37826_ (.A(_08459_),
    .B(_08462_),
    .Y(_08463_));
 INVx1_ASAP7_75t_R _37827_ (.A(_08463_),
    .Y(_08464_));
 AO21x1_ASAP7_75t_R _37828_ (.A1(_05360_),
    .A2(_05095_),
    .B(net3103),
    .Y(_08465_));
 AO21x1_ASAP7_75t_R _37829_ (.A1(net1402),
    .A2(net1945),
    .B(net3103),
    .Y(_08466_));
 AND2x2_ASAP7_75t_R _37830_ (.A(_08466_),
    .B(_08465_),
    .Y(_08467_));
 AOI21x1_ASAP7_75t_R _37831_ (.A1(_05218_),
    .A2(_05087_),
    .B(_08162_),
    .Y(_08468_));
 NAND2x2_ASAP7_75t_R _37832_ (.A(_08468_),
    .B(_08467_),
    .Y(_08469_));
 NOR2x2_ASAP7_75t_R _37833_ (.A(_08464_),
    .B(_08469_),
    .Y(_08470_));
 AO21x1_ASAP7_75t_R _37834_ (.A1(_05211_),
    .A2(net1836),
    .B(net3107),
    .Y(_08471_));
 INVx1_ASAP7_75t_R _37835_ (.A(_08471_),
    .Y(_08473_));
 AOI211x1_ASAP7_75t_R _37836_ (.A1(net3439),
    .A2(_05068_),
    .B(net2273),
    .C(net3107),
    .Y(_08474_));
 NOR3x2_ASAP7_75t_R _37837_ (.B(_08474_),
    .C(_07600_),
    .Y(_08475_),
    .A(_08473_));
 NAND2x1_ASAP7_75t_R _37838_ (.A(_05239_),
    .B(_05108_),
    .Y(_08476_));
 NAND2x1_ASAP7_75t_R _37839_ (.A(_05308_),
    .B(_05108_),
    .Y(_08477_));
 NAND2x1_ASAP7_75t_R _37840_ (.A(_05200_),
    .B(_05108_),
    .Y(_08478_));
 NAND3x1_ASAP7_75t_R _37841_ (.A(_08476_),
    .B(_08477_),
    .C(_08478_),
    .Y(_08479_));
 NOR2x1_ASAP7_75t_R _37842_ (.A(_05115_),
    .B(_08479_),
    .Y(_08480_));
 NAND2x2_ASAP7_75t_R _37843_ (.A(_08475_),
    .B(_08480_),
    .Y(_08481_));
 INVx1_ASAP7_75t_R _37844_ (.A(_08481_),
    .Y(_08482_));
 NAND2x1_ASAP7_75t_R _37845_ (.A(_08482_),
    .B(_08470_),
    .Y(_08484_));
 AO21x1_ASAP7_75t_R _37846_ (.A1(net2027),
    .A2(_05345_),
    .B(_05215_),
    .Y(_08485_));
 OAI21x1_ASAP7_75t_R _37847_ (.A1(net2146),
    .A2(_05215_),
    .B(_08485_),
    .Y(_08486_));
 AO21x1_ASAP7_75t_R _37848_ (.A1(net3452),
    .A2(net990),
    .B(_05186_),
    .Y(_08487_));
 NAND2x1_ASAP7_75t_R _37849_ (.A(net2224),
    .B(_05247_),
    .Y(_08488_));
 OAI21x1_ASAP7_75t_R _37850_ (.A1(_06321_),
    .A2(_06956_),
    .B(_05247_),
    .Y(_08489_));
 NAND3x1_ASAP7_75t_R _37851_ (.A(_08487_),
    .B(_08488_),
    .C(_08489_),
    .Y(_08490_));
 NOR2x1_ASAP7_75t_R _37852_ (.A(_08486_),
    .B(_08490_),
    .Y(_08491_));
 NOR2x1_ASAP7_75t_R _37853_ (.A(_06312_),
    .B(_08128_),
    .Y(_08492_));
 AO221x1_ASAP7_75t_R _37854_ (.A1(net1321),
    .A2(net3442),
    .B1(_05345_),
    .B2(_05090_),
    .C(_05153_),
    .Y(_08493_));
 NAND2x1_ASAP7_75t_R _37855_ (.A(_08492_),
    .B(_08493_),
    .Y(_08495_));
 NOR2x2_ASAP7_75t_R _37856_ (.A(_08133_),
    .B(_05411_),
    .Y(_08496_));
 AO21x1_ASAP7_75t_R _37857_ (.A1(_05211_),
    .A2(net1835),
    .B(_05306_),
    .Y(_08497_));
 AO21x1_ASAP7_75t_R _37858_ (.A1(net992),
    .A2(net1946),
    .B(_05306_),
    .Y(_08498_));
 NAND3x2_ASAP7_75t_R _37859_ (.B(_08497_),
    .C(_08498_),
    .Y(_08499_),
    .A(_08496_));
 NOR2x1_ASAP7_75t_R _37860_ (.A(_08495_),
    .B(_08499_),
    .Y(_08500_));
 NAND2x1_ASAP7_75t_R _37861_ (.A(_08491_),
    .B(_08500_),
    .Y(_08501_));
 NOR2x1_ASAP7_75t_R _37862_ (.A(_08501_),
    .B(_08484_),
    .Y(_08502_));
 NAND2x2_ASAP7_75t_R _37863_ (.A(_08457_),
    .B(_08502_),
    .Y(_08503_));
 NOR2x2_ASAP7_75t_R _37864_ (.A(_05717_),
    .B(_08503_),
    .Y(_08504_));
 NOR2x2_ASAP7_75t_R _37865_ (.A(net1860),
    .B(_08504_),
    .Y(_08506_));
 NOR2x2_ASAP7_75t_R _37866_ (.A(_08380_),
    .B(_08419_),
    .Y(_08507_));
 NAND2x2_ASAP7_75t_R _37867_ (.A(_05479_),
    .B(_08507_),
    .Y(_08508_));
 INVx1_ASAP7_75t_R _37868_ (.A(_08491_),
    .Y(_08509_));
 NOR3x1_ASAP7_75t_R _37869_ (.A(_08509_),
    .B(_08499_),
    .C(_08495_),
    .Y(_08510_));
 INVx1_ASAP7_75t_R _37870_ (.A(_08470_),
    .Y(_08511_));
 NOR2x1_ASAP7_75t_R _37871_ (.A(_08481_),
    .B(_08511_),
    .Y(_08512_));
 NAND2x1_ASAP7_75t_R _37872_ (.A(_08510_),
    .B(_08512_),
    .Y(_08513_));
 INVx1_ASAP7_75t_R _37873_ (.A(_08457_),
    .Y(_08514_));
 NOR2x1_ASAP7_75t_R _37874_ (.A(_08513_),
    .B(_08514_),
    .Y(_08515_));
 NAND2x2_ASAP7_75t_R _37875_ (.A(_05329_),
    .B(_08515_),
    .Y(_08517_));
 NOR2x2_ASAP7_75t_R _37876_ (.A(_08508_),
    .B(_08517_),
    .Y(_08518_));
 NOR2x2_ASAP7_75t_R _37877_ (.A(_08518_),
    .B(_08506_),
    .Y(_08519_));
 AO21x1_ASAP7_75t_R _37878_ (.A1(_08339_),
    .A2(_08341_),
    .B(_08519_),
    .Y(_08520_));
 NAND3x1_ASAP7_75t_R _37879_ (.A(_08519_),
    .B(_08339_),
    .C(_08341_),
    .Y(_08521_));
 AOI21x1_ASAP7_75t_R _37880_ (.A1(_08520_),
    .A2(_08521_),
    .B(net388),
    .Y(_08522_));
 NOR2x1_ASAP7_75t_R _37881_ (.A(_08185_),
    .B(_08522_),
    .Y(_08523_));
 XOR2x1_ASAP7_75t_R _37882_ (.A(_08523_),
    .Y(_00110_),
    .B(_00498_));
 NOR2x2_ASAP7_75t_R _37883_ (.A(net394),
    .B(_00845_),
    .Y(_08524_));
 NOR2x1_ASAP7_75t_R _37884_ (.A(_06061_),
    .B(net1591),
    .Y(_08525_));
 INVx1_ASAP7_75t_R _37885_ (.A(_08525_),
    .Y(_08527_));
 AO21x1_ASAP7_75t_R _37886_ (.A1(_08527_),
    .A2(net3231),
    .B(_06240_),
    .Y(_08528_));
 AO21x1_ASAP7_75t_R _37887_ (.A1(_06099_),
    .A2(_06052_),
    .B(_06240_),
    .Y(_08529_));
 NAND2x1_ASAP7_75t_R _37888_ (.A(_08528_),
    .B(_08529_),
    .Y(_08530_));
 OA21x2_ASAP7_75t_R _37889_ (.A1(_06109_),
    .A2(net3432),
    .B(_06775_),
    .Y(_08531_));
 OA21x2_ASAP7_75t_R _37890_ (.A1(net2744),
    .A2(_06799_),
    .B(_06775_),
    .Y(_08532_));
 OR3x1_ASAP7_75t_R _37891_ (.A(_08531_),
    .B(_08532_),
    .C(_06235_),
    .Y(_08533_));
 NOR2x1_ASAP7_75t_R _37892_ (.A(_08530_),
    .B(_08533_),
    .Y(_08534_));
 OA21x2_ASAP7_75t_R _37893_ (.A1(_06250_),
    .A2(net3330),
    .B(_06253_),
    .Y(_08535_));
 AO21x1_ASAP7_75t_R _37894_ (.A1(net1260),
    .A2(_06219_),
    .B(_06268_),
    .Y(_08536_));
 AO21x1_ASAP7_75t_R _37895_ (.A1(net2639),
    .A2(_06118_),
    .B(_06268_),
    .Y(_08538_));
 AND2x2_ASAP7_75t_R _37896_ (.A(_08536_),
    .B(_08538_),
    .Y(_08539_));
 AO31x2_ASAP7_75t_R _37897_ (.A1(_06078_),
    .A2(_06070_),
    .A3(net2234),
    .B(_06250_),
    .Y(_08540_));
 AND3x1_ASAP7_75t_R _37898_ (.A(_08535_),
    .B(_08539_),
    .C(_08540_),
    .Y(_08541_));
 NAND2x2_ASAP7_75t_R _37899_ (.A(_08534_),
    .B(_08541_),
    .Y(_08542_));
 AO21x1_ASAP7_75t_R _37900_ (.A1(_06190_),
    .A2(_06078_),
    .B(_06203_),
    .Y(_08543_));
 NAND2x1_ASAP7_75t_R _37901_ (.A(_06088_),
    .B(_06207_),
    .Y(_08544_));
 NAND2x1_ASAP7_75t_R _37902_ (.A(_06259_),
    .B(_06207_),
    .Y(_08545_));
 NAND2x1_ASAP7_75t_R _37903_ (.A(_06799_),
    .B(_06207_),
    .Y(_08546_));
 AND4x2_ASAP7_75t_R _37904_ (.A(_08543_),
    .B(_08544_),
    .C(_08545_),
    .D(_08546_),
    .Y(_08547_));
 AO21x1_ASAP7_75t_R _37905_ (.A1(_06036_),
    .A2(_06089_),
    .B(_06191_),
    .Y(_08549_));
 AO21x1_ASAP7_75t_R _37906_ (.A1(net3328),
    .A2(net1217),
    .B(_06191_),
    .Y(_08550_));
 NAND2x2_ASAP7_75t_R _37907_ (.A(_07461_),
    .B(_06194_),
    .Y(_08551_));
 NAND3x2_ASAP7_75t_R _37908_ (.B(_08550_),
    .C(_08551_),
    .Y(_08552_),
    .A(_08549_));
 NAND2x2_ASAP7_75t_R _37909_ (.A(net2857),
    .B(_06781_),
    .Y(_08553_));
 NAND3x2_ASAP7_75t_R _37910_ (.B(_07312_),
    .C(_08553_),
    .Y(_08554_),
    .A(_06179_));
 NOR2x2_ASAP7_75t_R _37911_ (.A(_08552_),
    .B(_08554_),
    .Y(_08555_));
 AOI211x1_ASAP7_75t_R _37912_ (.A1(net1276),
    .A2(_06061_),
    .B(net3235),
    .C(net3433),
    .Y(_08556_));
 INVx1_ASAP7_75t_R _37913_ (.A(_08556_),
    .Y(_08557_));
 AO21x1_ASAP7_75t_R _37914_ (.A1(_06863_),
    .A2(net2234),
    .B(net3235),
    .Y(_08558_));
 AO21x1_ASAP7_75t_R _37915_ (.A1(net2639),
    .A2(_06150_),
    .B(net3235),
    .Y(_08560_));
 AND3x2_ASAP7_75t_R _37916_ (.A(_08557_),
    .B(_08558_),
    .C(_08560_),
    .Y(_08561_));
 NAND3x2_ASAP7_75t_R _37917_ (.B(_08555_),
    .C(_08561_),
    .Y(_08562_),
    .A(_08547_));
 NOR2x2_ASAP7_75t_R _37918_ (.A(_08542_),
    .B(_08562_),
    .Y(_08563_));
 AO221x1_ASAP7_75t_R _37919_ (.A1(net1276),
    .A2(_06061_),
    .B1(net3329),
    .B2(net3433),
    .C(_06151_),
    .Y(_08564_));
 OA21x2_ASAP7_75t_R _37920_ (.A1(_06151_),
    .A2(_07345_),
    .B(_06884_),
    .Y(_08565_));
 AND2x2_ASAP7_75t_R _37921_ (.A(_08564_),
    .B(_08565_),
    .Y(_08566_));
 AO21x1_ASAP7_75t_R _37922_ (.A1(_06118_),
    .A2(net3329),
    .B(_06121_),
    .Y(_08567_));
 OAI21x1_ASAP7_75t_R _37923_ (.A1(_06121_),
    .A2(_06226_),
    .B(_08567_),
    .Y(_08568_));
 AO21x1_ASAP7_75t_R _37924_ (.A1(_07345_),
    .A2(_06841_),
    .B(_06710_),
    .Y(_08569_));
 AO21x1_ASAP7_75t_R _37925_ (.A1(net3328),
    .A2(net2639),
    .B(_06710_),
    .Y(_08571_));
 NAND3x2_ASAP7_75t_R _37926_ (.B(_08571_),
    .C(_08210_),
    .Y(_08572_),
    .A(_08569_));
 NOR2x2_ASAP7_75t_R _37927_ (.A(_08568_),
    .B(_08572_),
    .Y(_08573_));
 INVx1_ASAP7_75t_R _37928_ (.A(_06165_),
    .Y(_08574_));
 NOR2x1_ASAP7_75t_R _37929_ (.A(_07480_),
    .B(_08574_),
    .Y(_08575_));
 AOI211x1_ASAP7_75t_R _37930_ (.A1(net1276),
    .A2(_06061_),
    .B(net2346),
    .C(net1591),
    .Y(_08576_));
 OA21x2_ASAP7_75t_R _37931_ (.A1(net2813),
    .A2(net2084),
    .B(_06159_),
    .Y(_08577_));
 NOR2x1_ASAP7_75t_R _37932_ (.A(_08576_),
    .B(_08577_),
    .Y(_08578_));
 AND2x2_ASAP7_75t_R _37933_ (.A(_08575_),
    .B(_08578_),
    .Y(_08579_));
 NAND3x2_ASAP7_75t_R _37934_ (.B(_08573_),
    .C(_08579_),
    .Y(_08580_),
    .A(_08566_));
 AO21x1_ASAP7_75t_R _37935_ (.A1(_06181_),
    .A2(_06070_),
    .B(net2399),
    .Y(_08582_));
 AO21x1_ASAP7_75t_R _37936_ (.A1(_07475_),
    .A2(_06089_),
    .B(net2399),
    .Y(_08583_));
 NAND3x2_ASAP7_75t_R _37937_ (.B(_08583_),
    .C(_07843_),
    .Y(_08584_),
    .A(_08582_));
 AO21x1_ASAP7_75t_R _37938_ (.A1(net1216),
    .A2(net2234),
    .B(net2764),
    .Y(_08585_));
 OAI21x1_ASAP7_75t_R _37939_ (.A1(net2764),
    .A2(_06226_),
    .B(_08585_),
    .Y(_08586_));
 NOR3x2_ASAP7_75t_R _37940_ (.B(_06832_),
    .C(_08586_),
    .Y(_08587_),
    .A(_08584_));
 AOI22x1_ASAP7_75t_R _37941_ (.A1(_07351_),
    .A2(_06058_),
    .B1(_07455_),
    .B2(net3473),
    .Y(_08588_));
 AO21x1_ASAP7_75t_R _37942_ (.A1(net3231),
    .A2(net1217),
    .B(net2786),
    .Y(_08589_));
 NAND3x1_ASAP7_75t_R _37943_ (.A(_08588_),
    .B(_07825_),
    .C(_08589_),
    .Y(_08590_));
 AOI211x1_ASAP7_75t_R _37944_ (.A1(_06029_),
    .A2(net1551),
    .B(net1590),
    .C(_06064_),
    .Y(_08591_));
 NOR2x1_ASAP7_75t_R _37945_ (.A(_08591_),
    .B(_06818_),
    .Y(_08593_));
 NAND2x1_ASAP7_75t_R _37946_ (.A(_06256_),
    .B(_06816_),
    .Y(_08594_));
 AO21x1_ASAP7_75t_R _37947_ (.A1(_06181_),
    .A2(net2234),
    .B(_06064_),
    .Y(_08595_));
 NAND3x1_ASAP7_75t_R _37948_ (.A(_08593_),
    .B(_08594_),
    .C(_08595_),
    .Y(_08596_));
 NOR2x1_ASAP7_75t_R _37949_ (.A(_08590_),
    .B(_08596_),
    .Y(_08597_));
 NAND2x2_ASAP7_75t_R _37950_ (.A(_08587_),
    .B(_08597_),
    .Y(_08598_));
 NOR2x2_ASAP7_75t_R _37951_ (.A(_08580_),
    .B(_08598_),
    .Y(_08599_));
 NAND2x2_ASAP7_75t_R _37952_ (.A(_08563_),
    .B(_08599_),
    .Y(_08600_));
 NOR2x2_ASAP7_75t_R _37953_ (.A(_06890_),
    .B(_08600_),
    .Y(_08601_));
 NAND2x2_ASAP7_75t_R _37954_ (.A(_08601_),
    .B(_08504_),
    .Y(_08602_));
 OAI22x1_ASAP7_75t_R _37955_ (.A1(_08600_),
    .A2(_06890_),
    .B1(_08503_),
    .B2(_05717_),
    .Y(_08604_));
 AO21x1_ASAP7_75t_R _37956_ (.A1(_05833_),
    .A2(_05860_),
    .B(net3352),
    .Y(_08605_));
 AO21x1_ASAP7_75t_R _37957_ (.A1(net2423),
    .A2(net3355),
    .B(net3352),
    .Y(_08606_));
 NAND2x1_ASAP7_75t_R _37958_ (.A(_05930_),
    .B(_05953_),
    .Y(_08607_));
 AND3x1_ASAP7_75t_R _37959_ (.A(_08605_),
    .B(_08606_),
    .C(_08607_),
    .Y(_08608_));
 AO21x1_ASAP7_75t_R _37960_ (.A1(net1037),
    .A2(_05796_),
    .B(_05938_),
    .Y(_08609_));
 OAI21x1_ASAP7_75t_R _37961_ (.A1(_05807_),
    .A2(_05938_),
    .B(_08609_),
    .Y(_08610_));
 OR3x2_ASAP7_75t_R _37962_ (.A(_05938_),
    .B(net1226),
    .C(_05741_),
    .Y(_08611_));
 NAND2x1_ASAP7_75t_R _37963_ (.A(_07503_),
    .B(_08611_),
    .Y(_08612_));
 NOR2x1_ASAP7_75t_R _37964_ (.A(_08610_),
    .B(_08612_),
    .Y(_08613_));
 NAND2x1_ASAP7_75t_R _37965_ (.A(_08608_),
    .B(_08613_),
    .Y(_08615_));
 AND3x1_ASAP7_75t_R _37966_ (.A(_05762_),
    .B(_05753_),
    .C(_07237_),
    .Y(_08616_));
 AO21x1_ASAP7_75t_R _37967_ (.A1(net980),
    .A2(_05887_),
    .B(_05787_),
    .Y(_08617_));
 NAND2x1_ASAP7_75t_R _37968_ (.A(_08023_),
    .B(_08617_),
    .Y(_08618_));
 OA211x2_ASAP7_75t_R _37969_ (.A1(_05740_),
    .A2(_05757_),
    .B(_05926_),
    .C(net2705),
    .Y(_08619_));
 NOR2x1_ASAP7_75t_R _37970_ (.A(_08618_),
    .B(_08619_),
    .Y(_08620_));
 NAND2x1_ASAP7_75t_R _37971_ (.A(_08616_),
    .B(_08620_),
    .Y(_08621_));
 NOR2x2_ASAP7_75t_R _37972_ (.A(_08615_),
    .B(_08621_),
    .Y(_08622_));
 NOR2x1_ASAP7_75t_R _37973_ (.A(_05993_),
    .B(net1807),
    .Y(_08623_));
 AO21x1_ASAP7_75t_R _37974_ (.A1(_06541_),
    .A2(_05844_),
    .B(_08623_),
    .Y(_08624_));
 NOR2x2_ASAP7_75t_R _37975_ (.A(net2232),
    .B(net2525),
    .Y(_08626_));
 INVx2_ASAP7_75t_R _37976_ (.A(_08626_),
    .Y(_08627_));
 AO21x1_ASAP7_75t_R _37977_ (.A1(net2743),
    .A2(_05817_),
    .B(net2525),
    .Y(_08628_));
 NAND2x1_ASAP7_75t_R _37978_ (.A(_08627_),
    .B(_08628_),
    .Y(_08629_));
 NOR2x1_ASAP7_75t_R _37979_ (.A(_08624_),
    .B(_08629_),
    .Y(_08630_));
 OA21x2_ASAP7_75t_R _37980_ (.A1(net2519),
    .A2(_05897_),
    .B(_06017_),
    .Y(_08631_));
 NOR3x1_ASAP7_75t_R _37981_ (.A(_08631_),
    .B(_08043_),
    .C(_06011_),
    .Y(_08632_));
 AOI21x1_ASAP7_75t_R _37982_ (.A1(_05880_),
    .A2(_06017_),
    .B(_06018_),
    .Y(_08633_));
 NAND3x1_ASAP7_75t_R _37983_ (.A(_08630_),
    .B(_08632_),
    .C(_08633_),
    .Y(_08634_));
 OAI21x1_ASAP7_75t_R _37984_ (.A1(_05931_),
    .A2(_06494_),
    .B(net2636),
    .Y(_08635_));
 NAND2x1_ASAP7_75t_R _37985_ (.A(net2636),
    .B(_06521_),
    .Y(_08637_));
 OA211x2_ASAP7_75t_R _37986_ (.A1(_07522_),
    .A2(_05933_),
    .B(_08635_),
    .C(_08637_),
    .Y(_08638_));
 NAND2x1_ASAP7_75t_R _37987_ (.A(_05986_),
    .B(_05984_),
    .Y(_08639_));
 OA21x2_ASAP7_75t_R _37988_ (.A1(_06515_),
    .A2(net1178),
    .B(_05978_),
    .Y(_08640_));
 NOR2x1_ASAP7_75t_R _37989_ (.A(_05977_),
    .B(_07168_),
    .Y(_08641_));
 NOR3x1_ASAP7_75t_R _37990_ (.A(_08639_),
    .B(_08640_),
    .C(_08641_),
    .Y(_08642_));
 NAND2x1_ASAP7_75t_R _37991_ (.A(_08638_),
    .B(_08642_),
    .Y(_08643_));
 NOR2x1_ASAP7_75t_R _37992_ (.A(_08643_),
    .B(_08634_),
    .Y(_08644_));
 NAND2x2_ASAP7_75t_R _37993_ (.A(_08622_),
    .B(_08644_),
    .Y(_08645_));
 AO21x1_ASAP7_75t_R _37994_ (.A1(net3468),
    .A2(net2081),
    .B(_05800_),
    .Y(_08646_));
 AO21x1_ASAP7_75t_R _37995_ (.A1(net1807),
    .A2(net1695),
    .B(_05800_),
    .Y(_08648_));
 NAND2x1_ASAP7_75t_R _37996_ (.A(_05880_),
    .B(_05812_),
    .Y(_08649_));
 AND3x1_ASAP7_75t_R _37997_ (.A(_08646_),
    .B(_08648_),
    .C(_08649_),
    .Y(_08650_));
 AO21x1_ASAP7_75t_R _37998_ (.A1(net2743),
    .A2(net2485),
    .B(net3351),
    .Y(_08651_));
 AO21x1_ASAP7_75t_R _37999_ (.A1(net2098),
    .A2(_05850_),
    .B(net3351),
    .Y(_08652_));
 NAND2x1_ASAP7_75t_R _38000_ (.A(_08651_),
    .B(_08652_),
    .Y(_08653_));
 AO21x1_ASAP7_75t_R _38001_ (.A1(net1805),
    .A2(_06429_),
    .B(_05821_),
    .Y(_08654_));
 OAI21x1_ASAP7_75t_R _38002_ (.A1(net1118),
    .A2(net3351),
    .B(_08654_),
    .Y(_08655_));
 NOR2x1_ASAP7_75t_R _38003_ (.A(_08653_),
    .B(_08655_),
    .Y(_08656_));
 NAND2x2_ASAP7_75t_R _38004_ (.A(_08650_),
    .B(_08656_),
    .Y(_08657_));
 OA21x2_ASAP7_75t_R _38005_ (.A1(_07229_),
    .A2(net2679),
    .B(_05856_),
    .Y(_08659_));
 AO21x1_ASAP7_75t_R _38006_ (.A1(net1560),
    .A2(_07207_),
    .B(net2679),
    .Y(_08660_));
 AO21x1_ASAP7_75t_R _38007_ (.A1(net2270),
    .A2(_05918_),
    .B(_05839_),
    .Y(_08661_));
 AO21x1_ASAP7_75t_R _38008_ (.A1(net1805),
    .A2(net3372),
    .B(_05839_),
    .Y(_08662_));
 AND2x2_ASAP7_75t_R _38009_ (.A(_08661_),
    .B(_08662_),
    .Y(_08663_));
 NAND3x2_ASAP7_75t_R _38010_ (.B(_08660_),
    .C(_08663_),
    .Y(_08664_),
    .A(_08659_));
 NOR2x2_ASAP7_75t_R _38011_ (.A(_08657_),
    .B(_08664_),
    .Y(_08665_));
 AOI211x1_ASAP7_75t_R _38012_ (.A1(_05764_),
    .A2(net1776),
    .B(_05873_),
    .C(net1445),
    .Y(_08666_));
 OA21x2_ASAP7_75t_R _38013_ (.A1(_06481_),
    .A2(_06472_),
    .B(_05878_),
    .Y(_08667_));
 NOR2x1_ASAP7_75t_R _38014_ (.A(_08666_),
    .B(_08667_),
    .Y(_08668_));
 NAND2x1_ASAP7_75t_R _38015_ (.A(_05810_),
    .B(net1811),
    .Y(_08670_));
 AOI21x1_ASAP7_75t_R _38016_ (.A1(_05905_),
    .A2(_08670_),
    .B(_05884_),
    .Y(_08671_));
 AOI21x1_ASAP7_75t_R _38017_ (.A1(net2743),
    .A2(_07501_),
    .B(_05884_),
    .Y(_08672_));
 NOR2x1_ASAP7_75t_R _38018_ (.A(_08671_),
    .B(_08672_),
    .Y(_08673_));
 AO21x1_ASAP7_75t_R _38019_ (.A1(_05807_),
    .A2(net2541),
    .B(_05873_),
    .Y(_08674_));
 NAND3x1_ASAP7_75t_R _38020_ (.A(_08668_),
    .B(_08673_),
    .C(_08674_),
    .Y(_08675_));
 OA21x2_ASAP7_75t_R _38021_ (.A1(_05931_),
    .A2(_06494_),
    .B(_05898_),
    .Y(_08676_));
 NAND2x1_ASAP7_75t_R _38022_ (.A(_06461_),
    .B(_07190_),
    .Y(_08677_));
 NOR2x1_ASAP7_75t_R _38023_ (.A(_08676_),
    .B(_08677_),
    .Y(_08678_));
 AO21x1_ASAP7_75t_R _38024_ (.A1(_05850_),
    .A2(net1913),
    .B(_05894_),
    .Y(_08679_));
 AO21x1_ASAP7_75t_R _38025_ (.A1(_05857_),
    .A2(net2845),
    .B(_05894_),
    .Y(_08681_));
 AND2x2_ASAP7_75t_R _38026_ (.A(_08679_),
    .B(_08681_),
    .Y(_08682_));
 AO21x1_ASAP7_75t_R _38027_ (.A1(net2743),
    .A2(_05835_),
    .B(_05908_),
    .Y(_08683_));
 AO21x1_ASAP7_75t_R _38028_ (.A1(net1786),
    .A2(_07207_),
    .B(_05908_),
    .Y(_08684_));
 AND2x2_ASAP7_75t_R _38029_ (.A(_08683_),
    .B(_08684_),
    .Y(_08685_));
 NAND3x1_ASAP7_75t_R _38030_ (.A(_08678_),
    .B(_08682_),
    .C(_08685_),
    .Y(_08686_));
 NOR2x1_ASAP7_75t_R _38031_ (.A(_08675_),
    .B(_08686_),
    .Y(_08687_));
 NAND2x2_ASAP7_75t_R _38032_ (.A(_08665_),
    .B(_08687_),
    .Y(_08688_));
 NOR3x2_ASAP7_75t_R _38033_ (.B(_08645_),
    .C(_08688_),
    .Y(_08689_),
    .A(_06425_));
 NAND3x1_ASAP7_75t_R _38034_ (.A(_08602_),
    .B(_08604_),
    .C(_08689_),
    .Y(_08690_));
 INVx1_ASAP7_75t_R _38035_ (.A(_08690_),
    .Y(_08692_));
 AO21x1_ASAP7_75t_R _38036_ (.A1(_08602_),
    .A2(_08604_),
    .B(_08689_),
    .Y(_08693_));
 INVx1_ASAP7_75t_R _38037_ (.A(_08693_),
    .Y(_08694_));
 INVx1_ASAP7_75t_R _38038_ (.A(_05468_),
    .Y(_08695_));
 AO21x1_ASAP7_75t_R _38039_ (.A1(_05685_),
    .A2(net1667),
    .B(_05472_),
    .Y(_08696_));
 AO21x1_ASAP7_75t_R _38040_ (.A1(net2191),
    .A2(net3115),
    .B(_05472_),
    .Y(_08697_));
 NAND2x1_ASAP7_75t_R _38041_ (.A(_08696_),
    .B(_08697_),
    .Y(_08698_));
 OR3x1_ASAP7_75t_R _38042_ (.A(_07079_),
    .B(_08695_),
    .C(_08698_),
    .Y(_08699_));
 AO21x1_ASAP7_75t_R _38043_ (.A1(net2833),
    .A2(_05486_),
    .B(net2389),
    .Y(_08700_));
 NAND2x1_ASAP7_75t_R _38044_ (.A(_05568_),
    .B(_05564_),
    .Y(_08701_));
 OA211x2_ASAP7_75t_R _38045_ (.A1(net1124),
    .A2(net2389),
    .B(_08700_),
    .C(_08701_),
    .Y(_08703_));
 OA21x2_ASAP7_75t_R _38046_ (.A1(_06637_),
    .A2(_05561_),
    .B(_05577_),
    .Y(_08704_));
 INVx1_ASAP7_75t_R _38047_ (.A(_08704_),
    .Y(_08705_));
 AO21x1_ASAP7_75t_R _38048_ (.A1(net2833),
    .A2(net1085),
    .B(_05581_),
    .Y(_08706_));
 NAND2x1_ASAP7_75t_R _38049_ (.A(_05577_),
    .B(_05441_),
    .Y(_08707_));
 AND4x1_ASAP7_75t_R _38050_ (.A(_08705_),
    .B(_08706_),
    .C(_08707_),
    .D(_07699_),
    .Y(_08708_));
 NAND2x1_ASAP7_75t_R _38051_ (.A(_08703_),
    .B(_08708_),
    .Y(_08709_));
 NOR2x1_ASAP7_75t_R _38052_ (.A(_08699_),
    .B(_08709_),
    .Y(_08710_));
 AO21x1_ASAP7_75t_R _38053_ (.A1(_05447_),
    .A2(net2663),
    .B(_05492_),
    .Y(_08711_));
 OAI21x1_ASAP7_75t_R _38054_ (.A1(_05457_),
    .A2(_05492_),
    .B(_08711_),
    .Y(_08712_));
 NAND2x1_ASAP7_75t_R _38055_ (.A(_05499_),
    .B(_07718_),
    .Y(_08714_));
 OA21x2_ASAP7_75t_R _38056_ (.A1(net3106),
    .A2(_06647_),
    .B(net3373),
    .Y(_08715_));
 OA21x2_ASAP7_75t_R _38057_ (.A1(_07066_),
    .A2(net1528),
    .B(net3373),
    .Y(_08716_));
 OR4x1_ASAP7_75t_R _38058_ (.A(_08712_),
    .B(_08714_),
    .C(_08715_),
    .D(_08716_),
    .Y(_08717_));
 AO21x1_ASAP7_75t_R _38059_ (.A1(_06627_),
    .A2(_06626_),
    .B(_06631_),
    .Y(_08718_));
 OA21x2_ASAP7_75t_R _38060_ (.A1(net2834),
    .A2(_05566_),
    .B(_06627_),
    .Y(_08719_));
 AO21x1_ASAP7_75t_R _38061_ (.A1(_06627_),
    .A2(_06637_),
    .B(_08719_),
    .Y(_08720_));
 NOR2x1_ASAP7_75t_R _38062_ (.A(_08718_),
    .B(_08720_),
    .Y(_08721_));
 AO21x1_ASAP7_75t_R _38063_ (.A1(net1627),
    .A2(net2658),
    .B(_05548_),
    .Y(_08722_));
 AO21x1_ASAP7_75t_R _38064_ (.A1(_05496_),
    .A2(net2509),
    .B(_05548_),
    .Y(_08723_));
 AND2x2_ASAP7_75t_R _38065_ (.A(_08722_),
    .B(_08723_),
    .Y(_08725_));
 AOI21x1_ASAP7_75t_R _38066_ (.A1(_05682_),
    .A2(_05545_),
    .B(_05555_),
    .Y(_08726_));
 NAND3x1_ASAP7_75t_R _38067_ (.A(_08721_),
    .B(_08725_),
    .C(_08726_),
    .Y(_08727_));
 NOR2x1_ASAP7_75t_R _38068_ (.A(_08717_),
    .B(_08727_),
    .Y(_08728_));
 NAND2x1_ASAP7_75t_R _38069_ (.A(_08710_),
    .B(_08728_),
    .Y(_08729_));
 AO21x1_ASAP7_75t_R _38070_ (.A1(net3350),
    .A2(net2509),
    .B(net2447),
    .Y(_08730_));
 AO21x1_ASAP7_75t_R _38071_ (.A1(net2658),
    .A2(net1773),
    .B(net2447),
    .Y(_08731_));
 AO21x1_ASAP7_75t_R _38072_ (.A1(net1083),
    .A2(net2401),
    .B(net2447),
    .Y(_08732_));
 NAND2x1_ASAP7_75t_R _38073_ (.A(net3106),
    .B(_06613_),
    .Y(_08733_));
 AND4x1_ASAP7_75t_R _38074_ (.A(_08730_),
    .B(_08731_),
    .C(_08732_),
    .D(_08733_),
    .Y(_08734_));
 AO21x1_ASAP7_75t_R _38075_ (.A1(net3349),
    .A2(net1267),
    .B(net2411),
    .Y(_08736_));
 AO21x1_ASAP7_75t_R _38076_ (.A1(net2003),
    .A2(net2116),
    .B(net2411),
    .Y(_08737_));
 OA211x2_ASAP7_75t_R _38077_ (.A1(net2221),
    .A2(net2411),
    .B(_08736_),
    .C(_08737_),
    .Y(_08738_));
 NAND2x1_ASAP7_75t_R _38078_ (.A(_08734_),
    .B(_08738_),
    .Y(_08739_));
 AO21x1_ASAP7_75t_R _38079_ (.A1(net1124),
    .A2(_05676_),
    .B(net2616),
    .Y(_08740_));
 OA211x2_ASAP7_75t_R _38080_ (.A1(_05496_),
    .A2(net2616),
    .B(_05641_),
    .C(_08740_),
    .Y(_08741_));
 AO21x1_ASAP7_75t_R _38081_ (.A1(net1772),
    .A2(net1267),
    .B(net2461),
    .Y(_08742_));
 AO21x1_ASAP7_75t_R _38082_ (.A1(net2401),
    .A2(net2613),
    .B(net2461),
    .Y(_08743_));
 OA211x2_ASAP7_75t_R _38083_ (.A1(net2461),
    .A2(net1627),
    .B(_08742_),
    .C(_08743_),
    .Y(_08744_));
 NAND2x1_ASAP7_75t_R _38084_ (.A(_08741_),
    .B(_08744_),
    .Y(_08745_));
 NOR2x1_ASAP7_75t_R _38085_ (.A(_08739_),
    .B(_08745_),
    .Y(_08747_));
 AO21x1_ASAP7_75t_R _38086_ (.A1(net2703),
    .A2(net1772),
    .B(_05683_),
    .Y(_08748_));
 AO21x1_ASAP7_75t_R _38087_ (.A1(_05496_),
    .A2(net2509),
    .B(_05683_),
    .Y(_08749_));
 OA211x2_ASAP7_75t_R _38088_ (.A1(_05683_),
    .A2(_07112_),
    .B(_08748_),
    .C(_08749_),
    .Y(_08750_));
 NAND2x1_ASAP7_75t_R _38089_ (.A(_05675_),
    .B(_05665_),
    .Y(_08751_));
 NOR2x2_ASAP7_75t_R _38090_ (.A(_05677_),
    .B(net3356),
    .Y(_08752_));
 INVx1_ASAP7_75t_R _38091_ (.A(_08752_),
    .Y(_08753_));
 AND4x1_ASAP7_75t_R _38092_ (.A(_07788_),
    .B(_06563_),
    .C(_08751_),
    .D(_08753_),
    .Y(_08754_));
 AND2x2_ASAP7_75t_R _38093_ (.A(_08750_),
    .B(_08754_),
    .Y(_08755_));
 AO21x1_ASAP7_75t_R _38094_ (.A1(net1083),
    .A2(net2401),
    .B(_06576_),
    .Y(_08756_));
 AO21x1_ASAP7_75t_R _38095_ (.A1(net2567),
    .A2(net2612),
    .B(_06576_),
    .Y(_08758_));
 AND3x1_ASAP7_75t_R _38096_ (.A(_08756_),
    .B(_08758_),
    .C(_06581_),
    .Y(_08759_));
 AO21x1_ASAP7_75t_R _38097_ (.A1(net3356),
    .A2(net2815),
    .B(_06576_),
    .Y(_08760_));
 AO21x1_ASAP7_75t_R _38098_ (.A1(net2658),
    .A2(net1772),
    .B(_06576_),
    .Y(_08761_));
 AND2x2_ASAP7_75t_R _38099_ (.A(_08760_),
    .B(_08761_),
    .Y(_08762_));
 AO21x1_ASAP7_75t_R _38100_ (.A1(net3350),
    .A2(_05464_),
    .B(_05654_),
    .Y(_08763_));
 AO21x1_ASAP7_75t_R _38101_ (.A1(net2115),
    .A2(_05676_),
    .B(_05654_),
    .Y(_08764_));
 AND2x2_ASAP7_75t_R _38102_ (.A(_08763_),
    .B(_08764_),
    .Y(_08765_));
 AND3x1_ASAP7_75t_R _38103_ (.A(_08759_),
    .B(_08762_),
    .C(_08765_),
    .Y(_08766_));
 AND2x4_ASAP7_75t_R _38104_ (.A(_08755_),
    .B(_08766_),
    .Y(_08767_));
 NAND2x2_ASAP7_75t_R _38105_ (.A(_08747_),
    .B(_08767_),
    .Y(_08769_));
 NOR2x2_ASAP7_75t_R _38106_ (.A(_08729_),
    .B(_08769_),
    .Y(_08770_));
 NAND2x2_ASAP7_75t_R _38107_ (.A(_05479_),
    .B(_08770_),
    .Y(_08771_));
 AO21x1_ASAP7_75t_R _38108_ (.A1(net3101),
    .A2(net1237),
    .B(_05062_),
    .Y(_08772_));
 AO21x1_ASAP7_75t_R _38109_ (.A1(net1877),
    .A2(_05360_),
    .B(_05062_),
    .Y(_08773_));
 NOR2x1_ASAP7_75t_R _38110_ (.A(_05062_),
    .B(net3454),
    .Y(_08774_));
 INVx1_ASAP7_75t_R _38111_ (.A(_08774_),
    .Y(_08775_));
 NAND3x1_ASAP7_75t_R _38112_ (.A(_08772_),
    .B(_08773_),
    .C(_08775_),
    .Y(_08776_));
 INVx1_ASAP7_75t_R _38113_ (.A(_05128_),
    .Y(_08777_));
 AO21x1_ASAP7_75t_R _38114_ (.A1(_08777_),
    .A2(net1154),
    .B(_05219_),
    .Y(_08778_));
 AO21x1_ASAP7_75t_R _38115_ (.A1(net1921),
    .A2(net1091),
    .B(net3411),
    .Y(_08780_));
 AO21x1_ASAP7_75t_R _38116_ (.A1(_05206_),
    .A2(net1140),
    .B(net3411),
    .Y(_08781_));
 NAND2x1_ASAP7_75t_R _38117_ (.A(_08780_),
    .B(_08781_),
    .Y(_08782_));
 NOR3x1_ASAP7_75t_R _38118_ (.A(_08776_),
    .B(_08778_),
    .C(_08782_),
    .Y(_08783_));
 AO21x1_ASAP7_75t_R _38119_ (.A1(_05265_),
    .A2(net2149),
    .B(_05118_),
    .Y(_08784_));
 NAND3x1_ASAP7_75t_R _38120_ (.A(_05374_),
    .B(_08784_),
    .C(_07645_),
    .Y(_08785_));
 OA211x2_ASAP7_75t_R _38121_ (.A1(net3436),
    .A2(net3442),
    .B(_06394_),
    .C(_05066_),
    .Y(_08786_));
 OA21x2_ASAP7_75t_R _38122_ (.A1(_05106_),
    .A2(_05092_),
    .B(_06394_),
    .Y(_08787_));
 NOR3x1_ASAP7_75t_R _38123_ (.A(_08785_),
    .B(_08786_),
    .C(_08787_),
    .Y(_08788_));
 NAND2x1_ASAP7_75t_R _38124_ (.A(_08783_),
    .B(_08788_),
    .Y(_08789_));
 AO21x1_ASAP7_75t_R _38125_ (.A1(_05206_),
    .A2(_05143_),
    .B(_05198_),
    .Y(_08791_));
 NAND2x1_ASAP7_75t_R _38126_ (.A(_07646_),
    .B(_05199_),
    .Y(_08792_));
 NAND3x1_ASAP7_75t_R _38127_ (.A(_08791_),
    .B(_08102_),
    .C(_08792_),
    .Y(_08793_));
 AO21x1_ASAP7_75t_R _38128_ (.A1(net1921),
    .A2(net1091),
    .B(_05208_),
    .Y(_08794_));
 NAND2x1_ASAP7_75t_R _38129_ (.A(_08794_),
    .B(_05330_),
    .Y(_08795_));
 AO21x1_ASAP7_75t_R _38130_ (.A1(_05058_),
    .A2(net964),
    .B(_05208_),
    .Y(_08796_));
 AO21x1_ASAP7_75t_R _38131_ (.A1(net2139),
    .A2(net1877),
    .B(_05208_),
    .Y(_08797_));
 NAND2x1_ASAP7_75t_R _38132_ (.A(_08796_),
    .B(_08797_),
    .Y(_08798_));
 NOR3x1_ASAP7_75t_R _38133_ (.A(_08793_),
    .B(_08795_),
    .C(_08798_),
    .Y(_08799_));
 AO21x1_ASAP7_75t_R _38134_ (.A1(_05181_),
    .A2(_05205_),
    .B(_07680_),
    .Y(_08800_));
 AO21x1_ASAP7_75t_R _38135_ (.A1(net1768),
    .A2(net1091),
    .B(net3095),
    .Y(_08802_));
 AO21x1_ASAP7_75t_R _38136_ (.A1(_05265_),
    .A2(net1140),
    .B(net3095),
    .Y(_08803_));
 AO21x1_ASAP7_75t_R _38137_ (.A1(_05058_),
    .A2(_05090_),
    .B(net3095),
    .Y(_08804_));
 NAND3x1_ASAP7_75t_R _38138_ (.A(_08802_),
    .B(_08803_),
    .C(_08804_),
    .Y(_08805_));
 AO21x1_ASAP7_75t_R _38139_ (.A1(net990),
    .A2(net964),
    .B(_05256_),
    .Y(_08806_));
 NAND2x1_ASAP7_75t_R _38140_ (.A(_08806_),
    .B(_06378_),
    .Y(_08807_));
 NOR3x1_ASAP7_75t_R _38141_ (.A(_08800_),
    .B(_08805_),
    .C(_08807_),
    .Y(_08808_));
 NAND2x1_ASAP7_75t_R _38142_ (.A(_08799_),
    .B(_08808_),
    .Y(_08809_));
 NOR2x2_ASAP7_75t_R _38143_ (.A(_08789_),
    .B(_08809_),
    .Y(_08810_));
 AO21x1_ASAP7_75t_R _38144_ (.A1(net1835),
    .A2(_05058_),
    .B(_05186_),
    .Y(_08811_));
 INVx1_ASAP7_75t_R _38145_ (.A(_07635_),
    .Y(_08813_));
 NAND3x1_ASAP7_75t_R _38146_ (.A(_05417_),
    .B(_08811_),
    .C(_08813_),
    .Y(_08814_));
 AO21x1_ASAP7_75t_R _38147_ (.A1(_05202_),
    .A2(_05089_),
    .B(_05345_),
    .Y(_08815_));
 AO21x1_ASAP7_75t_R _38148_ (.A1(_08815_),
    .A2(net1794),
    .B(_05215_),
    .Y(_08816_));
 OAI21x1_ASAP7_75t_R _38149_ (.A1(_05215_),
    .A2(_05233_),
    .B(_08816_),
    .Y(_08817_));
 NOR2x1_ASAP7_75t_R _38150_ (.A(_08814_),
    .B(_08817_),
    .Y(_08818_));
 AO21x1_ASAP7_75t_R _38151_ (.A1(net1091),
    .A2(net2149),
    .B(_05306_),
    .Y(_08819_));
 AO21x1_ASAP7_75t_R _38152_ (.A1(net3426),
    .A2(_05259_),
    .B(_05306_),
    .Y(_08820_));
 NAND2x1_ASAP7_75t_R _38153_ (.A(_05100_),
    .B(net2161),
    .Y(_08821_));
 NAND2x1_ASAP7_75t_R _38154_ (.A(_05100_),
    .B(_06323_),
    .Y(_08822_));
 AND4x1_ASAP7_75t_R _38155_ (.A(_08819_),
    .B(_08820_),
    .C(_08821_),
    .D(_08822_),
    .Y(_08824_));
 NOR2x1_ASAP7_75t_R _38156_ (.A(_07036_),
    .B(_05323_),
    .Y(_08825_));
 NAND3x1_ASAP7_75t_R _38157_ (.A(_08818_),
    .B(_08824_),
    .C(_08825_),
    .Y(_08826_));
 OA21x2_ASAP7_75t_R _38158_ (.A1(net2493),
    .A2(_05345_),
    .B(_06341_),
    .Y(_08827_));
 AO21x1_ASAP7_75t_R _38159_ (.A1(net1867),
    .A2(net1091),
    .B(net2621),
    .Y(_08828_));
 AO21x1_ASAP7_75t_R _38160_ (.A1(_07609_),
    .A2(net992),
    .B(net2621),
    .Y(_08829_));
 AND2x2_ASAP7_75t_R _38161_ (.A(_08828_),
    .B(_08829_),
    .Y(_08830_));
 OAI21x1_ASAP7_75t_R _38162_ (.A1(net2493),
    .A2(_05122_),
    .B(_05266_),
    .Y(_08831_));
 INVx1_ASAP7_75t_R _38163_ (.A(_08831_),
    .Y(_08832_));
 AND3x1_ASAP7_75t_R _38164_ (.A(_08827_),
    .B(_08830_),
    .C(_08832_),
    .Y(_08833_));
 OA21x2_ASAP7_75t_R _38165_ (.A1(_05185_),
    .A2(net2529),
    .B(_05267_),
    .Y(_08835_));
 NOR2x1_ASAP7_75t_R _38166_ (.A(_05119_),
    .B(net2529),
    .Y(_08836_));
 AOI211x1_ASAP7_75t_R _38167_ (.A1(_06328_),
    .A2(net1322),
    .B(_05300_),
    .C(_08836_),
    .Y(_08837_));
 NAND2x1_ASAP7_75t_R _38168_ (.A(_08835_),
    .B(_08837_),
    .Y(_08838_));
 AO21x1_ASAP7_75t_R _38169_ (.A1(_05206_),
    .A2(net2146),
    .B(_05086_),
    .Y(_08839_));
 OA21x2_ASAP7_75t_R _38170_ (.A1(net1237),
    .A2(_05086_),
    .B(_08839_),
    .Y(_08840_));
 NAND2x1_ASAP7_75t_R _38171_ (.A(_05087_),
    .B(_06346_),
    .Y(_08841_));
 AND2x2_ASAP7_75t_R _38172_ (.A(_06333_),
    .B(_08841_),
    .Y(_08842_));
 NAND2x1_ASAP7_75t_R _38173_ (.A(_08840_),
    .B(_08842_),
    .Y(_08843_));
 NOR2x1_ASAP7_75t_R _38174_ (.A(_08838_),
    .B(_08843_),
    .Y(_08844_));
 NAND2x1_ASAP7_75t_R _38175_ (.A(_08833_),
    .B(_08844_),
    .Y(_08846_));
 NOR2x1_ASAP7_75t_R _38176_ (.A(_08826_),
    .B(_08846_),
    .Y(_08847_));
 NAND2x2_ASAP7_75t_R _38177_ (.A(_08810_),
    .B(_08847_),
    .Y(_08848_));
 NOR2x2_ASAP7_75t_R _38178_ (.A(_05717_),
    .B(_08848_),
    .Y(_08849_));
 XOR2x2_ASAP7_75t_R _38179_ (.A(_08771_),
    .B(_08849_),
    .Y(_08850_));
 OAI21x1_ASAP7_75t_R _38180_ (.A1(_08692_),
    .A2(_08694_),
    .B(net3347),
    .Y(_08851_));
 NOR2x2_ASAP7_75t_R _38181_ (.A(_08688_),
    .B(_08645_),
    .Y(_08852_));
 NAND2x2_ASAP7_75t_R _38182_ (.A(net1978),
    .B(_08852_),
    .Y(_08853_));
 AO21x1_ASAP7_75t_R _38183_ (.A1(_08602_),
    .A2(_08604_),
    .B(net1948),
    .Y(_08854_));
 NAND3x1_ASAP7_75t_R _38184_ (.A(_08602_),
    .B(_08604_),
    .C(net1948),
    .Y(_08855_));
 AOI21x1_ASAP7_75t_R _38185_ (.A1(_08854_),
    .A2(_08855_),
    .B(_08850_),
    .Y(_08856_));
 INVx1_ASAP7_75t_R _38186_ (.A(_08856_),
    .Y(_08857_));
 AOI21x1_ASAP7_75t_R _38187_ (.A1(_08851_),
    .A2(_08857_),
    .B(net388),
    .Y(_08858_));
 OAI21x1_ASAP7_75t_R _38188_ (.A1(_08524_),
    .A2(_08858_),
    .B(_00497_),
    .Y(_08859_));
 XNOR2x2_ASAP7_75t_R _38189_ (.A(_08849_),
    .B(_08771_),
    .Y(_08860_));
 AOI21x1_ASAP7_75t_R _38190_ (.A1(_08693_),
    .A2(_08690_),
    .B(_08860_),
    .Y(_08861_));
 OAI21x1_ASAP7_75t_R _38191_ (.A1(_08856_),
    .A2(_08861_),
    .B(net394),
    .Y(_08862_));
 INVx1_ASAP7_75t_R _38192_ (.A(_08524_),
    .Y(_08863_));
 NAND3x2_ASAP7_75t_R _38193_ (.B(_14360_),
    .C(_08863_),
    .Y(_08864_),
    .A(_08862_));
 NAND2x2_ASAP7_75t_R _38194_ (.A(_08864_),
    .B(_08859_),
    .Y(_00111_));
 NAND2x1_ASAP7_75t_R _38195_ (.A(_06481_),
    .B(_05898_),
    .Y(_08866_));
 NAND3x1_ASAP7_75t_R _38196_ (.A(_08681_),
    .B(_07191_),
    .C(_08866_),
    .Y(_08867_));
 AO31x2_ASAP7_75t_R _38197_ (.A1(net2845),
    .A2(_05918_),
    .A3(net3467),
    .B(_05908_),
    .Y(_08868_));
 AO21x1_ASAP7_75t_R _38198_ (.A1(net2423),
    .A2(net2736),
    .B(_05908_),
    .Y(_08869_));
 NAND3x1_ASAP7_75t_R _38199_ (.A(_08868_),
    .B(_07548_),
    .C(_08869_),
    .Y(_08870_));
 NOR2x1_ASAP7_75t_R _38200_ (.A(_08867_),
    .B(_08870_),
    .Y(_08871_));
 AO21x1_ASAP7_75t_R _38201_ (.A1(net3357),
    .A2(net3467),
    .B(_05873_),
    .Y(_08872_));
 AO21x1_ASAP7_75t_R _38202_ (.A1(_06490_),
    .A2(net2416),
    .B(_05873_),
    .Y(_08873_));
 AND3x1_ASAP7_75t_R _38203_ (.A(_08872_),
    .B(_05877_),
    .C(_08873_),
    .Y(_08874_));
 AO21x1_ASAP7_75t_R _38204_ (.A1(net3466),
    .A2(net1786),
    .B(_05884_),
    .Y(_08875_));
 AO21x1_ASAP7_75t_R _38205_ (.A1(net2416),
    .A2(_05807_),
    .B(_05884_),
    .Y(_08877_));
 NAND2x1_ASAP7_75t_R _38206_ (.A(_05897_),
    .B(_05885_),
    .Y(_08878_));
 AND3x1_ASAP7_75t_R _38207_ (.A(_08875_),
    .B(_08877_),
    .C(_08878_),
    .Y(_08879_));
 AND2x2_ASAP7_75t_R _38208_ (.A(_08874_),
    .B(_08879_),
    .Y(_08880_));
 NAND2x1_ASAP7_75t_R _38209_ (.A(_08871_),
    .B(_08880_),
    .Y(_08881_));
 AO21x1_ASAP7_75t_R _38210_ (.A1(_05817_),
    .A2(net2098),
    .B(_05821_),
    .Y(_08882_));
 NAND2x1_ASAP7_75t_R _38211_ (.A(_05930_),
    .B(_05829_),
    .Y(_08883_));
 AO21x1_ASAP7_75t_R _38212_ (.A1(_05807_),
    .A2(net2737),
    .B(_05821_),
    .Y(_08884_));
 AND3x1_ASAP7_75t_R _38213_ (.A(_08882_),
    .B(_08883_),
    .C(_08884_),
    .Y(_08885_));
 AOI211x1_ASAP7_75t_R _38214_ (.A1(net1224),
    .A2(net1779),
    .B(_05800_),
    .C(_05957_),
    .Y(_08886_));
 AOI21x1_ASAP7_75t_R _38215_ (.A1(_06427_),
    .A2(net3357),
    .B(_05800_),
    .Y(_08888_));
 NOR3x1_ASAP7_75t_R _38216_ (.A(_08886_),
    .B(_07569_),
    .C(_08888_),
    .Y(_08889_));
 AND2x2_ASAP7_75t_R _38217_ (.A(_08885_),
    .B(_08889_),
    .Y(_08890_));
 AO21x1_ASAP7_75t_R _38218_ (.A1(_06453_),
    .A2(_05865_),
    .B(net2679),
    .Y(_08891_));
 AO21x1_ASAP7_75t_R _38219_ (.A1(_05817_),
    .A2(_07229_),
    .B(net2679),
    .Y(_08892_));
 AO21x1_ASAP7_75t_R _38220_ (.A1(_05819_),
    .A2(_05918_),
    .B(net2679),
    .Y(_08893_));
 NAND3x1_ASAP7_75t_R _38221_ (.A(_08891_),
    .B(_08892_),
    .C(_08893_),
    .Y(_08894_));
 AOI211x1_ASAP7_75t_R _38222_ (.A1(_05764_),
    .A2(_05755_),
    .B(_05839_),
    .C(net1440),
    .Y(_08895_));
 NOR2x1_ASAP7_75t_R _38223_ (.A(_06447_),
    .B(_08895_),
    .Y(_08896_));
 NAND2x1_ASAP7_75t_R _38224_ (.A(_06523_),
    .B(_05846_),
    .Y(_08897_));
 NAND3x1_ASAP7_75t_R _38225_ (.A(_08896_),
    .B(_08897_),
    .C(_08297_),
    .Y(_08899_));
 NOR2x1_ASAP7_75t_R _38226_ (.A(_08894_),
    .B(_08899_),
    .Y(_08900_));
 NAND2x2_ASAP7_75t_R _38227_ (.A(_08890_),
    .B(_08900_),
    .Y(_08901_));
 NOR2x2_ASAP7_75t_R _38228_ (.A(_08881_),
    .B(_08901_),
    .Y(_08902_));
 AND2x2_ASAP7_75t_R _38229_ (.A(_08605_),
    .B(_06502_),
    .Y(_08903_));
 AO21x1_ASAP7_75t_R _38230_ (.A1(_06429_),
    .A2(_05796_),
    .B(net3352),
    .Y(_08904_));
 AO21x1_ASAP7_75t_R _38231_ (.A1(_05879_),
    .A2(_05805_),
    .B(net3352),
    .Y(_08905_));
 AND2x2_ASAP7_75t_R _38232_ (.A(_08904_),
    .B(_08905_),
    .Y(_08906_));
 NAND2x1_ASAP7_75t_R _38233_ (.A(_08903_),
    .B(_08906_),
    .Y(_08907_));
 AO21x1_ASAP7_75t_R _38234_ (.A1(_05921_),
    .A2(net3370),
    .B(net2520),
    .Y(_08908_));
 NAND3x1_ASAP7_75t_R _38235_ (.A(_05948_),
    .B(_08611_),
    .C(_08908_),
    .Y(_08910_));
 NOR2x1_ASAP7_75t_R _38236_ (.A(_08907_),
    .B(_08910_),
    .Y(_08911_));
 AO31x2_ASAP7_75t_R _38237_ (.A1(_05775_),
    .A2(_05807_),
    .A3(_05887_),
    .B(_05787_),
    .Y(_08912_));
 AO21x1_ASAP7_75t_R _38238_ (.A1(_05817_),
    .A2(_07229_),
    .B(_05787_),
    .Y(_08913_));
 NAND3x1_ASAP7_75t_R _38239_ (.A(_08912_),
    .B(_08328_),
    .C(_08913_),
    .Y(_08914_));
 OA21x2_ASAP7_75t_R _38240_ (.A1(_06517_),
    .A2(_05845_),
    .B(_05751_),
    .Y(_08915_));
 NOR2x1_ASAP7_75t_R _38241_ (.A(net2416),
    .B(_05752_),
    .Y(_08916_));
 NOR2x1_ASAP7_75t_R _38242_ (.A(_05764_),
    .B(_05780_),
    .Y(_08917_));
 OR3x1_ASAP7_75t_R _38243_ (.A(_08915_),
    .B(_08916_),
    .C(_08917_),
    .Y(_08918_));
 NOR2x1_ASAP7_75t_R _38244_ (.A(_08914_),
    .B(_08918_),
    .Y(_08919_));
 NAND2x1_ASAP7_75t_R _38245_ (.A(_08911_),
    .B(_08919_),
    .Y(_08921_));
 OA21x2_ASAP7_75t_R _38246_ (.A1(_06521_),
    .A2(_05976_),
    .B(_05966_),
    .Y(_08922_));
 NAND2x1_ASAP7_75t_R _38247_ (.A(_08305_),
    .B(_06530_),
    .Y(_08923_));
 AOI211x1_ASAP7_75t_R _38248_ (.A1(net2636),
    .A2(_05776_),
    .B(_08922_),
    .C(_08923_),
    .Y(_08924_));
 AO21x1_ASAP7_75t_R _38249_ (.A1(net2875),
    .A2(net3471),
    .B(_05977_),
    .Y(_08925_));
 NAND2x1_ASAP7_75t_R _38250_ (.A(_05979_),
    .B(_08925_),
    .Y(_08926_));
 AO21x1_ASAP7_75t_R _38251_ (.A1(_05833_),
    .A2(net2846),
    .B(_05977_),
    .Y(_08927_));
 AO21x1_ASAP7_75t_R _38252_ (.A1(net2098),
    .A2(_05819_),
    .B(_05977_),
    .Y(_08928_));
 NAND2x1_ASAP7_75t_R _38253_ (.A(_08927_),
    .B(_08928_),
    .Y(_08929_));
 NOR2x1_ASAP7_75t_R _38254_ (.A(_08926_),
    .B(_08929_),
    .Y(_08930_));
 AND2x2_ASAP7_75t_R _38255_ (.A(_08930_),
    .B(_08924_),
    .Y(_08932_));
 AND2x2_ASAP7_75t_R _38256_ (.A(_06542_),
    .B(_08037_),
    .Y(_08933_));
 AO21x1_ASAP7_75t_R _38257_ (.A1(_05876_),
    .A2(net2231),
    .B(_05993_),
    .Y(_08934_));
 OA21x2_ASAP7_75t_R _38258_ (.A1(_06426_),
    .A2(net2525),
    .B(_08934_),
    .Y(_08935_));
 NAND2x1_ASAP7_75t_R _38259_ (.A(_08933_),
    .B(_08935_),
    .Y(_08936_));
 NOR2x1_ASAP7_75t_R _38260_ (.A(_05835_),
    .B(_06007_),
    .Y(_08937_));
 NOR2x1_ASAP7_75t_R _38261_ (.A(_08937_),
    .B(_08631_),
    .Y(_08938_));
 NAND2x1_ASAP7_75t_R _38262_ (.A(_06017_),
    .B(net2404),
    .Y(_08939_));
 AO21x1_ASAP7_75t_R _38263_ (.A1(net2875),
    .A2(_05905_),
    .B(_06007_),
    .Y(_08940_));
 NAND3x1_ASAP7_75t_R _38264_ (.A(_08938_),
    .B(_08939_),
    .C(_08940_),
    .Y(_08941_));
 NOR2x1_ASAP7_75t_R _38265_ (.A(_08936_),
    .B(_08941_),
    .Y(_08943_));
 NAND2x1_ASAP7_75t_R _38266_ (.A(_08932_),
    .B(_08943_),
    .Y(_08944_));
 NOR2x1_ASAP7_75t_R _38267_ (.A(_08921_),
    .B(_08944_),
    .Y(_08945_));
 NAND2x2_ASAP7_75t_R _38268_ (.A(_08902_),
    .B(_08945_),
    .Y(_08946_));
 INVx3_ASAP7_75t_R _38269_ (.A(_08946_),
    .Y(_08947_));
 XOR2x1_ASAP7_75t_R _38270_ (.A(_08849_),
    .Y(_08948_),
    .B(_08947_));
 INVx1_ASAP7_75t_R _38271_ (.A(_08948_),
    .Y(_08949_));
 AO21x1_ASAP7_75t_R _38272_ (.A1(net3331),
    .A2(_06150_),
    .B(_06710_),
    .Y(_08950_));
 AND3x1_ASAP7_75t_R _38273_ (.A(_08950_),
    .B(_07849_),
    .C(_06713_),
    .Y(_08951_));
 AO21x1_ASAP7_75t_R _38274_ (.A1(net3328),
    .A2(net1217),
    .B(_06121_),
    .Y(_08952_));
 INVx1_ASAP7_75t_R _38275_ (.A(net2531),
    .Y(_08954_));
 NAND2x1_ASAP7_75t_R _38276_ (.A(_08954_),
    .B(_06764_),
    .Y(_08955_));
 NAND2x1_ASAP7_75t_R _38277_ (.A(_06817_),
    .B(_06764_),
    .Y(_08956_));
 AND3x1_ASAP7_75t_R _38278_ (.A(_08952_),
    .B(_08955_),
    .C(_08956_),
    .Y(_08957_));
 AND2x2_ASAP7_75t_R _38279_ (.A(_08951_),
    .B(_08957_),
    .Y(_08958_));
 AND4x1_ASAP7_75t_R _38280_ (.A(_06883_),
    .B(_07472_),
    .C(_06884_),
    .D(_06885_),
    .Y(_08959_));
 AO21x1_ASAP7_75t_R _38281_ (.A1(_06863_),
    .A2(_06098_),
    .B(net2345),
    .Y(_08960_));
 AO21x1_ASAP7_75t_R _38282_ (.A1(net2639),
    .A2(net1217),
    .B(net2345),
    .Y(_08961_));
 AND3x1_ASAP7_75t_R _38283_ (.A(_08960_),
    .B(_08961_),
    .C(_08254_),
    .Y(_08962_));
 AND3x1_ASAP7_75t_R _38284_ (.A(_08958_),
    .B(_08959_),
    .C(_08962_),
    .Y(_08963_));
 AO21x1_ASAP7_75t_R _38285_ (.A1(_08527_),
    .A2(net3231),
    .B(net2764),
    .Y(_08965_));
 OA21x2_ASAP7_75t_R _38286_ (.A1(net2764),
    .A2(_06099_),
    .B(_08965_),
    .Y(_08966_));
 AO21x1_ASAP7_75t_R _38287_ (.A1(_06196_),
    .A2(net3329),
    .B(net2399),
    .Y(_08967_));
 OA211x2_ASAP7_75t_R _38288_ (.A1(net2399),
    .A2(_06841_),
    .B(_07840_),
    .C(_08967_),
    .Y(_08968_));
 NAND2x1_ASAP7_75t_R _38289_ (.A(_08966_),
    .B(_08968_),
    .Y(_08969_));
 NAND2x1_ASAP7_75t_R _38290_ (.A(_06816_),
    .B(_06108_),
    .Y(_08970_));
 NAND2x1_ASAP7_75t_R _38291_ (.A(_08196_),
    .B(_06816_),
    .Y(_08971_));
 AO21x1_ASAP7_75t_R _38292_ (.A1(_06190_),
    .A2(_06226_),
    .B(_06064_),
    .Y(_08972_));
 AND4x1_ASAP7_75t_R _38293_ (.A(_07357_),
    .B(_08970_),
    .C(_08971_),
    .D(_08972_),
    .Y(_08973_));
 OA211x2_ASAP7_75t_R _38294_ (.A1(net1276),
    .A2(_06061_),
    .B(_07455_),
    .C(net2744),
    .Y(_08974_));
 AO21x1_ASAP7_75t_R _38295_ (.A1(_07455_),
    .A2(_06272_),
    .B(_06813_),
    .Y(_08976_));
 AO21x1_ASAP7_75t_R _38296_ (.A1(_07907_),
    .A2(_07455_),
    .B(_07822_),
    .Y(_08977_));
 NOR3x1_ASAP7_75t_R _38297_ (.A(_08974_),
    .B(_08976_),
    .C(_08977_),
    .Y(_08978_));
 NAND2x1_ASAP7_75t_R _38298_ (.A(_08973_),
    .B(_08978_),
    .Y(_08979_));
 NOR2x1_ASAP7_75t_R _38299_ (.A(_08969_),
    .B(_08979_),
    .Y(_08980_));
 AND2x4_ASAP7_75t_R _38300_ (.A(_08963_),
    .B(_08980_),
    .Y(_08981_));
 OA211x2_ASAP7_75t_R _38301_ (.A1(_06029_),
    .A2(_06061_),
    .B(_06251_),
    .C(net2507),
    .Y(_08982_));
 INVx1_ASAP7_75t_R _38302_ (.A(_08982_),
    .Y(_08983_));
 AO21x1_ASAP7_75t_R _38303_ (.A1(_06219_),
    .A2(_06070_),
    .B(_06268_),
    .Y(_08984_));
 AO21x1_ASAP7_75t_R _38304_ (.A1(_06118_),
    .A2(_06750_),
    .B(_06268_),
    .Y(_08985_));
 AND2x2_ASAP7_75t_R _38305_ (.A(_08984_),
    .B(_08985_),
    .Y(_08987_));
 AO21x1_ASAP7_75t_R _38306_ (.A1(_07475_),
    .A2(net3231),
    .B(_06250_),
    .Y(_08988_));
 NAND3x1_ASAP7_75t_R _38307_ (.A(_08983_),
    .B(_08987_),
    .C(_08988_),
    .Y(_08989_));
 INVx1_ASAP7_75t_R _38308_ (.A(_08989_),
    .Y(_08990_));
 AO21x1_ASAP7_75t_R _38309_ (.A1(_06078_),
    .A2(net2234),
    .B(_06240_),
    .Y(_08991_));
 AO21x1_ASAP7_75t_R _38310_ (.A1(net3330),
    .A2(_06196_),
    .B(_06240_),
    .Y(_08992_));
 NOR2x1_ASAP7_75t_R _38311_ (.A(_06240_),
    .B(net3328),
    .Y(_08993_));
 INVx1_ASAP7_75t_R _38312_ (.A(_08993_),
    .Y(_08994_));
 AND3x2_ASAP7_75t_R _38313_ (.A(_08991_),
    .B(_08992_),
    .C(_08994_),
    .Y(_08995_));
 AO21x1_ASAP7_75t_R _38314_ (.A1(_07475_),
    .A2(net3330),
    .B(net2412),
    .Y(_08996_));
 NAND2x1_ASAP7_75t_R _38315_ (.A(net3327),
    .B(_06775_),
    .Y(_08998_));
 AND2x2_ASAP7_75t_R _38316_ (.A(_08996_),
    .B(_08998_),
    .Y(_08999_));
 AO21x1_ASAP7_75t_R _38317_ (.A1(_06190_),
    .A2(net2590),
    .B(net2412),
    .Y(_09000_));
 AO21x1_ASAP7_75t_R _38318_ (.A1(net1260),
    .A2(_06181_),
    .B(net2412),
    .Y(_09001_));
 AND3x2_ASAP7_75t_R _38319_ (.A(_08999_),
    .B(_09000_),
    .C(_09001_),
    .Y(_09002_));
 NAND3x2_ASAP7_75t_R _38320_ (.B(_08995_),
    .C(_09002_),
    .Y(_09003_),
    .A(_08990_));
 NAND2x1_ASAP7_75t_R _38321_ (.A(_06208_),
    .B(_07876_),
    .Y(_09004_));
 NAND2x1_ASAP7_75t_R _38322_ (.A(net2756),
    .B(_06207_),
    .Y(_09005_));
 INVx1_ASAP7_75t_R _38323_ (.A(_09005_),
    .Y(_09006_));
 OR3x1_ASAP7_75t_R _38324_ (.A(_09004_),
    .B(_09006_),
    .C(_07323_),
    .Y(_09007_));
 OA21x2_ASAP7_75t_R _38325_ (.A1(_06193_),
    .A2(_06799_),
    .B(_06212_),
    .Y(_09009_));
 OA21x2_ASAP7_75t_R _38326_ (.A1(_07393_),
    .A2(net1600),
    .B(_06212_),
    .Y(_09010_));
 OR4x1_ASAP7_75t_R _38327_ (.A(_09009_),
    .B(_09010_),
    .C(_06220_),
    .D(_07885_),
    .Y(_09011_));
 NOR2x1_ASAP7_75t_R _38328_ (.A(_09007_),
    .B(_09011_),
    .Y(_09012_));
 OAI21x1_ASAP7_75t_R _38329_ (.A1(_06191_),
    .A2(_06853_),
    .B(_06192_),
    .Y(_09013_));
 OA31x2_ASAP7_75t_R _38330_ (.A1(_06270_),
    .A2(_07393_),
    .A3(_08525_),
    .B1(_06194_),
    .Y(_09014_));
 NOR2x1_ASAP7_75t_R _38331_ (.A(_09013_),
    .B(_09014_),
    .Y(_09015_));
 AO21x1_ASAP7_75t_R _38332_ (.A1(_06190_),
    .A2(_06794_),
    .B(_06176_),
    .Y(_09016_));
 AO21x1_ASAP7_75t_R _38333_ (.A1(_06196_),
    .A2(_06750_),
    .B(_06176_),
    .Y(_09017_));
 AND3x1_ASAP7_75t_R _38334_ (.A(_09015_),
    .B(_09016_),
    .C(_09017_),
    .Y(_09018_));
 NAND2x1_ASAP7_75t_R _38335_ (.A(_09012_),
    .B(_09018_),
    .Y(_09020_));
 NOR2x2_ASAP7_75t_R _38336_ (.A(_09003_),
    .B(_09020_),
    .Y(_09021_));
 NAND3x2_ASAP7_75t_R _38337_ (.B(_09021_),
    .C(_06920_),
    .Y(_09022_),
    .A(_08981_));
 OAI21x1_ASAP7_75t_R _38338_ (.A1(_05495_),
    .A2(_05669_),
    .B(_05684_),
    .Y(_09023_));
 AO21x1_ASAP7_75t_R _38339_ (.A1(_05605_),
    .A2(net2033),
    .B(_05683_),
    .Y(_09024_));
 NAND2x2_ASAP7_75t_R _38340_ (.A(_09023_),
    .B(_09024_),
    .Y(_09025_));
 AOI221x1_ASAP7_75t_R _38341_ (.A1(net2814),
    .A2(net3111),
    .B1(_05440_),
    .B2(_05457_),
    .C(_05677_),
    .Y(_09026_));
 NOR3x2_ASAP7_75t_R _38342_ (.B(_09026_),
    .C(_08752_),
    .Y(_09027_),
    .A(_09025_));
 AO21x1_ASAP7_75t_R _38343_ (.A1(net2698),
    .A2(net2401),
    .B(_06576_),
    .Y(_09028_));
 NAND2x1_ASAP7_75t_R _38344_ (.A(_05661_),
    .B(_07066_),
    .Y(_09029_));
 AND3x2_ASAP7_75t_R _38345_ (.A(_09028_),
    .B(_08760_),
    .C(_09029_),
    .Y(_09031_));
 AO21x1_ASAP7_75t_R _38346_ (.A1(net1772),
    .A2(_05503_),
    .B(_05654_),
    .Y(_09032_));
 AO21x1_ASAP7_75t_R _38347_ (.A1(_05462_),
    .A2(net2815),
    .B(_05654_),
    .Y(_09033_));
 NAND2x1_ASAP7_75t_R _38348_ (.A(_09032_),
    .B(_09033_),
    .Y(_09034_));
 AO21x1_ASAP7_75t_R _38349_ (.A1(_05598_),
    .A2(_05655_),
    .B(_07772_),
    .Y(_09035_));
 NOR2x2_ASAP7_75t_R _38350_ (.A(_09034_),
    .B(_09035_),
    .Y(_09036_));
 NAND3x2_ASAP7_75t_R _38351_ (.B(_09031_),
    .C(_09036_),
    .Y(_09037_),
    .A(_09027_));
 OA21x2_ASAP7_75t_R _38352_ (.A1(_05566_),
    .A2(_05561_),
    .B(_06613_),
    .Y(_09038_));
 AOI211x1_ASAP7_75t_R _38353_ (.A1(net3110),
    .A2(net1204),
    .B(_05616_),
    .C(_05457_),
    .Y(_09039_));
 NOR3x2_ASAP7_75t_R _38354_ (.B(_09039_),
    .C(_08347_),
    .Y(_09040_),
    .A(_09038_));
 INVx1_ASAP7_75t_R _38355_ (.A(_09040_),
    .Y(_09042_));
 OA21x2_ASAP7_75t_R _38356_ (.A1(_05664_),
    .A2(_05665_),
    .B(_05627_),
    .Y(_09043_));
 NOR2x2_ASAP7_75t_R _38357_ (.A(_07749_),
    .B(_09043_),
    .Y(_09044_));
 AOI211x1_ASAP7_75t_R _38358_ (.A1(net1313),
    .A2(net989),
    .B(_05626_),
    .C(net1670),
    .Y(_09045_));
 AOI21x1_ASAP7_75t_R _38359_ (.A1(_05642_),
    .A2(_05627_),
    .B(_09045_),
    .Y(_09046_));
 NAND2x1_ASAP7_75t_R _38360_ (.A(_09044_),
    .B(_09046_),
    .Y(_09047_));
 NOR2x1_ASAP7_75t_R _38361_ (.A(_09042_),
    .B(_09047_),
    .Y(_09048_));
 AOI21x1_ASAP7_75t_R _38362_ (.A1(_07919_),
    .A2(_05447_),
    .B(_05634_),
    .Y(_09049_));
 OAI21x1_ASAP7_75t_R _38363_ (.A1(_05495_),
    .A2(_05566_),
    .B(_06593_),
    .Y(_09050_));
 NAND2x1_ASAP7_75t_R _38364_ (.A(_07151_),
    .B(_09050_),
    .Y(_09051_));
 NOR2x1_ASAP7_75t_R _38365_ (.A(_09049_),
    .B(_09051_),
    .Y(_09053_));
 AOI211x1_ASAP7_75t_R _38366_ (.A1(net1000),
    .A2(net989),
    .B(_05640_),
    .C(net1666),
    .Y(_09054_));
 OA21x2_ASAP7_75t_R _38367_ (.A1(_05495_),
    .A2(_05566_),
    .B(_05647_),
    .Y(_09055_));
 NOR2x1_ASAP7_75t_R _38368_ (.A(_09054_),
    .B(_09055_),
    .Y(_09056_));
 AOI21x1_ASAP7_75t_R _38369_ (.A1(_05513_),
    .A2(_05648_),
    .B(_06590_),
    .Y(_09057_));
 NAND3x1_ASAP7_75t_R _38370_ (.A(_09053_),
    .B(_09056_),
    .C(_09057_),
    .Y(_09058_));
 INVx1_ASAP7_75t_R _38371_ (.A(_09058_),
    .Y(_09059_));
 NAND2x2_ASAP7_75t_R _38372_ (.A(_09059_),
    .B(_09048_),
    .Y(_09060_));
 NOR2x2_ASAP7_75t_R _38373_ (.A(_09037_),
    .B(_09060_),
    .Y(_09061_));
 AO21x1_ASAP7_75t_R _38374_ (.A1(_05447_),
    .A2(_06574_),
    .B(_05492_),
    .Y(_09062_));
 NAND2x1_ASAP7_75t_R _38375_ (.A(_05488_),
    .B(_09062_),
    .Y(_09064_));
 INVx1_ASAP7_75t_R _38376_ (.A(_09064_),
    .Y(_09065_));
 OA21x2_ASAP7_75t_R _38377_ (.A1(_05646_),
    .A2(_05441_),
    .B(net3373),
    .Y(_09066_));
 OA21x2_ASAP7_75t_R _38378_ (.A1(_06637_),
    .A2(_05656_),
    .B(net3373),
    .Y(_09067_));
 NOR2x2_ASAP7_75t_R _38379_ (.A(_09066_),
    .B(_09067_),
    .Y(_09068_));
 OA21x2_ASAP7_75t_R _38380_ (.A1(_07066_),
    .A2(_05561_),
    .B(_05484_),
    .Y(_09069_));
 OA21x2_ASAP7_75t_R _38381_ (.A1(_07152_),
    .A2(_05656_),
    .B(_05484_),
    .Y(_09070_));
 NOR2x2_ASAP7_75t_R _38382_ (.A(_09069_),
    .B(_09070_),
    .Y(_09071_));
 NAND3x2_ASAP7_75t_R _38383_ (.B(_09068_),
    .C(_09071_),
    .Y(_09072_),
    .A(_09065_));
 AOI211x1_ASAP7_75t_R _38384_ (.A1(net3110),
    .A2(net989),
    .B(net2755),
    .C(net1672),
    .Y(_09073_));
 AOI21x1_ASAP7_75t_R _38385_ (.A1(_06627_),
    .A2(_05568_),
    .B(_09073_),
    .Y(_09075_));
 AO21x1_ASAP7_75t_R _38386_ (.A1(_05447_),
    .A2(_05580_),
    .B(_05548_),
    .Y(_09076_));
 AO21x1_ASAP7_75t_R _38387_ (.A1(_05503_),
    .A2(net1213),
    .B(_05548_),
    .Y(_09077_));
 AND2x2_ASAP7_75t_R _38388_ (.A(_09076_),
    .B(_09077_),
    .Y(_09078_));
 INVx1_ASAP7_75t_R _38389_ (.A(_07947_),
    .Y(_09079_));
 NOR2x2_ASAP7_75t_R _38390_ (.A(_06631_),
    .B(_09079_),
    .Y(_09080_));
 NAND3x2_ASAP7_75t_R _38391_ (.B(_09078_),
    .C(_09080_),
    .Y(_09081_),
    .A(_09075_));
 NOR2x2_ASAP7_75t_R _38392_ (.A(_09072_),
    .B(_09081_),
    .Y(_09082_));
 INVx2_ASAP7_75t_R _38393_ (.A(_09082_),
    .Y(_09083_));
 NAND2x1_ASAP7_75t_R _38394_ (.A(_08701_),
    .B(_06668_),
    .Y(_09084_));
 AO21x1_ASAP7_75t_R _38395_ (.A1(_05579_),
    .A2(net2035),
    .B(net2389),
    .Y(_09086_));
 OAI21x1_ASAP7_75t_R _38396_ (.A1(net2389),
    .A2(_05605_),
    .B(_09086_),
    .Y(_09087_));
 NOR2x1_ASAP7_75t_R _38397_ (.A(_09084_),
    .B(_09087_),
    .Y(_09088_));
 NAND2x1_ASAP7_75t_R _38398_ (.A(_07700_),
    .B(_05578_),
    .Y(_09089_));
 NOR3x1_ASAP7_75t_R _38399_ (.A(_09089_),
    .B(_05586_),
    .C(_08704_),
    .Y(_09090_));
 NAND2x1_ASAP7_75t_R _38400_ (.A(_09088_),
    .B(_09090_),
    .Y(_09091_));
 INVx1_ASAP7_75t_R _38401_ (.A(_09091_),
    .Y(_09092_));
 AOI211x1_ASAP7_75t_R _38402_ (.A1(net3110),
    .A2(_05500_),
    .B(_05453_),
    .C(_05457_),
    .Y(_09093_));
 INVx1_ASAP7_75t_R _38403_ (.A(_09093_),
    .Y(_09094_));
 AO21x1_ASAP7_75t_R _38404_ (.A1(net3249),
    .A2(_05503_),
    .B(_05453_),
    .Y(_09095_));
 AND2x2_ASAP7_75t_R _38405_ (.A(_09094_),
    .B(_09095_),
    .Y(_09097_));
 INVx1_ASAP7_75t_R _38406_ (.A(_09097_),
    .Y(_09098_));
 AOI211x1_ASAP7_75t_R _38407_ (.A1(net3110),
    .A2(net989),
    .B(_05472_),
    .C(_05457_),
    .Y(_09099_));
 NOR2x2_ASAP7_75t_R _38408_ (.A(_05599_),
    .B(_09099_),
    .Y(_09100_));
 AO21x1_ASAP7_75t_R _38409_ (.A1(_05613_),
    .A2(_05496_),
    .B(_05472_),
    .Y(_09101_));
 OA21x2_ASAP7_75t_R _38410_ (.A1(_07760_),
    .A2(_05601_),
    .B(_09101_),
    .Y(_09102_));
 NAND2x1_ASAP7_75t_R _38411_ (.A(_09100_),
    .B(_09102_),
    .Y(_09103_));
 NOR2x1_ASAP7_75t_R _38412_ (.A(_09098_),
    .B(_09103_),
    .Y(_09104_));
 NAND2x1_ASAP7_75t_R _38413_ (.A(_09092_),
    .B(_09104_),
    .Y(_09105_));
 NOR2x2_ASAP7_75t_R _38414_ (.A(_09083_),
    .B(_09105_),
    .Y(_09106_));
 NAND2x2_ASAP7_75t_R _38415_ (.A(_09061_),
    .B(_09106_),
    .Y(_09108_));
 XOR2x2_ASAP7_75t_R _38416_ (.A(_09108_),
    .B(_05427_),
    .Y(_09109_));
 XOR2x2_ASAP7_75t_R _38417_ (.A(_09022_),
    .B(_09109_),
    .Y(_09110_));
 NAND2x1_ASAP7_75t_R _38418_ (.A(_08949_),
    .B(_09110_),
    .Y(_09111_));
 INVx2_ASAP7_75t_R _38419_ (.A(_09110_),
    .Y(_09112_));
 NAND2x1_ASAP7_75t_R _38420_ (.A(_08948_),
    .B(_09112_),
    .Y(_09113_));
 NAND2x1_ASAP7_75t_R _38421_ (.A(_09111_),
    .B(_09113_),
    .Y(_09114_));
 NOR2x1_ASAP7_75t_R _38422_ (.A(net394),
    .B(_00844_),
    .Y(_09115_));
 AOI21x1_ASAP7_75t_R _38423_ (.A1(net394),
    .A2(_09114_),
    .B(_09115_),
    .Y(_09116_));
 XOR2x1_ASAP7_75t_R _38424_ (.A(_09116_),
    .Y(_00112_),
    .B(_00388_));
 NAND2x1_ASAP7_75t_R _38425_ (.A(_00843_),
    .B(net388),
    .Y(_09118_));
 XOR2x1_ASAP7_75t_R _38426_ (.A(_06913_),
    .Y(_09119_),
    .B(net1964));
 OAI21x1_ASAP7_75t_R _38427_ (.A1(_06290_),
    .A2(_06291_),
    .B(_09119_),
    .Y(_09120_));
 XOR2x1_ASAP7_75t_R _38428_ (.A(_06913_),
    .Y(_09121_),
    .B(_08947_));
 OAI21x1_ASAP7_75t_R _38429_ (.A1(_06294_),
    .A2(_06295_),
    .B(_09121_),
    .Y(_09122_));
 AO21x1_ASAP7_75t_R _38430_ (.A1(_09120_),
    .A2(_09122_),
    .B(net388),
    .Y(_09123_));
 AOI21x1_ASAP7_75t_R _38431_ (.A1(_09118_),
    .A2(_09123_),
    .B(_14603_),
    .Y(_09124_));
 AOI21x1_ASAP7_75t_R _38432_ (.A1(_09120_),
    .A2(_09122_),
    .B(net388),
    .Y(_09125_));
 AND2x2_ASAP7_75t_R _38433_ (.A(net388),
    .B(_00843_),
    .Y(_09126_));
 NOR3x2_ASAP7_75t_R _38434_ (.B(_00496_),
    .C(_09126_),
    .Y(_09127_),
    .A(_09125_));
 NOR2x2_ASAP7_75t_R _38435_ (.A(_09127_),
    .B(_09124_),
    .Y(_00073_));
 TAPCELL_ASAP7_75t_R PHY_286 ();
 AND2x2_ASAP7_75t_R _38437_ (.A(net388),
    .B(_00842_),
    .Y(_09130_));
 AOI21x1_ASAP7_75t_R _38438_ (.A1(net1978),
    .A2(_06025_),
    .B(_08946_),
    .Y(_09131_));
 INVx1_ASAP7_75t_R _38439_ (.A(_09131_),
    .Y(_09132_));
 NAND3x2_ASAP7_75t_R _38440_ (.B(net2305),
    .C(net1978),
    .Y(_09133_),
    .A(_06025_));
 NAND2x2_ASAP7_75t_R _38441_ (.A(_09132_),
    .B(_09133_),
    .Y(_09134_));
 XOR2x2_ASAP7_75t_R _38442_ (.A(net3435),
    .B(_06679_),
    .Y(_09135_));
 NOR2x2_ASAP7_75t_R _38443_ (.A(_09134_),
    .B(_09135_),
    .Y(_09136_));
 XOR2x2_ASAP7_75t_R _38444_ (.A(net3435),
    .B(net1927),
    .Y(_09137_));
 INVx3_ASAP7_75t_R _38445_ (.A(_09134_),
    .Y(_09139_));
 NOR2x1_ASAP7_75t_R _38446_ (.A(_09137_),
    .B(_09139_),
    .Y(_09140_));
 INVx1_ASAP7_75t_R _38447_ (.A(_07381_),
    .Y(_09141_));
 XOR2x2_ASAP7_75t_R _38448_ (.A(_06913_),
    .B(_09141_),
    .Y(_09142_));
 OAI21x1_ASAP7_75t_R _38449_ (.A1(_09136_),
    .A2(_09140_),
    .B(_09142_),
    .Y(_09143_));
 NOR2x2_ASAP7_75t_R _38450_ (.A(_09134_),
    .B(_09137_),
    .Y(_09144_));
 NOR2x1_ASAP7_75t_R _38451_ (.A(_09135_),
    .B(_09139_),
    .Y(_09145_));
 INVx2_ASAP7_75t_R _38452_ (.A(_09142_),
    .Y(_09146_));
 OAI21x1_ASAP7_75t_R _38453_ (.A1(_09144_),
    .A2(_09145_),
    .B(_09146_),
    .Y(_09147_));
 AOI21x1_ASAP7_75t_R _38454_ (.A1(_09143_),
    .A2(_09147_),
    .B(net388),
    .Y(_09148_));
 OAI21x1_ASAP7_75t_R _38455_ (.A1(_09130_),
    .A2(_09148_),
    .B(_17184_),
    .Y(_09150_));
 NOR2x1_ASAP7_75t_R _38456_ (.A(net394),
    .B(_00842_),
    .Y(_09151_));
 OAI21x1_ASAP7_75t_R _38457_ (.A1(_09144_),
    .A2(_09145_),
    .B(_09142_),
    .Y(_09152_));
 OAI21x1_ASAP7_75t_R _38458_ (.A1(_09136_),
    .A2(_09140_),
    .B(_09146_),
    .Y(_09153_));
 TAPCELL_ASAP7_75t_R PHY_285 ();
 AOI21x1_ASAP7_75t_R _38460_ (.A1(_09152_),
    .A2(_09153_),
    .B(net388),
    .Y(_09155_));
 OAI21x1_ASAP7_75t_R _38461_ (.A1(_09151_),
    .A2(_09155_),
    .B(_00495_),
    .Y(_09156_));
 NAND2x2_ASAP7_75t_R _38462_ (.A(_09156_),
    .B(_09150_),
    .Y(_00074_));
 AND2x2_ASAP7_75t_R _38463_ (.A(net388),
    .B(_00841_),
    .Y(_09157_));
 INVx3_ASAP7_75t_R _38464_ (.A(net3382),
    .Y(_09158_));
 AOI21x1_ASAP7_75t_R _38465_ (.A1(_07160_),
    .A2(_07167_),
    .B(_09158_),
    .Y(_09160_));
 AOI21x1_ASAP7_75t_R _38466_ (.A1(_07274_),
    .A2(_07275_),
    .B(net3383),
    .Y(_09161_));
 XOR2x2_ASAP7_75t_R _38467_ (.A(_07381_),
    .B(_06697_),
    .Y(_09162_));
 OAI21x1_ASAP7_75t_R _38468_ (.A1(_09160_),
    .A2(_09161_),
    .B(_09162_),
    .Y(_09163_));
 AOI21x1_ASAP7_75t_R _38469_ (.A1(_07160_),
    .A2(_07167_),
    .B(net3383),
    .Y(_09164_));
 AOI21x1_ASAP7_75t_R _38470_ (.A1(_07274_),
    .A2(_07275_),
    .B(_09158_),
    .Y(_09165_));
 XOR2x2_ASAP7_75t_R _38471_ (.A(_07381_),
    .B(_06552_),
    .Y(_09166_));
 OAI21x1_ASAP7_75t_R _38472_ (.A1(_09164_),
    .A2(_09165_),
    .B(_09166_),
    .Y(_09167_));
 AOI21x1_ASAP7_75t_R _38473_ (.A1(_09163_),
    .A2(_09167_),
    .B(net388),
    .Y(_09168_));
 NOR2x1_ASAP7_75t_R _38474_ (.A(_09157_),
    .B(_09168_),
    .Y(_09169_));
 XNOR2x2_ASAP7_75t_R _38475_ (.A(_00389_),
    .B(_09169_),
    .Y(_00075_));
 XOR2x1_ASAP7_75t_R _38476_ (.A(_07500_),
    .Y(_09171_),
    .B(_07917_));
 XNOR2x2_ASAP7_75t_R _38477_ (.A(_08946_),
    .B(_07271_),
    .Y(_09172_));
 XOR2x1_ASAP7_75t_R _38478_ (.A(_07807_),
    .Y(_09173_),
    .B(_09172_));
 XOR2x2_ASAP7_75t_R _38479_ (.A(_09171_),
    .B(_09173_),
    .Y(_09174_));
 NOR2x2_ASAP7_75t_R _38480_ (.A(net391),
    .B(_00840_),
    .Y(_09175_));
 AOI21x1_ASAP7_75t_R _38481_ (.A1(net391),
    .A2(_09174_),
    .B(_09175_),
    .Y(_09176_));
 XOR2x1_ASAP7_75t_R _38482_ (.A(_09176_),
    .Y(_00076_),
    .B(_00390_));
 TAPCELL_ASAP7_75t_R PHY_284 ();
 NOR2x1_ASAP7_75t_R _38484_ (.A(net391),
    .B(_00839_),
    .Y(_09178_));
 INVx1_ASAP7_75t_R _38485_ (.A(_08222_),
    .Y(_09180_));
 NAND2x1_ASAP7_75t_R _38486_ (.A(_08233_),
    .B(_08206_),
    .Y(_09181_));
 NOR2x2_ASAP7_75t_R _38487_ (.A(_09180_),
    .B(_09181_),
    .Y(_09182_));
 INVx1_ASAP7_75t_R _38488_ (.A(_08250_),
    .Y(_09183_));
 NAND2x1_ASAP7_75t_R _38489_ (.A(_08264_),
    .B(_08240_),
    .Y(_09184_));
 NOR2x1_ASAP7_75t_R _38490_ (.A(_09183_),
    .B(_09184_),
    .Y(_09185_));
 NAND2x2_ASAP7_75t_R _38491_ (.A(_09182_),
    .B(_09185_),
    .Y(_09186_));
 XOR2x1_ASAP7_75t_R _38492_ (.A(_07918_),
    .Y(_09187_),
    .B(_09186_));
 XOR2x2_ASAP7_75t_R _38493_ (.A(_07593_),
    .B(_08947_),
    .Y(_09188_));
 XOR2x2_ASAP7_75t_R _38494_ (.A(_08005_),
    .B(_08169_),
    .Y(_09189_));
 XOR2x1_ASAP7_75t_R _38495_ (.A(_09188_),
    .Y(_09191_),
    .B(_09189_));
 NOR2x1_ASAP7_75t_R _38496_ (.A(_09187_),
    .B(_09191_),
    .Y(_09192_));
 XOR2x1_ASAP7_75t_R _38497_ (.A(_07918_),
    .Y(_09193_),
    .B(_08266_));
 XNOR2x1_ASAP7_75t_R _38498_ (.B(_09188_),
    .Y(_09194_),
    .A(_09189_));
 NOR2x1_ASAP7_75t_R _38499_ (.A(_09193_),
    .B(_09194_),
    .Y(_09195_));
 OAI21x1_ASAP7_75t_R _38500_ (.A1(_09192_),
    .A2(_09195_),
    .B(_00528_),
    .Y(_09196_));
 INVx1_ASAP7_75t_R _38501_ (.A(_09196_),
    .Y(_09197_));
 OAI21x1_ASAP7_75t_R _38502_ (.A1(_09178_),
    .A2(_09197_),
    .B(_00391_),
    .Y(_09198_));
 INVx1_ASAP7_75t_R _38503_ (.A(_09178_),
    .Y(_09199_));
 NAND3x1_ASAP7_75t_R _38504_ (.A(_09196_),
    .B(_17199_),
    .C(_09199_),
    .Y(_09200_));
 NAND2x1_ASAP7_75t_R _38505_ (.A(_09200_),
    .B(_09198_),
    .Y(_00077_));
 NOR2x2_ASAP7_75t_R _38506_ (.A(_00528_),
    .B(_00838_),
    .Y(_09202_));
 XOR2x2_ASAP7_75t_R _38507_ (.A(_08266_),
    .B(_08086_),
    .Y(_09203_));
 NAND2x1_ASAP7_75t_R _38508_ (.A(_08601_),
    .B(_09203_),
    .Y(_09204_));
 NAND2x1_ASAP7_75t_R _38509_ (.A(_08086_),
    .B(_08266_),
    .Y(_09205_));
 OAI22x1_ASAP7_75t_R _38510_ (.A1(_08265_),
    .A2(_08234_),
    .B1(_08085_),
    .B2(_08048_),
    .Y(_09206_));
 AO21x1_ASAP7_75t_R _38511_ (.A1(_09205_),
    .A2(_09206_),
    .B(_08601_),
    .Y(_09207_));
 AOI21x1_ASAP7_75t_R _38512_ (.A1(_09204_),
    .A2(_09207_),
    .B(_08519_),
    .Y(_09208_));
 NOR2x1_ASAP7_75t_R _38513_ (.A(_08508_),
    .B(_08504_),
    .Y(_09209_));
 NOR2x1_ASAP7_75t_R _38514_ (.A(net1860),
    .B(_08517_),
    .Y(_09210_));
 NOR2x1_ASAP7_75t_R _38515_ (.A(_09209_),
    .B(_09210_),
    .Y(_09212_));
 NAND3x2_ASAP7_75t_R _38516_ (.B(_08599_),
    .C(_08563_),
    .Y(_09213_),
    .A(net2156));
 XOR2x1_ASAP7_75t_R _38517_ (.A(_09203_),
    .Y(_09214_),
    .B(_09213_));
 NOR2x1_ASAP7_75t_R _38518_ (.A(_09212_),
    .B(_09214_),
    .Y(_09215_));
 OAI21x1_ASAP7_75t_R _38519_ (.A1(_09208_),
    .A2(_09215_),
    .B(net394),
    .Y(_09216_));
 INVx1_ASAP7_75t_R _38520_ (.A(_09216_),
    .Y(_09217_));
 OAI21x1_ASAP7_75t_R _38521_ (.A1(_09202_),
    .A2(_09217_),
    .B(_00494_),
    .Y(_09218_));
 INVx1_ASAP7_75t_R _38522_ (.A(_09202_),
    .Y(_09219_));
 NAND3x1_ASAP7_75t_R _38523_ (.A(_09216_),
    .B(_17206_),
    .C(_09219_),
    .Y(_09220_));
 NAND2x1_ASAP7_75t_R _38524_ (.A(_09220_),
    .B(_09218_),
    .Y(_00078_));
 AND2x2_ASAP7_75t_R _38525_ (.A(net388),
    .B(_00837_),
    .Y(_09222_));
 NAND3x2_ASAP7_75t_R _38526_ (.B(_08336_),
    .C(_08304_),
    .Y(_09223_),
    .A(_05794_));
 NOR2x2_ASAP7_75t_R _38527_ (.A(_09223_),
    .B(_09213_),
    .Y(_09224_));
 NOR2x2_ASAP7_75t_R _38528_ (.A(_08601_),
    .B(net2774),
    .Y(_09225_));
 NAND2x2_ASAP7_75t_R _38529_ (.A(_09021_),
    .B(_08981_),
    .Y(_09226_));
 NOR2x2_ASAP7_75t_R _38530_ (.A(_06890_),
    .B(_09226_),
    .Y(_09227_));
 OA21x2_ASAP7_75t_R _38531_ (.A1(_09224_),
    .A2(_09225_),
    .B(_09227_),
    .Y(_09228_));
 NOR2x2_ASAP7_75t_R _38532_ (.A(_09213_),
    .B(net2774),
    .Y(_09229_));
 NOR2x2_ASAP7_75t_R _38533_ (.A(_08601_),
    .B(_09223_),
    .Y(_09230_));
 OA21x2_ASAP7_75t_R _38534_ (.A1(_09229_),
    .A2(_09230_),
    .B(_09022_),
    .Y(_09231_));
 OAI21x1_ASAP7_75t_R _38535_ (.A1(_09228_),
    .A2(_09231_),
    .B(net3347),
    .Y(_09233_));
 OA21x2_ASAP7_75t_R _38536_ (.A1(_09224_),
    .A2(_09225_),
    .B(_09022_),
    .Y(_09234_));
 OA21x2_ASAP7_75t_R _38537_ (.A1(_09229_),
    .A2(_09230_),
    .B(_09227_),
    .Y(_09235_));
 OAI21x1_ASAP7_75t_R _38538_ (.A1(_09234_),
    .A2(_09235_),
    .B(_08860_),
    .Y(_09236_));
 TAPCELL_ASAP7_75t_R PHY_283 ();
 AOI21x1_ASAP7_75t_R _38540_ (.A1(_09233_),
    .A2(_09236_),
    .B(net388),
    .Y(_09238_));
 OAI21x1_ASAP7_75t_R _38541_ (.A1(_09222_),
    .A2(_09238_),
    .B(_17214_),
    .Y(_09239_));
 NOR2x1_ASAP7_75t_R _38542_ (.A(net394),
    .B(_00837_),
    .Y(_09240_));
 OAI21x1_ASAP7_75t_R _38543_ (.A1(_09228_),
    .A2(_09231_),
    .B(_08860_),
    .Y(_09241_));
 OAI21x1_ASAP7_75t_R _38544_ (.A1(_09234_),
    .A2(_09235_),
    .B(net3347),
    .Y(_09242_));
 AOI21x1_ASAP7_75t_R _38545_ (.A1(_09241_),
    .A2(_09242_),
    .B(net388),
    .Y(_09244_));
 OAI21x1_ASAP7_75t_R _38546_ (.A1(_09240_),
    .A2(_09244_),
    .B(_00493_),
    .Y(_09245_));
 NAND2x1_ASAP7_75t_R _38547_ (.A(_09239_),
    .B(_09245_),
    .Y(_00079_));
 AND2x2_ASAP7_75t_R _38548_ (.A(net388),
    .B(_00836_),
    .Y(_09246_));
 XOR2x2_ASAP7_75t_R _38549_ (.A(_08853_),
    .B(_06729_),
    .Y(_09247_));
 NAND2x1_ASAP7_75t_R _38550_ (.A(_09247_),
    .B(_09110_),
    .Y(_09248_));
 XOR2x2_ASAP7_75t_R _38551_ (.A(_08853_),
    .B(_06286_),
    .Y(_09249_));
 NAND2x1_ASAP7_75t_R _38552_ (.A(_09112_),
    .B(_09249_),
    .Y(_09250_));
 AOI21x1_ASAP7_75t_R _38553_ (.A1(_09248_),
    .A2(_09250_),
    .B(net388),
    .Y(_09251_));
 OAI21x1_ASAP7_75t_R _38554_ (.A1(_09246_),
    .A2(_09251_),
    .B(_17220_),
    .Y(_09252_));
 NOR2x1_ASAP7_75t_R _38555_ (.A(_09246_),
    .B(_09251_),
    .Y(_09254_));
 NAND2x1_ASAP7_75t_R _38556_ (.A(_00392_),
    .B(_09254_),
    .Y(_09255_));
 NAND2x1_ASAP7_75t_R _38557_ (.A(_09255_),
    .B(_09252_),
    .Y(_00080_));
 NOR2x1_ASAP7_75t_R _38558_ (.A(net394),
    .B(_00835_),
    .Y(_09256_));
 INVx1_ASAP7_75t_R _38559_ (.A(_09256_),
    .Y(_09257_));
 NAND3x1_ASAP7_75t_R _38560_ (.A(_09097_),
    .B(_09102_),
    .C(_09100_),
    .Y(_09258_));
 NOR2x1_ASAP7_75t_R _38561_ (.A(_09091_),
    .B(_09258_),
    .Y(_09259_));
 NAND2x2_ASAP7_75t_R _38562_ (.A(_09082_),
    .B(_09259_),
    .Y(_09260_));
 INVx1_ASAP7_75t_R _38563_ (.A(_09027_),
    .Y(_09261_));
 NAND2x1_ASAP7_75t_R _38564_ (.A(_09031_),
    .B(_09036_),
    .Y(_09262_));
 NOR2x1_ASAP7_75t_R _38565_ (.A(_09261_),
    .B(_09262_),
    .Y(_09264_));
 NAND3x1_ASAP7_75t_R _38566_ (.A(_09040_),
    .B(_09046_),
    .C(_09044_),
    .Y(_09265_));
 NOR2x1_ASAP7_75t_R _38567_ (.A(_09058_),
    .B(_09265_),
    .Y(_09266_));
 NAND2x1_ASAP7_75t_R _38568_ (.A(_09264_),
    .B(_09266_),
    .Y(_09267_));
 NOR2x2_ASAP7_75t_R _38569_ (.A(_09260_),
    .B(_09267_),
    .Y(_09268_));
 NAND2x1_ASAP7_75t_R _38570_ (.A(_09268_),
    .B(_05728_),
    .Y(_09269_));
 AO21x1_ASAP7_75t_R _38571_ (.A1(_05317_),
    .A2(net3428),
    .B(_09268_),
    .Y(_09270_));
 NAND2x2_ASAP7_75t_R _38572_ (.A(_06920_),
    .B(_06876_),
    .Y(_09271_));
 NAND3x1_ASAP7_75t_R _38573_ (.A(_09269_),
    .B(_09270_),
    .C(_09271_),
    .Y(_09272_));
 AO21x1_ASAP7_75t_R _38574_ (.A1(_09269_),
    .A2(_09270_),
    .B(_09271_),
    .Y(_09273_));
 AOI21x1_ASAP7_75t_R _38575_ (.A1(_09272_),
    .A2(_09273_),
    .B(_09139_),
    .Y(_09275_));
 TAPCELL_ASAP7_75t_R PHY_282 ();
 XOR2x1_ASAP7_75t_R _38577_ (.A(_05728_),
    .Y(_09277_),
    .B(_09271_));
 NAND2x1_ASAP7_75t_R _38578_ (.A(_09108_),
    .B(_09277_),
    .Y(_09278_));
 XNOR2x1_ASAP7_75t_R _38579_ (.B(_05728_),
    .Y(_09279_),
    .A(_09271_));
 NAND2x1_ASAP7_75t_R _38580_ (.A(_09268_),
    .B(_09279_),
    .Y(_09280_));
 AOI21x1_ASAP7_75t_R _38581_ (.A1(_09278_),
    .A2(_09280_),
    .B(_09134_),
    .Y(_09281_));
 OAI21x1_ASAP7_75t_R _38582_ (.A1(_09275_),
    .A2(_09281_),
    .B(net394),
    .Y(_09282_));
 NAND2x1_ASAP7_75t_R _38583_ (.A(_09257_),
    .B(_09282_),
    .Y(_09283_));
 INVx3_ASAP7_75t_R _38584_ (.A(_00492_),
    .Y(_09284_));
 XOR2x2_ASAP7_75t_R _38585_ (.A(_09283_),
    .B(_09284_),
    .Y(_00041_));
 AND2x2_ASAP7_75t_R _38586_ (.A(net388),
    .B(_00834_),
    .Y(_09286_));
 NOR2x1_ASAP7_75t_R _38587_ (.A(_09166_),
    .B(_09134_),
    .Y(_09287_));
 NOR2x1_ASAP7_75t_R _38588_ (.A(_09162_),
    .B(_09139_),
    .Y(_09288_));
 AO21x2_ASAP7_75t_R _38589_ (.A1(_05692_),
    .A2(_05479_),
    .B(_09108_),
    .Y(_09289_));
 NAND3x2_ASAP7_75t_R _38590_ (.B(_09108_),
    .C(net2350),
    .Y(_09290_),
    .A(_05692_));
 AOI21x1_ASAP7_75t_R _38591_ (.A1(_09289_),
    .A2(_09290_),
    .B(_06422_),
    .Y(_09291_));
 AO21x2_ASAP7_75t_R _38592_ (.A1(_05692_),
    .A2(_05479_),
    .B(_09268_),
    .Y(_09292_));
 NAND3x2_ASAP7_75t_R _38593_ (.B(_09268_),
    .C(_05479_),
    .Y(_09293_),
    .A(_05692_));
 AOI21x1_ASAP7_75t_R _38594_ (.A1(_09292_),
    .A2(_09293_),
    .B(net3435),
    .Y(_09294_));
 NOR2x2_ASAP7_75t_R _38595_ (.A(_09291_),
    .B(_09294_),
    .Y(_09296_));
 OAI21x1_ASAP7_75t_R _38596_ (.A1(_09287_),
    .A2(_09288_),
    .B(_09296_),
    .Y(_09297_));
 INVx1_ASAP7_75t_R _38597_ (.A(_09296_),
    .Y(_09298_));
 XOR2x1_ASAP7_75t_R _38598_ (.A(_09134_),
    .Y(_09299_),
    .B(_09166_));
 NAND2x1_ASAP7_75t_R _38599_ (.A(_09299_),
    .B(_09298_),
    .Y(_09300_));
 AOI21x1_ASAP7_75t_R _38600_ (.A1(_09297_),
    .A2(_09300_),
    .B(net388),
    .Y(_09301_));
 INVx1_ASAP7_75t_R _38601_ (.A(_00491_),
    .Y(_09302_));
 OAI21x1_ASAP7_75t_R _38602_ (.A1(_09286_),
    .A2(_09301_),
    .B(_09302_),
    .Y(_09303_));
 NOR2x1_ASAP7_75t_R _38603_ (.A(net394),
    .B(_00834_),
    .Y(_09304_));
 NAND2x2_ASAP7_75t_R _38604_ (.A(_09289_),
    .B(_09290_),
    .Y(_09305_));
 NOR2x1_ASAP7_75t_R _38605_ (.A(_09162_),
    .B(_09305_),
    .Y(_09307_));
 NAND2x2_ASAP7_75t_R _38606_ (.A(_09292_),
    .B(_09293_),
    .Y(_09308_));
 NOR2x1_ASAP7_75t_R _38607_ (.A(_09166_),
    .B(_09308_),
    .Y(_09309_));
 NOR2x1_ASAP7_75t_R _38608_ (.A(_06025_),
    .B(_08947_),
    .Y(_09310_));
 NOR2x1_ASAP7_75t_R _38609_ (.A(net1964),
    .B(_06026_),
    .Y(_09311_));
 OAI21x1_ASAP7_75t_R _38610_ (.A1(_09310_),
    .A2(_09311_),
    .B(net3419),
    .Y(_09312_));
 INVx1_ASAP7_75t_R _38611_ (.A(_09133_),
    .Y(_09313_));
 OAI21x1_ASAP7_75t_R _38612_ (.A1(_09131_),
    .A2(_09313_),
    .B(_06422_),
    .Y(_09314_));
 NAND2x2_ASAP7_75t_R _38613_ (.A(_09312_),
    .B(_09314_),
    .Y(_09315_));
 OAI21x1_ASAP7_75t_R _38614_ (.A1(_09307_),
    .A2(_09309_),
    .B(_09315_),
    .Y(_09316_));
 XOR2x1_ASAP7_75t_R _38615_ (.A(_09305_),
    .Y(_09318_),
    .B(_09162_));
 INVx1_ASAP7_75t_R _38616_ (.A(_09315_),
    .Y(_09319_));
 NAND2x1_ASAP7_75t_R _38617_ (.A(_09318_),
    .B(_09319_),
    .Y(_09320_));
 AOI21x1_ASAP7_75t_R _38618_ (.A1(_09316_),
    .A2(_09320_),
    .B(net388),
    .Y(_09321_));
 OAI21x1_ASAP7_75t_R _38619_ (.A1(_09304_),
    .A2(_09321_),
    .B(_00491_),
    .Y(_09322_));
 NAND2x2_ASAP7_75t_R _38620_ (.A(_09322_),
    .B(_09303_),
    .Y(_00042_));
 NOR2x1_ASAP7_75t_R _38621_ (.A(_00528_),
    .B(_00833_),
    .Y(_09323_));
 XOR2x2_ASAP7_75t_R _38622_ (.A(_06697_),
    .B(net1927),
    .Y(_09324_));
 XNOR2x2_ASAP7_75t_R _38623_ (.A(_07271_),
    .B(_07049_),
    .Y(_09325_));
 XOR2x1_ASAP7_75t_R _38624_ (.A(_09325_),
    .Y(_09326_),
    .B(net3382));
 NOR2x1_ASAP7_75t_R _38625_ (.A(_09324_),
    .B(_09326_),
    .Y(_09328_));
 INVx2_ASAP7_75t_R _38626_ (.A(_09324_),
    .Y(_09329_));
 XOR2x1_ASAP7_75t_R _38627_ (.A(_09325_),
    .Y(_09330_),
    .B(_09158_));
 NOR2x1_ASAP7_75t_R _38628_ (.A(_09329_),
    .B(_09330_),
    .Y(_09331_));
 OAI21x1_ASAP7_75t_R _38629_ (.A1(_09328_),
    .A2(_09331_),
    .B(net394),
    .Y(_09332_));
 INVx1_ASAP7_75t_R _38630_ (.A(_09332_),
    .Y(_09333_));
 OAI21x1_ASAP7_75t_R _38631_ (.A1(_09323_),
    .A2(_09333_),
    .B(_00393_),
    .Y(_09334_));
 INVx1_ASAP7_75t_R _38632_ (.A(_09323_),
    .Y(_09335_));
 NAND3x2_ASAP7_75t_R _38633_ (.B(_17369_),
    .C(_09335_),
    .Y(_09336_),
    .A(_09332_));
 NAND2x2_ASAP7_75t_R _38634_ (.A(_09334_),
    .B(_09336_),
    .Y(_00043_));
 AND2x2_ASAP7_75t_R _38635_ (.A(net388),
    .B(_00832_),
    .Y(_09338_));
 XNOR2x2_ASAP7_75t_R _38636_ (.A(_07917_),
    .B(_07593_),
    .Y(_09339_));
 NOR2x2_ASAP7_75t_R _38637_ (.A(_09172_),
    .B(_09339_),
    .Y(_09340_));
 AND2x4_ASAP7_75t_R _38638_ (.A(_09339_),
    .B(_09172_),
    .Y(_09341_));
 NOR2x2_ASAP7_75t_R _38639_ (.A(_09268_),
    .B(net3420),
    .Y(_09342_));
 NOR2x2_ASAP7_75t_R _38640_ (.A(net1739),
    .B(_07165_),
    .Y(_09343_));
 OAI21x1_ASAP7_75t_R _38641_ (.A1(_09342_),
    .A2(_09343_),
    .B(_07697_),
    .Y(_09344_));
 NOR2x2_ASAP7_75t_R _38642_ (.A(net1739),
    .B(net3420),
    .Y(_09345_));
 NOR2x2_ASAP7_75t_R _38643_ (.A(_09268_),
    .B(_07165_),
    .Y(_09346_));
 INVx1_ASAP7_75t_R _38644_ (.A(_07697_),
    .Y(_09347_));
 OAI21x1_ASAP7_75t_R _38645_ (.A1(_09345_),
    .A2(_09346_),
    .B(_09347_),
    .Y(_09349_));
 NAND2x2_ASAP7_75t_R _38646_ (.A(_09344_),
    .B(_09349_),
    .Y(_09350_));
 OAI21x1_ASAP7_75t_R _38647_ (.A1(_09340_),
    .A2(_09341_),
    .B(_09350_),
    .Y(_09351_));
 OAI21x1_ASAP7_75t_R _38648_ (.A1(_09342_),
    .A2(_09343_),
    .B(_09347_),
    .Y(_09352_));
 OAI21x1_ASAP7_75t_R _38649_ (.A1(_09345_),
    .A2(_09346_),
    .B(_07697_),
    .Y(_09353_));
 NAND2x2_ASAP7_75t_R _38650_ (.A(_09352_),
    .B(_09353_),
    .Y(_09354_));
 NOR2x1_ASAP7_75t_R _38651_ (.A(_09341_),
    .B(_09340_),
    .Y(_09355_));
 NAND2x1_ASAP7_75t_R _38652_ (.A(_09354_),
    .B(_09355_),
    .Y(_09356_));
 AOI21x1_ASAP7_75t_R _38653_ (.A1(_09351_),
    .A2(_09356_),
    .B(net388),
    .Y(_09357_));
 INVx1_ASAP7_75t_R _38654_ (.A(_00394_),
    .Y(_09358_));
 OAI21x1_ASAP7_75t_R _38655_ (.A1(_09338_),
    .A2(_09357_),
    .B(_09358_),
    .Y(_09360_));
 TAPCELL_ASAP7_75t_R PHY_281 ();
 NOR2x1_ASAP7_75t_R _38657_ (.A(_00528_),
    .B(_00832_),
    .Y(_09362_));
 OAI21x1_ASAP7_75t_R _38658_ (.A1(_09340_),
    .A2(_09341_),
    .B(_09354_),
    .Y(_09363_));
 NAND2x1_ASAP7_75t_R _38659_ (.A(_09355_),
    .B(_09350_),
    .Y(_09364_));
 AOI21x1_ASAP7_75t_R _38660_ (.A1(_09363_),
    .A2(_09364_),
    .B(net388),
    .Y(_09365_));
 OAI21x1_ASAP7_75t_R _38661_ (.A1(_09362_),
    .A2(_09365_),
    .B(_00394_),
    .Y(_09366_));
 NAND2x2_ASAP7_75t_R _38662_ (.A(_09366_),
    .B(_09360_),
    .Y(_00044_));
 OR2x2_ASAP7_75t_R _38663_ (.A(_00528_),
    .B(_00831_),
    .Y(_09367_));
 NOR2x1_ASAP7_75t_R _38664_ (.A(net1739),
    .B(_07806_),
    .Y(_09368_));
 INVx1_ASAP7_75t_R _38665_ (.A(_07717_),
    .Y(_09370_));
 INVx1_ASAP7_75t_R _38666_ (.A(_07728_),
    .Y(_09371_));
 NOR2x1_ASAP7_75t_R _38667_ (.A(_07741_),
    .B(_09371_),
    .Y(_09372_));
 NAND2x1_ASAP7_75t_R _38668_ (.A(_09370_),
    .B(_09372_),
    .Y(_09373_));
 NAND3x1_ASAP7_75t_R _38669_ (.A(_07790_),
    .B(_07800_),
    .C(_07796_),
    .Y(_09374_));
 INVx1_ASAP7_75t_R _38670_ (.A(_07785_),
    .Y(_09375_));
 NOR2x1_ASAP7_75t_R _38671_ (.A(_09374_),
    .B(_09375_),
    .Y(_09376_));
 INVx1_ASAP7_75t_R _38672_ (.A(_07771_),
    .Y(_09377_));
 NAND2x2_ASAP7_75t_R _38673_ (.A(_09376_),
    .B(_09377_),
    .Y(_09378_));
 NOR2x2_ASAP7_75t_R _38674_ (.A(_09373_),
    .B(_09378_),
    .Y(_09379_));
 NOR2x1_ASAP7_75t_R _38675_ (.A(_09268_),
    .B(_09379_),
    .Y(_09381_));
 OAI21x1_ASAP7_75t_R _38676_ (.A1(_09368_),
    .A2(_09381_),
    .B(_08170_),
    .Y(_09382_));
 NOR2x1_ASAP7_75t_R _38677_ (.A(_09268_),
    .B(_07806_),
    .Y(_09383_));
 NOR2x1_ASAP7_75t_R _38678_ (.A(net1739),
    .B(_09379_),
    .Y(_09384_));
 OAI21x1_ASAP7_75t_R _38679_ (.A1(_09383_),
    .A2(_09384_),
    .B(_08169_),
    .Y(_09385_));
 NAND2x2_ASAP7_75t_R _38680_ (.A(_09382_),
    .B(_09385_),
    .Y(_09386_));
 INVx1_ASAP7_75t_R _38681_ (.A(_09386_),
    .Y(_09387_));
 XOR2x1_ASAP7_75t_R _38682_ (.A(_09203_),
    .Y(_09388_),
    .B(_09188_));
 NAND2x1_ASAP7_75t_R _38683_ (.A(_09388_),
    .B(_09387_),
    .Y(_09389_));
 NOR2x1_ASAP7_75t_R _38684_ (.A(_09188_),
    .B(_09203_),
    .Y(_09390_));
 AND2x2_ASAP7_75t_R _38685_ (.A(_09203_),
    .B(_09188_),
    .Y(_09392_));
 OAI21x1_ASAP7_75t_R _38686_ (.A1(_09390_),
    .A2(_09392_),
    .B(_09386_),
    .Y(_09393_));
 NAND3x1_ASAP7_75t_R _38687_ (.A(_09389_),
    .B(_09393_),
    .C(_00528_),
    .Y(_09394_));
 AOI21x1_ASAP7_75t_R _38688_ (.A1(_09367_),
    .A2(_09394_),
    .B(_00395_),
    .Y(_09395_));
 NAND2x1_ASAP7_75t_R _38689_ (.A(_00831_),
    .B(net388),
    .Y(_09396_));
 AO21x1_ASAP7_75t_R _38690_ (.A1(_09389_),
    .A2(_09393_),
    .B(net388),
    .Y(_09397_));
 AOI21x1_ASAP7_75t_R _38691_ (.A1(_09396_),
    .A2(_09397_),
    .B(_17244_),
    .Y(_09398_));
 NOR2x1_ASAP7_75t_R _38692_ (.A(_09395_),
    .B(_09398_),
    .Y(_00045_));
 AND2x2_ASAP7_75t_R _38693_ (.A(net388),
    .B(_00830_),
    .Y(_09399_));
 NOR2x1_ASAP7_75t_R _38694_ (.A(_08338_),
    .B(_08504_),
    .Y(_09400_));
 NOR2x1_ASAP7_75t_R _38695_ (.A(_09223_),
    .B(_08517_),
    .Y(_09402_));
 OAI21x1_ASAP7_75t_R _38696_ (.A1(_09400_),
    .A2(_09402_),
    .B(_08601_),
    .Y(_09403_));
 INVx2_ASAP7_75t_R _38697_ (.A(_09403_),
    .Y(_09404_));
 NAND2x2_ASAP7_75t_R _38698_ (.A(_08504_),
    .B(_08338_),
    .Y(_09405_));
 OAI22x1_ASAP7_75t_R _38699_ (.A1(_08337_),
    .A2(_06425_),
    .B1(_08503_),
    .B2(_05717_),
    .Y(_09406_));
 NAND3x2_ASAP7_75t_R _38700_ (.B(_09406_),
    .C(_09213_),
    .Y(_09407_),
    .A(_09405_));
 INVx1_ASAP7_75t_R _38701_ (.A(_09407_),
    .Y(_09408_));
 INVx1_ASAP7_75t_R _38702_ (.A(_08087_),
    .Y(_09409_));
 OAI21x1_ASAP7_75t_R _38703_ (.A1(_09404_),
    .A2(_09408_),
    .B(_09409_),
    .Y(_09410_));
 NAND3x1_ASAP7_75t_R _38704_ (.A(_09407_),
    .B(_08087_),
    .C(_09403_),
    .Y(_09411_));
 AOI21x1_ASAP7_75t_R _38705_ (.A1(_09410_),
    .A2(_09411_),
    .B(net388),
    .Y(_09413_));
 OAI21x1_ASAP7_75t_R _38706_ (.A1(_09399_),
    .A2(_09413_),
    .B(_16062_),
    .Y(_09414_));
 NOR2x1_ASAP7_75t_R _38707_ (.A(_00528_),
    .B(_00830_),
    .Y(_09415_));
 OAI21x1_ASAP7_75t_R _38708_ (.A1(_09404_),
    .A2(_09408_),
    .B(_08087_),
    .Y(_09416_));
 NAND3x1_ASAP7_75t_R _38709_ (.A(_09407_),
    .B(_09409_),
    .C(_09403_),
    .Y(_09417_));
 AOI21x1_ASAP7_75t_R _38710_ (.A1(_09416_),
    .A2(_09417_),
    .B(net388),
    .Y(_09418_));
 OAI21x1_ASAP7_75t_R _38711_ (.A1(_09415_),
    .A2(_09418_),
    .B(_00490_),
    .Y(_09419_));
 NAND2x2_ASAP7_75t_R _38712_ (.A(_09419_),
    .B(_09414_),
    .Y(_00046_));
 NOR2x2_ASAP7_75t_R _38713_ (.A(net394),
    .B(_00829_),
    .Y(_09420_));
 INVx1_ASAP7_75t_R _38714_ (.A(_09420_),
    .Y(_09421_));
 NAND2x1_ASAP7_75t_R _38715_ (.A(_08420_),
    .B(net3448),
    .Y(_09423_));
 NOR2x1_ASAP7_75t_R _38716_ (.A(net1860),
    .B(net3448),
    .Y(_09424_));
 INVx1_ASAP7_75t_R _38717_ (.A(_09424_),
    .Y(_09425_));
 AOI21x1_ASAP7_75t_R _38718_ (.A1(_09423_),
    .A2(_09425_),
    .B(_09227_),
    .Y(_09426_));
 AOI22x1_ASAP7_75t_R _38719_ (.A1(_08852_),
    .A2(net1978),
    .B1(_08507_),
    .B2(_05479_),
    .Y(_09427_));
 NOR2x1_ASAP7_75t_R _38720_ (.A(_08508_),
    .B(_08853_),
    .Y(_09428_));
 OAI21x1_ASAP7_75t_R _38721_ (.A1(_09427_),
    .A2(_09428_),
    .B(_09227_),
    .Y(_09429_));
 INVx1_ASAP7_75t_R _38722_ (.A(_09429_),
    .Y(_09430_));
 XNOR2x1_ASAP7_75t_R _38723_ (.B(net2774),
    .Y(_09431_),
    .A(_08849_));
 INVx1_ASAP7_75t_R _38724_ (.A(_09431_),
    .Y(_09432_));
 OAI21x1_ASAP7_75t_R _38725_ (.A1(_09426_),
    .A2(_09430_),
    .B(_09432_),
    .Y(_09434_));
 NOR2x1_ASAP7_75t_R _38726_ (.A(_08508_),
    .B(_08689_),
    .Y(_09435_));
 OAI21x1_ASAP7_75t_R _38727_ (.A1(_09424_),
    .A2(_09435_),
    .B(_09022_),
    .Y(_09436_));
 NAND3x1_ASAP7_75t_R _38728_ (.A(_09436_),
    .B(_09429_),
    .C(_09431_),
    .Y(_09437_));
 AOI21x1_ASAP7_75t_R _38729_ (.A1(_09434_),
    .A2(_09437_),
    .B(net388),
    .Y(_09438_));
 INVx1_ASAP7_75t_R _38730_ (.A(_09438_),
    .Y(_09439_));
 AOI21x1_ASAP7_75t_R _38731_ (.A1(_09421_),
    .A2(_09439_),
    .B(_00489_),
    .Y(_09440_));
 NOR3x1_ASAP7_75t_R _38732_ (.A(_09438_),
    .B(_16132_),
    .C(_09420_),
    .Y(_09441_));
 NOR2x1_ASAP7_75t_R _38733_ (.A(_09441_),
    .B(_09440_),
    .Y(_00047_));
 AND2x2_ASAP7_75t_R _38734_ (.A(net388),
    .B(_00828_),
    .Y(_09442_));
 NOR2x2_ASAP7_75t_R _38735_ (.A(net2471),
    .B(_09247_),
    .Y(_09444_));
 AND2x4_ASAP7_75t_R _38736_ (.A(_09247_),
    .B(net2471),
    .Y(_09445_));
 XOR2x2_ASAP7_75t_R _38737_ (.A(_08946_),
    .B(_05715_),
    .Y(_09446_));
 OAI21x1_ASAP7_75t_R _38738_ (.A1(_09444_),
    .A2(_09445_),
    .B(_09446_),
    .Y(_09447_));
 NOR2x2_ASAP7_75t_R _38739_ (.A(net2471),
    .B(_09249_),
    .Y(_09448_));
 AND2x4_ASAP7_75t_R _38740_ (.A(_09249_),
    .B(net2471),
    .Y(_09449_));
 INVx1_ASAP7_75t_R _38741_ (.A(_09446_),
    .Y(_09450_));
 OAI21x1_ASAP7_75t_R _38742_ (.A1(_09448_),
    .A2(_09449_),
    .B(_09450_),
    .Y(_09451_));
 AOI21x1_ASAP7_75t_R _38743_ (.A1(_09447_),
    .A2(_09451_),
    .B(net388),
    .Y(_09452_));
 INVx1_ASAP7_75t_R _38744_ (.A(_00396_),
    .Y(_09453_));
 OAI21x1_ASAP7_75t_R _38745_ (.A1(_09442_),
    .A2(_09452_),
    .B(_09453_),
    .Y(_09455_));
 NOR2x1_ASAP7_75t_R _38746_ (.A(net394),
    .B(_00828_),
    .Y(_09456_));
 OAI21x1_ASAP7_75t_R _38747_ (.A1(_09444_),
    .A2(_09445_),
    .B(_09450_),
    .Y(_09457_));
 OAI21x1_ASAP7_75t_R _38748_ (.A1(_09448_),
    .A2(_09449_),
    .B(_09446_),
    .Y(_09458_));
 AOI21x1_ASAP7_75t_R _38749_ (.A1(_09457_),
    .A2(_09458_),
    .B(net388),
    .Y(_09459_));
 OAI21x1_ASAP7_75t_R _38750_ (.A1(_09456_),
    .A2(_09459_),
    .B(_00396_),
    .Y(_09460_));
 NAND2x2_ASAP7_75t_R _38751_ (.A(_09455_),
    .B(_09460_),
    .Y(_00048_));
 XOR2x1_ASAP7_75t_R _38752_ (.A(net3119),
    .Y(_09461_),
    .B(_09271_));
 XOR2x1_ASAP7_75t_R _38753_ (.A(_06026_),
    .Y(_09462_),
    .B(_05693_));
 XOR2x1_ASAP7_75t_R _38754_ (.A(_09461_),
    .Y(_09463_),
    .B(_09462_));
 NOR2x1_ASAP7_75t_R _38755_ (.A(net394),
    .B(_00827_),
    .Y(_09465_));
 AO21x1_ASAP7_75t_R _38756_ (.A1(_09463_),
    .A2(net394),
    .B(_09465_),
    .Y(_09466_));
 XOR2x1_ASAP7_75t_R _38757_ (.A(_09466_),
    .Y(_00009_),
    .B(_17386_));
 AND2x2_ASAP7_75t_R _38758_ (.A(net388),
    .B(_00826_),
    .Y(_09467_));
 NOR2x1_ASAP7_75t_R _38759_ (.A(_09324_),
    .B(_09308_),
    .Y(_09468_));
 NOR2x2_ASAP7_75t_R _38760_ (.A(_09305_),
    .B(_09329_),
    .Y(_09469_));
 AOI21x1_ASAP7_75t_R _38761_ (.A1(_05430_),
    .A2(_05428_),
    .B(_07381_),
    .Y(_09470_));
 AOI21x1_ASAP7_75t_R _38762_ (.A1(_05731_),
    .A2(_05729_),
    .B(_09141_),
    .Y(_09471_));
 NOR2x2_ASAP7_75t_R _38763_ (.A(_09471_),
    .B(_09470_),
    .Y(_09472_));
 OAI21x1_ASAP7_75t_R _38764_ (.A1(_09468_),
    .A2(_09469_),
    .B(_09472_),
    .Y(_09473_));
 INVx2_ASAP7_75t_R _38765_ (.A(_09472_),
    .Y(_09475_));
 XOR2x1_ASAP7_75t_R _38766_ (.A(_09308_),
    .Y(_09476_),
    .B(_09324_));
 NAND2x1_ASAP7_75t_R _38767_ (.A(_09476_),
    .B(_09475_),
    .Y(_09477_));
 AOI21x1_ASAP7_75t_R _38768_ (.A1(_09473_),
    .A2(_09477_),
    .B(net388),
    .Y(_09478_));
 INVx1_ASAP7_75t_R _38769_ (.A(_00400_),
    .Y(_09479_));
 OAI21x1_ASAP7_75t_R _38770_ (.A1(_09467_),
    .A2(_09478_),
    .B(_09479_),
    .Y(_09480_));
 NOR2x1_ASAP7_75t_R _38771_ (.A(net394),
    .B(_00826_),
    .Y(_09481_));
 NAND2x1_ASAP7_75t_R _38772_ (.A(_09472_),
    .B(_09476_),
    .Y(_09482_));
 OAI21x1_ASAP7_75t_R _38773_ (.A1(_09469_),
    .A2(_09468_),
    .B(_09475_),
    .Y(_09483_));
 AOI21x1_ASAP7_75t_R _38774_ (.A1(_09482_),
    .A2(_09483_),
    .B(net388),
    .Y(_09484_));
 OAI21x1_ASAP7_75t_R _38775_ (.A1(_09481_),
    .A2(_09484_),
    .B(_00400_),
    .Y(_09486_));
 NAND2x1_ASAP7_75t_R _38776_ (.A(_09486_),
    .B(_09480_),
    .Y(_00010_));
 NOR2x1_ASAP7_75t_R _38777_ (.A(_06679_),
    .B(net3419),
    .Y(_09487_));
 NOR2x1_ASAP7_75t_R _38778_ (.A(net1927),
    .B(_06422_),
    .Y(_09488_));
 OAI21x1_ASAP7_75t_R _38779_ (.A1(_09487_),
    .A2(_09488_),
    .B(_07499_),
    .Y(_09489_));
 NOR2x1_ASAP7_75t_R _38780_ (.A(net1927),
    .B(net3419),
    .Y(_09490_));
 NOR2x1_ASAP7_75t_R _38781_ (.A(_06679_),
    .B(_06422_),
    .Y(_09491_));
 OAI21x1_ASAP7_75t_R _38782_ (.A1(_09490_),
    .A2(_09491_),
    .B(_09158_),
    .Y(_09492_));
 XOR2x1_ASAP7_75t_R _38783_ (.A(_07159_),
    .Y(_09493_),
    .B(_07272_));
 INVx1_ASAP7_75t_R _38784_ (.A(_09493_),
    .Y(_09494_));
 NAND3x1_ASAP7_75t_R _38785_ (.A(_09489_),
    .B(_09492_),
    .C(_09494_),
    .Y(_09496_));
 NAND2x1_ASAP7_75t_R _38786_ (.A(_09489_),
    .B(_09492_),
    .Y(_09497_));
 AOI21x1_ASAP7_75t_R _38787_ (.A1(_09493_),
    .A2(_09497_),
    .B(net388),
    .Y(_09498_));
 AND2x2_ASAP7_75t_R _38788_ (.A(net388),
    .B(_00825_),
    .Y(_09499_));
 AOI21x1_ASAP7_75t_R _38789_ (.A1(_09496_),
    .A2(_09498_),
    .B(_09499_),
    .Y(_09500_));
 XOR2x1_ASAP7_75t_R _38790_ (.A(_09500_),
    .Y(_00011_),
    .B(_17275_));
 AND2x2_ASAP7_75t_R _38791_ (.A(net388),
    .B(_00824_),
    .Y(_09501_));
 NOR2x2_ASAP7_75t_R _38792_ (.A(_09345_),
    .B(_09346_),
    .Y(_09502_));
 NOR2x2_ASAP7_75t_R _38793_ (.A(_07812_),
    .B(_09502_),
    .Y(_09503_));
 NOR2x1_ASAP7_75t_R _38794_ (.A(_09343_),
    .B(_09342_),
    .Y(_09504_));
 NOR2x1_ASAP7_75t_R _38795_ (.A(_07596_),
    .B(_09504_),
    .Y(_09506_));
 XOR2x2_ASAP7_75t_R _38796_ (.A(_09339_),
    .B(_09379_),
    .Y(_09507_));
 OAI21x1_ASAP7_75t_R _38797_ (.A1(_09503_),
    .A2(_09506_),
    .B(_09507_),
    .Y(_09508_));
 NOR2x2_ASAP7_75t_R _38798_ (.A(_07596_),
    .B(_09502_),
    .Y(_09509_));
 NOR2x1_ASAP7_75t_R _38799_ (.A(_07812_),
    .B(_09504_),
    .Y(_09510_));
 XOR2x2_ASAP7_75t_R _38800_ (.A(_09339_),
    .B(_07806_),
    .Y(_09511_));
 OAI21x1_ASAP7_75t_R _38801_ (.A1(_09509_),
    .A2(_09510_),
    .B(_09511_),
    .Y(_09512_));
 AOI21x1_ASAP7_75t_R _38802_ (.A1(_09508_),
    .A2(_09512_),
    .B(net388),
    .Y(_09513_));
 OAI21x1_ASAP7_75t_R _38803_ (.A1(_09501_),
    .A2(_09513_),
    .B(_17284_),
    .Y(_09514_));
 NOR2x1_ASAP7_75t_R _38804_ (.A(net394),
    .B(_00824_),
    .Y(_09515_));
 OAI21x1_ASAP7_75t_R _38805_ (.A1(_09509_),
    .A2(_09510_),
    .B(_09507_),
    .Y(_09517_));
 OAI21x1_ASAP7_75t_R _38806_ (.A1(_09503_),
    .A2(_09506_),
    .B(_09511_),
    .Y(_09518_));
 AOI21x1_ASAP7_75t_R _38807_ (.A1(_09517_),
    .A2(_09518_),
    .B(net388),
    .Y(_09519_));
 OAI21x1_ASAP7_75t_R _38808_ (.A1(_09515_),
    .A2(_09519_),
    .B(_00487_),
    .Y(_09520_));
 NAND2x1_ASAP7_75t_R _38809_ (.A(_09514_),
    .B(_09520_),
    .Y(_00012_));
 NOR2x2_ASAP7_75t_R _38810_ (.A(net394),
    .B(_00823_),
    .Y(_09521_));
 INVx1_ASAP7_75t_R _38811_ (.A(_09521_),
    .Y(_09522_));
 XOR2x1_ASAP7_75t_R _38812_ (.A(_08087_),
    .Y(_09523_),
    .B(_08266_));
 XOR2x2_ASAP7_75t_R _38813_ (.A(_07806_),
    .B(net1739),
    .Y(_09524_));
 XOR2x1_ASAP7_75t_R _38814_ (.A(_08090_),
    .Y(_09525_),
    .B(_09524_));
 NAND2x1_ASAP7_75t_R _38815_ (.A(_09525_),
    .B(_09523_),
    .Y(_09527_));
 NOR2x1_ASAP7_75t_R _38816_ (.A(_09524_),
    .B(_08090_),
    .Y(_09528_));
 AND2x2_ASAP7_75t_R _38817_ (.A(_08090_),
    .B(_09524_),
    .Y(_09529_));
 INVx1_ASAP7_75t_R _38818_ (.A(_08005_),
    .Y(_09530_));
 AOI21x1_ASAP7_75t_R _38819_ (.A1(_09206_),
    .A2(_09205_),
    .B(_09530_),
    .Y(_09531_));
 OAI21x1_ASAP7_75t_R _38820_ (.A1(_08085_),
    .A2(_08048_),
    .B(_08266_),
    .Y(_09532_));
 NAND2x1_ASAP7_75t_R _38821_ (.A(_08086_),
    .B(_09186_),
    .Y(_09533_));
 AOI21x1_ASAP7_75t_R _38822_ (.A1(_09532_),
    .A2(_09533_),
    .B(_08005_),
    .Y(_09534_));
 NOR2x1_ASAP7_75t_R _38823_ (.A(_09531_),
    .B(_09534_),
    .Y(_09535_));
 OAI21x1_ASAP7_75t_R _38824_ (.A1(_09528_),
    .A2(_09529_),
    .B(_09535_),
    .Y(_09536_));
 AOI21x1_ASAP7_75t_R _38825_ (.A1(_09527_),
    .A2(_09536_),
    .B(net388),
    .Y(_09538_));
 INVx1_ASAP7_75t_R _38826_ (.A(_09538_),
    .Y(_09539_));
 AOI21x1_ASAP7_75t_R _38827_ (.A1(_09522_),
    .A2(_09539_),
    .B(_00486_),
    .Y(_09540_));
 NOR3x1_ASAP7_75t_R _38828_ (.A(_09538_),
    .B(_17293_),
    .C(_09521_),
    .Y(_09541_));
 NOR2x1_ASAP7_75t_R _38829_ (.A(_09540_),
    .B(_09541_),
    .Y(_00013_));
 OAI21x1_ASAP7_75t_R _38830_ (.A1(_09230_),
    .A2(_09229_),
    .B(net1860),
    .Y(_09542_));
 OAI21x1_ASAP7_75t_R _38831_ (.A1(_09225_),
    .A2(_09224_),
    .B(_08508_),
    .Y(_09543_));
 AOI21x1_ASAP7_75t_R _38832_ (.A1(_09542_),
    .A2(_09543_),
    .B(_09189_),
    .Y(_09544_));
 AO31x2_ASAP7_75t_R _38833_ (.A1(_09542_),
    .A2(_09543_),
    .A3(_09189_),
    .B(net388),
    .Y(_09545_));
 NAND2x1_ASAP7_75t_R _38834_ (.A(_00822_),
    .B(net388),
    .Y(_09546_));
 OAI21x1_ASAP7_75t_R _38835_ (.A1(_09544_),
    .A2(_09545_),
    .B(_09546_),
    .Y(_09548_));
 XOR2x1_ASAP7_75t_R _38836_ (.A(_09548_),
    .Y(_00014_),
    .B(_00405_));
 XOR2x1_ASAP7_75t_R _38837_ (.A(_08771_),
    .Y(_09549_),
    .B(_09022_));
 OAI21x1_ASAP7_75t_R _38838_ (.A1(_08506_),
    .A2(_08518_),
    .B(_08689_),
    .Y(_09550_));
 OAI21x1_ASAP7_75t_R _38839_ (.A1(_09209_),
    .A2(_09210_),
    .B(net1948),
    .Y(_09551_));
 NAND2x1_ASAP7_75t_R _38840_ (.A(_09551_),
    .B(_09550_),
    .Y(_09552_));
 OAI21x1_ASAP7_75t_R _38841_ (.A1(_09549_),
    .A2(_09552_),
    .B(net394),
    .Y(_09553_));
 AND2x2_ASAP7_75t_R _38842_ (.A(_09549_),
    .B(_09552_),
    .Y(_09554_));
 NAND2x1_ASAP7_75t_R _38843_ (.A(_00821_),
    .B(net388),
    .Y(_09555_));
 OAI21x1_ASAP7_75t_R _38844_ (.A1(_09553_),
    .A2(_09554_),
    .B(_09555_),
    .Y(_09556_));
 XOR2x1_ASAP7_75t_R _38845_ (.A(_09556_),
    .Y(_00015_),
    .B(_00407_));
 NOR2x2_ASAP7_75t_R _38846_ (.A(net394),
    .B(_00820_),
    .Y(_09558_));
 XOR2x1_ASAP7_75t_R _38847_ (.A(_09108_),
    .Y(_09559_),
    .B(_06729_));
 XOR2x1_ASAP7_75t_R _38848_ (.A(_09559_),
    .Y(_09560_),
    .B(net1964));
 NOR2x1_ASAP7_75t_R _38849_ (.A(_09560_),
    .B(_08850_),
    .Y(_09561_));
 AND2x2_ASAP7_75t_R _38850_ (.A(_08850_),
    .B(_09560_),
    .Y(_09562_));
 OAI21x1_ASAP7_75t_R _38851_ (.A1(_09561_),
    .A2(_09562_),
    .B(net394),
    .Y(_09563_));
 INVx1_ASAP7_75t_R _38852_ (.A(_09563_),
    .Y(_09564_));
 OAI21x1_ASAP7_75t_R _38853_ (.A1(_09558_),
    .A2(_09564_),
    .B(_00485_),
    .Y(_09565_));
 INVx1_ASAP7_75t_R _38854_ (.A(_09558_),
    .Y(_09566_));
 NAND3x1_ASAP7_75t_R _38855_ (.A(_09563_),
    .B(_17312_),
    .C(_09566_),
    .Y(_09568_));
 NAND2x1_ASAP7_75t_R _38856_ (.A(_09565_),
    .B(_09568_),
    .Y(_00016_));
 NOR2x2_ASAP7_75t_R _38857_ (.A(net393),
    .B(_00819_),
    .Y(_09569_));
 TAPCELL_ASAP7_75t_R PHY_280 ();
 TAPCELL_ASAP7_75t_R PHY_279 ();
 TAPCELL_ASAP7_75t_R PHY_278 ();
 CKINVDCx20_ASAP7_75t_R _38861_ (.A(net1278),
    .Y(_09573_));
 NAND2x2_ASAP7_75t_R _38862_ (.A(net1105),
    .B(_09573_),
    .Y(_09574_));
 TAPCELL_ASAP7_75t_R PHY_277 ();
 TAPCELL_ASAP7_75t_R PHY_276 ();
 INVx4_ASAP7_75t_R _38865_ (.A(net1625),
    .Y(_09578_));
 NAND2x2_ASAP7_75t_R _38866_ (.A(net1723),
    .B(_09578_),
    .Y(_09579_));
 NOR2x2_ASAP7_75t_R _38867_ (.A(_09574_),
    .B(_09579_),
    .Y(_09580_));
 NAND2x2_ASAP7_75t_R _38868_ (.A(net1106),
    .B(net1283),
    .Y(_09581_));
 NOR2x1_ASAP7_75t_R _38869_ (.A(_09581_),
    .B(net1476),
    .Y(_09582_));
 NAND2x2_ASAP7_75t_R _38870_ (.A(_00611_),
    .B(net2173),
    .Y(_09583_));
 TAPCELL_ASAP7_75t_R PHY_275 ();
 NAND2x2_ASAP7_75t_R _38872_ (.A(_00609_),
    .B(_00610_),
    .Y(_09585_));
 NOR2x2_ASAP7_75t_R _38873_ (.A(_09583_),
    .B(_09585_),
    .Y(_09586_));
 OA21x2_ASAP7_75t_R _38874_ (.A1(_09580_),
    .A2(_09582_),
    .B(net1218),
    .Y(_09587_));
 CKINVDCx20_ASAP7_75t_R _38875_ (.A(net1111),
    .Y(_09589_));
 INVx2_ASAP7_75t_R _38876_ (.A(_00614_),
    .Y(_09590_));
 NOR2x2_ASAP7_75t_R _38877_ (.A(net1625),
    .B(_09590_),
    .Y(_09591_));
 NAND2x2_ASAP7_75t_R _38878_ (.A(_09589_),
    .B(_09591_),
    .Y(_09592_));
 TAPCELL_ASAP7_75t_R PHY_274 ();
 CKINVDCx10_ASAP7_75t_R _38880_ (.A(net2927),
    .Y(_09594_));
 NOR2x2_ASAP7_75t_R _38881_ (.A(_09592_),
    .B(net2656),
    .Y(_09595_));
 NOR2x2_ASAP7_75t_R _38882_ (.A(net1625),
    .B(net1722),
    .Y(_09596_));
 CKINVDCx20_ASAP7_75t_R _38883_ (.A(net1099),
    .Y(_09597_));
 TAPCELL_ASAP7_75t_R PHY_273 ();
 TAPCELL_ASAP7_75t_R PHY_272 ();
 NOR2x2_ASAP7_75t_R _38886_ (.A(_09597_),
    .B(net2656),
    .Y(_09601_));
 NOR3x2_ASAP7_75t_R _38887_ (.B(_09595_),
    .C(_09601_),
    .Y(_09602_),
    .A(_09587_));
 NOR2x2_ASAP7_75t_R _38888_ (.A(net1723),
    .B(_09578_),
    .Y(_09603_));
 TAPCELL_ASAP7_75t_R PHY_271 ();
 NAND2x2_ASAP7_75t_R _38890_ (.A(net1930),
    .B(net1218),
    .Y(_09605_));
 NOR2x2_ASAP7_75t_R _38891_ (.A(_09589_),
    .B(net1282),
    .Y(_09606_));
 NAND2x2_ASAP7_75t_R _38892_ (.A(net1625),
    .B(_00614_),
    .Y(_09607_));
 CKINVDCx10_ASAP7_75t_R _38893_ (.A(net981),
    .Y(_09608_));
 TAPCELL_ASAP7_75t_R PHY_270 ();
 NAND2x2_ASAP7_75t_R _38895_ (.A(_09606_),
    .B(_09608_),
    .Y(_09611_));
 NOR2x2_ASAP7_75t_R _38896_ (.A(net1111),
    .B(net2798),
    .Y(_09612_));
 INVx4_ASAP7_75t_R _38897_ (.A(_09612_),
    .Y(_09613_));
 AO21x2_ASAP7_75t_R _38898_ (.A1(_09611_),
    .A2(_09613_),
    .B(_09594_),
    .Y(_09614_));
 NAND2x2_ASAP7_75t_R _38899_ (.A(_09614_),
    .B(_09605_),
    .Y(_09615_));
 INVx2_ASAP7_75t_R _38900_ (.A(_09615_),
    .Y(_09616_));
 INVx2_ASAP7_75t_R _38901_ (.A(_00611_),
    .Y(_09617_));
 NOR2x2_ASAP7_75t_R _38902_ (.A(net2173),
    .B(_09617_),
    .Y(_09618_));
 INVx4_ASAP7_75t_R _38903_ (.A(net2481),
    .Y(_09619_));
 NAND2x2_ASAP7_75t_R _38904_ (.A(_09618_),
    .B(_09619_),
    .Y(_09620_));
 TAPCELL_ASAP7_75t_R PHY_269 ();
 NAND3x2_ASAP7_75t_R _38906_ (.B(_09616_),
    .C(net2289),
    .Y(_09623_),
    .A(_09602_));
 INVx3_ASAP7_75t_R _38907_ (.A(net1760),
    .Y(_09624_));
 NOR2x2_ASAP7_75t_R _38908_ (.A(net1842),
    .B(_09624_),
    .Y(_09625_));
 AND3x2_ASAP7_75t_R _38909_ (.A(_09617_),
    .B(net1760),
    .C(_00610_),
    .Y(_09626_));
 NOR3x2_ASAP7_75t_R _38910_ (.B(net2931),
    .C(_09626_),
    .Y(_09627_),
    .A(_09623_));
 NAND2x2_ASAP7_75t_R _38911_ (.A(net1761),
    .B(_09627_),
    .Y(_09628_));
 NOR2x2_ASAP7_75t_R _38912_ (.A(net1105),
    .B(net1282),
    .Y(_09629_));
 TAPCELL_ASAP7_75t_R PHY_268 ();
 NAND2x2_ASAP7_75t_R _38914_ (.A(net2068),
    .B(_09629_),
    .Y(_09631_));
 INVx1_ASAP7_75t_R _38915_ (.A(_09631_),
    .Y(_09633_));
 TAPCELL_ASAP7_75t_R PHY_267 ();
 NAND2x2_ASAP7_75t_R _38917_ (.A(net1107),
    .B(net2068),
    .Y(_09635_));
 NAND2x2_ASAP7_75t_R _38918_ (.A(_09606_),
    .B(_09591_),
    .Y(_09636_));
 NAND2x1_ASAP7_75t_R _38919_ (.A(_09635_),
    .B(net1289),
    .Y(_09637_));
 NAND2x2_ASAP7_75t_R _38920_ (.A(net2174),
    .B(_09617_),
    .Y(_09638_));
 NAND2x2_ASAP7_75t_R _38921_ (.A(net1842),
    .B(_09624_),
    .Y(_09639_));
 NOR2x2_ASAP7_75t_R _38922_ (.A(_09638_),
    .B(_09639_),
    .Y(_09640_));
 OAI21x1_ASAP7_75t_R _38923_ (.A1(_09633_),
    .A2(_09637_),
    .B(_09640_),
    .Y(_09641_));
 NAND2x2_ASAP7_75t_R _38924_ (.A(net2068),
    .B(_09606_),
    .Y(_09642_));
 NAND2x2_ASAP7_75t_R _38925_ (.A(_09589_),
    .B(net2068),
    .Y(_09644_));
 TAPCELL_ASAP7_75t_R PHY_266 ();
 INVx2_ASAP7_75t_R _38927_ (.A(net2287),
    .Y(_09646_));
 NOR2x2_ASAP7_75t_R _38928_ (.A(net1760),
    .B(_09646_),
    .Y(_09647_));
 INVx3_ASAP7_75t_R _38929_ (.A(_09583_),
    .Y(_09648_));
 NAND2x2_ASAP7_75t_R _38930_ (.A(_09647_),
    .B(_09648_),
    .Y(_09649_));
 AO21x2_ASAP7_75t_R _38931_ (.A1(_09642_),
    .A2(_09644_),
    .B(_09649_),
    .Y(_09650_));
 AND2x2_ASAP7_75t_R _38932_ (.A(_09641_),
    .B(_09650_),
    .Y(_09651_));
 TAPCELL_ASAP7_75t_R PHY_265 ();
 NAND2x2_ASAP7_75t_R _38934_ (.A(_09629_),
    .B(_09591_),
    .Y(_09653_));
 NAND2x2_ASAP7_75t_R _38935_ (.A(_09625_),
    .B(_09648_),
    .Y(_09655_));
 AO21x2_ASAP7_75t_R _38936_ (.A1(net2771),
    .A2(_09653_),
    .B(_09655_),
    .Y(_09656_));
 AND2x4_ASAP7_75t_R _38937_ (.A(net1108),
    .B(net1284),
    .Y(_09657_));
 NAND2x2_ASAP7_75t_R _38938_ (.A(net2068),
    .B(_09657_),
    .Y(_09658_));
 AO21x1_ASAP7_75t_R _38939_ (.A1(_09658_),
    .A2(_09642_),
    .B(net3241),
    .Y(_09659_));
 NAND2x2_ASAP7_75t_R _38940_ (.A(net1763),
    .B(_09646_),
    .Y(_09660_));
 NOR2x2_ASAP7_75t_R _38941_ (.A(net1843),
    .B(_09660_),
    .Y(_09661_));
 NAND2x2_ASAP7_75t_R _38942_ (.A(net1282),
    .B(_09589_),
    .Y(_09662_));
 TAPCELL_ASAP7_75t_R PHY_264 ();
 NOR2x2_ASAP7_75t_R _38944_ (.A(_09662_),
    .B(_09597_),
    .Y(_09664_));
 NAND2x1_ASAP7_75t_R _38945_ (.A(_09661_),
    .B(_09664_),
    .Y(_09666_));
 AND3x2_ASAP7_75t_R _38946_ (.A(_09656_),
    .B(_09659_),
    .C(_09666_),
    .Y(_09667_));
 NAND2x1_ASAP7_75t_R _38947_ (.A(_09651_),
    .B(_09667_),
    .Y(_09668_));
 TAPCELL_ASAP7_75t_R PHY_263 ();
 INVx2_ASAP7_75t_R _38949_ (.A(net2173),
    .Y(_09670_));
 NOR2x2_ASAP7_75t_R _38950_ (.A(net2929),
    .B(_09670_),
    .Y(_09671_));
 NAND2x2_ASAP7_75t_R _38951_ (.A(_09625_),
    .B(_09671_),
    .Y(_09672_));
 TAPCELL_ASAP7_75t_R PHY_262 ();
 NAND2x2_ASAP7_75t_R _38953_ (.A(_09590_),
    .B(net1625),
    .Y(_09674_));
 TAPCELL_ASAP7_75t_R PHY_261 ();
 NOR2x2_ASAP7_75t_R _38955_ (.A(_00609_),
    .B(net3060),
    .Y(_09677_));
 NAND2x2_ASAP7_75t_R _38956_ (.A(_09677_),
    .B(_09618_),
    .Y(_09678_));
 TAPCELL_ASAP7_75t_R PHY_260 ();
 TAPCELL_ASAP7_75t_R PHY_259 ();
 OAI22x1_ASAP7_75t_R _38959_ (.A1(net2775),
    .A2(_09674_),
    .B1(_09678_),
    .B2(net3066),
    .Y(_09681_));
 NAND2x2_ASAP7_75t_R _38960_ (.A(_09671_),
    .B(_09647_),
    .Y(_09682_));
 TAPCELL_ASAP7_75t_R PHY_258 ();
 NAND2x2_ASAP7_75t_R _38962_ (.A(net1933),
    .B(_09657_),
    .Y(_09684_));
 TAPCELL_ASAP7_75t_R PHY_257 ();
 NOR2x1_ASAP7_75t_R _38964_ (.A(_09682_),
    .B(net2724),
    .Y(_09686_));
 AOI211x1_ASAP7_75t_R _38965_ (.A1(net1218),
    .A2(_09580_),
    .B(_09681_),
    .C(_09686_),
    .Y(_09688_));
 NAND2x2_ASAP7_75t_R _38966_ (.A(_09591_),
    .B(_09657_),
    .Y(_09689_));
 TAPCELL_ASAP7_75t_R PHY_256 ();
 NOR2x2_ASAP7_75t_R _38968_ (.A(_00611_),
    .B(net2173),
    .Y(_09691_));
 NAND2x2_ASAP7_75t_R _38969_ (.A(_09691_),
    .B(_09619_),
    .Y(_09692_));
 TAPCELL_ASAP7_75t_R PHY_255 ();
 AO21x1_ASAP7_75t_R _38971_ (.A1(_09689_),
    .A2(_09631_),
    .B(_09692_),
    .Y(_09694_));
 NAND2x2_ASAP7_75t_R _38972_ (.A(_09625_),
    .B(_09618_),
    .Y(_09695_));
 INVx2_ASAP7_75t_R _38973_ (.A(_09695_),
    .Y(_09696_));
 NAND2x1_ASAP7_75t_R _38974_ (.A(_09633_),
    .B(_09696_),
    .Y(_09697_));
 TAPCELL_ASAP7_75t_R PHY_254 ();
 NOR2x2_ASAP7_75t_R _38976_ (.A(net2799),
    .B(_09574_),
    .Y(_09700_));
 NOR2x2_ASAP7_75t_R _38977_ (.A(_09660_),
    .B(_09638_),
    .Y(_09701_));
 TAPCELL_ASAP7_75t_R PHY_253 ();
 NAND2x1_ASAP7_75t_R _38979_ (.A(_09700_),
    .B(_09701_),
    .Y(_09703_));
 AND3x2_ASAP7_75t_R _38980_ (.A(_09694_),
    .B(_09697_),
    .C(_09703_),
    .Y(_09704_));
 NAND2x1_ASAP7_75t_R _38981_ (.A(_09688_),
    .B(_09704_),
    .Y(_09705_));
 NOR2x1_ASAP7_75t_R _38982_ (.A(_09668_),
    .B(_09705_),
    .Y(_09706_));
 NAND2x2_ASAP7_75t_R _38983_ (.A(_09671_),
    .B(_09619_),
    .Y(_09707_));
 TAPCELL_ASAP7_75t_R PHY_252 ();
 NOR2x2_ASAP7_75t_R _38985_ (.A(net1107),
    .B(_09573_),
    .Y(_09710_));
 NAND2x2_ASAP7_75t_R _38986_ (.A(net1933),
    .B(_09710_),
    .Y(_09711_));
 TAPCELL_ASAP7_75t_R PHY_251 ();
 OAI22x1_ASAP7_75t_R _38988_ (.A1(_09605_),
    .A2(net1113),
    .B1(_09707_),
    .B2(net1387),
    .Y(_09713_));
 NAND2x2_ASAP7_75t_R _38989_ (.A(_09710_),
    .B(_09608_),
    .Y(_09714_));
 NAND2x2_ASAP7_75t_R _38990_ (.A(net1105),
    .B(_09608_),
    .Y(_09715_));
 AO21x2_ASAP7_75t_R _38991_ (.A1(_09714_),
    .A2(_09715_),
    .B(_09707_),
    .Y(_09716_));
 NAND2x2_ASAP7_75t_R _38992_ (.A(net2068),
    .B(_09710_),
    .Y(_09717_));
 NAND2x2_ASAP7_75t_R _38993_ (.A(_09691_),
    .B(_09677_),
    .Y(_09718_));
 AO21x1_ASAP7_75t_R _38994_ (.A1(net1384),
    .A2(net2558),
    .B(net2959),
    .Y(_09719_));
 NAND2x1_ASAP7_75t_R _38995_ (.A(_09716_),
    .B(_09719_),
    .Y(_09721_));
 NOR2x1_ASAP7_75t_R _38996_ (.A(_09713_),
    .B(_09721_),
    .Y(_09722_));
 NOR2x1_ASAP7_75t_R _38997_ (.A(_09597_),
    .B(_09692_),
    .Y(_09723_));
 NOR2x1_ASAP7_75t_R _38998_ (.A(net3241),
    .B(net1384),
    .Y(_09724_));
 AO21x1_ASAP7_75t_R _38999_ (.A1(net1113),
    .A2(_09723_),
    .B(_09724_),
    .Y(_09725_));
 NOR2x2_ASAP7_75t_R _39000_ (.A(net2100),
    .B(_09638_),
    .Y(_09726_));
 NAND2x2_ASAP7_75t_R _39001_ (.A(net1100),
    .B(_09726_),
    .Y(_09727_));
 TAPCELL_ASAP7_75t_R PHY_250 ();
 TAPCELL_ASAP7_75t_R PHY_249 ();
 NAND2x2_ASAP7_75t_R _39004_ (.A(_09618_),
    .B(_09647_),
    .Y(_09730_));
 TAPCELL_ASAP7_75t_R PHY_248 ();
 AO21x1_ASAP7_75t_R _39006_ (.A1(_09714_),
    .A2(net1925),
    .B(_09730_),
    .Y(_09733_));
 OAI21x1_ASAP7_75t_R _39007_ (.A1(net1113),
    .A2(_09727_),
    .B(_09733_),
    .Y(_09734_));
 NOR2x1_ASAP7_75t_R _39008_ (.A(_09725_),
    .B(_09734_),
    .Y(_09735_));
 NAND2x1_ASAP7_75t_R _39009_ (.A(_09722_),
    .B(_09735_),
    .Y(_09736_));
 OAI22x1_ASAP7_75t_R _39010_ (.A1(_09727_),
    .A2(_09581_),
    .B1(net1387),
    .B2(net2547),
    .Y(_09737_));
 NAND2x2_ASAP7_75t_R _39011_ (.A(_09606_),
    .B(net1933),
    .Y(_09738_));
 NAND2x2_ASAP7_75t_R _39012_ (.A(_09629_),
    .B(_09608_),
    .Y(_09739_));
 AO21x1_ASAP7_75t_R _39013_ (.A1(net1562),
    .A2(net2047),
    .B(_09594_),
    .Y(_09740_));
 NOR2x2_ASAP7_75t_R _39014_ (.A(net1279),
    .B(net982),
    .Y(_09741_));
 INVx1_ASAP7_75t_R _39015_ (.A(_09741_),
    .Y(_09743_));
 AO21x1_ASAP7_75t_R _39016_ (.A1(_09714_),
    .A2(_09743_),
    .B(net2268),
    .Y(_09744_));
 NAND2x1_ASAP7_75t_R _39017_ (.A(_09740_),
    .B(_09744_),
    .Y(_09745_));
 NOR2x1_ASAP7_75t_R _39018_ (.A(_09737_),
    .B(_09745_),
    .Y(_09746_));
 AO21x1_ASAP7_75t_R _39019_ (.A1(net2771),
    .A2(_09592_),
    .B(_09707_),
    .Y(_09747_));
 NAND2x2_ASAP7_75t_R _39020_ (.A(_09677_),
    .B(_09648_),
    .Y(_09748_));
 NOR2x1_ASAP7_75t_R _39021_ (.A(_09592_),
    .B(net1502),
    .Y(_09749_));
 NAND2x2_ASAP7_75t_R _39022_ (.A(_09573_),
    .B(_09749_),
    .Y(_09750_));
 NAND2x1_ASAP7_75t_R _39023_ (.A(_09747_),
    .B(_09750_),
    .Y(_09751_));
 NAND2x2_ASAP7_75t_R _39024_ (.A(net1107),
    .B(net1933),
    .Y(_09752_));
 INVx2_ASAP7_75t_R _39025_ (.A(_09752_),
    .Y(_09754_));
 NAND2x2_ASAP7_75t_R _39026_ (.A(_09677_),
    .B(_09671_),
    .Y(_09755_));
 TAPCELL_ASAP7_75t_R PHY_247 ();
 CKINVDCx6p67_ASAP7_75t_R _39028_ (.A(_09755_),
    .Y(_09757_));
 NAND2x2_ASAP7_75t_R _39029_ (.A(_09754_),
    .B(_09757_),
    .Y(_09758_));
 INVx6_ASAP7_75t_R _39030_ (.A(net2959),
    .Y(_09759_));
 NAND2x2_ASAP7_75t_R _39031_ (.A(net2686),
    .B(_09759_),
    .Y(_09760_));
 NOR2x2_ASAP7_75t_R _39032_ (.A(net988),
    .B(net2817),
    .Y(_09761_));
 NAND2x1_ASAP7_75t_R _39033_ (.A(net2927),
    .B(_09761_),
    .Y(_09762_));
 NAND3x1_ASAP7_75t_R _39034_ (.A(_09758_),
    .B(_09760_),
    .C(_09762_),
    .Y(_09763_));
 NOR2x1_ASAP7_75t_R _39035_ (.A(_09751_),
    .B(_09763_),
    .Y(_09765_));
 NAND2x1_ASAP7_75t_R _39036_ (.A(_09746_),
    .B(_09765_),
    .Y(_09766_));
 NOR2x1_ASAP7_75t_R _39037_ (.A(_09766_),
    .B(_09736_),
    .Y(_09767_));
 NAND2x1_ASAP7_75t_R _39038_ (.A(_09706_),
    .B(_09767_),
    .Y(_09768_));
 NAND2x2_ASAP7_75t_R _39039_ (.A(_09662_),
    .B(net1933),
    .Y(_09769_));
 NAND2x2_ASAP7_75t_R _39040_ (.A(_09691_),
    .B(_09647_),
    .Y(_09770_));
 TAPCELL_ASAP7_75t_R PHY_246 ();
 NAND2x1_ASAP7_75t_R _39042_ (.A(net2551),
    .B(net2152),
    .Y(_09772_));
 OAI22x1_ASAP7_75t_R _39043_ (.A1(_09769_),
    .A2(net2339),
    .B1(_09772_),
    .B2(net1942),
    .Y(_09773_));
 TAPCELL_ASAP7_75t_R PHY_245 ();
 NAND2x1_ASAP7_75t_R _39045_ (.A(_09573_),
    .B(net1218),
    .Y(_09776_));
 AOI21x1_ASAP7_75t_R _39046_ (.A1(net1506),
    .A2(_09776_),
    .B(_09635_),
    .Y(_09777_));
 NOR2x1_ASAP7_75t_R _39047_ (.A(_09773_),
    .B(_09777_),
    .Y(_09778_));
 INVx6_ASAP7_75t_R _39048_ (.A(_09629_),
    .Y(_09779_));
 NAND2x1_ASAP7_75t_R _39049_ (.A(_09581_),
    .B(_09779_),
    .Y(_09780_));
 INVx1_ASAP7_75t_R _39050_ (.A(_09780_),
    .Y(_09781_));
 OAI22x1_ASAP7_75t_R _39051_ (.A1(net2291),
    .A2(_09674_),
    .B1(_09678_),
    .B2(_09597_),
    .Y(_09782_));
 NOR2x2_ASAP7_75t_R _39052_ (.A(net982),
    .B(_09779_),
    .Y(_09783_));
 OA21x2_ASAP7_75t_R _39053_ (.A1(_09783_),
    .A2(_09664_),
    .B(_09701_),
    .Y(_09784_));
 AOI21x1_ASAP7_75t_R _39054_ (.A1(_09781_),
    .A2(_09782_),
    .B(_09784_),
    .Y(_09785_));
 NAND2x1_ASAP7_75t_R _39055_ (.A(_09778_),
    .B(_09785_),
    .Y(_09787_));
 TAPCELL_ASAP7_75t_R PHY_244 ();
 TAPCELL_ASAP7_75t_R PHY_243 ();
 TAPCELL_ASAP7_75t_R PHY_242 ();
 TAPCELL_ASAP7_75t_R PHY_241 ();
 AO211x2_ASAP7_75t_R _39060_ (.A1(net2942),
    .A2(net1743),
    .B(net1282),
    .C(net3066),
    .Y(_09792_));
 NOR2x1_ASAP7_75t_R _39061_ (.A(net981),
    .B(net2914),
    .Y(_09793_));
 NOR2x1_ASAP7_75t_R _39062_ (.A(net3066),
    .B(net2775),
    .Y(_09794_));
 OAI21x1_ASAP7_75t_R _39063_ (.A1(_09793_),
    .A2(_09794_),
    .B(_09662_),
    .Y(_09795_));
 TAPCELL_ASAP7_75t_R PHY_240 ();
 NAND2x2_ASAP7_75t_R _39065_ (.A(_09629_),
    .B(net1932),
    .Y(_09798_));
 TAPCELL_ASAP7_75t_R PHY_239 ();
 TAPCELL_ASAP7_75t_R PHY_238 ();
 NAND2x2_ASAP7_75t_R _39068_ (.A(_09691_),
    .B(_09625_),
    .Y(_09801_));
 TAPCELL_ASAP7_75t_R PHY_237 ();
 AO21x2_ASAP7_75t_R _39070_ (.A1(net1246),
    .A2(net1102),
    .B(_09801_),
    .Y(_09803_));
 NAND3x2_ASAP7_75t_R _39071_ (.B(_09795_),
    .C(_09803_),
    .Y(_09804_),
    .A(_09792_));
 NOR2x2_ASAP7_75t_R _39072_ (.A(_09787_),
    .B(_09804_),
    .Y(_09805_));
 CKINVDCx6p67_ASAP7_75t_R _39073_ (.A(net1507),
    .Y(_09806_));
 CKINVDCx5p33_ASAP7_75t_R _39074_ (.A(_09770_),
    .Y(_09807_));
 NOR2x2_ASAP7_75t_R _39075_ (.A(_09581_),
    .B(_09597_),
    .Y(_09809_));
 TAPCELL_ASAP7_75t_R PHY_236 ();
 AOI22x1_ASAP7_75t_R _39077_ (.A1(_09806_),
    .A2(_09664_),
    .B1(_09807_),
    .B2(net2956),
    .Y(_09811_));
 NAND2x2_ASAP7_75t_R _39078_ (.A(_09573_),
    .B(net1100),
    .Y(_09812_));
 NOR2x1_ASAP7_75t_R _39079_ (.A(_09812_),
    .B(net1942),
    .Y(_09813_));
 AOI21x1_ASAP7_75t_R _39080_ (.A1(net2919),
    .A2(_09806_),
    .B(_09813_),
    .Y(_09814_));
 NAND2x2_ASAP7_75t_R _39081_ (.A(_09811_),
    .B(_09814_),
    .Y(_09815_));
 NOR2x2_ASAP7_75t_R _39082_ (.A(net984),
    .B(_09581_),
    .Y(_09816_));
 INVx5_ASAP7_75t_R _39083_ (.A(_09816_),
    .Y(_09817_));
 TAPCELL_ASAP7_75t_R PHY_235 ();
 TAPCELL_ASAP7_75t_R PHY_234 ();
 AO21x1_ASAP7_75t_R _39086_ (.A1(_09817_),
    .A2(net2048),
    .B(net1942),
    .Y(_09821_));
 NOR2x2_ASAP7_75t_R _39087_ (.A(_09579_),
    .B(_09779_),
    .Y(_09822_));
 TAPCELL_ASAP7_75t_R PHY_233 ();
 TAPCELL_ASAP7_75t_R PHY_232 ();
 NAND2x2_ASAP7_75t_R _39090_ (.A(net3069),
    .B(net2453),
    .Y(_09825_));
 INVx8_ASAP7_75t_R _39091_ (.A(_09801_),
    .Y(_09826_));
 TAPCELL_ASAP7_75t_R PHY_231 ();
 OAI21x1_ASAP7_75t_R _39093_ (.A1(net2941),
    .A2(_09825_),
    .B(_09826_),
    .Y(_09828_));
 NAND2x2_ASAP7_75t_R _39094_ (.A(_09821_),
    .B(_09828_),
    .Y(_09829_));
 AO21x1_ASAP7_75t_R _39095_ (.A1(_09748_),
    .A2(_09678_),
    .B(net2732),
    .Y(_09831_));
 NOR2x2_ASAP7_75t_R _39096_ (.A(_09674_),
    .B(net2552),
    .Y(_09832_));
 TAPCELL_ASAP7_75t_R PHY_230 ();
 AOI22x1_ASAP7_75t_R _39098_ (.A1(_09832_),
    .A2(_09726_),
    .B1(_09664_),
    .B2(net2927),
    .Y(_09834_));
 NAND2x2_ASAP7_75t_R _39099_ (.A(_09831_),
    .B(_09834_),
    .Y(_09835_));
 NOR3x2_ASAP7_75t_R _39100_ (.B(_09829_),
    .C(_09835_),
    .Y(_09836_),
    .A(_09815_));
 NAND2x2_ASAP7_75t_R _39101_ (.A(net2930),
    .B(_09670_),
    .Y(_09837_));
 NOR2x2_ASAP7_75t_R _39102_ (.A(_09585_),
    .B(_09837_),
    .Y(_09838_));
 OA21x2_ASAP7_75t_R _39103_ (.A1(_09822_),
    .A2(_09582_),
    .B(_09838_),
    .Y(_09839_));
 TAPCELL_ASAP7_75t_R PHY_229 ();
 TAPCELL_ASAP7_75t_R PHY_228 ();
 OAI22x1_ASAP7_75t_R _39106_ (.A1(_09613_),
    .A2(net3016),
    .B1(net3241),
    .B2(net2103),
    .Y(_09843_));
 NOR2x1_ASAP7_75t_R _39107_ (.A(_09839_),
    .B(_09843_),
    .Y(_09844_));
 AND4x1_ASAP7_75t_R _39108_ (.A(_09608_),
    .B(_09625_),
    .C(_09662_),
    .D(_09691_),
    .Y(_09845_));
 NOR2x2_ASAP7_75t_R _39109_ (.A(net1843),
    .B(_09639_),
    .Y(_09846_));
 AND3x1_ASAP7_75t_R _39110_ (.A(_09846_),
    .B(net1282),
    .C(_09608_),
    .Y(_09847_));
 NOR2x1_ASAP7_75t_R _39111_ (.A(_09845_),
    .B(_09847_),
    .Y(_09848_));
 NAND2x1_ASAP7_75t_R _39112_ (.A(_09844_),
    .B(_09848_),
    .Y(_09849_));
 TAPCELL_ASAP7_75t_R PHY_227 ();
 TAPCELL_ASAP7_75t_R PHY_226 ();
 OAI22x1_ASAP7_75t_R _39115_ (.A1(net1246),
    .A2(net1998),
    .B1(net1477),
    .B2(net1868),
    .Y(_09853_));
 NAND2x2_ASAP7_75t_R _39116_ (.A(_09589_),
    .B(net1933),
    .Y(_09854_));
 OAI22x1_ASAP7_75t_R _39117_ (.A1(net2656),
    .A2(net1577),
    .B1(net1743),
    .B2(_09854_),
    .Y(_09855_));
 NOR2x1_ASAP7_75t_R _39118_ (.A(_09853_),
    .B(_09855_),
    .Y(_09856_));
 OAI22x1_ASAP7_75t_R _39119_ (.A1(_09649_),
    .A2(_09769_),
    .B1(_09730_),
    .B2(_09644_),
    .Y(_09857_));
 NAND2x2_ASAP7_75t_R _39120_ (.A(net2550),
    .B(_09608_),
    .Y(_09858_));
 NAND2x2_ASAP7_75t_R _39121_ (.A(_09700_),
    .B(_09759_),
    .Y(_09859_));
 OAI21x1_ASAP7_75t_R _39122_ (.A1(net2085),
    .A2(_09858_),
    .B(_09859_),
    .Y(_09860_));
 NOR2x1_ASAP7_75t_R _39123_ (.A(_09857_),
    .B(_09860_),
    .Y(_09861_));
 NAND2x2_ASAP7_75t_R _39124_ (.A(_09856_),
    .B(_09861_),
    .Y(_09862_));
 NOR2x2_ASAP7_75t_R _39125_ (.A(_09849_),
    .B(_09862_),
    .Y(_09864_));
 NAND3x2_ASAP7_75t_R _39126_ (.B(_09836_),
    .C(_09864_),
    .Y(_09865_),
    .A(_09805_));
 NOR2x2_ASAP7_75t_R _39127_ (.A(_09768_),
    .B(_09865_),
    .Y(_09866_));
 NAND2x2_ASAP7_75t_R _39128_ (.A(net1493),
    .B(_09866_),
    .Y(_09867_));
 TAPCELL_ASAP7_75t_R PHY_225 ();
 TAPCELL_ASAP7_75t_R PHY_224 ();
 INVx3_ASAP7_75t_R _39131_ (.A(net2830),
    .Y(_09870_));
 NAND2x2_ASAP7_75t_R _39132_ (.A(_00649_),
    .B(_09870_),
    .Y(_09871_));
 TAPCELL_ASAP7_75t_R PHY_223 ();
 INVx2_ASAP7_75t_R _39134_ (.A(_00652_),
    .Y(_09873_));
 NAND2x2_ASAP7_75t_R _39135_ (.A(net3159),
    .B(_09873_),
    .Y(_09875_));
 NOR2x2_ASAP7_75t_R _39136_ (.A(_09871_),
    .B(_09875_),
    .Y(_09876_));
 TAPCELL_ASAP7_75t_R PHY_222 ();
 NOR2x2_ASAP7_75t_R _39138_ (.A(_00653_),
    .B(_00654_),
    .Y(_09878_));
 TAPCELL_ASAP7_75t_R PHY_221 ();
 TAPCELL_ASAP7_75t_R PHY_220 ();
 NOR2x2_ASAP7_75t_R _39141_ (.A(net1015),
    .B(net1161),
    .Y(_09881_));
 NAND2x2_ASAP7_75t_R _39142_ (.A(net1247),
    .B(_09881_),
    .Y(_09882_));
 INVx3_ASAP7_75t_R _39143_ (.A(_09882_),
    .Y(_09883_));
 NAND2x2_ASAP7_75t_R _39144_ (.A(_09876_),
    .B(_09883_),
    .Y(_09884_));
 INVx3_ASAP7_75t_R _39145_ (.A(_00654_),
    .Y(_09886_));
 NOR2x2_ASAP7_75t_R _39146_ (.A(net2564),
    .B(_09886_),
    .Y(_09887_));
 CKINVDCx20_ASAP7_75t_R _39147_ (.A(net1017),
    .Y(_09888_));
 NOR2x2_ASAP7_75t_R _39148_ (.A(net1159),
    .B(_09888_),
    .Y(_09889_));
 NAND2x2_ASAP7_75t_R _39149_ (.A(net1699),
    .B(net2470),
    .Y(_09890_));
 TAPCELL_ASAP7_75t_R PHY_219 ();
 CKINVDCx16_ASAP7_75t_R _39151_ (.A(net1159),
    .Y(_09892_));
 NOR2x2_ASAP7_75t_R _39152_ (.A(net1019),
    .B(_09892_),
    .Y(_09893_));
 TAPCELL_ASAP7_75t_R PHY_218 ();
 NAND2x2_ASAP7_75t_R _39154_ (.A(net1699),
    .B(_09893_),
    .Y(_09895_));
 INVx2_ASAP7_75t_R _39155_ (.A(_00649_),
    .Y(_09897_));
 NOR2x2_ASAP7_75t_R _39156_ (.A(net2831),
    .B(_09897_),
    .Y(_09898_));
 INVx2_ASAP7_75t_R _39157_ (.A(_00651_),
    .Y(_09899_));
 NOR2x2_ASAP7_75t_R _39158_ (.A(_00652_),
    .B(_09899_),
    .Y(_09900_));
 NAND2x2_ASAP7_75t_R _39159_ (.A(_09898_),
    .B(_09900_),
    .Y(_09901_));
 AO21x1_ASAP7_75t_R _39160_ (.A1(net945),
    .A2(_09895_),
    .B(_09901_),
    .Y(_09902_));
 NAND2x1_ASAP7_75t_R _39161_ (.A(_09884_),
    .B(_09902_),
    .Y(_09903_));
 NAND2x2_ASAP7_75t_R _39162_ (.A(_00653_),
    .B(_00654_),
    .Y(_09904_));
 CKINVDCx8_ASAP7_75t_R _39163_ (.A(net1353),
    .Y(_09905_));
 NAND2x2_ASAP7_75t_R _39164_ (.A(net1028),
    .B(_09905_),
    .Y(_09906_));
 NAND2x2_ASAP7_75t_R _39165_ (.A(net976),
    .B(_09905_),
    .Y(_09908_));
 AO21x1_ASAP7_75t_R _39166_ (.A1(_09906_),
    .A2(net2444),
    .B(_09901_),
    .Y(_09909_));
 INVx3_ASAP7_75t_R _39167_ (.A(net3074),
    .Y(_09910_));
 NOR2x2_ASAP7_75t_R _39168_ (.A(net2838),
    .B(_09910_),
    .Y(_09911_));
 TAPCELL_ASAP7_75t_R PHY_217 ();
 NAND2x2_ASAP7_75t_R _39170_ (.A(_09893_),
    .B(net2282),
    .Y(_09913_));
 NAND2x2_ASAP7_75t_R _39171_ (.A(net2049),
    .B(_09911_),
    .Y(_09914_));
 AO21x1_ASAP7_75t_R _39172_ (.A1(_09913_),
    .A2(net2356),
    .B(_09901_),
    .Y(_09915_));
 NAND2x1_ASAP7_75t_R _39173_ (.A(_09909_),
    .B(_09915_),
    .Y(_09916_));
 NOR2x1_ASAP7_75t_R _39174_ (.A(_09903_),
    .B(_09916_),
    .Y(_09917_));
 NAND2x2_ASAP7_75t_R _39175_ (.A(net2192),
    .B(net1699),
    .Y(_09919_));
 NAND2x2_ASAP7_75t_R _39176_ (.A(_00651_),
    .B(_00652_),
    .Y(_09920_));
 INVx3_ASAP7_75t_R _39177_ (.A(_09920_),
    .Y(_09921_));
 NAND2x2_ASAP7_75t_R _39178_ (.A(_09898_),
    .B(_09921_),
    .Y(_09922_));
 AO21x1_ASAP7_75t_R _39179_ (.A1(net2213),
    .A2(net2936),
    .B(net2660),
    .Y(_09923_));
 TAPCELL_ASAP7_75t_R PHY_216 ();
 NAND2x2_ASAP7_75t_R _39181_ (.A(net2192),
    .B(_09911_),
    .Y(_09925_));
 AO21x1_ASAP7_75t_R _39182_ (.A1(_09906_),
    .A2(net3059),
    .B(_09922_),
    .Y(_09926_));
 TAPCELL_ASAP7_75t_R PHY_215 ();
 NAND2x2_ASAP7_75t_R _39184_ (.A(net1250),
    .B(net2470),
    .Y(_09928_));
 AO21x1_ASAP7_75t_R _39185_ (.A1(_09928_),
    .A2(net3245),
    .B(_09922_),
    .Y(_09930_));
 AND3x1_ASAP7_75t_R _39186_ (.A(_09923_),
    .B(_09926_),
    .C(_09930_),
    .Y(_09931_));
 NAND2x1_ASAP7_75t_R _39187_ (.A(_09917_),
    .B(_09931_),
    .Y(_09932_));
 NAND2x2_ASAP7_75t_R _39188_ (.A(net1013),
    .B(net1159),
    .Y(_09933_));
 CKINVDCx12_ASAP7_75t_R _39189_ (.A(net1249),
    .Y(_09934_));
 TAPCELL_ASAP7_75t_R PHY_214 ();
 NOR2x2_ASAP7_75t_R _39191_ (.A(_00651_),
    .B(_00652_),
    .Y(_09936_));
 NAND2x2_ASAP7_75t_R _39192_ (.A(_09936_),
    .B(_09898_),
    .Y(_09937_));
 NOR2x2_ASAP7_75t_R _39193_ (.A(_09934_),
    .B(_09937_),
    .Y(_09938_));
 NAND2x2_ASAP7_75t_R _39194_ (.A(net2837),
    .B(_09910_),
    .Y(_09939_));
 NOR2x2_ASAP7_75t_R _39195_ (.A(_09888_),
    .B(_09939_),
    .Y(_09941_));
 INVx4_ASAP7_75t_R _39196_ (.A(_09936_),
    .Y(_09942_));
 NOR2x2_ASAP7_75t_R _39197_ (.A(_09871_),
    .B(_09942_),
    .Y(_09943_));
 NAND2x2_ASAP7_75t_R _39198_ (.A(_09941_),
    .B(_09943_),
    .Y(_09944_));
 NAND2x2_ASAP7_75t_R _39199_ (.A(net1160),
    .B(_09888_),
    .Y(_09945_));
 NOR2x2_ASAP7_75t_R _39200_ (.A(_09939_),
    .B(_09945_),
    .Y(_09946_));
 NAND2x2_ASAP7_75t_R _39201_ (.A(_09946_),
    .B(net1951),
    .Y(_09947_));
 NAND2x2_ASAP7_75t_R _39202_ (.A(_09944_),
    .B(_09947_),
    .Y(_09948_));
 AOI21x1_ASAP7_75t_R _39203_ (.A1(net1065),
    .A2(_09938_),
    .B(_09948_),
    .Y(_09949_));
 NAND2x2_ASAP7_75t_R _39204_ (.A(net3017),
    .B(net1248),
    .Y(_09950_));
 NOR2x2_ASAP7_75t_R _39205_ (.A(_00651_),
    .B(_09873_),
    .Y(_09952_));
 NAND2x2_ASAP7_75t_R _39206_ (.A(_09898_),
    .B(_09952_),
    .Y(_09953_));
 AO21x1_ASAP7_75t_R _39207_ (.A1(net947),
    .A2(_09950_),
    .B(_09953_),
    .Y(_09954_));
 TAPCELL_ASAP7_75t_R PHY_213 ();
 AO21x1_ASAP7_75t_R _39209_ (.A1(net3059),
    .A2(net1351),
    .B(_09953_),
    .Y(_09956_));
 AND2x2_ASAP7_75t_R _39210_ (.A(_09954_),
    .B(_09956_),
    .Y(_09957_));
 NAND2x2_ASAP7_75t_R _39211_ (.A(net2564),
    .B(_09886_),
    .Y(_09958_));
 NOR2x2_ASAP7_75t_R _39212_ (.A(net3017),
    .B(net1703),
    .Y(_09959_));
 TAPCELL_ASAP7_75t_R PHY_212 ();
 NOR2x2_ASAP7_75t_R _39214_ (.A(net1162),
    .B(net1353),
    .Y(_09961_));
 INVx3_ASAP7_75t_R _39215_ (.A(_09961_),
    .Y(_09963_));
 NOR2x1_ASAP7_75t_R _39216_ (.A(_09937_),
    .B(_09963_),
    .Y(_09964_));
 NOR2x1_ASAP7_75t_R _39217_ (.A(net3059),
    .B(_09937_),
    .Y(_09965_));
 AOI211x1_ASAP7_75t_R _39218_ (.A1(_09959_),
    .A2(net1951),
    .B(_09964_),
    .C(_09965_),
    .Y(_09966_));
 NAND3x1_ASAP7_75t_R _39219_ (.A(_09949_),
    .B(_09957_),
    .C(_09966_),
    .Y(_09967_));
 NOR2x1_ASAP7_75t_R _39220_ (.A(_09932_),
    .B(_09967_),
    .Y(_09968_));
 NAND2x2_ASAP7_75t_R _39221_ (.A(_00655_),
    .B(_09892_),
    .Y(_09969_));
 NOR2x2_ASAP7_75t_R _39222_ (.A(_09969_),
    .B(_09934_),
    .Y(_09970_));
 NAND2x2_ASAP7_75t_R _39223_ (.A(_00649_),
    .B(net2830),
    .Y(_09971_));
 NAND2x2_ASAP7_75t_R _39224_ (.A(_00652_),
    .B(_09899_),
    .Y(_09972_));
 NOR2x2_ASAP7_75t_R _39225_ (.A(net2584),
    .B(_09972_),
    .Y(_09974_));
 TAPCELL_ASAP7_75t_R PHY_211 ();
 TAPCELL_ASAP7_75t_R PHY_210 ();
 TAPCELL_ASAP7_75t_R PHY_209 ();
 NOR2x2_ASAP7_75t_R _39229_ (.A(net1016),
    .B(net1703),
    .Y(_09978_));
 NOR2x2_ASAP7_75t_R _39230_ (.A(net1353),
    .B(net979),
    .Y(_09979_));
 OA21x2_ASAP7_75t_R _39231_ (.A1(_09978_),
    .A2(_09979_),
    .B(net2430),
    .Y(_09980_));
 NOR2x2_ASAP7_75t_R _39232_ (.A(_09939_),
    .B(_09969_),
    .Y(_09981_));
 NOR2x2_ASAP7_75t_R _39233_ (.A(net1015),
    .B(_09939_),
    .Y(_09982_));
 OA21x2_ASAP7_75t_R _39234_ (.A1(_09981_),
    .A2(_09982_),
    .B(net2430),
    .Y(_09983_));
 AOI211x1_ASAP7_75t_R _39235_ (.A1(_09970_),
    .A2(net2430),
    .B(_09980_),
    .C(_09983_),
    .Y(_09985_));
 TAPCELL_ASAP7_75t_R PHY_208 ();
 NOR2x2_ASAP7_75t_R _39237_ (.A(net1162),
    .B(net1704),
    .Y(_09987_));
 INVx2_ASAP7_75t_R _39238_ (.A(_09987_),
    .Y(_09988_));
 INVx3_ASAP7_75t_R _39239_ (.A(_09971_),
    .Y(_09989_));
 NAND2x2_ASAP7_75t_R _39240_ (.A(net2866),
    .B(_09989_),
    .Y(_09990_));
 AO21x1_ASAP7_75t_R _39241_ (.A1(_09988_),
    .A2(_09963_),
    .B(_09990_),
    .Y(_09991_));
 NOR2x2_ASAP7_75t_R _39242_ (.A(_09971_),
    .B(_09942_),
    .Y(_09992_));
 NAND2x1_ASAP7_75t_R _39243_ (.A(_09982_),
    .B(_09992_),
    .Y(_09993_));
 AND2x6_ASAP7_75t_R _39244_ (.A(net1164),
    .B(net1018),
    .Y(_09994_));
 NAND2x2_ASAP7_75t_R _39245_ (.A(net1247),
    .B(_09994_),
    .Y(_09996_));
 TAPCELL_ASAP7_75t_R PHY_207 ();
 NAND2x2_ASAP7_75t_R _39247_ (.A(net1250),
    .B(_09893_),
    .Y(_09998_));
 TAPCELL_ASAP7_75t_R PHY_206 ();
 AO21x1_ASAP7_75t_R _39249_ (.A1(net2409),
    .A2(_09998_),
    .B(_09990_),
    .Y(_10000_));
 AND3x1_ASAP7_75t_R _39250_ (.A(_09991_),
    .B(_09993_),
    .C(_10000_),
    .Y(_10001_));
 NAND2x1_ASAP7_75t_R _39251_ (.A(_09985_),
    .B(_10001_),
    .Y(_10002_));
 NAND2x2_ASAP7_75t_R _39252_ (.A(net1017),
    .B(net1247),
    .Y(_10003_));
 NOR2x2_ASAP7_75t_R _39253_ (.A(_09920_),
    .B(_09971_),
    .Y(_10004_));
 CKINVDCx10_ASAP7_75t_R _39254_ (.A(_10004_),
    .Y(_10005_));
 AO21x1_ASAP7_75t_R _39255_ (.A1(_10003_),
    .A2(net2235),
    .B(_10005_),
    .Y(_10007_));
 NAND2x2_ASAP7_75t_R _39256_ (.A(_09911_),
    .B(_09994_),
    .Y(_10008_));
 AO21x1_ASAP7_75t_R _39257_ (.A1(_10008_),
    .A2(net3059),
    .B(_10005_),
    .Y(_10009_));
 NAND2x1_ASAP7_75t_R _39258_ (.A(_10007_),
    .B(_10009_),
    .Y(_10010_));
 NAND2x2_ASAP7_75t_R _39259_ (.A(_09900_),
    .B(_09989_),
    .Y(_10011_));
 AO21x2_ASAP7_75t_R _39260_ (.A1(_10008_),
    .A2(net3059),
    .B(_10011_),
    .Y(_10012_));
 NAND2x2_ASAP7_75t_R _39261_ (.A(_09893_),
    .B(_09905_),
    .Y(_10013_));
 NOR2x2_ASAP7_75t_R _39262_ (.A(net3017),
    .B(net1353),
    .Y(_10014_));
 INVx4_ASAP7_75t_R _39263_ (.A(_10014_),
    .Y(_10015_));
 AO21x1_ASAP7_75t_R _39264_ (.A1(net1962),
    .A2(_10015_),
    .B(_10011_),
    .Y(_10016_));
 NAND2x1_ASAP7_75t_R _39265_ (.A(_10012_),
    .B(_10016_),
    .Y(_10018_));
 TAPCELL_ASAP7_75t_R PHY_205 ();
 NOR2x1_ASAP7_75t_R _39267_ (.A(net1796),
    .B(_10011_),
    .Y(_10020_));
 INVx1_ASAP7_75t_R _39268_ (.A(_10020_),
    .Y(_10021_));
 AO21x1_ASAP7_75t_R _39269_ (.A1(_10003_),
    .A2(net3245),
    .B(_10011_),
    .Y(_10022_));
 NAND2x1_ASAP7_75t_R _39270_ (.A(_10021_),
    .B(_10022_),
    .Y(_10023_));
 OR3x1_ASAP7_75t_R _39271_ (.A(_10010_),
    .B(_10018_),
    .C(_10023_),
    .Y(_10024_));
 NOR2x1_ASAP7_75t_R _39272_ (.A(_10024_),
    .B(_10002_),
    .Y(_10025_));
 NAND2x1_ASAP7_75t_R _39273_ (.A(_09968_),
    .B(_10025_),
    .Y(_10026_));
 NOR2x2_ASAP7_75t_R _39274_ (.A(_09933_),
    .B(net1354),
    .Y(_10027_));
 NAND2x2_ASAP7_75t_R _39275_ (.A(net2830),
    .B(_09897_),
    .Y(_10029_));
 NOR2x2_ASAP7_75t_R _39276_ (.A(_09972_),
    .B(_10029_),
    .Y(_10030_));
 NAND2x1_ASAP7_75t_R _39277_ (.A(_10027_),
    .B(_10030_),
    .Y(_10031_));
 INVx2_ASAP7_75t_R _39278_ (.A(_10031_),
    .Y(_10032_));
 TAPCELL_ASAP7_75t_R PHY_204 ();
 NOR2x2_ASAP7_75t_R _39280_ (.A(_00649_),
    .B(_09870_),
    .Y(_10034_));
 NAND2x2_ASAP7_75t_R _39281_ (.A(_09952_),
    .B(_10034_),
    .Y(_10035_));
 AOI221x1_ASAP7_75t_R _39282_ (.A1(net3015),
    .A2(_09892_),
    .B1(net1801),
    .B2(_09934_),
    .C(_10035_),
    .Y(_10036_));
 NOR2x1_ASAP7_75t_R _39283_ (.A(_10032_),
    .B(_10036_),
    .Y(_10037_));
 NAND2x2_ASAP7_75t_R _39284_ (.A(net1021),
    .B(net2284),
    .Y(_10038_));
 NAND2x2_ASAP7_75t_R _39285_ (.A(net2867),
    .B(_10034_),
    .Y(_10040_));
 AO21x1_ASAP7_75t_R _39286_ (.A1(_10038_),
    .A2(_09925_),
    .B(_10040_),
    .Y(_10041_));
 NAND2x2_ASAP7_75t_R _39287_ (.A(net3017),
    .B(net1699),
    .Y(_10042_));
 AO21x1_ASAP7_75t_R _39288_ (.A1(_09998_),
    .A2(_10042_),
    .B(_10040_),
    .Y(_10043_));
 NOR2x2_ASAP7_75t_R _39289_ (.A(_10029_),
    .B(_09942_),
    .Y(_10044_));
 NAND2x1_ASAP7_75t_R _39290_ (.A(_10014_),
    .B(_10044_),
    .Y(_10045_));
 AND3x1_ASAP7_75t_R _39291_ (.A(_10041_),
    .B(_10043_),
    .C(_10045_),
    .Y(_10046_));
 NAND2x1_ASAP7_75t_R _39292_ (.A(_10037_),
    .B(_10046_),
    .Y(_10047_));
 NAND2x2_ASAP7_75t_R _39293_ (.A(_09900_),
    .B(_10034_),
    .Y(_10048_));
 TAPCELL_ASAP7_75t_R PHY_203 ();
 AO21x1_ASAP7_75t_R _39295_ (.A1(net2397),
    .A2(_09882_),
    .B(_10048_),
    .Y(_10051_));
 AO21x2_ASAP7_75t_R _39296_ (.A1(net2037),
    .A2(_09895_),
    .B(_10048_),
    .Y(_10052_));
 NAND2x1_ASAP7_75t_R _39297_ (.A(_10051_),
    .B(_10052_),
    .Y(_10053_));
 AO21x1_ASAP7_75t_R _39298_ (.A1(_09906_),
    .A2(net2444),
    .B(_10048_),
    .Y(_10054_));
 AO21x1_ASAP7_75t_R _39299_ (.A1(_09913_),
    .A2(_09925_),
    .B(_10048_),
    .Y(_10055_));
 NAND2x1_ASAP7_75t_R _39300_ (.A(_10054_),
    .B(_10055_),
    .Y(_10056_));
 NOR2x1_ASAP7_75t_R _39301_ (.A(_10053_),
    .B(_10056_),
    .Y(_10057_));
 INVx6_ASAP7_75t_R _39302_ (.A(net977),
    .Y(_10058_));
 AO21x2_ASAP7_75t_R _39303_ (.A1(_10058_),
    .A2(net1066),
    .B(_09904_),
    .Y(_10059_));
 NAND2x2_ASAP7_75t_R _39304_ (.A(_10034_),
    .B(_09921_),
    .Y(_10060_));
 AO21x1_ASAP7_75t_R _39305_ (.A1(_10059_),
    .A2(net2357),
    .B(_10060_),
    .Y(_10062_));
 NAND2x2_ASAP7_75t_R _39306_ (.A(net1699),
    .B(_09994_),
    .Y(_10063_));
 AO21x1_ASAP7_75t_R _39307_ (.A1(_10063_),
    .A2(_09890_),
    .B(_10060_),
    .Y(_10064_));
 AND2x2_ASAP7_75t_R _39308_ (.A(_10062_),
    .B(_10064_),
    .Y(_10065_));
 NAND2x2_ASAP7_75t_R _39309_ (.A(_10057_),
    .B(_10065_),
    .Y(_10066_));
 NOR2x2_ASAP7_75t_R _39310_ (.A(_10047_),
    .B(_10066_),
    .Y(_10067_));
 TAPCELL_ASAP7_75t_R PHY_202 ();
 NOR2x2_ASAP7_75t_R _39312_ (.A(_00649_),
    .B(net2830),
    .Y(_10069_));
 NAND2x2_ASAP7_75t_R _39313_ (.A(_10069_),
    .B(_09936_),
    .Y(_10070_));
 CKINVDCx8_ASAP7_75t_R _39314_ (.A(_10070_),
    .Y(_10071_));
 NAND2x2_ASAP7_75t_R _39315_ (.A(net1247),
    .B(_10071_),
    .Y(_10073_));
 NOR2x2_ASAP7_75t_R _39316_ (.A(net2252),
    .B(net2374),
    .Y(_10074_));
 INVx1_ASAP7_75t_R _39317_ (.A(_10074_),
    .Y(_10075_));
 OAI21x1_ASAP7_75t_R _39318_ (.A1(net3309),
    .A2(_10073_),
    .B(_10075_),
    .Y(_10076_));
 NOR2x2_ASAP7_75t_R _39319_ (.A(net1355),
    .B(_09969_),
    .Y(_10077_));
 OAI21x1_ASAP7_75t_R _39320_ (.A1(_10027_),
    .A2(_10077_),
    .B(_10071_),
    .Y(_10078_));
 NAND2x2_ASAP7_75t_R _39321_ (.A(_09959_),
    .B(_10071_),
    .Y(_10079_));
 NOR2x2_ASAP7_75t_R _39322_ (.A(net1354),
    .B(_09945_),
    .Y(_10080_));
 NAND2x1_ASAP7_75t_R _39323_ (.A(_10080_),
    .B(_10071_),
    .Y(_10081_));
 NAND3x1_ASAP7_75t_R _39324_ (.A(_10078_),
    .B(_10079_),
    .C(_10081_),
    .Y(_10082_));
 NOR2x1_ASAP7_75t_R _39325_ (.A(_10076_),
    .B(_10082_),
    .Y(_10084_));
 NAND2x2_ASAP7_75t_R _39326_ (.A(net3017),
    .B(net2285),
    .Y(_10085_));
 NAND2x2_ASAP7_75t_R _39327_ (.A(_10069_),
    .B(_09952_),
    .Y(_10086_));
 AO21x1_ASAP7_75t_R _39328_ (.A1(_09914_),
    .A2(_10085_),
    .B(net3244),
    .Y(_10087_));
 TAPCELL_ASAP7_75t_R PHY_201 ();
 AO21x1_ASAP7_75t_R _39330_ (.A1(_10013_),
    .A2(_10015_),
    .B(net3244),
    .Y(_10089_));
 NAND2x1_ASAP7_75t_R _39331_ (.A(_10087_),
    .B(_10089_),
    .Y(_10090_));
 AO21x1_ASAP7_75t_R _39332_ (.A1(net2408),
    .A2(_09882_),
    .B(_10086_),
    .Y(_10091_));
 OR3x1_ASAP7_75t_R _39333_ (.A(_10086_),
    .B(net1798),
    .C(net2049),
    .Y(_10092_));
 NAND2x1_ASAP7_75t_R _39334_ (.A(_10091_),
    .B(_10092_),
    .Y(_10093_));
 NOR2x1_ASAP7_75t_R _39335_ (.A(_10090_),
    .B(_10093_),
    .Y(_10095_));
 NAND2x1_ASAP7_75t_R _39336_ (.A(_10084_),
    .B(_10095_),
    .Y(_10096_));
 NOR2x2_ASAP7_75t_R _39337_ (.A(_09945_),
    .B(net1703),
    .Y(_10097_));
 NAND2x2_ASAP7_75t_R _39338_ (.A(_10069_),
    .B(_09900_),
    .Y(_10098_));
 INVx8_ASAP7_75t_R _39339_ (.A(_10098_),
    .Y(_10099_));
 OA21x2_ASAP7_75t_R _39340_ (.A1(net2583),
    .A2(_10080_),
    .B(_10099_),
    .Y(_10100_));
 TAPCELL_ASAP7_75t_R PHY_200 ();
 AOI21x1_ASAP7_75t_R _39342_ (.A1(_09882_),
    .A2(_10003_),
    .B(net2535),
    .Y(_10102_));
 NOR2x1_ASAP7_75t_R _39343_ (.A(net3093),
    .B(net1660),
    .Y(_10103_));
 NOR3x1_ASAP7_75t_R _39344_ (.A(_10100_),
    .B(_10102_),
    .C(_10103_),
    .Y(_10104_));
 NAND2x2_ASAP7_75t_R _39345_ (.A(_10069_),
    .B(_09921_),
    .Y(_10106_));
 INVx4_ASAP7_75t_R _39346_ (.A(_10027_),
    .Y(_10107_));
 NOR2x1_ASAP7_75t_R _39347_ (.A(net2628),
    .B(_10107_),
    .Y(_10108_));
 AOI211x1_ASAP7_75t_R _39348_ (.A1(net1023),
    .A2(net1166),
    .B(net1703),
    .C(net2628),
    .Y(_10109_));
 NOR2x1_ASAP7_75t_R _39349_ (.A(_10108_),
    .B(_10109_),
    .Y(_10110_));
 NAND2x2_ASAP7_75t_R _39350_ (.A(net1017),
    .B(net1699),
    .Y(_10111_));
 NOR2x2_ASAP7_75t_R _39351_ (.A(_10111_),
    .B(net2629),
    .Y(_10112_));
 INVx2_ASAP7_75t_R _39352_ (.A(_09950_),
    .Y(_10113_));
 INVx3_ASAP7_75t_R _39353_ (.A(net3064),
    .Y(_10114_));
 OA21x2_ASAP7_75t_R _39354_ (.A1(_10113_),
    .A2(_09970_),
    .B(_10114_),
    .Y(_10115_));
 NOR2x1_ASAP7_75t_R _39355_ (.A(_10112_),
    .B(_10115_),
    .Y(_10117_));
 NAND3x1_ASAP7_75t_R _39356_ (.A(_10104_),
    .B(_10110_),
    .C(_10117_),
    .Y(_10118_));
 NOR2x1_ASAP7_75t_R _39357_ (.A(_10118_),
    .B(_10096_),
    .Y(_10119_));
 NAND2x2_ASAP7_75t_R _39358_ (.A(_10067_),
    .B(_10119_),
    .Y(_10120_));
 NOR2x2_ASAP7_75t_R _39359_ (.A(_10026_),
    .B(_10120_),
    .Y(_10121_));
 NOR2x2_ASAP7_75t_R _39360_ (.A(_09871_),
    .B(_09972_),
    .Y(_10122_));
 NAND2x1_ASAP7_75t_R _39361_ (.A(net2382),
    .B(_10113_),
    .Y(_10123_));
 NAND2x1_ASAP7_75t_R _39362_ (.A(_09941_),
    .B(_09992_),
    .Y(_10124_));
 AO21x2_ASAP7_75t_R _39363_ (.A1(_10123_),
    .A2(_10124_),
    .B(net3309),
    .Y(_10125_));
 NOR2x2_ASAP7_75t_R _39364_ (.A(net1065),
    .B(net1704),
    .Y(_10126_));
 TAPCELL_ASAP7_75t_R PHY_199 ();
 OAI21x1_ASAP7_75t_R _39366_ (.A1(_10126_),
    .A2(net2222),
    .B(net2382),
    .Y(_10129_));
 NAND2x2_ASAP7_75t_R _39367_ (.A(_09987_),
    .B(net2280),
    .Y(_10130_));
 NAND3x2_ASAP7_75t_R _39368_ (.B(_10129_),
    .C(_10130_),
    .Y(_10131_),
    .A(_10125_));
 NAND2x1_ASAP7_75t_R _39369_ (.A(_09978_),
    .B(_09876_),
    .Y(_10132_));
 NOR2x2_ASAP7_75t_R _39370_ (.A(_09920_),
    .B(_09871_),
    .Y(_10133_));
 NAND2x1_ASAP7_75t_R _39371_ (.A(_10014_),
    .B(_10133_),
    .Y(_10134_));
 NAND2x1_ASAP7_75t_R _39372_ (.A(net1893),
    .B(_09978_),
    .Y(_10135_));
 AND3x1_ASAP7_75t_R _39373_ (.A(_10132_),
    .B(_10134_),
    .C(_10135_),
    .Y(_10136_));
 NAND2x2_ASAP7_75t_R _39374_ (.A(_09892_),
    .B(net1247),
    .Y(_10137_));
 INVx1_ASAP7_75t_R _39375_ (.A(_10137_),
    .Y(_10139_));
 CKINVDCx6p67_ASAP7_75t_R _39376_ (.A(_10086_),
    .Y(_10140_));
 NAND2x1_ASAP7_75t_R _39377_ (.A(_10139_),
    .B(_10140_),
    .Y(_10141_));
 OAI21x1_ASAP7_75t_R _39378_ (.A1(_09950_),
    .A2(_10048_),
    .B(_10141_),
    .Y(_10142_));
 INVx2_ASAP7_75t_R _39379_ (.A(_09919_),
    .Y(_10143_));
 NOR2x2_ASAP7_75t_R _39380_ (.A(_09920_),
    .B(_10029_),
    .Y(_10144_));
 TAPCELL_ASAP7_75t_R PHY_198 ();
 AO21x1_ASAP7_75t_R _39382_ (.A1(_10143_),
    .A2(net2805),
    .B(_09964_),
    .Y(_10146_));
 NOR2x1_ASAP7_75t_R _39383_ (.A(_10142_),
    .B(_10146_),
    .Y(_10147_));
 NAND2x1_ASAP7_75t_R _39384_ (.A(_10136_),
    .B(_10147_),
    .Y(_10148_));
 NOR2x2_ASAP7_75t_R _39385_ (.A(_10131_),
    .B(_10148_),
    .Y(_10150_));
 AOI22x1_ASAP7_75t_R _39386_ (.A1(_09992_),
    .A2(net2222),
    .B1(_10027_),
    .B2(net2804),
    .Y(_10151_));
 NOR2x2_ASAP7_75t_R _39387_ (.A(net1014),
    .B(net1355),
    .Y(_10152_));
 INVx3_ASAP7_75t_R _39388_ (.A(_10152_),
    .Y(_10153_));
 TAPCELL_ASAP7_75t_R PHY_197 ();
 AO21x1_ASAP7_75t_R _39390_ (.A1(_10153_),
    .A2(net2958),
    .B(_10070_),
    .Y(_10155_));
 AND2x2_ASAP7_75t_R _39391_ (.A(_10151_),
    .B(_10155_),
    .Y(_10156_));
 NOR2x2_ASAP7_75t_R _39392_ (.A(_09875_),
    .B(_10029_),
    .Y(_10157_));
 TAPCELL_ASAP7_75t_R PHY_196 ();
 OAI21x1_ASAP7_75t_R _39394_ (.A1(_10077_),
    .A2(_10080_),
    .B(_10157_),
    .Y(_10159_));
 NOR2x2_ASAP7_75t_R _39395_ (.A(_09945_),
    .B(_09934_),
    .Y(_10161_));
 TAPCELL_ASAP7_75t_R PHY_195 ();
 NAND2x1_ASAP7_75t_R _39397_ (.A(_10161_),
    .B(_10099_),
    .Y(_10163_));
 NOR2x2_ASAP7_75t_R _39398_ (.A(_09904_),
    .B(_10058_),
    .Y(_10164_));
 NAND2x2_ASAP7_75t_R _39399_ (.A(net2382),
    .B(_10164_),
    .Y(_10165_));
 AND3x1_ASAP7_75t_R _39400_ (.A(_10159_),
    .B(_10163_),
    .C(_10165_),
    .Y(_10166_));
 NAND2x1_ASAP7_75t_R _39401_ (.A(_10156_),
    .B(_10166_),
    .Y(_10167_));
 NAND2x2_ASAP7_75t_R _39402_ (.A(net2804),
    .B(_09981_),
    .Y(_10168_));
 NOR2x2_ASAP7_75t_R _39403_ (.A(net1356),
    .B(net1027),
    .Y(_10169_));
 NAND2x2_ASAP7_75t_R _39404_ (.A(_10169_),
    .B(_10044_),
    .Y(_10170_));
 NAND2x1_ASAP7_75t_R _39405_ (.A(_10168_),
    .B(_10170_),
    .Y(_10172_));
 NAND2x1_ASAP7_75t_R _39406_ (.A(_10077_),
    .B(_10071_),
    .Y(_10173_));
 TAPCELL_ASAP7_75t_R PHY_194 ();
 NOR2x1_ASAP7_75t_R _39408_ (.A(net1963),
    .B(_10060_),
    .Y(_10175_));
 INVx2_ASAP7_75t_R _39409_ (.A(_10175_),
    .Y(_10176_));
 NAND2x1_ASAP7_75t_R _39410_ (.A(_10173_),
    .B(_10176_),
    .Y(_10177_));
 NOR2x1_ASAP7_75t_R _39411_ (.A(_10172_),
    .B(_10177_),
    .Y(_10178_));
 AO22x1_ASAP7_75t_R _39412_ (.A1(_10030_),
    .A2(_10126_),
    .B1(_10113_),
    .B2(net2431),
    .Y(_10179_));
 NOR2x2_ASAP7_75t_R _39413_ (.A(net3063),
    .B(net1660),
    .Y(_10180_));
 AO21x1_ASAP7_75t_R _39414_ (.A1(net1699),
    .A2(_10071_),
    .B(_10180_),
    .Y(_10181_));
 NOR2x1_ASAP7_75t_R _39415_ (.A(_10179_),
    .B(_10181_),
    .Y(_10183_));
 NAND2x1_ASAP7_75t_R _39416_ (.A(_10178_),
    .B(_10183_),
    .Y(_10184_));
 NOR2x2_ASAP7_75t_R _39417_ (.A(_10167_),
    .B(_10184_),
    .Y(_10185_));
 AO21x1_ASAP7_75t_R _39418_ (.A1(_09969_),
    .A2(_09945_),
    .B(_09934_),
    .Y(_10186_));
 AO21x1_ASAP7_75t_R _39419_ (.A1(_10186_),
    .A2(_09919_),
    .B(_09937_),
    .Y(_10187_));
 NAND2x1_ASAP7_75t_R _39420_ (.A(_09987_),
    .B(net1951),
    .Y(_10188_));
 NAND2x1_ASAP7_75t_R _39421_ (.A(_10077_),
    .B(net2382),
    .Y(_10189_));
 AND3x4_ASAP7_75t_R _39422_ (.A(_09884_),
    .B(_10188_),
    .C(_10189_),
    .Y(_10190_));
 NAND2x1_ASAP7_75t_R _39423_ (.A(_10187_),
    .B(_10190_),
    .Y(_10191_));
 AO21x1_ASAP7_75t_R _39424_ (.A1(_09939_),
    .A2(net1703),
    .B(_09969_),
    .Y(_10192_));
 TAPCELL_ASAP7_75t_R PHY_193 ();
 AO21x1_ASAP7_75t_R _39426_ (.A1(_10186_),
    .A2(_10192_),
    .B(_10005_),
    .Y(_10195_));
 NOR2x1_ASAP7_75t_R _39427_ (.A(net1797),
    .B(_09953_),
    .Y(_10196_));
 INVx1_ASAP7_75t_R _39428_ (.A(_10196_),
    .Y(_10197_));
 TAPCELL_ASAP7_75t_R PHY_192 ();
 TAPCELL_ASAP7_75t_R PHY_191 ();
 AO21x1_ASAP7_75t_R _39431_ (.A1(_10015_),
    .A2(_09908_),
    .B(_09901_),
    .Y(_10200_));
 OA21x2_ASAP7_75t_R _39432_ (.A1(net2373),
    .A2(_10197_),
    .B(_10200_),
    .Y(_10201_));
 NAND2x1_ASAP7_75t_R _39433_ (.A(_10195_),
    .B(_10201_),
    .Y(_10202_));
 NOR2x2_ASAP7_75t_R _39434_ (.A(_10191_),
    .B(_10202_),
    .Y(_10203_));
 NAND3x2_ASAP7_75t_R _39435_ (.B(_10185_),
    .C(_10203_),
    .Y(_10205_),
    .A(_10150_));
 TAPCELL_ASAP7_75t_R PHY_190 ();
 NAND2x2_ASAP7_75t_R _39437_ (.A(net1251),
    .B(net2667),
    .Y(_10207_));
 TAPCELL_ASAP7_75t_R PHY_189 ();
 AO21x1_ASAP7_75t_R _39439_ (.A1(net949),
    .A2(_10207_),
    .B(_10035_),
    .Y(_10209_));
 AO21x1_ASAP7_75t_R _39440_ (.A1(_09998_),
    .A2(_09928_),
    .B(_10060_),
    .Y(_10210_));
 NAND2x2_ASAP7_75t_R _39441_ (.A(net2804),
    .B(_09883_),
    .Y(_10211_));
 AND3x4_ASAP7_75t_R _39442_ (.A(_10209_),
    .B(_10210_),
    .C(_10211_),
    .Y(_10212_));
 AO21x2_ASAP7_75t_R _39443_ (.A1(net942),
    .A2(_09919_),
    .B(_09922_),
    .Y(_10213_));
 TAPCELL_ASAP7_75t_R PHY_188 ();
 AO21x1_ASAP7_75t_R _39445_ (.A1(net2409),
    .A2(_09998_),
    .B(_09922_),
    .Y(_10216_));
 NOR2x1_ASAP7_75t_R _39446_ (.A(_09928_),
    .B(_09922_),
    .Y(_10217_));
 INVx1_ASAP7_75t_R _39447_ (.A(_10217_),
    .Y(_10218_));
 AND3x4_ASAP7_75t_R _39448_ (.A(_10213_),
    .B(_10216_),
    .C(_10218_),
    .Y(_10219_));
 NAND2x2_ASAP7_75t_R _39449_ (.A(_10219_),
    .B(_10212_),
    .Y(_10220_));
 TAPCELL_ASAP7_75t_R PHY_187 ();
 AO21x1_ASAP7_75t_R _39451_ (.A1(net2397),
    .A2(net2734),
    .B(_09990_),
    .Y(_10222_));
 AO21x1_ASAP7_75t_R _39452_ (.A1(_10013_),
    .A2(_09963_),
    .B(_09990_),
    .Y(_10223_));
 NAND2x1_ASAP7_75t_R _39453_ (.A(_10222_),
    .B(_10223_),
    .Y(_10224_));
 NAND2x2_ASAP7_75t_R _39454_ (.A(net1701),
    .B(_09876_),
    .Y(_10225_));
 TAPCELL_ASAP7_75t_R PHY_186 ();
 OAI22x1_ASAP7_75t_R _39456_ (.A1(_10225_),
    .A2(net1163),
    .B1(net2353),
    .B2(_10038_),
    .Y(_10228_));
 NOR2x1_ASAP7_75t_R _39457_ (.A(_10224_),
    .B(_10228_),
    .Y(_10229_));
 AOI22x1_ASAP7_75t_R _39458_ (.A1(_09981_),
    .A2(net2430),
    .B1(_10044_),
    .B2(_09959_),
    .Y(_10230_));
 AND2x2_ASAP7_75t_R _39459_ (.A(_10092_),
    .B(_10230_),
    .Y(_10231_));
 TAPCELL_ASAP7_75t_R PHY_185 ();
 TAPCELL_ASAP7_75t_R PHY_184 ();
 NOR2x1_ASAP7_75t_R _39462_ (.A(net1757),
    .B(_10040_),
    .Y(_10234_));
 OA21x2_ASAP7_75t_R _39463_ (.A1(_09982_),
    .A2(_09979_),
    .B(net2430),
    .Y(_10235_));
 NOR2x1_ASAP7_75t_R _39464_ (.A(_10234_),
    .B(_10235_),
    .Y(_10236_));
 NAND3x1_ASAP7_75t_R _39465_ (.A(_10229_),
    .B(_10231_),
    .C(_10236_),
    .Y(_10238_));
 NOR2x1_ASAP7_75t_R _39466_ (.A(_10238_),
    .B(_10220_),
    .Y(_10239_));
 NAND2x2_ASAP7_75t_R _39467_ (.A(net2281),
    .B(net2804),
    .Y(_10240_));
 NAND2x2_ASAP7_75t_R _39468_ (.A(_09992_),
    .B(_09883_),
    .Y(_10241_));
 OAI21x1_ASAP7_75t_R _39469_ (.A1(net2591),
    .A2(_10240_),
    .B(_10241_),
    .Y(_10242_));
 TAPCELL_ASAP7_75t_R PHY_183 ();
 AO21x1_ASAP7_75t_R _39471_ (.A1(net1963),
    .A2(net2958),
    .B(net2925),
    .Y(_10244_));
 TAPCELL_ASAP7_75t_R PHY_182 ();
 NAND2x2_ASAP7_75t_R _39473_ (.A(_09952_),
    .B(_09989_),
    .Y(_10246_));
 OAI21x1_ASAP7_75t_R _39474_ (.A1(net2470),
    .A2(_09893_),
    .B(net2282),
    .Y(_10247_));
 AO21x1_ASAP7_75t_R _39475_ (.A1(_10011_),
    .A2(_10246_),
    .B(_10247_),
    .Y(_10249_));
 NAND2x1_ASAP7_75t_R _39476_ (.A(_10244_),
    .B(_10249_),
    .Y(_10250_));
 NOR2x1_ASAP7_75t_R _39477_ (.A(_10242_),
    .B(_10250_),
    .Y(_10251_));
 NOR2x2_ASAP7_75t_R _39478_ (.A(net2408),
    .B(_10246_),
    .Y(_10252_));
 AO21x1_ASAP7_75t_R _39479_ (.A1(_10126_),
    .A2(_10133_),
    .B(_10252_),
    .Y(_10253_));
 NAND2x2_ASAP7_75t_R _39480_ (.A(net1065),
    .B(_10058_),
    .Y(_10254_));
 NOR2x2_ASAP7_75t_R _39481_ (.A(net2584),
    .B(_09875_),
    .Y(_10255_));
 TAPCELL_ASAP7_75t_R PHY_181 ();
 AND3x4_ASAP7_75t_R _39483_ (.A(_10254_),
    .B(_10255_),
    .C(net1701),
    .Y(_10257_));
 NOR2x1_ASAP7_75t_R _39484_ (.A(net3244),
    .B(_10059_),
    .Y(_10258_));
 NOR3x1_ASAP7_75t_R _39485_ (.A(_10253_),
    .B(_10257_),
    .C(_10258_),
    .Y(_10259_));
 NAND2x1_ASAP7_75t_R _39486_ (.A(_10251_),
    .B(_10259_),
    .Y(_10260_));
 NOR2x1_ASAP7_75t_R _39487_ (.A(_09934_),
    .B(_10106_),
    .Y(_10261_));
 INVx1_ASAP7_75t_R _39488_ (.A(_10261_),
    .Y(_10262_));
 OAI22x1_ASAP7_75t_R _39489_ (.A1(_10262_),
    .A2(net3015),
    .B1(net3309),
    .B2(_10079_),
    .Y(_10263_));
 INVx4_ASAP7_75t_R _39490_ (.A(net2408),
    .Y(_10264_));
 TAPCELL_ASAP7_75t_R PHY_180 ();
 NOR2x1_ASAP7_75t_R _39492_ (.A(_10003_),
    .B(net3093),
    .Y(_10266_));
 AO22x1_ASAP7_75t_R _39493_ (.A1(_10264_),
    .A2(_10044_),
    .B1(_10266_),
    .B2(_09892_),
    .Y(_10267_));
 NOR2x1_ASAP7_75t_R _39494_ (.A(_10263_),
    .B(_10267_),
    .Y(_10268_));
 AOI22x1_ASAP7_75t_R _39495_ (.A1(_10099_),
    .A2(net1700),
    .B1(_10152_),
    .B2(_10255_),
    .Y(_10270_));
 TAPCELL_ASAP7_75t_R PHY_179 ();
 NAND2x1_ASAP7_75t_R _39497_ (.A(net1893),
    .B(_09982_),
    .Y(_10272_));
 OA21x2_ASAP7_75t_R _39498_ (.A1(net3093),
    .A2(_09914_),
    .B(_10272_),
    .Y(_10273_));
 NAND2x1_ASAP7_75t_R _39499_ (.A(_10270_),
    .B(_10273_),
    .Y(_10274_));
 NAND2x1_ASAP7_75t_R _39500_ (.A(_10152_),
    .B(net1890),
    .Y(_10275_));
 OA21x2_ASAP7_75t_R _39501_ (.A1(_09890_),
    .A2(net2925),
    .B(_10275_),
    .Y(_10276_));
 NAND2x1_ASAP7_75t_R _39502_ (.A(_10080_),
    .B(_10099_),
    .Y(_10277_));
 NAND2x2_ASAP7_75t_R _39503_ (.A(_10027_),
    .B(net1949),
    .Y(_10278_));
 AND2x2_ASAP7_75t_R _39504_ (.A(_10277_),
    .B(_10278_),
    .Y(_10279_));
 NAND2x1_ASAP7_75t_R _39505_ (.A(_10276_),
    .B(_10279_),
    .Y(_10281_));
 NOR2x1_ASAP7_75t_R _39506_ (.A(_10274_),
    .B(_10281_),
    .Y(_10282_));
 NAND2x1_ASAP7_75t_R _39507_ (.A(_10268_),
    .B(_10282_),
    .Y(_10283_));
 NOR2x1_ASAP7_75t_R _39508_ (.A(_10260_),
    .B(_10283_),
    .Y(_10284_));
 NAND2x1_ASAP7_75t_R _39509_ (.A(_10239_),
    .B(_10284_),
    .Y(_10285_));
 NOR2x2_ASAP7_75t_R _39510_ (.A(_10205_),
    .B(_10285_),
    .Y(_10286_));
 NOR2x2_ASAP7_75t_R _39511_ (.A(_10286_),
    .B(_10121_),
    .Y(_10287_));
 INVx3_ASAP7_75t_R _39512_ (.A(_10287_),
    .Y(_10288_));
 OAI21x1_ASAP7_75t_R _39513_ (.A1(_09881_),
    .A2(_09994_),
    .B(net2282),
    .Y(_10289_));
 AOI21x1_ASAP7_75t_R _39514_ (.A1(_10013_),
    .A2(_10289_),
    .B(_10005_),
    .Y(_10290_));
 AOI21x1_ASAP7_75t_R _39515_ (.A1(_09963_),
    .A2(_10247_),
    .B(_10005_),
    .Y(_10292_));
 NOR2x2_ASAP7_75t_R _39516_ (.A(_10290_),
    .B(_10292_),
    .Y(_10293_));
 NOR2x1_ASAP7_75t_R _39517_ (.A(_09934_),
    .B(_10005_),
    .Y(_10294_));
 TAPCELL_ASAP7_75t_R PHY_178 ();
 AOI21x1_ASAP7_75t_R _39519_ (.A1(_10111_),
    .A2(_10042_),
    .B(_10005_),
    .Y(_10296_));
 NOR2x1_ASAP7_75t_R _39520_ (.A(_10294_),
    .B(_10296_),
    .Y(_10297_));
 OR3x1_ASAP7_75t_R _39521_ (.A(_09897_),
    .B(_09870_),
    .C(net3160),
    .Y(_10298_));
 AND4x2_ASAP7_75t_R _39522_ (.A(_10293_),
    .B(_10011_),
    .C(_10297_),
    .D(_10298_),
    .Y(_10299_));
 NAND3x2_ASAP7_75t_R _39523_ (.B(_00649_),
    .C(net2832),
    .Y(_10300_),
    .A(_10299_));
 TAPCELL_ASAP7_75t_R PHY_177 ();
 NAND3x2_ASAP7_75t_R _39525_ (.B(_10121_),
    .C(net2681),
    .Y(_10303_),
    .A(_10286_));
 NAND2x2_ASAP7_75t_R _39526_ (.A(_10288_),
    .B(_10303_),
    .Y(_10304_));
 NOR2x1_ASAP7_75t_R _39527_ (.A(_09867_),
    .B(_10304_),
    .Y(_10305_));
 INVx2_ASAP7_75t_R _39528_ (.A(_09867_),
    .Y(_10306_));
 AO21x1_ASAP7_75t_R _39529_ (.A1(_10303_),
    .A2(_10288_),
    .B(_10306_),
    .Y(_10307_));
 INVx1_ASAP7_75t_R _39530_ (.A(_10307_),
    .Y(_10308_));
 TAPCELL_ASAP7_75t_R PHY_176 ();
 NAND2x2_ASAP7_75t_R _39532_ (.A(net1374),
    .B(net1582),
    .Y(_10310_));
 INVx6_ASAP7_75t_R _39533_ (.A(net1960),
    .Y(_10311_));
 NAND2x2_ASAP7_75t_R _39534_ (.A(net2311),
    .B(_10311_),
    .Y(_10312_));
 TAPCELL_ASAP7_75t_R PHY_175 ();
 NOR2x2_ASAP7_75t_R _39536_ (.A(net960),
    .B(net1513),
    .Y(_10315_));
 CKINVDCx16_ASAP7_75t_R _39537_ (.A(net1582),
    .Y(_10316_));
 NAND2x2_ASAP7_75t_R _39538_ (.A(net1374),
    .B(_10316_),
    .Y(_10317_));
 NOR2x2_ASAP7_75t_R _39539_ (.A(_10317_),
    .B(_10312_),
    .Y(_10318_));
 TAPCELL_ASAP7_75t_R PHY_174 ();
 TAPCELL_ASAP7_75t_R PHY_173 ();
 NAND2x2_ASAP7_75t_R _39542_ (.A(net3361),
    .B(net2741),
    .Y(_10321_));
 NAND2x2_ASAP7_75t_R _39543_ (.A(_00569_),
    .B(_00570_),
    .Y(_10322_));
 NOR2x2_ASAP7_75t_R _39544_ (.A(_10321_),
    .B(_10322_),
    .Y(_10323_));
 OAI21x1_ASAP7_75t_R _39545_ (.A1(_10315_),
    .A2(_10318_),
    .B(_10323_),
    .Y(_10325_));
 NOR2x2_ASAP7_75t_R _39546_ (.A(net1374),
    .B(_10316_),
    .Y(_10326_));
 INVx3_ASAP7_75t_R _39547_ (.A(_00574_),
    .Y(_10327_));
 NOR2x2_ASAP7_75t_R _39548_ (.A(net1960),
    .B(_10327_),
    .Y(_10328_));
 NAND2x2_ASAP7_75t_R _39549_ (.A(_10326_),
    .B(net3035),
    .Y(_10329_));
 TAPCELL_ASAP7_75t_R PHY_172 ();
 TAPCELL_ASAP7_75t_R PHY_171 ();
 NOR2x2_ASAP7_75t_R _39552_ (.A(net1374),
    .B(net1582),
    .Y(_10332_));
 NAND2x2_ASAP7_75t_R _39553_ (.A(_10332_),
    .B(net2745),
    .Y(_10333_));
 TAPCELL_ASAP7_75t_R PHY_170 ();
 CKINVDCx8_ASAP7_75t_R _39555_ (.A(_10323_),
    .Y(_10336_));
 AO21x1_ASAP7_75t_R _39556_ (.A1(_10329_),
    .A2(_10333_),
    .B(_10336_),
    .Y(_10337_));
 NAND2x2_ASAP7_75t_R _39557_ (.A(_10325_),
    .B(_10337_),
    .Y(_10338_));
 NOR2x2_ASAP7_75t_R _39558_ (.A(net1960),
    .B(_00574_),
    .Y(_10339_));
 TAPCELL_ASAP7_75t_R PHY_169 ();
 INVx11_ASAP7_75t_R _39560_ (.A(net1273),
    .Y(_10341_));
 NOR2x2_ASAP7_75t_R _39561_ (.A(_10341_),
    .B(_10336_),
    .Y(_10342_));
 NOR2x2_ASAP7_75t_R _39562_ (.A(net2311),
    .B(_10311_),
    .Y(_10343_));
 TAPCELL_ASAP7_75t_R PHY_168 ();
 NAND2x2_ASAP7_75t_R _39564_ (.A(net1885),
    .B(_10323_),
    .Y(_10345_));
 TAPCELL_ASAP7_75t_R PHY_167 ();
 NAND2x2_ASAP7_75t_R _39566_ (.A(net1960),
    .B(_00574_),
    .Y(_10348_));
 NOR2x2_ASAP7_75t_R _39567_ (.A(net1379),
    .B(net972),
    .Y(_10349_));
 NOR2x2_ASAP7_75t_R _39568_ (.A(net968),
    .B(_10317_),
    .Y(_10350_));
 OAI21x1_ASAP7_75t_R _39569_ (.A1(_10349_),
    .A2(_10350_),
    .B(_10323_),
    .Y(_10351_));
 NAND2x2_ASAP7_75t_R _39570_ (.A(_10345_),
    .B(_10351_),
    .Y(_10352_));
 NOR3x2_ASAP7_75t_R _39571_ (.B(_10342_),
    .C(_10352_),
    .Y(_10353_),
    .A(_10338_));
 INVx3_ASAP7_75t_R _39572_ (.A(net3361),
    .Y(_10354_));
 NOR2x2_ASAP7_75t_R _39573_ (.A(net2741),
    .B(_10354_),
    .Y(_10355_));
 INVx3_ASAP7_75t_R _39574_ (.A(_10322_),
    .Y(_10356_));
 NAND2x2_ASAP7_75t_R _39575_ (.A(_10355_),
    .B(_10356_),
    .Y(_10358_));
 TAPCELL_ASAP7_75t_R PHY_166 ();
 INVx4_ASAP7_75t_R _39577_ (.A(_00569_),
    .Y(_10360_));
 INVx3_ASAP7_75t_R _39578_ (.A(_00570_),
    .Y(_10361_));
 OR3x2_ASAP7_75t_R _39579_ (.A(_10360_),
    .B(_10361_),
    .C(net3362),
    .Y(_10362_));
 NAND3x2_ASAP7_75t_R _39580_ (.B(net2241),
    .C(_10362_),
    .Y(_10363_),
    .A(_10353_));
 NOR3x2_ASAP7_75t_R _39581_ (.B(_10360_),
    .C(_10361_),
    .Y(_10364_),
    .A(_10363_));
 NAND2x2_ASAP7_75t_R _39582_ (.A(_10326_),
    .B(_10343_),
    .Y(_10365_));
 TAPCELL_ASAP7_75t_R PHY_165 ();
 CKINVDCx20_ASAP7_75t_R _39584_ (.A(net1374),
    .Y(_10367_));
 NOR2x2_ASAP7_75t_R _39585_ (.A(net1582),
    .B(_10367_),
    .Y(_10369_));
 NAND2x2_ASAP7_75t_R _39586_ (.A(net3293),
    .B(net3038),
    .Y(_10370_));
 TAPCELL_ASAP7_75t_R PHY_164 ();
 AOI21x1_ASAP7_75t_R _39588_ (.A1(net1494),
    .A2(net1414),
    .B(_10358_),
    .Y(_10372_));
 TAPCELL_ASAP7_75t_R PHY_163 ();
 INVx4_ASAP7_75t_R _39590_ (.A(_10310_),
    .Y(_10374_));
 NAND2x2_ASAP7_75t_R _39591_ (.A(net1742),
    .B(_10374_),
    .Y(_10375_));
 AOI21x1_ASAP7_75t_R _39592_ (.A1(net2333),
    .A2(_10375_),
    .B(_10358_),
    .Y(_10376_));
 INVx1_ASAP7_75t_R _39593_ (.A(_10349_),
    .Y(_10377_));
 NOR2x2_ASAP7_75t_R _39594_ (.A(_10377_),
    .B(_10358_),
    .Y(_10378_));
 NOR3x2_ASAP7_75t_R _39595_ (.B(_10376_),
    .C(_10378_),
    .Y(_10380_),
    .A(_10372_));
 INVx1_ASAP7_75t_R _39596_ (.A(_10380_),
    .Y(_10381_));
 CKINVDCx5p33_ASAP7_75t_R _39597_ (.A(_10332_),
    .Y(_10382_));
 NOR2x2_ASAP7_75t_R _39598_ (.A(net968),
    .B(_10382_),
    .Y(_10383_));
 NAND2x2_ASAP7_75t_R _39599_ (.A(net1584),
    .B(_10367_),
    .Y(_10384_));
 NOR2x2_ASAP7_75t_R _39600_ (.A(net969),
    .B(_10384_),
    .Y(_10385_));
 TAPCELL_ASAP7_75t_R PHY_162 ();
 OA21x2_ASAP7_75t_R _39602_ (.A1(_10383_),
    .A2(_10385_),
    .B(_10323_),
    .Y(_10387_));
 TAPCELL_ASAP7_75t_R PHY_161 ();
 NAND2x2_ASAP7_75t_R _39604_ (.A(net1960),
    .B(_10327_),
    .Y(_10389_));
 TAPCELL_ASAP7_75t_R PHY_160 ();
 AOI211x1_ASAP7_75t_R _39606_ (.A1(net975),
    .A2(net1318),
    .B(_10336_),
    .C(_10389_),
    .Y(_10392_));
 NOR2x2_ASAP7_75t_R _39607_ (.A(_10387_),
    .B(_10392_),
    .Y(_10393_));
 NAND2x2_ASAP7_75t_R _39608_ (.A(net3032),
    .B(_10369_),
    .Y(_10394_));
 TAPCELL_ASAP7_75t_R PHY_159 ();
 NAND2x2_ASAP7_75t_R _39610_ (.A(net2566),
    .B(_10326_),
    .Y(_10396_));
 TAPCELL_ASAP7_75t_R PHY_158 ();
 AO21x1_ASAP7_75t_R _39612_ (.A1(net1079),
    .A2(net1090),
    .B(_10336_),
    .Y(_10398_));
 NOR2x2_ASAP7_75t_R _39613_ (.A(net1510),
    .B(_10374_),
    .Y(_10399_));
 NAND2x1_ASAP7_75t_R _39614_ (.A(_10323_),
    .B(_10399_),
    .Y(_10400_));
 AND2x2_ASAP7_75t_R _39615_ (.A(_10398_),
    .B(_10400_),
    .Y(_10402_));
 NAND2x1_ASAP7_75t_R _39616_ (.A(_10393_),
    .B(_10402_),
    .Y(_10403_));
 NOR2x1_ASAP7_75t_R _39617_ (.A(_10381_),
    .B(_10403_),
    .Y(_10404_));
 NAND2x2_ASAP7_75t_R _39618_ (.A(net2742),
    .B(_10354_),
    .Y(_10405_));
 NOR2x2_ASAP7_75t_R _39619_ (.A(net2355),
    .B(_10405_),
    .Y(_10406_));
 NAND2x1_ASAP7_75t_R _39620_ (.A(_10406_),
    .B(_10399_),
    .Y(_10407_));
 NAND2x2_ASAP7_75t_R _39621_ (.A(net3032),
    .B(_10374_),
    .Y(_10408_));
 TAPCELL_ASAP7_75t_R PHY_157 ();
 NAND2x2_ASAP7_75t_R _39623_ (.A(_10367_),
    .B(net1268),
    .Y(_10410_));
 TAPCELL_ASAP7_75t_R PHY_156 ();
 INVx2_ASAP7_75t_R _39625_ (.A(net2741),
    .Y(_10413_));
 NOR2x2_ASAP7_75t_R _39626_ (.A(net3361),
    .B(_10413_),
    .Y(_10414_));
 NAND2x2_ASAP7_75t_R _39627_ (.A(_10414_),
    .B(_10356_),
    .Y(_10415_));
 TAPCELL_ASAP7_75t_R PHY_155 ();
 AO21x1_ASAP7_75t_R _39629_ (.A1(net2954),
    .A2(_10410_),
    .B(_10415_),
    .Y(_10417_));
 NAND2x1_ASAP7_75t_R _39630_ (.A(_10407_),
    .B(_10417_),
    .Y(_10418_));
 INVx11_ASAP7_75t_R _39631_ (.A(net968),
    .Y(_10419_));
 NAND2x2_ASAP7_75t_R _39632_ (.A(_10326_),
    .B(_10419_),
    .Y(_10420_));
 NAND2x2_ASAP7_75t_R _39633_ (.A(_10419_),
    .B(net1377),
    .Y(_10421_));
 AO21x2_ASAP7_75t_R _39634_ (.A1(_10420_),
    .A2(_10421_),
    .B(_10415_),
    .Y(_10422_));
 TAPCELL_ASAP7_75t_R PHY_154 ();
 TAPCELL_ASAP7_75t_R PHY_153 ();
 AO21x1_ASAP7_75t_R _39637_ (.A1(net1494),
    .A2(_10370_),
    .B(_10415_),
    .Y(_10426_));
 NAND2x1_ASAP7_75t_R _39638_ (.A(_10426_),
    .B(_10422_),
    .Y(_10427_));
 NOR2x2_ASAP7_75t_R _39639_ (.A(_10418_),
    .B(_10427_),
    .Y(_10428_));
 INVx1_ASAP7_75t_R _39640_ (.A(_10428_),
    .Y(_10429_));
 NOR2x2_ASAP7_75t_R _39641_ (.A(net3361),
    .B(net2741),
    .Y(_10430_));
 NAND2x2_ASAP7_75t_R _39642_ (.A(net2491),
    .B(_10356_),
    .Y(_10431_));
 TAPCELL_ASAP7_75t_R PHY_152 ();
 TAPCELL_ASAP7_75t_R PHY_151 ();
 NOR2x1_ASAP7_75t_R _39645_ (.A(net1881),
    .B(net1494),
    .Y(_10435_));
 TAPCELL_ASAP7_75t_R PHY_150 ();
 AOI211x1_ASAP7_75t_R _39647_ (.A1(net1376),
    .A2(net1583),
    .B(_10431_),
    .C(net965),
    .Y(_10437_));
 NOR2x2_ASAP7_75t_R _39648_ (.A(_10435_),
    .B(_10437_),
    .Y(_10438_));
 NOR2x2_ASAP7_75t_R _39649_ (.A(_10341_),
    .B(_10431_),
    .Y(_10439_));
 TAPCELL_ASAP7_75t_R PHY_149 ();
 NOR2x1_ASAP7_75t_R _39651_ (.A(_10431_),
    .B(_10375_),
    .Y(_10441_));
 NAND2x2_ASAP7_75t_R _39652_ (.A(_10332_),
    .B(net3032),
    .Y(_10442_));
 NOR2x1_ASAP7_75t_R _39653_ (.A(_10442_),
    .B(_10431_),
    .Y(_10443_));
 AOI211x1_ASAP7_75t_R _39654_ (.A1(_10439_),
    .A2(net1376),
    .B(_10441_),
    .C(_10443_),
    .Y(_10444_));
 NAND2x1_ASAP7_75t_R _39655_ (.A(_10438_),
    .B(_10444_),
    .Y(_10446_));
 NOR2x1_ASAP7_75t_R _39656_ (.A(_10429_),
    .B(_10446_),
    .Y(_10447_));
 NAND2x2_ASAP7_75t_R _39657_ (.A(_10447_),
    .B(_10404_),
    .Y(_10448_));
 NAND2x2_ASAP7_75t_R _39658_ (.A(net3038),
    .B(_10419_),
    .Y(_10449_));
 TAPCELL_ASAP7_75t_R PHY_148 ();
 NAND2x2_ASAP7_75t_R _39660_ (.A(_10332_),
    .B(_10419_),
    .Y(_10451_));
 TAPCELL_ASAP7_75t_R PHY_147 ();
 NOR2x2_ASAP7_75t_R _39662_ (.A(_00570_),
    .B(_10360_),
    .Y(_10453_));
 NAND2x2_ASAP7_75t_R _39663_ (.A(_10453_),
    .B(_10414_),
    .Y(_10454_));
 TAPCELL_ASAP7_75t_R PHY_146 ();
 TAPCELL_ASAP7_75t_R PHY_145 ();
 AO21x1_ASAP7_75t_R _39666_ (.A1(net2463),
    .A2(net1125),
    .B(net2020),
    .Y(_10458_));
 NAND2x2_ASAP7_75t_R _39667_ (.A(_10384_),
    .B(net1741),
    .Y(_10459_));
 TAPCELL_ASAP7_75t_R PHY_144 ();
 AO21x1_ASAP7_75t_R _39669_ (.A1(_10459_),
    .A2(net1090),
    .B(net2020),
    .Y(_10461_));
 INVx3_ASAP7_75t_R _39670_ (.A(_10454_),
    .Y(_10462_));
 NAND2x1_ASAP7_75t_R _39671_ (.A(net1499),
    .B(_10462_),
    .Y(_10463_));
 NAND3x1_ASAP7_75t_R _39672_ (.A(_10458_),
    .B(_10461_),
    .C(_10463_),
    .Y(_10464_));
 TAPCELL_ASAP7_75t_R PHY_143 ();
 AO21x1_ASAP7_75t_R _39674_ (.A1(net2962),
    .A2(_10317_),
    .B(_10341_),
    .Y(_10466_));
 NAND2x2_ASAP7_75t_R _39675_ (.A(_10430_),
    .B(_10453_),
    .Y(_10468_));
 TAPCELL_ASAP7_75t_R PHY_142 ();
 AO21x1_ASAP7_75t_R _39677_ (.A1(_10466_),
    .A2(net3161),
    .B(net2233),
    .Y(_10470_));
 NAND2x2_ASAP7_75t_R _39678_ (.A(_10332_),
    .B(_10343_),
    .Y(_10471_));
 TAPCELL_ASAP7_75t_R PHY_141 ();
 AOI21x1_ASAP7_75t_R _39680_ (.A1(net3292),
    .A2(net2851),
    .B(net1979),
    .Y(_10473_));
 TAPCELL_ASAP7_75t_R PHY_140 ();
 TAPCELL_ASAP7_75t_R PHY_139 ();
 AOI211x1_ASAP7_75t_R _39683_ (.A1(_10367_),
    .A2(net1318),
    .B(net2233),
    .C(net968),
    .Y(_10476_));
 NOR2x1_ASAP7_75t_R _39684_ (.A(_10473_),
    .B(_10476_),
    .Y(_10477_));
 NAND2x1_ASAP7_75t_R _39685_ (.A(_10470_),
    .B(_10477_),
    .Y(_10479_));
 NOR2x1_ASAP7_75t_R _39686_ (.A(_10464_),
    .B(_10479_),
    .Y(_10480_));
 INVx2_ASAP7_75t_R _39687_ (.A(_10442_),
    .Y(_10481_));
 NAND2x2_ASAP7_75t_R _39688_ (.A(_10355_),
    .B(_10453_),
    .Y(_10482_));
 INVx4_ASAP7_75t_R _39689_ (.A(_10482_),
    .Y(_10483_));
 NAND2x1_ASAP7_75t_R _39690_ (.A(_10481_),
    .B(_10483_),
    .Y(_10484_));
 NAND2x2_ASAP7_75t_R _39691_ (.A(net3038),
    .B(net1740),
    .Y(_10485_));
 TAPCELL_ASAP7_75t_R PHY_138 ();
 AO21x1_ASAP7_75t_R _39693_ (.A1(net2957),
    .A2(net1114),
    .B(net2070),
    .Y(_10487_));
 NAND2x1_ASAP7_75t_R _39694_ (.A(_10484_),
    .B(_10487_),
    .Y(_10488_));
 NAND2x2_ASAP7_75t_R _39695_ (.A(_10384_),
    .B(_10419_),
    .Y(_10490_));
 INVx1_ASAP7_75t_R _39696_ (.A(_10490_),
    .Y(_10491_));
 NAND2x1_ASAP7_75t_R _39697_ (.A(_10491_),
    .B(_10483_),
    .Y(_10492_));
 TAPCELL_ASAP7_75t_R PHY_137 ();
 AO21x1_ASAP7_75t_R _39699_ (.A1(net1494),
    .A2(_10471_),
    .B(_10482_),
    .Y(_10494_));
 NAND2x1_ASAP7_75t_R _39700_ (.A(_10492_),
    .B(_10494_),
    .Y(_10495_));
 NOR2x1_ASAP7_75t_R _39701_ (.A(_10488_),
    .B(_10495_),
    .Y(_10496_));
 INVx4_ASAP7_75t_R _39702_ (.A(_10321_),
    .Y(_10497_));
 NAND2x2_ASAP7_75t_R _39703_ (.A(_10453_),
    .B(_10497_),
    .Y(_10498_));
 TAPCELL_ASAP7_75t_R PHY_136 ();
 AO21x1_ASAP7_75t_R _39705_ (.A1(_10485_),
    .A2(net2333),
    .B(net2249),
    .Y(_10501_));
 NAND2x2_ASAP7_75t_R _39706_ (.A(net1841),
    .B(_10374_),
    .Y(_10502_));
 TAPCELL_ASAP7_75t_R PHY_135 ();
 AO21x1_ASAP7_75t_R _39708_ (.A1(_10502_),
    .A2(_10421_),
    .B(net2249),
    .Y(_10504_));
 NAND2x2_ASAP7_75t_R _39709_ (.A(net1375),
    .B(net2566),
    .Y(_10505_));
 TAPCELL_ASAP7_75t_R PHY_134 ();
 AO21x1_ASAP7_75t_R _39711_ (.A1(net2441),
    .A2(_10505_),
    .B(net2249),
    .Y(_10507_));
 AND3x1_ASAP7_75t_R _39712_ (.A(_10501_),
    .B(_10504_),
    .C(_10507_),
    .Y(_10508_));
 NAND2x1_ASAP7_75t_R _39713_ (.A(_10496_),
    .B(_10508_),
    .Y(_10509_));
 INVx1_ASAP7_75t_R _39714_ (.A(_10509_),
    .Y(_10510_));
 NAND2x1_ASAP7_75t_R _39715_ (.A(_10510_),
    .B(_10480_),
    .Y(_10512_));
 NOR2x2_ASAP7_75t_R _39716_ (.A(_10448_),
    .B(_10512_),
    .Y(_10513_));
 NOR2x2_ASAP7_75t_R _39717_ (.A(net2727),
    .B(_10361_),
    .Y(_10514_));
 NAND2x2_ASAP7_75t_R _39718_ (.A(_10430_),
    .B(_10514_),
    .Y(_10515_));
 TAPCELL_ASAP7_75t_R PHY_133 ();
 TAPCELL_ASAP7_75t_R PHY_132 ();
 AO21x1_ASAP7_75t_R _39721_ (.A1(_10367_),
    .A2(net1585),
    .B(net3011),
    .Y(_10518_));
 NOR2x1_ASAP7_75t_R _39722_ (.A(net2228),
    .B(_10518_),
    .Y(_10519_));
 NOR2x2_ASAP7_75t_R _39723_ (.A(_10316_),
    .B(net970),
    .Y(_10520_));
 INVx1_ASAP7_75t_R _39724_ (.A(_10520_),
    .Y(_10521_));
 AOI21x1_ASAP7_75t_R _39725_ (.A1(net1125),
    .A2(_10521_),
    .B(net2228),
    .Y(_10523_));
 NOR2x1_ASAP7_75t_R _39726_ (.A(net2228),
    .B(net1143),
    .Y(_10524_));
 NOR3x1_ASAP7_75t_R _39727_ (.A(_10519_),
    .B(_10523_),
    .C(_10524_),
    .Y(_10525_));
 INVx1_ASAP7_75t_R _39728_ (.A(_10505_),
    .Y(_10526_));
 NAND2x2_ASAP7_75t_R _39729_ (.A(_00570_),
    .B(_10360_),
    .Y(_10527_));
 NOR2x2_ASAP7_75t_R _39730_ (.A(_10405_),
    .B(_10527_),
    .Y(_10528_));
 OAI21x1_ASAP7_75t_R _39731_ (.A1(_10526_),
    .A2(_10481_),
    .B(_10528_),
    .Y(_10529_));
 NAND2x1_ASAP7_75t_R _39732_ (.A(_10318_),
    .B(_10528_),
    .Y(_10530_));
 NOR2x2_ASAP7_75t_R _39733_ (.A(net957),
    .B(net3010),
    .Y(_10531_));
 NAND2x1_ASAP7_75t_R _39734_ (.A(_10531_),
    .B(_10528_),
    .Y(_10532_));
 AND3x1_ASAP7_75t_R _39735_ (.A(_10529_),
    .B(_10530_),
    .C(_10532_),
    .Y(_10534_));
 NAND2x1_ASAP7_75t_R _39736_ (.A(_10525_),
    .B(_10534_),
    .Y(_10535_));
 NAND2x2_ASAP7_75t_R _39737_ (.A(net2839),
    .B(_10413_),
    .Y(_10536_));
 NOR2x2_ASAP7_75t_R _39738_ (.A(_10536_),
    .B(_10527_),
    .Y(_10537_));
 AND3x1_ASAP7_75t_R _39739_ (.A(_10537_),
    .B(_10367_),
    .C(net1270),
    .Y(_10538_));
 TAPCELL_ASAP7_75t_R PHY_131 ();
 NAND2x2_ASAP7_75t_R _39741_ (.A(_10355_),
    .B(_10514_),
    .Y(_10540_));
 AO21x1_ASAP7_75t_R _39742_ (.A1(net2695),
    .A2(net2463),
    .B(_10540_),
    .Y(_10541_));
 INVx1_ASAP7_75t_R _39743_ (.A(_10541_),
    .Y(_10542_));
 NOR2x1_ASAP7_75t_R _39744_ (.A(_10538_),
    .B(_10542_),
    .Y(_10543_));
 NOR2x2_ASAP7_75t_R _39745_ (.A(net1512),
    .B(_10382_),
    .Y(_10545_));
 NAND2x2_ASAP7_75t_R _39746_ (.A(_10514_),
    .B(_10497_),
    .Y(_10546_));
 INVx11_ASAP7_75t_R _39747_ (.A(_10546_),
    .Y(_10547_));
 TAPCELL_ASAP7_75t_R PHY_130 ();
 OAI21x1_ASAP7_75t_R _39749_ (.A1(net1264),
    .A2(_10545_),
    .B(_10547_),
    .Y(_10549_));
 INVx1_ASAP7_75t_R _39750_ (.A(_10410_),
    .Y(_10550_));
 INVx6_ASAP7_75t_R _39751_ (.A(_10394_),
    .Y(_10551_));
 OAI21x1_ASAP7_75t_R _39752_ (.A1(_10550_),
    .A2(_10551_),
    .B(_10547_),
    .Y(_10552_));
 NAND2x1_ASAP7_75t_R _39753_ (.A(_10549_),
    .B(_10552_),
    .Y(_10553_));
 NOR2x2_ASAP7_75t_R _39754_ (.A(net956),
    .B(net973),
    .Y(_10554_));
 OAI21x1_ASAP7_75t_R _39755_ (.A1(_10554_),
    .A2(_10385_),
    .B(_10547_),
    .Y(_10556_));
 OA21x2_ASAP7_75t_R _39756_ (.A1(net1377),
    .A2(_10316_),
    .B(net1498),
    .Y(_10557_));
 NAND2x2_ASAP7_75t_R _39757_ (.A(_10547_),
    .B(_10557_),
    .Y(_10558_));
 NAND2x1_ASAP7_75t_R _39758_ (.A(_10556_),
    .B(_10558_),
    .Y(_10559_));
 NOR2x1_ASAP7_75t_R _39759_ (.A(_10553_),
    .B(_10559_),
    .Y(_10560_));
 NAND2x1_ASAP7_75t_R _39760_ (.A(_10543_),
    .B(_10560_),
    .Y(_10561_));
 NOR2x2_ASAP7_75t_R _39761_ (.A(_10535_),
    .B(_10561_),
    .Y(_10562_));
 INVx1_ASAP7_75t_R _39762_ (.A(_10562_),
    .Y(_10563_));
 TAPCELL_ASAP7_75t_R PHY_129 ();
 NOR2x2_ASAP7_75t_R _39764_ (.A(net2727),
    .B(_00570_),
    .Y(_10565_));
 NAND2x2_ASAP7_75t_R _39765_ (.A(_10565_),
    .B(_10497_),
    .Y(_10567_));
 TAPCELL_ASAP7_75t_R PHY_128 ();
 TAPCELL_ASAP7_75t_R PHY_127 ();
 AOI211x1_ASAP7_75t_R _39768_ (.A1(_10367_),
    .A2(net3338),
    .B(net2211),
    .C(_10341_),
    .Y(_10570_));
 INVx1_ASAP7_75t_R _39769_ (.A(_10570_),
    .Y(_10571_));
 INVx3_ASAP7_75t_R _39770_ (.A(_10567_),
    .Y(_10572_));
 NAND2x2_ASAP7_75t_R _39771_ (.A(net2454),
    .B(_10572_),
    .Y(_10573_));
 AO21x2_ASAP7_75t_R _39772_ (.A1(net2854),
    .A2(net3161),
    .B(net2211),
    .Y(_10574_));
 NAND3x2_ASAP7_75t_R _39773_ (.B(_10573_),
    .C(_10574_),
    .Y(_10575_),
    .A(_10571_));
 NOR2x2_ASAP7_75t_R _39774_ (.A(net2188),
    .B(net3296),
    .Y(_10576_));
 NAND2x2_ASAP7_75t_R _39775_ (.A(_10565_),
    .B(_10355_),
    .Y(_10578_));
 INVx3_ASAP7_75t_R _39776_ (.A(_10578_),
    .Y(_10579_));
 OA21x2_ASAP7_75t_R _39777_ (.A1(net2454),
    .A2(_10576_),
    .B(_10579_),
    .Y(_10580_));
 TAPCELL_ASAP7_75t_R PHY_126 ();
 NOR2x1_ASAP7_75t_R _39779_ (.A(net1515),
    .B(net1840),
    .Y(_10582_));
 AOI21x1_ASAP7_75t_R _39780_ (.A1(net1078),
    .A2(net1090),
    .B(net1840),
    .Y(_10583_));
 OR3x1_ASAP7_75t_R _39781_ (.A(_10580_),
    .B(_10582_),
    .C(_10583_),
    .Y(_10584_));
 NOR2x2_ASAP7_75t_R _39782_ (.A(_10575_),
    .B(_10584_),
    .Y(_10585_));
 NAND2x2_ASAP7_75t_R _39783_ (.A(_10565_),
    .B(_10430_),
    .Y(_10586_));
 AO21x2_ASAP7_75t_R _39784_ (.A1(_10329_),
    .A2(_10333_),
    .B(_10586_),
    .Y(_10587_));
 CKINVDCx6p67_ASAP7_75t_R _39785_ (.A(_10586_),
    .Y(_10589_));
 TAPCELL_ASAP7_75t_R PHY_125 ();
 OAI21x1_ASAP7_75t_R _39787_ (.A1(_10315_),
    .A2(net3018),
    .B(_10589_),
    .Y(_10591_));
 NOR2x1_ASAP7_75t_R _39788_ (.A(_10586_),
    .B(net2441),
    .Y(_10592_));
 INVx1_ASAP7_75t_R _39789_ (.A(_10592_),
    .Y(_10593_));
 NAND3x2_ASAP7_75t_R _39790_ (.B(_10591_),
    .C(_10593_),
    .Y(_10594_),
    .A(_10587_));
 AOI211x1_ASAP7_75t_R _39791_ (.A1(net975),
    .A2(net1318),
    .B(net2227),
    .C(net967),
    .Y(_10595_));
 AO21x1_ASAP7_75t_R _39792_ (.A1(_10589_),
    .A2(_10531_),
    .B(_10595_),
    .Y(_10596_));
 NOR2x2_ASAP7_75t_R _39793_ (.A(_10367_),
    .B(net3011),
    .Y(_10597_));
 NOR2x1_ASAP7_75t_R _39794_ (.A(net3039),
    .B(_10490_),
    .Y(_10598_));
 NAND2x2_ASAP7_75t_R _39795_ (.A(_10565_),
    .B(_10414_),
    .Y(_10600_));
 INVx3_ASAP7_75t_R _39796_ (.A(_10600_),
    .Y(_10601_));
 OAI21x1_ASAP7_75t_R _39797_ (.A1(_10597_),
    .A2(_10598_),
    .B(_10601_),
    .Y(_10602_));
 TAPCELL_ASAP7_75t_R PHY_124 ();
 NAND2x2_ASAP7_75t_R _39799_ (.A(_10317_),
    .B(net1740),
    .Y(_10604_));
 NOR2x1_ASAP7_75t_R _39800_ (.A(net2180),
    .B(_10604_),
    .Y(_10605_));
 TAPCELL_ASAP7_75t_R PHY_123 ();
 AOI21x1_ASAP7_75t_R _39802_ (.A1(net1051),
    .A2(net1077),
    .B(net2180),
    .Y(_10607_));
 NOR2x1_ASAP7_75t_R _39803_ (.A(_10605_),
    .B(_10607_),
    .Y(_10608_));
 NAND2x2_ASAP7_75t_R _39804_ (.A(_10602_),
    .B(_10608_),
    .Y(_10609_));
 NOR3x2_ASAP7_75t_R _39805_ (.B(_10596_),
    .C(_10609_),
    .Y(_10611_),
    .A(_10594_));
 NAND2x1_ASAP7_75t_R _39806_ (.A(_10585_),
    .B(_10611_),
    .Y(_10612_));
 NOR2x1_ASAP7_75t_R _39807_ (.A(_10563_),
    .B(_10612_),
    .Y(_10613_));
 NAND2x2_ASAP7_75t_R _39808_ (.A(_10513_),
    .B(_10613_),
    .Y(_10614_));
 NOR2x2_ASAP7_75t_R _39809_ (.A(_10364_),
    .B(_10614_),
    .Y(_10615_));
 TAPCELL_ASAP7_75t_R PHY_122 ();
 TAPCELL_ASAP7_75t_R PHY_121 ();
 NOR2x2_ASAP7_75t_R _39812_ (.A(net2933),
    .B(net3028),
    .Y(_10618_));
 TAPCELL_ASAP7_75t_R PHY_120 ();
 TAPCELL_ASAP7_75t_R PHY_119 ();
 NAND2x2_ASAP7_75t_R _39815_ (.A(net1716),
    .B(net1421),
    .Y(_10622_));
 INVx3_ASAP7_75t_R _39816_ (.A(_10622_),
    .Y(_10623_));
 NAND2x2_ASAP7_75t_R _39817_ (.A(net1336),
    .B(_10623_),
    .Y(_10624_));
 TAPCELL_ASAP7_75t_R PHY_118 ();
 CKINVDCx16_ASAP7_75t_R _39819_ (.A(net1716),
    .Y(_10626_));
 NOR2x2_ASAP7_75t_R _39820_ (.A(net1416),
    .B(_10626_),
    .Y(_10627_));
 NAND2x2_ASAP7_75t_R _39821_ (.A(net1338),
    .B(_10627_),
    .Y(_10628_));
 TAPCELL_ASAP7_75t_R PHY_117 ();
 TAPCELL_ASAP7_75t_R PHY_116 ();
 INVx2_ASAP7_75t_R _39824_ (.A(_00531_),
    .Y(_10631_));
 NOR2x2_ASAP7_75t_R _39825_ (.A(_00532_),
    .B(_10631_),
    .Y(_10633_));
 TAPCELL_ASAP7_75t_R PHY_115 ();
 TAPCELL_ASAP7_75t_R PHY_114 ();
 AND2x6_ASAP7_75t_R _39828_ (.A(_00529_),
    .B(_00530_),
    .Y(_10636_));
 NAND2x2_ASAP7_75t_R _39829_ (.A(_10633_),
    .B(_10636_),
    .Y(_10637_));
 AO21x1_ASAP7_75t_R _39830_ (.A1(_10624_),
    .A2(_10628_),
    .B(_10637_),
    .Y(_10638_));
 NAND2x2_ASAP7_75t_R _39831_ (.A(_00529_),
    .B(_00530_),
    .Y(_10639_));
 INVx2_ASAP7_75t_R _39832_ (.A(_00532_),
    .Y(_10640_));
 NAND2x1_ASAP7_75t_R _39833_ (.A(_00531_),
    .B(_10640_),
    .Y(_10641_));
 NOR2x2_ASAP7_75t_R _39834_ (.A(_10639_),
    .B(_10641_),
    .Y(_10642_));
 NOR2x2_ASAP7_75t_R _39835_ (.A(_00535_),
    .B(net1415),
    .Y(_10644_));
 NAND2x2_ASAP7_75t_R _39836_ (.A(_10618_),
    .B(_10644_),
    .Y(_10645_));
 TAPCELL_ASAP7_75t_R PHY_113 ();
 INVx1_ASAP7_75t_R _39838_ (.A(_10645_),
    .Y(_10647_));
 NAND2x1_ASAP7_75t_R _39839_ (.A(_10642_),
    .B(_10647_),
    .Y(_10648_));
 INVx2_ASAP7_75t_R _39840_ (.A(_00534_),
    .Y(_10649_));
 NOR2x2_ASAP7_75t_R _39841_ (.A(net2933),
    .B(_10649_),
    .Y(_10650_));
 TAPCELL_ASAP7_75t_R PHY_112 ();
 NAND2x2_ASAP7_75t_R _39843_ (.A(net1347),
    .B(_10642_),
    .Y(_10652_));
 NAND3x1_ASAP7_75t_R _39844_ (.A(_10638_),
    .B(_10648_),
    .C(_10652_),
    .Y(_10653_));
 TAPCELL_ASAP7_75t_R PHY_111 ();
 NAND2x2_ASAP7_75t_R _39846_ (.A(net1721),
    .B(net1336),
    .Y(_10656_));
 TAPCELL_ASAP7_75t_R PHY_110 ();
 CKINVDCx20_ASAP7_75t_R _39848_ (.A(net1416),
    .Y(_10658_));
 NOR2x2_ASAP7_75t_R _39849_ (.A(net1716),
    .B(_10658_),
    .Y(_10659_));
 NAND2x2_ASAP7_75t_R _39850_ (.A(net1336),
    .B(_10659_),
    .Y(_10660_));
 TAPCELL_ASAP7_75t_R PHY_109 ();
 NAND2x2_ASAP7_75t_R _39852_ (.A(_00531_),
    .B(_00532_),
    .Y(_10662_));
 INVx3_ASAP7_75t_R _39853_ (.A(_10662_),
    .Y(_10663_));
 NAND2x2_ASAP7_75t_R _39854_ (.A(_10636_),
    .B(_10663_),
    .Y(_10664_));
 TAPCELL_ASAP7_75t_R PHY_108 ();
 AO21x1_ASAP7_75t_R _39856_ (.A1(_10656_),
    .A2(_10660_),
    .B(_10664_),
    .Y(_10667_));
 INVx3_ASAP7_75t_R _39857_ (.A(net2933),
    .Y(_10668_));
 NOR2x2_ASAP7_75t_R _39858_ (.A(net3025),
    .B(_10668_),
    .Y(_10669_));
 TAPCELL_ASAP7_75t_R PHY_107 ();
 NAND2x2_ASAP7_75t_R _39860_ (.A(_10669_),
    .B(_10623_),
    .Y(_10671_));
 NAND2x2_ASAP7_75t_R _39861_ (.A(_10644_),
    .B(_10669_),
    .Y(_10672_));
 TAPCELL_ASAP7_75t_R PHY_106 ();
 AO21x1_ASAP7_75t_R _39863_ (.A1(_10671_),
    .A2(_10672_),
    .B(_10664_),
    .Y(_10674_));
 NAND2x1_ASAP7_75t_R _39864_ (.A(_10667_),
    .B(_10674_),
    .Y(_10675_));
 AND2x6_ASAP7_75t_R _39865_ (.A(net2933),
    .B(_00534_),
    .Y(_10677_));
 NAND2x2_ASAP7_75t_R _39866_ (.A(_10659_),
    .B(_10677_),
    .Y(_10678_));
 TAPCELL_ASAP7_75t_R PHY_105 ();
 NAND2x2_ASAP7_75t_R _39868_ (.A(net2934),
    .B(net3024),
    .Y(_10680_));
 NOR2x2_ASAP7_75t_R _39869_ (.A(_10626_),
    .B(net1995),
    .Y(_10681_));
 INVx2_ASAP7_75t_R _39870_ (.A(_10681_),
    .Y(_10682_));
 AO21x1_ASAP7_75t_R _39871_ (.A1(_10678_),
    .A2(_10682_),
    .B(_10637_),
    .Y(_10683_));
 INVx3_ASAP7_75t_R _39872_ (.A(_10644_),
    .Y(_10684_));
 NAND2x2_ASAP7_75t_R _39873_ (.A(net2933),
    .B(_10649_),
    .Y(_10685_));
 AO21x1_ASAP7_75t_R _39874_ (.A1(_10684_),
    .A2(_10622_),
    .B(net2026),
    .Y(_10686_));
 NOR2x2_ASAP7_75t_R _39875_ (.A(_10637_),
    .B(_10686_),
    .Y(_10688_));
 INVx1_ASAP7_75t_R _39876_ (.A(_10688_),
    .Y(_10689_));
 NAND2x1_ASAP7_75t_R _39877_ (.A(_10683_),
    .B(_10689_),
    .Y(_10690_));
 NOR3x1_ASAP7_75t_R _39878_ (.A(_10653_),
    .B(_10675_),
    .C(_10690_),
    .Y(_10691_));
 TAPCELL_ASAP7_75t_R PHY_104 ();
 NAND2x2_ASAP7_75t_R _39880_ (.A(_10658_),
    .B(_10677_),
    .Y(_10693_));
 NAND2x2_ASAP7_75t_R _39881_ (.A(_10658_),
    .B(_10669_),
    .Y(_10694_));
 NOR2x2_ASAP7_75t_R _39882_ (.A(_00531_),
    .B(_00532_),
    .Y(_10695_));
 NAND2x2_ASAP7_75t_R _39883_ (.A(_10695_),
    .B(_10636_),
    .Y(_10696_));
 TAPCELL_ASAP7_75t_R PHY_103 ();
 AO21x1_ASAP7_75t_R _39885_ (.A1(_10693_),
    .A2(_10694_),
    .B(_10696_),
    .Y(_10699_));
 NAND2x2_ASAP7_75t_R _39886_ (.A(_10626_),
    .B(net2147),
    .Y(_10700_));
 NAND2x2_ASAP7_75t_R _39887_ (.A(net1417),
    .B(net1339),
    .Y(_10701_));
 AO21x1_ASAP7_75t_R _39888_ (.A1(_10700_),
    .A2(_10701_),
    .B(_10696_),
    .Y(_10702_));
 AND2x2_ASAP7_75t_R _39889_ (.A(_10699_),
    .B(_10702_),
    .Y(_10703_));
 NOR2x2_ASAP7_75t_R _39890_ (.A(_00531_),
    .B(_10640_),
    .Y(_10704_));
 NAND2x2_ASAP7_75t_R _39891_ (.A(_10704_),
    .B(_10636_),
    .Y(_10705_));
 NAND2x1_ASAP7_75t_R _39892_ (.A(_10677_),
    .B(_10684_),
    .Y(_10706_));
 NOR2x2_ASAP7_75t_R _39893_ (.A(_10705_),
    .B(_10706_),
    .Y(_10707_));
 NOR2x2_ASAP7_75t_R _39894_ (.A(net2021),
    .B(_10684_),
    .Y(_10708_));
 NAND2x2_ASAP7_75t_R _39895_ (.A(net1421),
    .B(_10626_),
    .Y(_10710_));
 NOR2x2_ASAP7_75t_R _39896_ (.A(_10710_),
    .B(_10685_),
    .Y(_10711_));
 NAND2x2_ASAP7_75t_R _39897_ (.A(_00532_),
    .B(_10631_),
    .Y(_10712_));
 NOR2x2_ASAP7_75t_R _39898_ (.A(_10639_),
    .B(_10712_),
    .Y(_10713_));
 OA21x2_ASAP7_75t_R _39899_ (.A1(_10708_),
    .A2(_10711_),
    .B(_10713_),
    .Y(_10714_));
 NOR2x1_ASAP7_75t_R _39900_ (.A(_10707_),
    .B(_10714_),
    .Y(_10715_));
 TAPCELL_ASAP7_75t_R PHY_102 ();
 NAND2x2_ASAP7_75t_R _39902_ (.A(_10622_),
    .B(net1343),
    .Y(_10717_));
 TAPCELL_ASAP7_75t_R PHY_101 ();
 AO21x1_ASAP7_75t_R _39904_ (.A1(net3048),
    .A2(_10717_),
    .B(_10705_),
    .Y(_10719_));
 AND3x1_ASAP7_75t_R _39905_ (.A(_10703_),
    .B(_10715_),
    .C(_10719_),
    .Y(_10721_));
 NAND2x1_ASAP7_75t_R _39906_ (.A(_10691_),
    .B(_10721_),
    .Y(_10722_));
 INVx4_ASAP7_75t_R _39907_ (.A(_00529_),
    .Y(_10723_));
 NOR2x2_ASAP7_75t_R _39908_ (.A(_00530_),
    .B(_10723_),
    .Y(_10724_));
 NAND2x2_ASAP7_75t_R _39909_ (.A(_10704_),
    .B(_10724_),
    .Y(_10725_));
 AO21x1_ASAP7_75t_R _39910_ (.A1(_10660_),
    .A2(_10645_),
    .B(_10725_),
    .Y(_10726_));
 TAPCELL_ASAP7_75t_R PHY_100 ();
 TAPCELL_ASAP7_75t_R PHY_99 ();
 AO21x1_ASAP7_75t_R _39913_ (.A1(_10672_),
    .A2(net1996),
    .B(_10725_),
    .Y(_10729_));
 NAND2x2_ASAP7_75t_R _39914_ (.A(net1718),
    .B(_10658_),
    .Y(_10730_));
 NAND2x2_ASAP7_75t_R _39915_ (.A(net3026),
    .B(_10668_),
    .Y(_10732_));
 NOR2x2_ASAP7_75t_R _39916_ (.A(_10730_),
    .B(_10732_),
    .Y(_10733_));
 INVx4_ASAP7_75t_R _39917_ (.A(_00530_),
    .Y(_10734_));
 NAND2x2_ASAP7_75t_R _39918_ (.A(_00529_),
    .B(_10734_),
    .Y(_10735_));
 NOR2x2_ASAP7_75t_R _39919_ (.A(_10712_),
    .B(_10735_),
    .Y(_10736_));
 NAND2x1_ASAP7_75t_R _39920_ (.A(_10733_),
    .B(_10736_),
    .Y(_10737_));
 NAND3x1_ASAP7_75t_R _39921_ (.A(_10726_),
    .B(_10729_),
    .C(_10737_),
    .Y(_10738_));
 NAND2x2_ASAP7_75t_R _39922_ (.A(_10695_),
    .B(_10724_),
    .Y(_10739_));
 CKINVDCx14_ASAP7_75t_R _39923_ (.A(net1338),
    .Y(_10740_));
 AOI211x1_ASAP7_75t_R _39924_ (.A1(net1720),
    .A2(net1422),
    .B(_10739_),
    .C(_10740_),
    .Y(_10741_));
 INVx1_ASAP7_75t_R _39925_ (.A(_10741_),
    .Y(_10743_));
 NAND2x2_ASAP7_75t_R _39926_ (.A(_10627_),
    .B(net2147),
    .Y(_10744_));
 NAND2x2_ASAP7_75t_R _39927_ (.A(net1422),
    .B(net1344),
    .Y(_10745_));
 AO21x1_ASAP7_75t_R _39928_ (.A1(_10744_),
    .A2(_10745_),
    .B(_10739_),
    .Y(_10746_));
 NAND2x2_ASAP7_75t_R _39929_ (.A(_10710_),
    .B(net2118),
    .Y(_10747_));
 AO21x1_ASAP7_75t_R _39930_ (.A1(_10747_),
    .A2(_10693_),
    .B(_10739_),
    .Y(_10748_));
 NAND3x1_ASAP7_75t_R _39931_ (.A(_10743_),
    .B(_10746_),
    .C(_10748_),
    .Y(_10749_));
 NOR2x1_ASAP7_75t_R _39932_ (.A(_10738_),
    .B(_10749_),
    .Y(_10750_));
 NAND2x2_ASAP7_75t_R _39933_ (.A(_10627_),
    .B(_10677_),
    .Y(_10751_));
 TAPCELL_ASAP7_75t_R PHY_98 ();
 NOR2x2_ASAP7_75t_R _39935_ (.A(_10662_),
    .B(_10735_),
    .Y(_10754_));
 CKINVDCx5p33_ASAP7_75t_R _39936_ (.A(_10754_),
    .Y(_10755_));
 AO21x1_ASAP7_75t_R _39937_ (.A1(net3053),
    .A2(net2061),
    .B(_10755_),
    .Y(_10756_));
 NAND2x2_ASAP7_75t_R _39938_ (.A(_10659_),
    .B(net2147),
    .Y(_10757_));
 TAPCELL_ASAP7_75t_R PHY_97 ();
 NAND2x2_ASAP7_75t_R _39940_ (.A(_10644_),
    .B(net2147),
    .Y(_10759_));
 TAPCELL_ASAP7_75t_R PHY_96 ();
 TAPCELL_ASAP7_75t_R PHY_95 ();
 AO21x1_ASAP7_75t_R _39943_ (.A1(_10757_),
    .A2(_10759_),
    .B(_10755_),
    .Y(_10762_));
 TAPCELL_ASAP7_75t_R PHY_94 ();
 AO21x1_ASAP7_75t_R _39945_ (.A1(net3048),
    .A2(net3058),
    .B(_10755_),
    .Y(_10765_));
 AND3x1_ASAP7_75t_R _39946_ (.A(_10756_),
    .B(_10762_),
    .C(_10765_),
    .Y(_10766_));
 NAND2x2_ASAP7_75t_R _39947_ (.A(_10669_),
    .B(_10627_),
    .Y(_10767_));
 NAND2x2_ASAP7_75t_R _39948_ (.A(_10659_),
    .B(_10669_),
    .Y(_10768_));
 NAND2x2_ASAP7_75t_R _39949_ (.A(_10633_),
    .B(_10724_),
    .Y(_10769_));
 AO21x1_ASAP7_75t_R _39950_ (.A1(_10767_),
    .A2(net2781),
    .B(net3040),
    .Y(_10770_));
 NAND2x2_ASAP7_75t_R _39951_ (.A(_10644_),
    .B(_10677_),
    .Y(_10771_));
 AO21x1_ASAP7_75t_R _39952_ (.A1(_10751_),
    .A2(_10771_),
    .B(net3040),
    .Y(_10772_));
 AND2x2_ASAP7_75t_R _39953_ (.A(_10770_),
    .B(_10772_),
    .Y(_10773_));
 INVx3_ASAP7_75t_R _39954_ (.A(net3040),
    .Y(_10774_));
 NOR2x1_ASAP7_75t_R _39955_ (.A(net3040),
    .B(_10757_),
    .Y(_10776_));
 NOR2x1_ASAP7_75t_R _39956_ (.A(_10645_),
    .B(net3040),
    .Y(_10777_));
 AOI211x1_ASAP7_75t_R _39957_ (.A1(_10774_),
    .A2(_10733_),
    .B(_10776_),
    .C(_10777_),
    .Y(_10778_));
 AND2x2_ASAP7_75t_R _39958_ (.A(_10773_),
    .B(_10778_),
    .Y(_10779_));
 NAND3x1_ASAP7_75t_R _39959_ (.A(_10750_),
    .B(_10766_),
    .C(_10779_),
    .Y(_10780_));
 NOR2x1_ASAP7_75t_R _39960_ (.A(_10722_),
    .B(_10780_),
    .Y(_10781_));
 NOR2x2_ASAP7_75t_R _39961_ (.A(_10622_),
    .B(_10680_),
    .Y(_10782_));
 CKINVDCx9p33_ASAP7_75t_R _39962_ (.A(_10782_),
    .Y(_10783_));
 NOR2x2_ASAP7_75t_R _39963_ (.A(_00529_),
    .B(_10734_),
    .Y(_10784_));
 NAND2x2_ASAP7_75t_R _39964_ (.A(_10784_),
    .B(_10663_),
    .Y(_10785_));
 AO21x1_ASAP7_75t_R _39965_ (.A1(_10783_),
    .A2(_10771_),
    .B(_10785_),
    .Y(_10787_));
 NAND2x2_ASAP7_75t_R _39966_ (.A(net1343),
    .B(_10623_),
    .Y(_10788_));
 AO21x1_ASAP7_75t_R _39967_ (.A1(_10744_),
    .A2(_10788_),
    .B(_10785_),
    .Y(_10789_));
 NAND2x2_ASAP7_75t_R _39968_ (.A(_00530_),
    .B(_10723_),
    .Y(_10790_));
 NOR2x2_ASAP7_75t_R _39969_ (.A(_10662_),
    .B(_10790_),
    .Y(_10791_));
 NOR2x2_ASAP7_75t_R _39970_ (.A(_10730_),
    .B(net2021),
    .Y(_10792_));
 NAND2x1_ASAP7_75t_R _39971_ (.A(_10791_),
    .B(_10792_),
    .Y(_10793_));
 NAND3x1_ASAP7_75t_R _39972_ (.A(_10787_),
    .B(_10789_),
    .C(_10793_),
    .Y(_10794_));
 TAPCELL_ASAP7_75t_R PHY_93 ();
 NAND2x2_ASAP7_75t_R _39974_ (.A(_10633_),
    .B(_10784_),
    .Y(_10796_));
 TAPCELL_ASAP7_75t_R PHY_92 ();
 AO21x1_ASAP7_75t_R _39976_ (.A1(net2781),
    .A2(_10672_),
    .B(_10796_),
    .Y(_10799_));
 TAPCELL_ASAP7_75t_R PHY_91 ();
 AO21x1_ASAP7_75t_R _39978_ (.A1(_10751_),
    .A2(_10771_),
    .B(_10796_),
    .Y(_10801_));
 NAND2x1_ASAP7_75t_R _39979_ (.A(_10799_),
    .B(_10801_),
    .Y(_10802_));
 AO21x1_ASAP7_75t_R _39980_ (.A1(_10624_),
    .A2(_10645_),
    .B(_10796_),
    .Y(_10803_));
 AO21x1_ASAP7_75t_R _39981_ (.A1(_10744_),
    .A2(_10757_),
    .B(_10796_),
    .Y(_10804_));
 NAND2x1_ASAP7_75t_R _39982_ (.A(_10803_),
    .B(_10804_),
    .Y(_10805_));
 NOR3x1_ASAP7_75t_R _39983_ (.A(_10794_),
    .B(_10802_),
    .C(_10805_),
    .Y(_10806_));
 NAND2x2_ASAP7_75t_R _39984_ (.A(net1716),
    .B(net1342),
    .Y(_10807_));
 NOR2x2_ASAP7_75t_R _39985_ (.A(_10712_),
    .B(_10790_),
    .Y(_10809_));
 INVx3_ASAP7_75t_R _39986_ (.A(_10809_),
    .Y(_10810_));
 AO21x1_ASAP7_75t_R _39987_ (.A1(_10807_),
    .A2(_10757_),
    .B(_10810_),
    .Y(_10811_));
 AO21x1_ASAP7_75t_R _39988_ (.A1(_10660_),
    .A2(_10656_),
    .B(_10810_),
    .Y(_10812_));
 AND2x2_ASAP7_75t_R _39989_ (.A(_10811_),
    .B(_10812_),
    .Y(_10813_));
 NOR2x1_ASAP7_75t_R _39990_ (.A(_10783_),
    .B(_10810_),
    .Y(_10814_));
 INVx1_ASAP7_75t_R _39991_ (.A(_10814_),
    .Y(_10815_));
 NAND2x2_ASAP7_75t_R _39992_ (.A(_10695_),
    .B(_10784_),
    .Y(_10816_));
 TAPCELL_ASAP7_75t_R PHY_90 ();
 AO21x1_ASAP7_75t_R _39994_ (.A1(_10682_),
    .A2(_10747_),
    .B(_10816_),
    .Y(_10818_));
 TAPCELL_ASAP7_75t_R PHY_89 ();
 AO21x1_ASAP7_75t_R _39996_ (.A1(_10660_),
    .A2(_10700_),
    .B(_10816_),
    .Y(_10821_));
 AND2x2_ASAP7_75t_R _39997_ (.A(_10818_),
    .B(_10821_),
    .Y(_10822_));
 AND3x1_ASAP7_75t_R _39998_ (.A(_10813_),
    .B(_10815_),
    .C(_10822_),
    .Y(_10823_));
 NAND2x1_ASAP7_75t_R _39999_ (.A(_10806_),
    .B(_10823_),
    .Y(_10824_));
 NOR2x2_ASAP7_75t_R _40000_ (.A(_00529_),
    .B(_00530_),
    .Y(_10825_));
 NAND2x2_ASAP7_75t_R _40001_ (.A(_10825_),
    .B(_10663_),
    .Y(_10826_));
 INVx3_ASAP7_75t_R _40002_ (.A(_10826_),
    .Y(_10827_));
 NOR2x1_ASAP7_75t_R _40003_ (.A(_10807_),
    .B(_10826_),
    .Y(_10828_));
 INVx1_ASAP7_75t_R _40004_ (.A(_10828_),
    .Y(_10829_));
 NOR2x2_ASAP7_75t_R _40005_ (.A(net1719),
    .B(_10740_),
    .Y(_10831_));
 INVx4_ASAP7_75t_R _40006_ (.A(_10831_),
    .Y(_10832_));
 TAPCELL_ASAP7_75t_R PHY_88 ();
 AO21x1_ASAP7_75t_R _40008_ (.A1(_10832_),
    .A2(net3047),
    .B(_10826_),
    .Y(_10834_));
 NAND2x1_ASAP7_75t_R _40009_ (.A(_10829_),
    .B(_10834_),
    .Y(_10835_));
 TAPCELL_ASAP7_75t_R PHY_87 ();
 TAPCELL_ASAP7_75t_R PHY_86 ();
 TAPCELL_ASAP7_75t_R PHY_85 ();
 AOI211x1_ASAP7_75t_R _40013_ (.A1(net1501),
    .A2(net1420),
    .B(_10826_),
    .C(net2023),
    .Y(_10839_));
 AOI211x1_ASAP7_75t_R _40014_ (.A1(net3068),
    .A2(_10827_),
    .B(_10835_),
    .C(_10839_),
    .Y(_10840_));
 TAPCELL_ASAP7_75t_R PHY_84 ();
 NAND2x2_ASAP7_75t_R _40016_ (.A(_10825_),
    .B(_10695_),
    .Y(_10843_));
 AOI211x1_ASAP7_75t_R _40017_ (.A1(_10626_),
    .A2(_10658_),
    .B(_10843_),
    .C(net1991),
    .Y(_10844_));
 INVx1_ASAP7_75t_R _40018_ (.A(_10844_),
    .Y(_10845_));
 NOR2x2_ASAP7_75t_R _40019_ (.A(_10626_),
    .B(net2022),
    .Y(_10846_));
 INVx2_ASAP7_75t_R _40020_ (.A(_10843_),
    .Y(_10847_));
 NAND2x2_ASAP7_75t_R _40021_ (.A(_10846_),
    .B(_10847_),
    .Y(_10848_));
 AO21x1_ASAP7_75t_R _40022_ (.A1(_10744_),
    .A2(_10701_),
    .B(_10843_),
    .Y(_10849_));
 NAND3x2_ASAP7_75t_R _40023_ (.B(_10848_),
    .C(_10849_),
    .Y(_10850_),
    .A(_10845_));
 NAND2x2_ASAP7_75t_R _40024_ (.A(_10825_),
    .B(_10704_),
    .Y(_10851_));
 TAPCELL_ASAP7_75t_R PHY_83 ();
 NAND2x2_ASAP7_75t_R _40026_ (.A(_10730_),
    .B(net1344),
    .Y(_10854_));
 NOR2x1_ASAP7_75t_R _40027_ (.A(_10851_),
    .B(_10854_),
    .Y(_10855_));
 AOI21x1_ASAP7_75t_R _40028_ (.A1(_10645_),
    .A2(_10624_),
    .B(_10851_),
    .Y(_10856_));
 NOR2x1_ASAP7_75t_R _40029_ (.A(_10855_),
    .B(_10856_),
    .Y(_10857_));
 AOI211x1_ASAP7_75t_R _40030_ (.A1(_10626_),
    .A2(_10658_),
    .B(net1992),
    .C(_10851_),
    .Y(_10858_));
 AOI211x1_ASAP7_75t_R _40031_ (.A1(net1717),
    .A2(net1418),
    .B(net2022),
    .C(_10851_),
    .Y(_10859_));
 NOR2x1_ASAP7_75t_R _40032_ (.A(_10858_),
    .B(_10859_),
    .Y(_10860_));
 NAND2x1_ASAP7_75t_R _40033_ (.A(_10857_),
    .B(_10860_),
    .Y(_10861_));
 NOR2x2_ASAP7_75t_R _40034_ (.A(_10850_),
    .B(_10861_),
    .Y(_10862_));
 NAND2x2_ASAP7_75t_R _40035_ (.A(_10825_),
    .B(_10633_),
    .Y(_10864_));
 TAPCELL_ASAP7_75t_R PHY_82 ();
 TAPCELL_ASAP7_75t_R PHY_81 ();
 AOI211x1_ASAP7_75t_R _40038_ (.A1(_10626_),
    .A2(net1418),
    .B(_10864_),
    .C(_10740_),
    .Y(_10867_));
 INVx1_ASAP7_75t_R _40039_ (.A(_10867_),
    .Y(_10868_));
 INVx4_ASAP7_75t_R _40040_ (.A(_10759_),
    .Y(_10869_));
 INVx3_ASAP7_75t_R _40041_ (.A(_10864_),
    .Y(_10870_));
 NAND2x1_ASAP7_75t_R _40042_ (.A(_10869_),
    .B(_10870_),
    .Y(_10871_));
 AO21x1_ASAP7_75t_R _40043_ (.A1(_10678_),
    .A2(_10768_),
    .B(_10864_),
    .Y(_10872_));
 AND3x2_ASAP7_75t_R _40044_ (.A(_10868_),
    .B(_10871_),
    .C(_10872_),
    .Y(_10873_));
 NAND3x2_ASAP7_75t_R _40045_ (.B(_10862_),
    .C(_10873_),
    .Y(_10875_),
    .A(_10840_));
 NOR2x2_ASAP7_75t_R _40046_ (.A(_10824_),
    .B(_10875_),
    .Y(_10876_));
 NAND2x2_ASAP7_75t_R _40047_ (.A(_10781_),
    .B(_10876_),
    .Y(_10877_));
 INVx2_ASAP7_75t_R _40048_ (.A(_10877_),
    .Y(_10878_));
 XOR2x1_ASAP7_75t_R _40049_ (.A(_10615_),
    .Y(_10879_),
    .B(_10878_));
 INVx1_ASAP7_75t_R _40050_ (.A(_10879_),
    .Y(_10880_));
 OAI21x1_ASAP7_75t_R _40051_ (.A1(_10305_),
    .A2(_10308_),
    .B(_10880_),
    .Y(_10881_));
 AO21x1_ASAP7_75t_R _40052_ (.A1(_10303_),
    .A2(_10288_),
    .B(_09867_),
    .Y(_10882_));
 INVx3_ASAP7_75t_R _40053_ (.A(_10121_),
    .Y(_10883_));
 NAND2x2_ASAP7_75t_R _40054_ (.A(net2681),
    .B(_10286_),
    .Y(_10884_));
 NOR2x2_ASAP7_75t_R _40055_ (.A(_10883_),
    .B(_10884_),
    .Y(_10886_));
 NOR2x1_ASAP7_75t_R _40056_ (.A(_10287_),
    .B(_10886_),
    .Y(_10887_));
 NAND2x1_ASAP7_75t_R _40057_ (.A(_09867_),
    .B(_10887_),
    .Y(_10888_));
 AOI21x1_ASAP7_75t_R _40058_ (.A1(_10882_),
    .A2(_10888_),
    .B(_10880_),
    .Y(_10889_));
 INVx1_ASAP7_75t_R _40059_ (.A(_10889_),
    .Y(_10890_));
 AOI21x1_ASAP7_75t_R _40060_ (.A1(_10881_),
    .A2(_10890_),
    .B(net389),
    .Y(_10891_));
 OAI21x1_ASAP7_75t_R _40061_ (.A1(_09569_),
    .A2(_10891_),
    .B(_00409_),
    .Y(_10892_));
 NAND2x1_ASAP7_75t_R _40062_ (.A(_10306_),
    .B(_10887_),
    .Y(_10893_));
 AOI21x1_ASAP7_75t_R _40063_ (.A1(_10307_),
    .A2(_10893_),
    .B(_10879_),
    .Y(_10894_));
 OAI21x1_ASAP7_75t_R _40064_ (.A1(_10894_),
    .A2(_10889_),
    .B(net392),
    .Y(_10895_));
 INVx2_ASAP7_75t_R _40065_ (.A(_00409_),
    .Y(_10897_));
 INVx1_ASAP7_75t_R _40066_ (.A(_09569_),
    .Y(_10898_));
 NAND3x2_ASAP7_75t_R _40067_ (.B(_10897_),
    .C(_10898_),
    .Y(_10899_),
    .A(_10895_));
 NAND2x2_ASAP7_75t_R _40068_ (.A(_10892_),
    .B(_10899_),
    .Y(_00097_));
 AND2x2_ASAP7_75t_R _40069_ (.A(net389),
    .B(_00818_),
    .Y(_10900_));
 NAND2x1_ASAP7_75t_R _40070_ (.A(_10622_),
    .B(_10684_),
    .Y(_10901_));
 INVx2_ASAP7_75t_R _40071_ (.A(_10901_),
    .Y(_10902_));
 NOR2x2_ASAP7_75t_R _40072_ (.A(_10902_),
    .B(_10652_),
    .Y(_10903_));
 OA21x2_ASAP7_75t_R _40073_ (.A1(_10792_),
    .A2(_10711_),
    .B(_10642_),
    .Y(_10904_));
 NAND2x2_ASAP7_75t_R _40074_ (.A(_10626_),
    .B(_10677_),
    .Y(_10905_));
 TAPCELL_ASAP7_75t_R PHY_80 ();
 NOR2x1_ASAP7_75t_R _40076_ (.A(_10905_),
    .B(_10637_),
    .Y(_10908_));
 OR3x1_ASAP7_75t_R _40077_ (.A(_10903_),
    .B(_10904_),
    .C(_10908_),
    .Y(_10909_));
 TAPCELL_ASAP7_75t_R PHY_79 ();
 AOI211x1_ASAP7_75t_R _40079_ (.A1(net1501),
    .A2(net1425),
    .B(net3021),
    .C(_10685_),
    .Y(_10911_));
 AO21x1_ASAP7_75t_R _40080_ (.A1(_10678_),
    .A2(_10771_),
    .B(_10664_),
    .Y(_10912_));
 INVx1_ASAP7_75t_R _40081_ (.A(_10912_),
    .Y(_10913_));
 NOR2x1_ASAP7_75t_R _40082_ (.A(_10911_),
    .B(_10913_),
    .Y(_10914_));
 AO21x1_ASAP7_75t_R _40083_ (.A1(net1288),
    .A2(_10660_),
    .B(net3021),
    .Y(_10915_));
 OA21x2_ASAP7_75t_R _40084_ (.A1(_10717_),
    .A2(net3021),
    .B(_10915_),
    .Y(_10916_));
 NAND2x1_ASAP7_75t_R _40085_ (.A(_10914_),
    .B(_10916_),
    .Y(_10918_));
 NOR2x1_ASAP7_75t_R _40086_ (.A(_10909_),
    .B(_10918_),
    .Y(_10919_));
 TAPCELL_ASAP7_75t_R PHY_78 ();
 AO21x1_ASAP7_75t_R _40088_ (.A1(net1501),
    .A2(net1421),
    .B(_10680_),
    .Y(_10921_));
 TAPCELL_ASAP7_75t_R PHY_77 ();
 AOI21x1_ASAP7_75t_R _40090_ (.A1(net1862),
    .A2(_10921_),
    .B(_10696_),
    .Y(_10923_));
 TAPCELL_ASAP7_75t_R PHY_76 ();
 NOR2x1_ASAP7_75t_R _40092_ (.A(_10696_),
    .B(_10788_),
    .Y(_10925_));
 AOI21x1_ASAP7_75t_R _40093_ (.A1(net3058),
    .A2(_10656_),
    .B(_10696_),
    .Y(_10926_));
 OR3x1_ASAP7_75t_R _40094_ (.A(_10923_),
    .B(_10925_),
    .C(_10926_),
    .Y(_10927_));
 OA21x2_ASAP7_75t_R _40095_ (.A1(_10792_),
    .A2(_10711_),
    .B(_10713_),
    .Y(_10929_));
 NOR2x1_ASAP7_75t_R _40096_ (.A(_10707_),
    .B(_10929_),
    .Y(_10930_));
 TAPCELL_ASAP7_75t_R PHY_75 ();
 AO21x1_ASAP7_75t_R _40098_ (.A1(net3022),
    .A2(_10700_),
    .B(_10705_),
    .Y(_10932_));
 TAPCELL_ASAP7_75t_R PHY_74 ();
 AO21x1_ASAP7_75t_R _40100_ (.A1(_10832_),
    .A2(net3020),
    .B(_10705_),
    .Y(_10934_));
 NAND3x1_ASAP7_75t_R _40101_ (.A(_10930_),
    .B(_10932_),
    .C(_10934_),
    .Y(_10935_));
 NOR2x1_ASAP7_75t_R _40102_ (.A(_10927_),
    .B(_10935_),
    .Y(_10936_));
 NAND2x1_ASAP7_75t_R _40103_ (.A(_10919_),
    .B(_10936_),
    .Y(_10937_));
 NAND2x2_ASAP7_75t_R _40104_ (.A(_10710_),
    .B(_10677_),
    .Y(_10938_));
 TAPCELL_ASAP7_75t_R PHY_73 ();
 NOR2x1_ASAP7_75t_R _40106_ (.A(_10938_),
    .B(net3040),
    .Y(_10941_));
 AOI21x1_ASAP7_75t_R _40107_ (.A1(net2061),
    .A2(net2053),
    .B(net3040),
    .Y(_10942_));
 NOR2x2_ASAP7_75t_R _40108_ (.A(_10941_),
    .B(_10942_),
    .Y(_10943_));
 INVx1_ASAP7_75t_R _40109_ (.A(_10777_),
    .Y(_10944_));
 AO21x1_ASAP7_75t_R _40110_ (.A1(_10744_),
    .A2(net1492),
    .B(net3040),
    .Y(_10945_));
 NAND3x2_ASAP7_75t_R _40111_ (.B(_10944_),
    .C(_10945_),
    .Y(_10946_),
    .A(_10943_));
 TAPCELL_ASAP7_75t_R PHY_72 ();
 TAPCELL_ASAP7_75t_R PHY_71 ();
 TAPCELL_ASAP7_75t_R PHY_70 ();
 TAPCELL_ASAP7_75t_R PHY_69 ();
 AO31x2_ASAP7_75t_R _40116_ (.A1(_10783_),
    .A2(net3053),
    .A3(_10671_),
    .B(_10755_),
    .Y(_10952_));
 OA21x2_ASAP7_75t_R _40117_ (.A1(_10869_),
    .A2(_10733_),
    .B(_10754_),
    .Y(_10953_));
 TAPCELL_ASAP7_75t_R PHY_68 ();
 AOI211x1_ASAP7_75t_R _40119_ (.A1(_10626_),
    .A2(_10658_),
    .B(_10755_),
    .C(_10740_),
    .Y(_10955_));
 NOR2x2_ASAP7_75t_R _40120_ (.A(_10953_),
    .B(_10955_),
    .Y(_10956_));
 NAND2x1_ASAP7_75t_R _40121_ (.A(_10952_),
    .B(_10956_),
    .Y(_10957_));
 NOR2x2_ASAP7_75t_R _40122_ (.A(_10946_),
    .B(_10957_),
    .Y(_10958_));
 AO21x2_ASAP7_75t_R _40123_ (.A1(_10768_),
    .A2(_10671_),
    .B(_10725_),
    .Y(_10959_));
 TAPCELL_ASAP7_75t_R PHY_67 ();
 AO21x2_ASAP7_75t_R _40125_ (.A1(_10767_),
    .A2(_10672_),
    .B(_10725_),
    .Y(_10962_));
 TAPCELL_ASAP7_75t_R PHY_66 ();
 AO21x1_ASAP7_75t_R _40127_ (.A1(net3065),
    .A2(net1475),
    .B(_10725_),
    .Y(_10964_));
 NAND3x2_ASAP7_75t_R _40128_ (.B(_10962_),
    .C(_10964_),
    .Y(_10965_),
    .A(_10959_));
 OR3x4_ASAP7_75t_R _40129_ (.A(_10725_),
    .B(net2935),
    .C(_10649_),
    .Y(_10966_));
 NOR2x2_ASAP7_75t_R _40130_ (.A(_10710_),
    .B(_10740_),
    .Y(_10967_));
 NAND2x2_ASAP7_75t_R _40131_ (.A(_10736_),
    .B(_10967_),
    .Y(_10968_));
 OAI21x1_ASAP7_75t_R _40132_ (.A1(_10659_),
    .A2(_10966_),
    .B(_10968_),
    .Y(_10969_));
 TAPCELL_ASAP7_75t_R PHY_65 ();
 NOR2x1_ASAP7_75t_R _40134_ (.A(_10759_),
    .B(_10739_),
    .Y(_10971_));
 TAPCELL_ASAP7_75t_R PHY_64 ();
 AOI21x1_ASAP7_75t_R _40136_ (.A1(net3046),
    .A2(_10660_),
    .B(_10739_),
    .Y(_10974_));
 NOR2x1_ASAP7_75t_R _40137_ (.A(_10971_),
    .B(_10974_),
    .Y(_10975_));
 AO31x2_ASAP7_75t_R _40138_ (.A1(_10694_),
    .A2(_10783_),
    .A3(_10693_),
    .B(_10739_),
    .Y(_10976_));
 NAND2x2_ASAP7_75t_R _40139_ (.A(_10975_),
    .B(_10976_),
    .Y(_10977_));
 NOR3x2_ASAP7_75t_R _40140_ (.B(_10969_),
    .C(_10977_),
    .Y(_10978_),
    .A(_10965_));
 NAND2x2_ASAP7_75t_R _40141_ (.A(_10958_),
    .B(_10978_),
    .Y(_10979_));
 NOR2x2_ASAP7_75t_R _40142_ (.A(_10937_),
    .B(_10979_),
    .Y(_10980_));
 AO21x1_ASAP7_75t_R _40143_ (.A1(_10740_),
    .A2(_10732_),
    .B(_10664_),
    .Y(_10981_));
 OR3x1_ASAP7_75t_R _40144_ (.A(_10685_),
    .B(_10639_),
    .C(_10662_),
    .Y(_10982_));
 AO21x1_ASAP7_75t_R _40145_ (.A1(_10693_),
    .A2(_10905_),
    .B(_10664_),
    .Y(_10984_));
 NAND2x1_ASAP7_75t_R _40146_ (.A(_10982_),
    .B(_10984_),
    .Y(_10985_));
 INVx1_ASAP7_75t_R _40147_ (.A(_10985_),
    .Y(_10986_));
 NAND2x2_ASAP7_75t_R _40148_ (.A(_10981_),
    .B(_10986_),
    .Y(_10987_));
 OR3x2_ASAP7_75t_R _40149_ (.A(_10723_),
    .B(_10734_),
    .C(_00531_),
    .Y(_10988_));
 INVx1_ASAP7_75t_R _40150_ (.A(_10988_),
    .Y(_10989_));
 NOR3x2_ASAP7_75t_R _40151_ (.B(_10642_),
    .C(_10989_),
    .Y(_10990_),
    .A(_10987_));
 NAND3x2_ASAP7_75t_R _40152_ (.B(_00529_),
    .C(_00530_),
    .Y(_10991_),
    .A(_10990_));
 INVx4_ASAP7_75t_R _40153_ (.A(_10816_),
    .Y(_10992_));
 INVx1_ASAP7_75t_R _40154_ (.A(_10624_),
    .Y(_10993_));
 NAND2x1_ASAP7_75t_R _40155_ (.A(_10992_),
    .B(_10993_),
    .Y(_10995_));
 NOR2x2_ASAP7_75t_R _40156_ (.A(net1990),
    .B(_10627_),
    .Y(_10996_));
 INVx1_ASAP7_75t_R _40157_ (.A(_10747_),
    .Y(_10997_));
 OAI21x1_ASAP7_75t_R _40158_ (.A1(_10996_),
    .A2(_10997_),
    .B(_10992_),
    .Y(_10998_));
 NAND2x1_ASAP7_75t_R _40159_ (.A(_10995_),
    .B(_10998_),
    .Y(_10999_));
 OAI21x1_ASAP7_75t_R _40160_ (.A1(net1501),
    .A2(_10658_),
    .B(net1337),
    .Y(_11000_));
 INVx1_ASAP7_75t_R _40161_ (.A(_11000_),
    .Y(_11001_));
 TAPCELL_ASAP7_75t_R PHY_63 ();
 OAI21x1_ASAP7_75t_R _40163_ (.A1(_10733_),
    .A2(_11001_),
    .B(_10809_),
    .Y(_11003_));
 OAI21x1_ASAP7_75t_R _40164_ (.A1(_10671_),
    .A2(_10810_),
    .B(_11003_),
    .Y(_11004_));
 NOR2x2_ASAP7_75t_R _40165_ (.A(_10999_),
    .B(_11004_),
    .Y(_11006_));
 NAND2x2_ASAP7_75t_R _40166_ (.A(net2119),
    .B(_10791_),
    .Y(_11007_));
 NOR2x2_ASAP7_75t_R _40167_ (.A(net1993),
    .B(_10710_),
    .Y(_11008_));
 OAI21x1_ASAP7_75t_R _40168_ (.A1(net3068),
    .A2(_11008_),
    .B(_10791_),
    .Y(_11009_));
 OAI21x1_ASAP7_75t_R _40169_ (.A1(_10659_),
    .A2(_11007_),
    .B(_11009_),
    .Y(_11010_));
 OAI21x1_ASAP7_75t_R _40170_ (.A1(_10733_),
    .A2(_10869_),
    .B(_10791_),
    .Y(_11011_));
 INVx2_ASAP7_75t_R _40171_ (.A(_10628_),
    .Y(_11012_));
 OAI21x1_ASAP7_75t_R _40172_ (.A1(_10831_),
    .A2(_11012_),
    .B(_10791_),
    .Y(_11013_));
 NAND2x1_ASAP7_75t_R _40173_ (.A(_11011_),
    .B(_11013_),
    .Y(_11014_));
 NOR2x2_ASAP7_75t_R _40174_ (.A(_11010_),
    .B(_11014_),
    .Y(_11015_));
 AO21x1_ASAP7_75t_R _40175_ (.A1(net3065),
    .A2(_10678_),
    .B(_10796_),
    .Y(_11017_));
 AO21x1_ASAP7_75t_R _40176_ (.A1(net3049),
    .A2(_10645_),
    .B(_10796_),
    .Y(_11018_));
 AND2x2_ASAP7_75t_R _40177_ (.A(_11017_),
    .B(_11018_),
    .Y(_11019_));
 NAND3x2_ASAP7_75t_R _40178_ (.B(_11015_),
    .C(_11019_),
    .Y(_11020_),
    .A(_11006_));
 AOI211x1_ASAP7_75t_R _40179_ (.A1(_10626_),
    .A2(_10658_),
    .B(_10826_),
    .C(_10740_),
    .Y(_11021_));
 OA21x2_ASAP7_75t_R _40180_ (.A1(_10869_),
    .A2(_10733_),
    .B(_10827_),
    .Y(_11022_));
 AOI211x1_ASAP7_75t_R _40181_ (.A1(_10827_),
    .A2(_11008_),
    .B(_11021_),
    .C(_11022_),
    .Y(_11023_));
 OA21x2_ASAP7_75t_R _40182_ (.A1(_10792_),
    .A2(_11008_),
    .B(_10870_),
    .Y(_11024_));
 OA211x2_ASAP7_75t_R _40183_ (.A1(net3027),
    .A2(_10902_),
    .B(_10870_),
    .C(_10668_),
    .Y(_11025_));
 NOR2x1_ASAP7_75t_R _40184_ (.A(_11024_),
    .B(_11025_),
    .Y(_11026_));
 NAND2x2_ASAP7_75t_R _40185_ (.A(_11023_),
    .B(_11026_),
    .Y(_11028_));
 TAPCELL_ASAP7_75t_R PHY_62 ();
 AOI21x1_ASAP7_75t_R _40187_ (.A1(net3057),
    .A2(_10788_),
    .B(_10843_),
    .Y(_11030_));
 TAPCELL_ASAP7_75t_R PHY_61 ();
 AOI21x1_ASAP7_75t_R _40189_ (.A1(net1492),
    .A2(net1446),
    .B(_10843_),
    .Y(_11032_));
 AOI211x1_ASAP7_75t_R _40190_ (.A1(_10967_),
    .A2(_10847_),
    .B(_11030_),
    .C(_11032_),
    .Y(_11033_));
 TAPCELL_ASAP7_75t_R PHY_60 ();
 AOI21x1_ASAP7_75t_R _40192_ (.A1(net1475),
    .A2(_10783_),
    .B(_10851_),
    .Y(_11035_));
 NAND2x2_ASAP7_75t_R _40193_ (.A(_10658_),
    .B(net1340),
    .Y(_11036_));
 AOI21x1_ASAP7_75t_R _40194_ (.A1(_11036_),
    .A2(_10854_),
    .B(_10851_),
    .Y(_11037_));
 NAND2x2_ASAP7_75t_R _40195_ (.A(net1718),
    .B(net2118),
    .Y(_11039_));
 NOR2x2_ASAP7_75t_R _40196_ (.A(_10851_),
    .B(_11039_),
    .Y(_11040_));
 NOR3x2_ASAP7_75t_R _40197_ (.B(_11037_),
    .C(_11040_),
    .Y(_11041_),
    .A(_11035_));
 AO21x1_ASAP7_75t_R _40198_ (.A1(net3065),
    .A2(_10905_),
    .B(_10843_),
    .Y(_11042_));
 NOR2x2_ASAP7_75t_R _40199_ (.A(_10622_),
    .B(_10685_),
    .Y(_11043_));
 NAND2x1_ASAP7_75t_R _40200_ (.A(_11043_),
    .B(_10847_),
    .Y(_11044_));
 AND2x2_ASAP7_75t_R _40201_ (.A(_11042_),
    .B(_11044_),
    .Y(_11045_));
 NAND3x2_ASAP7_75t_R _40202_ (.B(_11041_),
    .C(_11045_),
    .Y(_11046_),
    .A(_11033_));
 NOR3x2_ASAP7_75t_R _40203_ (.B(_11028_),
    .C(_11046_),
    .Y(_11047_),
    .A(_11020_));
 NAND3x2_ASAP7_75t_R _40204_ (.B(_10991_),
    .C(_11047_),
    .Y(_11048_),
    .A(_10980_));
 XOR2x2_ASAP7_75t_R _40205_ (.A(_11048_),
    .B(_10878_),
    .Y(_11050_));
 AO21x1_ASAP7_75t_R _40206_ (.A1(_09738_),
    .A2(_09798_),
    .B(_09692_),
    .Y(_11051_));
 TAPCELL_ASAP7_75t_R PHY_59 ();
 AO21x1_ASAP7_75t_R _40208_ (.A1(_09658_),
    .A2(_09631_),
    .B(_09755_),
    .Y(_11053_));
 NAND2x1_ASAP7_75t_R _40209_ (.A(_09741_),
    .B(_09826_),
    .Y(_11054_));
 AND3x1_ASAP7_75t_R _40210_ (.A(_11051_),
    .B(_11053_),
    .C(_11054_),
    .Y(_11055_));
 INVx6_ASAP7_75t_R _40211_ (.A(_09692_),
    .Y(_11056_));
 NAND2x2_ASAP7_75t_R _40212_ (.A(net3177),
    .B(_11056_),
    .Y(_11057_));
 AO21x1_ASAP7_75t_R _40213_ (.A1(net2453),
    .A2(_09631_),
    .B(net2960),
    .Y(_11058_));
 NAND2x1_ASAP7_75t_R _40214_ (.A(_11058_),
    .B(_11057_),
    .Y(_11059_));
 TAPCELL_ASAP7_75t_R PHY_58 ();
 AO21x1_ASAP7_75t_R _40216_ (.A1(_09674_),
    .A2(net1476),
    .B(_09730_),
    .Y(_11062_));
 NAND2x1_ASAP7_75t_R _40217_ (.A(_09816_),
    .B(_09807_),
    .Y(_11063_));
 OAI21x1_ASAP7_75t_R _40218_ (.A1(_09589_),
    .A2(_11062_),
    .B(_11063_),
    .Y(_11064_));
 NOR2x1_ASAP7_75t_R _40219_ (.A(_11064_),
    .B(_11059_),
    .Y(_11065_));
 NAND2x1_ASAP7_75t_R _40220_ (.A(_11055_),
    .B(_11065_),
    .Y(_11066_));
 NAND2x2_ASAP7_75t_R _40221_ (.A(net2686),
    .B(_09661_),
    .Y(_11067_));
 OAI22x1_ASAP7_75t_R _40222_ (.A1(_11067_),
    .A2(net1281),
    .B1(net1102),
    .B2(net1743),
    .Y(_11068_));
 NOR2x2_ASAP7_75t_R _40223_ (.A(net2915),
    .B(_09674_),
    .Y(_11069_));
 OAI21x1_ASAP7_75t_R _40224_ (.A1(_11069_),
    .A2(net3177),
    .B(_09759_),
    .Y(_11070_));
 OR4x2_ASAP7_75t_R _40225_ (.A(_09674_),
    .B(net1844),
    .C(_09629_),
    .D(_09585_),
    .Y(_11072_));
 NAND2x1_ASAP7_75t_R _40226_ (.A(_11070_),
    .B(_11072_),
    .Y(_11073_));
 NOR2x1_ASAP7_75t_R _40227_ (.A(_11068_),
    .B(_11073_),
    .Y(_11074_));
 NOR2x2_ASAP7_75t_R _40228_ (.A(net1109),
    .B(net1476),
    .Y(_11075_));
 AO22x1_ASAP7_75t_R _40229_ (.A1(_09726_),
    .A2(_09816_),
    .B1(_09701_),
    .B2(_11075_),
    .Y(_11076_));
 OAI22x1_ASAP7_75t_R _40230_ (.A1(net2046),
    .A2(net1504),
    .B1(net1923),
    .B2(net2000),
    .Y(_11077_));
 NOR2x1_ASAP7_75t_R _40231_ (.A(_09644_),
    .B(net1502),
    .Y(_11078_));
 NOR3x1_ASAP7_75t_R _40232_ (.A(_11076_),
    .B(_11077_),
    .C(_11078_),
    .Y(_11079_));
 NAND2x1_ASAP7_75t_R _40233_ (.A(_11074_),
    .B(_11079_),
    .Y(_11080_));
 NOR2x1_ASAP7_75t_R _40234_ (.A(_11080_),
    .B(_11066_),
    .Y(_11081_));
 NAND2x1_ASAP7_75t_R _40235_ (.A(_09631_),
    .B(_09658_),
    .Y(_11083_));
 TAPCELL_ASAP7_75t_R PHY_57 ();
 TAPCELL_ASAP7_75t_R PHY_56 ();
 AOI211x1_ASAP7_75t_R _40238_ (.A1(_09854_),
    .A2(_09644_),
    .B(net2339),
    .C(_09573_),
    .Y(_11086_));
 AO21x2_ASAP7_75t_R _40239_ (.A1(_09714_),
    .A2(_09769_),
    .B(_09649_),
    .Y(_11087_));
 INVx1_ASAP7_75t_R _40240_ (.A(_11087_),
    .Y(_11088_));
 AOI211x1_ASAP7_75t_R _40241_ (.A1(_09696_),
    .A2(_11083_),
    .B(_11086_),
    .C(_11088_),
    .Y(_11089_));
 CKINVDCx10_ASAP7_75t_R _40242_ (.A(net2002),
    .Y(_11090_));
 NAND2x1_ASAP7_75t_R _40243_ (.A(_09608_),
    .B(_11090_),
    .Y(_11091_));
 TAPCELL_ASAP7_75t_R PHY_55 ();
 AO21x1_ASAP7_75t_R _40245_ (.A1(net2771),
    .A2(_09689_),
    .B(net2691),
    .Y(_11094_));
 OAI21x1_ASAP7_75t_R _40246_ (.A1(_09779_),
    .A2(_11091_),
    .B(_11094_),
    .Y(_11095_));
 INVx4_ASAP7_75t_R _40247_ (.A(_09854_),
    .Y(_11096_));
 NAND2x2_ASAP7_75t_R _40248_ (.A(_11096_),
    .B(_09757_),
    .Y(_11097_));
 OAI22x1_ASAP7_75t_R _40249_ (.A1(_11097_),
    .A2(_09573_),
    .B1(_09631_),
    .B2(net2942),
    .Y(_11098_));
 NOR2x1_ASAP7_75t_R _40250_ (.A(_11095_),
    .B(_11098_),
    .Y(_11099_));
 NAND2x1_ASAP7_75t_R _40251_ (.A(_11089_),
    .B(_11099_),
    .Y(_11100_));
 TAPCELL_ASAP7_75t_R PHY_54 ();
 NAND2x1_ASAP7_75t_R _40253_ (.A(net2771),
    .B(net1384),
    .Y(_11102_));
 NOR2x2_ASAP7_75t_R _40254_ (.A(_09642_),
    .B(_09655_),
    .Y(_11103_));
 AO21x1_ASAP7_75t_R _40255_ (.A1(_11102_),
    .A2(_09826_),
    .B(_11103_),
    .Y(_11105_));
 INVx1_ASAP7_75t_R _40256_ (.A(_09723_),
    .Y(_11106_));
 AO21x1_ASAP7_75t_R _40257_ (.A1(_09658_),
    .A2(_09631_),
    .B(net2002),
    .Y(_11107_));
 OAI21x1_ASAP7_75t_R _40258_ (.A1(_09589_),
    .A2(_11106_),
    .B(_11107_),
    .Y(_11108_));
 NOR2x1_ASAP7_75t_R _40259_ (.A(_11105_),
    .B(_11108_),
    .Y(_11109_));
 NAND2x1_ASAP7_75t_R _40260_ (.A(_09744_),
    .B(_09750_),
    .Y(_11110_));
 NOR2x2_ASAP7_75t_R _40261_ (.A(_09589_),
    .B(_09579_),
    .Y(_11111_));
 TAPCELL_ASAP7_75t_R PHY_53 ();
 AOI22x1_ASAP7_75t_R _40263_ (.A1(_11056_),
    .A2(_11111_),
    .B1(_11090_),
    .B2(_09832_),
    .Y(_11113_));
 NOR2x2_ASAP7_75t_R _40264_ (.A(_09597_),
    .B(_09730_),
    .Y(_11114_));
 AOI21x1_ASAP7_75t_R _40265_ (.A1(net2928),
    .A2(net2686),
    .B(_11114_),
    .Y(_11116_));
 NAND2x1_ASAP7_75t_R _40266_ (.A(_11116_),
    .B(_11113_),
    .Y(_11117_));
 NOR2x1_ASAP7_75t_R _40267_ (.A(_11117_),
    .B(_11110_),
    .Y(_11118_));
 NAND2x1_ASAP7_75t_R _40268_ (.A(_11109_),
    .B(_11118_),
    .Y(_11119_));
 NOR2x1_ASAP7_75t_R _40269_ (.A(_11100_),
    .B(_11119_),
    .Y(_11120_));
 NAND2x2_ASAP7_75t_R _40270_ (.A(_11081_),
    .B(_11120_),
    .Y(_11121_));
 NOR2x1_ASAP7_75t_R _40271_ (.A(net2104),
    .B(_09695_),
    .Y(_11122_));
 INVx2_ASAP7_75t_R _40272_ (.A(_11122_),
    .Y(_11123_));
 NAND2x2_ASAP7_75t_R _40273_ (.A(_09846_),
    .B(_11075_),
    .Y(_11124_));
 AO21x1_ASAP7_75t_R _40274_ (.A1(_11123_),
    .A2(_11124_),
    .B(_09573_),
    .Y(_11125_));
 OA21x2_ASAP7_75t_R _40275_ (.A1(_09832_),
    .A2(_09816_),
    .B(_09806_),
    .Y(_11127_));
 NOR2x2_ASAP7_75t_R _40276_ (.A(_09674_),
    .B(net2817),
    .Y(_11128_));
 NOR2x2_ASAP7_75t_R _40277_ (.A(_09717_),
    .B(_09672_),
    .Y(_11129_));
 AOI21x1_ASAP7_75t_R _40278_ (.A1(_09838_),
    .A2(_11128_),
    .B(_11129_),
    .Y(_11130_));
 INVx1_ASAP7_75t_R _40279_ (.A(_11130_),
    .Y(_11131_));
 NOR2x1_ASAP7_75t_R _40280_ (.A(_11127_),
    .B(_11131_),
    .Y(_11132_));
 NAND2x1_ASAP7_75t_R _40281_ (.A(_11125_),
    .B(_11132_),
    .Y(_11133_));
 NOR2x2_ASAP7_75t_R _40282_ (.A(_09674_),
    .B(_09779_),
    .Y(_11134_));
 OA21x2_ASAP7_75t_R _40283_ (.A1(_11134_),
    .A2(_09809_),
    .B(_09806_),
    .Y(_11135_));
 NAND2x1_ASAP7_75t_R _40284_ (.A(net2152),
    .B(_09757_),
    .Y(_11136_));
 NAND2x1_ASAP7_75t_R _40285_ (.A(net2919),
    .B(_09807_),
    .Y(_11138_));
 OAI21x1_ASAP7_75t_R _40286_ (.A1(_09589_),
    .A2(_11136_),
    .B(_11138_),
    .Y(_11139_));
 NOR2x1_ASAP7_75t_R _40287_ (.A(_11135_),
    .B(_11139_),
    .Y(_11140_));
 AO21x2_ASAP7_75t_R _40288_ (.A1(_09642_),
    .A2(_09653_),
    .B(net2339),
    .Y(_11141_));
 INVx1_ASAP7_75t_R _40289_ (.A(_11141_),
    .Y(_11142_));
 AO21x1_ASAP7_75t_R _40290_ (.A1(_09592_),
    .A2(net2216),
    .B(_09620_),
    .Y(_11143_));
 AO21x2_ASAP7_75t_R _40291_ (.A1(_09611_),
    .A2(_09613_),
    .B(_09672_),
    .Y(_11144_));
 NAND2x1_ASAP7_75t_R _40292_ (.A(_11143_),
    .B(_11144_),
    .Y(_11145_));
 NOR2x1_ASAP7_75t_R _40293_ (.A(_11145_),
    .B(_11142_),
    .Y(_11146_));
 NAND2x2_ASAP7_75t_R _40294_ (.A(_11140_),
    .B(_11146_),
    .Y(_11147_));
 NOR2x2_ASAP7_75t_R _40295_ (.A(_11133_),
    .B(_11147_),
    .Y(_11149_));
 OAI22x1_ASAP7_75t_R _40296_ (.A1(net1518),
    .A2(_09682_),
    .B1(net2917),
    .B2(_09597_),
    .Y(_11150_));
 NAND2x2_ASAP7_75t_R _40297_ (.A(net2687),
    .B(_09640_),
    .Y(_11151_));
 OAI21x1_ASAP7_75t_R _40298_ (.A1(_09854_),
    .A2(net2000),
    .B(_11151_),
    .Y(_11152_));
 NOR2x1_ASAP7_75t_R _40299_ (.A(_11150_),
    .B(_11152_),
    .Y(_11153_));
 OAI22x1_ASAP7_75t_R _40300_ (.A1(net1925),
    .A2(_09682_),
    .B1(net2453),
    .B2(net2547),
    .Y(_11154_));
 OAI21x1_ASAP7_75t_R _40301_ (.A1(net2732),
    .A2(net2339),
    .B(_09666_),
    .Y(_11155_));
 NOR2x1_ASAP7_75t_R _40302_ (.A(_11154_),
    .B(_11155_),
    .Y(_11156_));
 NAND2x1_ASAP7_75t_R _40303_ (.A(_11153_),
    .B(_11156_),
    .Y(_11157_));
 OA21x2_ASAP7_75t_R _40304_ (.A1(_09661_),
    .A2(_09726_),
    .B(_11069_),
    .Y(_11158_));
 NAND2x1_ASAP7_75t_R _40305_ (.A(_09662_),
    .B(_09591_),
    .Y(_11160_));
 NAND2x2_ASAP7_75t_R _40306_ (.A(_09591_),
    .B(_09710_),
    .Y(_11161_));
 TAPCELL_ASAP7_75t_R PHY_52 ();
 OAI22x1_ASAP7_75t_R _40308_ (.A1(_09682_),
    .A2(_11160_),
    .B1(_11161_),
    .B2(net1942),
    .Y(_11163_));
 NOR2x1_ASAP7_75t_R _40309_ (.A(_11158_),
    .B(_11163_),
    .Y(_11164_));
 NAND2x2_ASAP7_75t_R _40310_ (.A(net1286),
    .B(net1934),
    .Y(_11165_));
 OAI22x1_ASAP7_75t_R _40311_ (.A1(_11161_),
    .A2(net2914),
    .B1(_09672_),
    .B2(_11165_),
    .Y(_11166_));
 NOR2x2_ASAP7_75t_R _40312_ (.A(_09581_),
    .B(_09674_),
    .Y(_11167_));
 NOR2x2_ASAP7_75t_R _40313_ (.A(_09837_),
    .B(_09639_),
    .Y(_11168_));
 AO22x1_ASAP7_75t_R _40314_ (.A1(_09838_),
    .A2(_11167_),
    .B1(_11168_),
    .B2(_09761_),
    .Y(_11169_));
 NOR2x1_ASAP7_75t_R _40315_ (.A(_11166_),
    .B(_11169_),
    .Y(_11171_));
 NAND2x1_ASAP7_75t_R _40316_ (.A(_11164_),
    .B(_11171_),
    .Y(_11172_));
 NOR2x2_ASAP7_75t_R _40317_ (.A(_11157_),
    .B(_11172_),
    .Y(_11173_));
 NOR2x1_ASAP7_75t_R _40318_ (.A(_09613_),
    .B(_09707_),
    .Y(_11174_));
 NOR2x1_ASAP7_75t_R _40319_ (.A(net2103),
    .B(_09620_),
    .Y(_11175_));
 OR3x2_ASAP7_75t_R _40320_ (.A(_09595_),
    .B(_11174_),
    .C(_11175_),
    .Y(_11176_));
 NAND2x2_ASAP7_75t_R _40321_ (.A(net1285),
    .B(net2151),
    .Y(_11177_));
 NOR2x2_ASAP7_75t_R _40322_ (.A(_11177_),
    .B(_09655_),
    .Y(_11178_));
 INVx3_ASAP7_75t_R _40323_ (.A(_11178_),
    .Y(_11179_));
 NOR2x2_ASAP7_75t_R _40324_ (.A(net1480),
    .B(_09662_),
    .Y(_11180_));
 AND2x2_ASAP7_75t_R _40325_ (.A(net1100),
    .B(_09581_),
    .Y(_11182_));
 OAI21x1_ASAP7_75t_R _40326_ (.A1(_11180_),
    .A2(_11182_),
    .B(_09826_),
    .Y(_11183_));
 NAND3x2_ASAP7_75t_R _40327_ (.B(_11179_),
    .C(_11183_),
    .Y(_11184_),
    .A(_09656_));
 NAND2x2_ASAP7_75t_R _40328_ (.A(_11180_),
    .B(_11090_),
    .Y(_11185_));
 NAND2x2_ASAP7_75t_R _40329_ (.A(_09661_),
    .B(_09700_),
    .Y(_11186_));
 NAND2x2_ASAP7_75t_R _40330_ (.A(_09846_),
    .B(net2918),
    .Y(_11187_));
 NAND3x2_ASAP7_75t_R _40331_ (.B(_11186_),
    .C(_11187_),
    .Y(_11188_),
    .A(_11185_));
 NOR3x2_ASAP7_75t_R _40332_ (.B(_11184_),
    .C(_11188_),
    .Y(_11189_),
    .A(_11176_));
 NAND3x2_ASAP7_75t_R _40333_ (.B(_11173_),
    .C(_11189_),
    .Y(_11190_),
    .A(_11149_));
 NOR2x2_ASAP7_75t_R _40334_ (.A(_11121_),
    .B(_11190_),
    .Y(_11191_));
 NAND2x2_ASAP7_75t_R _40335_ (.A(_09628_),
    .B(_11191_),
    .Y(_11193_));
 TAPCELL_ASAP7_75t_R PHY_51 ();
 AO21x1_ASAP7_75t_R _40337_ (.A1(_10111_),
    .A2(net1661),
    .B(_09990_),
    .Y(_11195_));
 NOR2x1_ASAP7_75t_R _40338_ (.A(_09934_),
    .B(_09990_),
    .Y(_11196_));
 OAI21x1_ASAP7_75t_R _40339_ (.A1(net1020),
    .A2(net1163),
    .B(_11196_),
    .Y(_11197_));
 NAND2x1_ASAP7_75t_R _40340_ (.A(_11195_),
    .B(_11197_),
    .Y(_11198_));
 OAI21x1_ASAP7_75t_R _40341_ (.A1(_09988_),
    .A2(_09990_),
    .B(_10223_),
    .Y(_11199_));
 NOR2x2_ASAP7_75t_R _40342_ (.A(net976),
    .B(net1704),
    .Y(_11200_));
 NAND2x2_ASAP7_75t_R _40343_ (.A(_11200_),
    .B(_09974_),
    .Y(_11201_));
 AO21x1_ASAP7_75t_R _40344_ (.A1(_10107_),
    .A2(_10153_),
    .B(_10246_),
    .Y(_11202_));
 NAND2x1_ASAP7_75t_R _40345_ (.A(_11201_),
    .B(_11202_),
    .Y(_11204_));
 NOR3x1_ASAP7_75t_R _40346_ (.A(_11198_),
    .B(_11199_),
    .C(_11204_),
    .Y(_11205_));
 TAPCELL_ASAP7_75t_R PHY_50 ();
 TAPCELL_ASAP7_75t_R PHY_49 ();
 AO21x1_ASAP7_75t_R _40349_ (.A1(_09913_),
    .A2(_10008_),
    .B(_10011_),
    .Y(_11208_));
 AO21x1_ASAP7_75t_R _40350_ (.A1(net2958),
    .A2(_10042_),
    .B(_10011_),
    .Y(_11209_));
 NAND2x1_ASAP7_75t_R _40351_ (.A(_10014_),
    .B(_10255_),
    .Y(_11210_));
 NAND3x1_ASAP7_75t_R _40352_ (.A(_11208_),
    .B(_11209_),
    .C(_11210_),
    .Y(_11211_));
 NOR2x2_ASAP7_75t_R _40353_ (.A(_09969_),
    .B(net1703),
    .Y(_11212_));
 OAI21x1_ASAP7_75t_R _40354_ (.A1(_10126_),
    .A2(_11212_),
    .B(net1892),
    .Y(_11213_));
 NAND2x1_ASAP7_75t_R _40355_ (.A(net1891),
    .B(net2222),
    .Y(_11215_));
 NAND3x1_ASAP7_75t_R _40356_ (.A(_11213_),
    .B(_10275_),
    .C(_11215_),
    .Y(_11216_));
 AO21x1_ASAP7_75t_R _40357_ (.A1(_09934_),
    .A2(_10042_),
    .B(_10005_),
    .Y(_11217_));
 INVx1_ASAP7_75t_R _40358_ (.A(_11217_),
    .Y(_11218_));
 NOR3x1_ASAP7_75t_R _40359_ (.A(_11211_),
    .B(_11216_),
    .C(_11218_),
    .Y(_11219_));
 NAND2x1_ASAP7_75t_R _40360_ (.A(_11205_),
    .B(_11219_),
    .Y(_11220_));
 NOR2x1_ASAP7_75t_R _40361_ (.A(_09892_),
    .B(net1798),
    .Y(_11221_));
 NAND2x2_ASAP7_75t_R _40362_ (.A(_11221_),
    .B(_10133_),
    .Y(_11222_));
 NAND2x2_ASAP7_75t_R _40363_ (.A(_11222_),
    .B(_10213_),
    .Y(_11223_));
 NAND2x2_ASAP7_75t_R _40364_ (.A(_11200_),
    .B(_10133_),
    .Y(_11224_));
 AO21x1_ASAP7_75t_R _40365_ (.A1(_09906_),
    .A2(net2444),
    .B(net2660),
    .Y(_11226_));
 NAND2x2_ASAP7_75t_R _40366_ (.A(_11224_),
    .B(_11226_),
    .Y(_11227_));
 NAND2x2_ASAP7_75t_R _40367_ (.A(_10133_),
    .B(_10161_),
    .Y(_11228_));
 NAND2x2_ASAP7_75t_R _40368_ (.A(_11228_),
    .B(_10218_),
    .Y(_11229_));
 NOR3x2_ASAP7_75t_R _40369_ (.B(_11227_),
    .C(_11229_),
    .Y(_11230_),
    .A(_11223_));
 NAND3x2_ASAP7_75t_R _40370_ (.B(net1067),
    .C(_09905_),
    .Y(_11231_),
    .A(net2382));
 OAI21x1_ASAP7_75t_R _40371_ (.A1(_09982_),
    .A2(_10161_),
    .B(net2382),
    .Y(_11232_));
 NAND3x2_ASAP7_75t_R _40372_ (.B(_10129_),
    .C(_11232_),
    .Y(_11233_),
    .A(_11231_));
 NAND3x2_ASAP7_75t_R _40373_ (.B(net1067),
    .C(net1252),
    .Y(_11234_),
    .A(net1952));
 OAI21x1_ASAP7_75t_R _40374_ (.A1(_09961_),
    .A2(_10126_),
    .B(net1953),
    .Y(_11235_));
 OAI21x1_ASAP7_75t_R _40375_ (.A1(_09981_),
    .A2(_09946_),
    .B(net1951),
    .Y(_11237_));
 NAND3x2_ASAP7_75t_R _40376_ (.B(_11235_),
    .C(_11237_),
    .Y(_11238_),
    .A(_11234_));
 NOR2x2_ASAP7_75t_R _40377_ (.A(_11233_),
    .B(_11238_),
    .Y(_11239_));
 AOI211x1_ASAP7_75t_R _40378_ (.A1(net3015),
    .A2(_09892_),
    .B(_09901_),
    .C(net1798),
    .Y(_11240_));
 INVx1_ASAP7_75t_R _40379_ (.A(_11240_),
    .Y(_11241_));
 AO21x1_ASAP7_75t_R _40380_ (.A1(net2397),
    .A2(_09882_),
    .B(_09901_),
    .Y(_11242_));
 AO21x1_ASAP7_75t_R _40381_ (.A1(_10107_),
    .A2(net1757),
    .B(_09901_),
    .Y(_11243_));
 AND3x1_ASAP7_75t_R _40382_ (.A(_11241_),
    .B(_11242_),
    .C(_11243_),
    .Y(_11244_));
 NAND3x2_ASAP7_75t_R _40383_ (.B(_11239_),
    .C(_11244_),
    .Y(_11245_),
    .A(_11230_));
 NOR2x2_ASAP7_75t_R _40384_ (.A(_11220_),
    .B(_11245_),
    .Y(_11246_));
 AO21x1_ASAP7_75t_R _40385_ (.A1(_09906_),
    .A2(_10153_),
    .B(_10035_),
    .Y(_11248_));
 NAND2x1_ASAP7_75t_R _40386_ (.A(_10030_),
    .B(_11212_),
    .Y(_11249_));
 NOR2x1_ASAP7_75t_R _40387_ (.A(net1798),
    .B(net2591),
    .Y(_11250_));
 NAND2x1_ASAP7_75t_R _40388_ (.A(_10030_),
    .B(_11250_),
    .Y(_11251_));
 NAND3x1_ASAP7_75t_R _40389_ (.A(_11248_),
    .B(_11249_),
    .C(_11251_),
    .Y(_11252_));
 NAND2x1_ASAP7_75t_R _40390_ (.A(net1163),
    .B(_09905_),
    .Y(_11253_));
 TAPCELL_ASAP7_75t_R PHY_48 ();
 AO21x1_ASAP7_75t_R _40392_ (.A1(_09913_),
    .A2(_11253_),
    .B(net2662),
    .Y(_11255_));
 AO21x1_ASAP7_75t_R _40393_ (.A1(net942),
    .A2(net1661),
    .B(net2662),
    .Y(_11256_));
 AO21x1_ASAP7_75t_R _40394_ (.A1(_09998_),
    .A2(_09928_),
    .B(net2662),
    .Y(_11257_));
 NAND3x1_ASAP7_75t_R _40395_ (.A(_11255_),
    .B(_11256_),
    .C(_11257_),
    .Y(_11259_));
 NOR2x1_ASAP7_75t_R _40396_ (.A(_11252_),
    .B(_11259_),
    .Y(_11260_));
 NAND2x2_ASAP7_75t_R _40397_ (.A(net2805),
    .B(_09946_),
    .Y(_11261_));
 NAND3x1_ASAP7_75t_R _40398_ (.A(_10211_),
    .B(_10168_),
    .C(_11261_),
    .Y(_11262_));
 AO21x1_ASAP7_75t_R _40399_ (.A1(_10111_),
    .A2(_09934_),
    .B(_10048_),
    .Y(_11263_));
 AO21x1_ASAP7_75t_R _40400_ (.A1(net2160),
    .A2(_10038_),
    .B(_10048_),
    .Y(_11264_));
 NAND2x1_ASAP7_75t_R _40401_ (.A(_11263_),
    .B(_11264_),
    .Y(_11265_));
 OAI21x1_ASAP7_75t_R _40402_ (.A1(net2591),
    .A2(_10240_),
    .B(_10176_),
    .Y(_11266_));
 NOR3x1_ASAP7_75t_R _40403_ (.A(_11262_),
    .B(_11265_),
    .C(_11266_),
    .Y(_11267_));
 NAND2x1_ASAP7_75t_R _40404_ (.A(_11260_),
    .B(_11267_),
    .Y(_11268_));
 TAPCELL_ASAP7_75t_R PHY_47 ();
 AO21x1_ASAP7_75t_R _40406_ (.A1(_09913_),
    .A2(_10038_),
    .B(net2253),
    .Y(_11271_));
 AO21x1_ASAP7_75t_R _40407_ (.A1(net2235),
    .A2(_09882_),
    .B(net2253),
    .Y(_11272_));
 NAND2x1_ASAP7_75t_R _40408_ (.A(_10071_),
    .B(_10143_),
    .Y(_11273_));
 NAND3x1_ASAP7_75t_R _40409_ (.A(_11271_),
    .B(_11272_),
    .C(_11273_),
    .Y(_11274_));
 TAPCELL_ASAP7_75t_R PHY_46 ();
 AO21x1_ASAP7_75t_R _40411_ (.A1(net2214),
    .A2(_10111_),
    .B(net2353),
    .Y(_11276_));
 NAND2x1_ASAP7_75t_R _40412_ (.A(net2222),
    .B(_10140_),
    .Y(_11277_));
 NAND3x1_ASAP7_75t_R _40413_ (.A(_11276_),
    .B(_10091_),
    .C(_11277_),
    .Y(_11278_));
 NOR2x1_ASAP7_75t_R _40414_ (.A(_11274_),
    .B(_11278_),
    .Y(_11279_));
 AO31x2_ASAP7_75t_R _40415_ (.A1(_09882_),
    .A2(net2214),
    .A3(net2397),
    .B(net2535),
    .Y(_11281_));
 NOR2x2_ASAP7_75t_R _40416_ (.A(net2351),
    .B(_09963_),
    .Y(_11282_));
 OA21x2_ASAP7_75t_R _40417_ (.A1(_09978_),
    .A2(_11212_),
    .B(_10099_),
    .Y(_11283_));
 NOR2x1_ASAP7_75t_R _40418_ (.A(_11282_),
    .B(_11283_),
    .Y(_11284_));
 NAND2x1_ASAP7_75t_R _40419_ (.A(_11281_),
    .B(_11284_),
    .Y(_11285_));
 NOR2x1_ASAP7_75t_R _40420_ (.A(net2408),
    .B(net2925),
    .Y(_11286_));
 AOI211x1_ASAP7_75t_R _40421_ (.A1(_10114_),
    .A2(_10113_),
    .B(_11286_),
    .C(_10180_),
    .Y(_11287_));
 AO21x1_ASAP7_75t_R _40422_ (.A1(_10107_),
    .A2(net2445),
    .B(net2628),
    .Y(_11288_));
 AO21x1_ASAP7_75t_R _40423_ (.A1(net2358),
    .A2(net1756),
    .B(net2628),
    .Y(_11289_));
 AND2x2_ASAP7_75t_R _40424_ (.A(_11288_),
    .B(_11289_),
    .Y(_11290_));
 NAND2x1_ASAP7_75t_R _40425_ (.A(_11290_),
    .B(_11287_),
    .Y(_11292_));
 NOR2x1_ASAP7_75t_R _40426_ (.A(_11285_),
    .B(_11292_),
    .Y(_11293_));
 NAND2x2_ASAP7_75t_R _40427_ (.A(_11279_),
    .B(_11293_),
    .Y(_11294_));
 NOR2x2_ASAP7_75t_R _40428_ (.A(_11268_),
    .B(_11294_),
    .Y(_11295_));
 NAND3x2_ASAP7_75t_R _40429_ (.B(_10300_),
    .C(_11295_),
    .Y(_11296_),
    .A(_11246_));
 XOR2x2_ASAP7_75t_R _40430_ (.A(_11193_),
    .B(_11296_),
    .Y(_11297_));
 NOR2x2_ASAP7_75t_R _40431_ (.A(_11050_),
    .B(_11297_),
    .Y(_11298_));
 TAPCELL_ASAP7_75t_R PHY_45 ();
 XOR2x2_ASAP7_75t_R _40433_ (.A(_11048_),
    .B(net2514),
    .Y(_11300_));
 INVx1_ASAP7_75t_R _40434_ (.A(_11296_),
    .Y(_11301_));
 XOR2x1_ASAP7_75t_R _40435_ (.A(_11301_),
    .Y(_11303_),
    .B(_11193_));
 NOR2x1_ASAP7_75t_R _40436_ (.A(_11300_),
    .B(_11303_),
    .Y(_11304_));
 TAPCELL_ASAP7_75t_R PHY_44 ();
 NAND2x2_ASAP7_75t_R _40438_ (.A(net1378),
    .B(net1497),
    .Y(_11306_));
 AO21x1_ASAP7_75t_R _40439_ (.A1(net1115),
    .A2(_11306_),
    .B(net2227),
    .Y(_11307_));
 AO21x1_ASAP7_75t_R _40440_ (.A1(net1090),
    .A2(net1051),
    .B(net2227),
    .Y(_11308_));
 NAND2x1_ASAP7_75t_R _40441_ (.A(_10545_),
    .B(_10589_),
    .Y(_11309_));
 NAND3x1_ASAP7_75t_R _40442_ (.A(_11307_),
    .B(_11308_),
    .C(_11309_),
    .Y(_11310_));
 TAPCELL_ASAP7_75t_R PHY_43 ();
 NAND2x2_ASAP7_75t_R _40444_ (.A(net3084),
    .B(net1740),
    .Y(_11312_));
 AO21x1_ASAP7_75t_R _40445_ (.A1(net2841),
    .A2(_11312_),
    .B(net2180),
    .Y(_11314_));
 TAPCELL_ASAP7_75t_R PHY_42 ();
 AO21x1_ASAP7_75t_R _40447_ (.A1(net1143),
    .A2(net1051),
    .B(net2180),
    .Y(_11316_));
 NOR2x2_ASAP7_75t_R _40448_ (.A(_10384_),
    .B(net2188),
    .Y(_11317_));
 NAND2x1_ASAP7_75t_R _40449_ (.A(_11317_),
    .B(_10601_),
    .Y(_11318_));
 NAND3x1_ASAP7_75t_R _40450_ (.A(_11314_),
    .B(_11316_),
    .C(_11318_),
    .Y(_11319_));
 NOR2x1_ASAP7_75t_R _40451_ (.A(_11310_),
    .B(_11319_),
    .Y(_11320_));
 AOI21x1_ASAP7_75t_R _40452_ (.A1(net1306),
    .A2(net1414),
    .B(_10567_),
    .Y(_11321_));
 TAPCELL_ASAP7_75t_R PHY_41 ();
 INVx8_ASAP7_75t_R _40454_ (.A(_10554_),
    .Y(_11323_));
 TAPCELL_ASAP7_75t_R PHY_40 ();
 AOI21x1_ASAP7_75t_R _40456_ (.A1(net1856),
    .A2(_11323_),
    .B(_10567_),
    .Y(_11325_));
 NOR2x1_ASAP7_75t_R _40457_ (.A(_11321_),
    .B(_11325_),
    .Y(_11326_));
 AO31x2_ASAP7_75t_R _40458_ (.A1(net1144),
    .A2(_10410_),
    .A3(net3161),
    .B(_10567_),
    .Y(_11327_));
 NAND2x1_ASAP7_75t_R _40459_ (.A(_11326_),
    .B(_11327_),
    .Y(_11328_));
 AO31x2_ASAP7_75t_R _40460_ (.A1(net1144),
    .A2(net1052),
    .A3(net1659),
    .B(net2313),
    .Y(_11329_));
 AOI21x1_ASAP7_75t_R _40461_ (.A1(net3335),
    .A2(net2463),
    .B(net2313),
    .Y(_11330_));
 AOI211x1_ASAP7_75t_R _40462_ (.A1(net975),
    .A2(net1586),
    .B(_10578_),
    .C(net3013),
    .Y(_11331_));
 NOR2x1_ASAP7_75t_R _40463_ (.A(_11330_),
    .B(_11331_),
    .Y(_11332_));
 NAND2x1_ASAP7_75t_R _40464_ (.A(_11332_),
    .B(_11329_),
    .Y(_11333_));
 NOR2x1_ASAP7_75t_R _40465_ (.A(_11328_),
    .B(_11333_),
    .Y(_11335_));
 NAND2x1_ASAP7_75t_R _40466_ (.A(_11335_),
    .B(_11320_),
    .Y(_11336_));
 NAND2x1_ASAP7_75t_R _40467_ (.A(_10481_),
    .B(_10547_),
    .Y(_11337_));
 NOR2x2_ASAP7_75t_R _40468_ (.A(_10384_),
    .B(_10312_),
    .Y(_11338_));
 OAI21x1_ASAP7_75t_R _40469_ (.A1(net1264),
    .A2(_11338_),
    .B(_10547_),
    .Y(_11339_));
 NAND2x1_ASAP7_75t_R _40470_ (.A(_11337_),
    .B(_11339_),
    .Y(_11340_));
 NOR2x2_ASAP7_75t_R _40471_ (.A(_10367_),
    .B(_10312_),
    .Y(_11341_));
 OAI21x1_ASAP7_75t_R _40472_ (.A1(net1272),
    .A2(_11341_),
    .B(_10537_),
    .Y(_11342_));
 OAI21x1_ASAP7_75t_R _40473_ (.A1(_10385_),
    .A2(_10597_),
    .B(_10537_),
    .Y(_11343_));
 NAND2x1_ASAP7_75t_R _40474_ (.A(_11342_),
    .B(_11343_),
    .Y(_11344_));
 TAPCELL_ASAP7_75t_R PHY_39 ();
 AOI21x1_ASAP7_75t_R _40476_ (.A1(net2695),
    .A2(_10518_),
    .B(net3043),
    .Y(_11347_));
 NOR3x1_ASAP7_75t_R _40477_ (.A(_11340_),
    .B(_11344_),
    .C(_11347_),
    .Y(_11348_));
 INVx2_ASAP7_75t_R _40478_ (.A(_10396_),
    .Y(_11349_));
 INVx3_ASAP7_75t_R _40479_ (.A(_10515_),
    .Y(_11350_));
 OA21x2_ASAP7_75t_R _40480_ (.A1(net3034),
    .A2(_11349_),
    .B(_11350_),
    .Y(_11351_));
 OA21x2_ASAP7_75t_R _40481_ (.A1(net1265),
    .A2(_10545_),
    .B(_11350_),
    .Y(_11352_));
 OA21x2_ASAP7_75t_R _40482_ (.A1(_11317_),
    .A2(_10520_),
    .B(_11350_),
    .Y(_11353_));
 NOR3x1_ASAP7_75t_R _40483_ (.A(_11351_),
    .B(_11352_),
    .C(_11353_),
    .Y(_11354_));
 NAND2x2_ASAP7_75t_R _40484_ (.A(_10414_),
    .B(_10514_),
    .Y(_11355_));
 TAPCELL_ASAP7_75t_R PHY_38 ();
 AOI211x1_ASAP7_75t_R _40486_ (.A1(net975),
    .A2(net1318),
    .B(_11355_),
    .C(net970),
    .Y(_11358_));
 NOR2x1_ASAP7_75t_R _40487_ (.A(_10459_),
    .B(_11355_),
    .Y(_11359_));
 AOI211x1_ASAP7_75t_R _40488_ (.A1(_10576_),
    .A2(_10528_),
    .B(_11358_),
    .C(_11359_),
    .Y(_11360_));
 NAND3x1_ASAP7_75t_R _40489_ (.A(_11348_),
    .B(_11354_),
    .C(_11360_),
    .Y(_11361_));
 NOR2x1_ASAP7_75t_R _40490_ (.A(_11336_),
    .B(_11361_),
    .Y(_11362_));
 AO21x1_ASAP7_75t_R _40491_ (.A1(net1115),
    .A2(_10502_),
    .B(_10358_),
    .Y(_11363_));
 NAND2x2_ASAP7_75t_R _40492_ (.A(_10367_),
    .B(_10328_),
    .Y(_11364_));
 TAPCELL_ASAP7_75t_R PHY_37 ();
 AO21x1_ASAP7_75t_R _40494_ (.A1(_11364_),
    .A2(net1090),
    .B(_10358_),
    .Y(_11366_));
 NOR2x2_ASAP7_75t_R _40495_ (.A(_10322_),
    .B(_10536_),
    .Y(_11368_));
 OAI21x1_ASAP7_75t_R _40496_ (.A1(_10554_),
    .A2(_10350_),
    .B(_11368_),
    .Y(_11369_));
 NAND3x1_ASAP7_75t_R _40497_ (.A(_11363_),
    .B(_11366_),
    .C(_11369_),
    .Y(_11370_));
 OA21x2_ASAP7_75t_R _40498_ (.A1(_10545_),
    .A2(_11338_),
    .B(_10323_),
    .Y(_11371_));
 NOR2x1_ASAP7_75t_R _40499_ (.A(_10342_),
    .B(_11371_),
    .Y(_11372_));
 NOR2x1_ASAP7_75t_R _40500_ (.A(_10332_),
    .B(_10345_),
    .Y(_11373_));
 NOR2x1_ASAP7_75t_R _40501_ (.A(_11373_),
    .B(_10387_),
    .Y(_11374_));
 NAND2x1_ASAP7_75t_R _40502_ (.A(_11372_),
    .B(_11374_),
    .Y(_11375_));
 NOR2x1_ASAP7_75t_R _40503_ (.A(_11370_),
    .B(_11375_),
    .Y(_11376_));
 AO21x1_ASAP7_75t_R _40504_ (.A1(net2695),
    .A2(net1125),
    .B(net2536),
    .Y(_11377_));
 NAND2x2_ASAP7_75t_R _40505_ (.A(net1500),
    .B(_10382_),
    .Y(_11379_));
 OR2x6_ASAP7_75t_R _40506_ (.A(net2329),
    .B(_11379_),
    .Y(_11380_));
 NAND2x1_ASAP7_75t_R _40507_ (.A(_10554_),
    .B(_10406_),
    .Y(_11381_));
 NAND3x1_ASAP7_75t_R _40508_ (.A(_11377_),
    .B(_11380_),
    .C(_11381_),
    .Y(_11382_));
 NAND2x1_ASAP7_75t_R _40509_ (.A(_10316_),
    .B(net1885),
    .Y(_11383_));
 NOR2x1_ASAP7_75t_R _40510_ (.A(_11383_),
    .B(net2448),
    .Y(_11384_));
 NOR2x1_ASAP7_75t_R _40511_ (.A(_11384_),
    .B(_10437_),
    .Y(_11385_));
 AOI211x1_ASAP7_75t_R _40512_ (.A1(_10367_),
    .A2(net1582),
    .B(net1510),
    .C(net1881),
    .Y(_11386_));
 AOI211x1_ASAP7_75t_R _40513_ (.A1(_10367_),
    .A2(net3338),
    .B(net1881),
    .C(_10341_),
    .Y(_11387_));
 NOR2x1_ASAP7_75t_R _40514_ (.A(_11386_),
    .B(_11387_),
    .Y(_11388_));
 NAND2x1_ASAP7_75t_R _40515_ (.A(_11385_),
    .B(_11388_),
    .Y(_11390_));
 NOR2x1_ASAP7_75t_R _40516_ (.A(_11382_),
    .B(_11390_),
    .Y(_11391_));
 NAND2x1_ASAP7_75t_R _40517_ (.A(_11376_),
    .B(_11391_),
    .Y(_11392_));
 NAND3x2_ASAP7_75t_R _40518_ (.B(net959),
    .C(net2951),
    .Y(_11393_),
    .A(_10462_));
 AO21x1_ASAP7_75t_R _40519_ (.A1(net2952),
    .A2(net2442),
    .B(_10454_),
    .Y(_11394_));
 AO21x1_ASAP7_75t_R _40520_ (.A1(net1115),
    .A2(_10502_),
    .B(_10454_),
    .Y(_11395_));
 NAND3x1_ASAP7_75t_R _40521_ (.A(_11393_),
    .B(_11394_),
    .C(_11395_),
    .Y(_11396_));
 INVx3_ASAP7_75t_R _40522_ (.A(_10468_),
    .Y(_11397_));
 AOI21x1_ASAP7_75t_R _40523_ (.A1(net2354),
    .A2(_10449_),
    .B(_10468_),
    .Y(_11398_));
 AOI21x1_ASAP7_75t_R _40524_ (.A1(_11397_),
    .A2(_10531_),
    .B(_11398_),
    .Y(_11399_));
 AOI21x1_ASAP7_75t_R _40525_ (.A1(_10485_),
    .A2(net1659),
    .B(net2233),
    .Y(_11401_));
 AOI211x1_ASAP7_75t_R _40526_ (.A1(net975),
    .A2(net1586),
    .B(_10468_),
    .C(_10341_),
    .Y(_11402_));
 NOR2x1_ASAP7_75t_R _40527_ (.A(_11401_),
    .B(_11402_),
    .Y(_11403_));
 NAND2x1_ASAP7_75t_R _40528_ (.A(_11399_),
    .B(_11403_),
    .Y(_11404_));
 NOR2x1_ASAP7_75t_R _40529_ (.A(_11396_),
    .B(_11404_),
    .Y(_11405_));
 TAPCELL_ASAP7_75t_R PHY_36 ();
 AO21x1_ASAP7_75t_R _40531_ (.A1(_11323_),
    .A2(net1306),
    .B(net2069),
    .Y(_11407_));
 AO21x1_ASAP7_75t_R _40532_ (.A1(net2841),
    .A2(_11312_),
    .B(net2069),
    .Y(_11408_));
 AO21x1_ASAP7_75t_R _40533_ (.A1(net1143),
    .A2(net1053),
    .B(net2069),
    .Y(_11409_));
 NAND3x1_ASAP7_75t_R _40534_ (.A(_11407_),
    .B(_11408_),
    .C(_11409_),
    .Y(_11410_));
 NOR2x1_ASAP7_75t_R _40535_ (.A(net2247),
    .B(_11379_),
    .Y(_11412_));
 INVx3_ASAP7_75t_R _40536_ (.A(_10498_),
    .Y(_11413_));
 OA21x2_ASAP7_75t_R _40537_ (.A1(net2806),
    .A2(net2715),
    .B(_11413_),
    .Y(_11414_));
 NOR2x1_ASAP7_75t_R _40538_ (.A(_11412_),
    .B(_11414_),
    .Y(_11415_));
 AO21x1_ASAP7_75t_R _40539_ (.A1(_10394_),
    .A2(net2442),
    .B(net2248),
    .Y(_11416_));
 NOR2x1_ASAP7_75t_R _40540_ (.A(net1516),
    .B(net2247),
    .Y(_11417_));
 INVx1_ASAP7_75t_R _40541_ (.A(_11417_),
    .Y(_11418_));
 AND2x2_ASAP7_75t_R _40542_ (.A(_11416_),
    .B(_11418_),
    .Y(_11419_));
 NAND2x1_ASAP7_75t_R _40543_ (.A(_11415_),
    .B(_11419_),
    .Y(_11420_));
 NOR2x1_ASAP7_75t_R _40544_ (.A(_11410_),
    .B(_11420_),
    .Y(_11421_));
 NAND2x1_ASAP7_75t_R _40545_ (.A(_11405_),
    .B(_11421_),
    .Y(_11423_));
 NOR2x1_ASAP7_75t_R _40546_ (.A(_11392_),
    .B(_11423_),
    .Y(_11424_));
 NAND2x2_ASAP7_75t_R _40547_ (.A(_11362_),
    .B(_11424_),
    .Y(_11425_));
 NOR2x2_ASAP7_75t_R _40548_ (.A(_10364_),
    .B(_11425_),
    .Y(_11426_));
 INVx3_ASAP7_75t_R _40549_ (.A(net3336),
    .Y(_11427_));
 OAI21x1_ASAP7_75t_R _40550_ (.A1(_10287_),
    .A2(_10886_),
    .B(_11427_),
    .Y(_11428_));
 NAND3x2_ASAP7_75t_R _40551_ (.B(_10288_),
    .C(net3336),
    .Y(_11429_),
    .A(_10303_));
 NAND2x2_ASAP7_75t_R _40552_ (.A(_11428_),
    .B(_11429_),
    .Y(_11430_));
 OAI21x1_ASAP7_75t_R _40553_ (.A1(_11298_),
    .A2(_11304_),
    .B(_11430_),
    .Y(_11431_));
 XOR2x2_ASAP7_75t_R _40554_ (.A(_10304_),
    .B(_11427_),
    .Y(_11432_));
 XOR2x1_ASAP7_75t_R _40555_ (.A(_11297_),
    .Y(_11434_),
    .B(_11050_));
 NAND2x1_ASAP7_75t_R _40556_ (.A(_11434_),
    .B(_11432_),
    .Y(_11435_));
 AOI21x1_ASAP7_75t_R _40557_ (.A1(_11431_),
    .A2(_11435_),
    .B(net389),
    .Y(_11436_));
 OAI21x1_ASAP7_75t_R _40558_ (.A1(_10900_),
    .A2(_11436_),
    .B(_17435_),
    .Y(_11437_));
 NOR2x1_ASAP7_75t_R _40559_ (.A(net392),
    .B(_00818_),
    .Y(_11438_));
 NAND2x1_ASAP7_75t_R _40560_ (.A(_11430_),
    .B(_11434_),
    .Y(_11439_));
 XOR2x1_ASAP7_75t_R _40561_ (.A(_11297_),
    .Y(_11440_),
    .B(_11300_));
 NAND2x1_ASAP7_75t_R _40562_ (.A(_11432_),
    .B(_11440_),
    .Y(_11441_));
 AOI21x1_ASAP7_75t_R _40563_ (.A1(_11439_),
    .A2(_11441_),
    .B(net389),
    .Y(_11442_));
 OAI21x1_ASAP7_75t_R _40564_ (.A1(_11438_),
    .A2(_11442_),
    .B(_00410_),
    .Y(_11443_));
 NAND2x2_ASAP7_75t_R _40565_ (.A(_11437_),
    .B(_11443_),
    .Y(_00098_));
 AND2x2_ASAP7_75t_R _40566_ (.A(net389),
    .B(_00817_),
    .Y(_11445_));
 AO21x1_ASAP7_75t_R _40567_ (.A1(net1659),
    .A2(_10410_),
    .B(net2248),
    .Y(_11446_));
 NAND2x1_ASAP7_75t_R _40568_ (.A(_10576_),
    .B(_11413_),
    .Y(_11447_));
 NAND2x2_ASAP7_75t_R _40569_ (.A(net2456),
    .B(_11413_),
    .Y(_11448_));
 AND3x1_ASAP7_75t_R _40570_ (.A(_11446_),
    .B(_11447_),
    .C(_11448_),
    .Y(_11449_));
 AO21x1_ASAP7_75t_R _40571_ (.A1(net2851),
    .A2(net1125),
    .B(net2070),
    .Y(_11450_));
 AO21x1_ASAP7_75t_R _40572_ (.A1(_10394_),
    .A2(net1056),
    .B(net2070),
    .Y(_11451_));
 NOR2x1_ASAP7_75t_R _40573_ (.A(net2070),
    .B(net1659),
    .Y(_11452_));
 INVx1_ASAP7_75t_R _40574_ (.A(_11452_),
    .Y(_11453_));
 AND3x1_ASAP7_75t_R _40575_ (.A(_11450_),
    .B(_11451_),
    .C(_11453_),
    .Y(_11455_));
 AND2x2_ASAP7_75t_R _40576_ (.A(_11449_),
    .B(_11455_),
    .Y(_11456_));
 AO21x1_ASAP7_75t_R _40577_ (.A1(_10375_),
    .A2(net1114),
    .B(net2464),
    .Y(_11457_));
 AO21x1_ASAP7_75t_R _40578_ (.A1(net1876),
    .A2(net2441),
    .B(net2464),
    .Y(_11458_));
 AND2x2_ASAP7_75t_R _40579_ (.A(_11457_),
    .B(_11458_),
    .Y(_11459_));
 AO21x1_ASAP7_75t_R _40580_ (.A1(net2851),
    .A2(net1306),
    .B(net2465),
    .Y(_11460_));
 OA21x2_ASAP7_75t_R _40581_ (.A1(net2463),
    .A2(net2020),
    .B(_11460_),
    .Y(_11461_));
 NAND2x1_ASAP7_75t_R _40582_ (.A(_11459_),
    .B(_11461_),
    .Y(_11462_));
 NAND2x2_ASAP7_75t_R _40583_ (.A(_11341_),
    .B(_11397_),
    .Y(_11463_));
 NAND2x1_ASAP7_75t_R _40584_ (.A(net3034),
    .B(_11397_),
    .Y(_11464_));
 NAND2x1_ASAP7_75t_R _40585_ (.A(_11463_),
    .B(_11464_),
    .Y(_11466_));
 NOR2x1_ASAP7_75t_R _40586_ (.A(net1979),
    .B(net2354),
    .Y(_11467_));
 OR3x1_ASAP7_75t_R _40587_ (.A(_11466_),
    .B(_11467_),
    .C(_10473_),
    .Y(_11468_));
 NOR2x1_ASAP7_75t_R _40588_ (.A(_11462_),
    .B(_11468_),
    .Y(_11469_));
 NAND2x1_ASAP7_75t_R _40589_ (.A(_11456_),
    .B(_11469_),
    .Y(_11470_));
 OA21x2_ASAP7_75t_R _40590_ (.A1(_10383_),
    .A2(_11317_),
    .B(_11368_),
    .Y(_11471_));
 OA21x2_ASAP7_75t_R _40591_ (.A1(_10545_),
    .A2(_11341_),
    .B(_11368_),
    .Y(_11472_));
 NOR2x1_ASAP7_75t_R _40592_ (.A(_10505_),
    .B(_10358_),
    .Y(_11473_));
 OR3x1_ASAP7_75t_R _40593_ (.A(_11471_),
    .B(_11472_),
    .C(_11473_),
    .Y(_11474_));
 AOI22x1_ASAP7_75t_R _40594_ (.A1(_10342_),
    .A2(net2962),
    .B1(_10323_),
    .B2(_11338_),
    .Y(_11475_));
 AO21x1_ASAP7_75t_R _40595_ (.A1(net1115),
    .A2(net1306),
    .B(_10336_),
    .Y(_11477_));
 AO21x1_ASAP7_75t_R _40596_ (.A1(net2695),
    .A2(net2463),
    .B(_10336_),
    .Y(_11478_));
 NAND3x1_ASAP7_75t_R _40597_ (.A(_11475_),
    .B(_11477_),
    .C(_11478_),
    .Y(_11479_));
 NOR2x1_ASAP7_75t_R _40598_ (.A(_11474_),
    .B(_11479_),
    .Y(_11480_));
 INVx1_ASAP7_75t_R _40599_ (.A(_10431_),
    .Y(_11481_));
 AOI211x1_ASAP7_75t_R _40600_ (.A1(_10551_),
    .A2(_11481_),
    .B(_10441_),
    .C(_10443_),
    .Y(_11482_));
 AO21x1_ASAP7_75t_R _40601_ (.A1(net1494),
    .A2(net2851),
    .B(net1881),
    .Y(_11483_));
 OA21x2_ASAP7_75t_R _40602_ (.A1(_10421_),
    .A2(net1881),
    .B(_11483_),
    .Y(_11484_));
 NAND2x1_ASAP7_75t_R _40603_ (.A(_11482_),
    .B(_11484_),
    .Y(_11485_));
 NAND2x1_ASAP7_75t_R _40604_ (.A(net2951),
    .B(_10406_),
    .Y(_11486_));
 NOR2x2_ASAP7_75t_R _40605_ (.A(net2190),
    .B(_10415_),
    .Y(_11488_));
 INVx1_ASAP7_75t_R _40606_ (.A(_11488_),
    .Y(_11489_));
 OA21x2_ASAP7_75t_R _40607_ (.A1(net2868),
    .A2(_11486_),
    .B(_11489_),
    .Y(_11490_));
 NAND2x1_ASAP7_75t_R _40608_ (.A(_10406_),
    .B(_10481_),
    .Y(_11491_));
 AO21x1_ASAP7_75t_R _40609_ (.A1(net1659),
    .A2(_11312_),
    .B(net2536),
    .Y(_11492_));
 NAND3x1_ASAP7_75t_R _40610_ (.A(_11490_),
    .B(_11491_),
    .C(_11492_),
    .Y(_11493_));
 NOR2x1_ASAP7_75t_R _40611_ (.A(_11485_),
    .B(_11493_),
    .Y(_11494_));
 NAND2x2_ASAP7_75t_R _40612_ (.A(_11480_),
    .B(_11494_),
    .Y(_11495_));
 NOR2x2_ASAP7_75t_R _40613_ (.A(_11470_),
    .B(_11495_),
    .Y(_11496_));
 AO21x1_ASAP7_75t_R _40614_ (.A1(_11312_),
    .A2(net3161),
    .B(_10540_),
    .Y(_11497_));
 NAND2x2_ASAP7_75t_R _40615_ (.A(net3290),
    .B(_10537_),
    .Y(_11499_));
 NAND2x1_ASAP7_75t_R _40616_ (.A(_10537_),
    .B(_10526_),
    .Y(_11500_));
 NAND3x1_ASAP7_75t_R _40617_ (.A(_11497_),
    .B(_11499_),
    .C(_11500_),
    .Y(_11501_));
 AO21x1_ASAP7_75t_R _40618_ (.A1(net2952),
    .A2(_10505_),
    .B(net3043),
    .Y(_11502_));
 NAND2x1_ASAP7_75t_R _40619_ (.A(_10491_),
    .B(_10547_),
    .Y(_11503_));
 NAND2x1_ASAP7_75t_R _40620_ (.A(net1264),
    .B(_10547_),
    .Y(_11504_));
 NAND3x1_ASAP7_75t_R _40621_ (.A(_11502_),
    .B(_11503_),
    .C(_11504_),
    .Y(_11505_));
 TAPCELL_ASAP7_75t_R PHY_35 ();
 AO21x1_ASAP7_75t_R _40623_ (.A1(net1115),
    .A2(net3051),
    .B(net3043),
    .Y(_11507_));
 NAND2x1_ASAP7_75t_R _40624_ (.A(_10558_),
    .B(_11507_),
    .Y(_11508_));
 NOR3x1_ASAP7_75t_R _40625_ (.A(_11501_),
    .B(_11505_),
    .C(_11508_),
    .Y(_11510_));
 AO21x1_ASAP7_75t_R _40626_ (.A1(net2841),
    .A2(_11312_),
    .B(_10515_),
    .Y(_11511_));
 AO21x1_ASAP7_75t_R _40627_ (.A1(net1143),
    .A2(net2442),
    .B(_10515_),
    .Y(_11512_));
 AND2x2_ASAP7_75t_R _40628_ (.A(_11511_),
    .B(_11512_),
    .Y(_11513_));
 AO21x1_ASAP7_75t_R _40629_ (.A1(net1494),
    .A2(_11306_),
    .B(_10515_),
    .Y(_11514_));
 OAI21x1_ASAP7_75t_R _40630_ (.A1(net2806),
    .A2(_10520_),
    .B(_11350_),
    .Y(_11515_));
 AND2x2_ASAP7_75t_R _40631_ (.A(_11514_),
    .B(_11515_),
    .Y(_11516_));
 NAND2x1_ASAP7_75t_R _40632_ (.A(_11513_),
    .B(_11516_),
    .Y(_11517_));
 OA21x2_ASAP7_75t_R _40633_ (.A1(net3034),
    .A2(_11349_),
    .B(_10528_),
    .Y(_11518_));
 NOR2x1_ASAP7_75t_R _40634_ (.A(_11355_),
    .B(net1659),
    .Y(_11519_));
 AOI211x1_ASAP7_75t_R _40635_ (.A1(net975),
    .A2(net1318),
    .B(_11355_),
    .C(net2189),
    .Y(_11521_));
 OR3x1_ASAP7_75t_R _40636_ (.A(_11518_),
    .B(_11519_),
    .C(_11521_),
    .Y(_11522_));
 NOR2x1_ASAP7_75t_R _40637_ (.A(_11517_),
    .B(_11522_),
    .Y(_11523_));
 NAND2x1_ASAP7_75t_R _40638_ (.A(_11510_),
    .B(_11523_),
    .Y(_11524_));
 NAND2x1_ASAP7_75t_R _40639_ (.A(net1269),
    .B(_10589_),
    .Y(_11525_));
 OA21x2_ASAP7_75t_R _40640_ (.A1(net1318),
    .A2(_11525_),
    .B(_10587_),
    .Y(_11526_));
 AO21x1_ASAP7_75t_R _40641_ (.A1(_11323_),
    .A2(net3335),
    .B(_10586_),
    .Y(_11527_));
 OA21x2_ASAP7_75t_R _40642_ (.A1(net2227),
    .A2(_11306_),
    .B(_11527_),
    .Y(_11528_));
 NAND2x1_ASAP7_75t_R _40643_ (.A(_11526_),
    .B(_11528_),
    .Y(_11529_));
 AND3x1_ASAP7_75t_R _40644_ (.A(_10601_),
    .B(net2962),
    .C(net1269),
    .Y(_11530_));
 NOR2x1_ASAP7_75t_R _40645_ (.A(net3011),
    .B(_10382_),
    .Y(_11532_));
 OA21x2_ASAP7_75t_R _40646_ (.A1(_11317_),
    .A2(_11532_),
    .B(_10601_),
    .Y(_11533_));
 OA21x2_ASAP7_75t_R _40647_ (.A1(net3018),
    .A2(_11338_),
    .B(_10601_),
    .Y(_11534_));
 OR3x1_ASAP7_75t_R _40648_ (.A(_11530_),
    .B(_11533_),
    .C(_11534_),
    .Y(_11535_));
 NOR2x1_ASAP7_75t_R _40649_ (.A(_11529_),
    .B(_11535_),
    .Y(_11536_));
 AO21x1_ASAP7_75t_R _40650_ (.A1(net2854),
    .A2(net2952),
    .B(_10567_),
    .Y(_11537_));
 NAND2x1_ASAP7_75t_R _40651_ (.A(_10551_),
    .B(_10572_),
    .Y(_11538_));
 AND2x2_ASAP7_75t_R _40652_ (.A(_11537_),
    .B(_11538_),
    .Y(_11539_));
 AO21x1_ASAP7_75t_R _40653_ (.A1(net2695),
    .A2(net1125),
    .B(net2211),
    .Y(_11540_));
 NAND2x1_ASAP7_75t_R _40654_ (.A(net1496),
    .B(_10572_),
    .Y(_11541_));
 NAND3x1_ASAP7_75t_R _40655_ (.A(_11539_),
    .B(_11540_),
    .C(_11541_),
    .Y(_11543_));
 TAPCELL_ASAP7_75t_R PHY_34 ();
 AO21x1_ASAP7_75t_R _40657_ (.A1(net2957),
    .A2(net2841),
    .B(net1840),
    .Y(_11545_));
 AO21x1_ASAP7_75t_R _40658_ (.A1(net1144),
    .A2(_10410_),
    .B(net1840),
    .Y(_11546_));
 AND2x2_ASAP7_75t_R _40659_ (.A(_11545_),
    .B(_11546_),
    .Y(_11547_));
 AO21x1_ASAP7_75t_R _40660_ (.A1(net2561),
    .A2(net3292),
    .B(net2312),
    .Y(_11548_));
 AO21x1_ASAP7_75t_R _40661_ (.A1(net2695),
    .A2(net3335),
    .B(net2312),
    .Y(_11549_));
 NAND2x1_ASAP7_75t_R _40662_ (.A(net2715),
    .B(_10579_),
    .Y(_11550_));
 AND3x1_ASAP7_75t_R _40663_ (.A(_11548_),
    .B(_11549_),
    .C(_11550_),
    .Y(_11551_));
 NAND2x1_ASAP7_75t_R _40664_ (.A(_11547_),
    .B(_11551_),
    .Y(_11552_));
 NOR2x1_ASAP7_75t_R _40665_ (.A(_11543_),
    .B(_11552_),
    .Y(_11554_));
 NAND2x1_ASAP7_75t_R _40666_ (.A(_11536_),
    .B(_11554_),
    .Y(_11555_));
 NOR2x1_ASAP7_75t_R _40667_ (.A(_11524_),
    .B(_11555_),
    .Y(_11556_));
 NAND2x2_ASAP7_75t_R _40668_ (.A(_11496_),
    .B(_11556_),
    .Y(_11557_));
 INVx3_ASAP7_75t_R _40669_ (.A(_10003_),
    .Y(_11558_));
 NAND2x1_ASAP7_75t_R _40670_ (.A(net2804),
    .B(_11558_),
    .Y(_11559_));
 OA21x2_ASAP7_75t_R _40671_ (.A1(_10111_),
    .A2(net2662),
    .B(_11559_),
    .Y(_11560_));
 NAND2x1_ASAP7_75t_R _40672_ (.A(_09886_),
    .B(net2049),
    .Y(_11561_));
 NAND2x1_ASAP7_75t_R _40673_ (.A(_10077_),
    .B(_10099_),
    .Y(_11562_));
 OA21x2_ASAP7_75t_R _40674_ (.A1(_10035_),
    .A2(_11561_),
    .B(_11562_),
    .Y(_11563_));
 NAND2x1_ASAP7_75t_R _40675_ (.A(_11560_),
    .B(_11563_),
    .Y(_11565_));
 NOR2x2_ASAP7_75t_R _40676_ (.A(net1706),
    .B(_10058_),
    .Y(_11566_));
 AO22x1_ASAP7_75t_R _40677_ (.A1(_10157_),
    .A2(_10152_),
    .B1(_11566_),
    .B2(net2429),
    .Y(_11567_));
 AO22x1_ASAP7_75t_R _40678_ (.A1(_10097_),
    .A2(_10030_),
    .B1(net2382),
    .B2(_09970_),
    .Y(_11568_));
 OR2x2_ASAP7_75t_R _40679_ (.A(_11567_),
    .B(_11568_),
    .Y(_11569_));
 NOR2x1_ASAP7_75t_R _40680_ (.A(_11565_),
    .B(_11569_),
    .Y(_11570_));
 NOR2x2_ASAP7_75t_R _40681_ (.A(_09933_),
    .B(net1796),
    .Y(_11571_));
 AOI22x1_ASAP7_75t_R _40682_ (.A1(_09970_),
    .A2(_09992_),
    .B1(_11571_),
    .B2(net2429),
    .Y(_11572_));
 NAND2x1_ASAP7_75t_R _40683_ (.A(_09943_),
    .B(_09970_),
    .Y(_11573_));
 OA21x2_ASAP7_75t_R _40684_ (.A1(_10070_),
    .A2(_10137_),
    .B(_11573_),
    .Y(_11574_));
 NAND2x1_ASAP7_75t_R _40685_ (.A(_11572_),
    .B(_11574_),
    .Y(_11576_));
 NAND2x1_ASAP7_75t_R _40686_ (.A(_11201_),
    .B(_11228_),
    .Y(_11577_));
 NAND2x1_ASAP7_75t_R _40687_ (.A(_09941_),
    .B(_10157_),
    .Y(_11578_));
 INVx1_ASAP7_75t_R _40688_ (.A(_11578_),
    .Y(_11579_));
 NOR2x1_ASAP7_75t_R _40689_ (.A(_10040_),
    .B(_09913_),
    .Y(_11580_));
 OR3x2_ASAP7_75t_R _40690_ (.A(_11577_),
    .B(_11579_),
    .C(_11580_),
    .Y(_11581_));
 NOR2x1_ASAP7_75t_R _40691_ (.A(_11576_),
    .B(_11581_),
    .Y(_11582_));
 NAND2x2_ASAP7_75t_R _40692_ (.A(_11570_),
    .B(_11582_),
    .Y(_11583_));
 AO21x1_ASAP7_75t_R _40693_ (.A1(_10247_),
    .A2(_10015_),
    .B(_09990_),
    .Y(_11584_));
 AND2x2_ASAP7_75t_R _40694_ (.A(_10125_),
    .B(_11584_),
    .Y(_11585_));
 NOR2x1_ASAP7_75t_R _40695_ (.A(_09982_),
    .B(_09970_),
    .Y(_11587_));
 AO21x2_ASAP7_75t_R _40696_ (.A1(_11587_),
    .A2(net2375),
    .B(net2925),
    .Y(_11588_));
 NAND3x2_ASAP7_75t_R _40697_ (.B(_10190_),
    .C(_11588_),
    .Y(_11589_),
    .A(_11585_));
 AO21x2_ASAP7_75t_R _40698_ (.A1(net2925),
    .A2(net3093),
    .B(_09904_),
    .Y(_11590_));
 AO21x1_ASAP7_75t_R _40699_ (.A1(_09895_),
    .A2(_10207_),
    .B(_10005_),
    .Y(_11591_));
 OAI21x1_ASAP7_75t_R _40700_ (.A1(_00655_),
    .A2(_11590_),
    .B(_11591_),
    .Y(_11592_));
 NOR2x2_ASAP7_75t_R _40701_ (.A(_09934_),
    .B(_10246_),
    .Y(_11593_));
 OA21x2_ASAP7_75t_R _40702_ (.A1(_10020_),
    .A2(_11593_),
    .B(net978),
    .Y(_11594_));
 NOR2x1_ASAP7_75t_R _40703_ (.A(net1352),
    .B(_10070_),
    .Y(_11595_));
 OA21x2_ASAP7_75t_R _40704_ (.A1(_10196_),
    .A2(_11595_),
    .B(_10254_),
    .Y(_11596_));
 OR3x2_ASAP7_75t_R _40705_ (.A(_11592_),
    .B(_11594_),
    .C(_11596_),
    .Y(_11598_));
 NOR3x2_ASAP7_75t_R _40706_ (.B(_11589_),
    .C(_11598_),
    .Y(_11599_),
    .A(_11583_));
 AO21x2_ASAP7_75t_R _40707_ (.A1(_09914_),
    .A2(_09908_),
    .B(_09901_),
    .Y(_11600_));
 NAND2x2_ASAP7_75t_R _40708_ (.A(_10255_),
    .B(_11558_),
    .Y(_11601_));
 NAND2x2_ASAP7_75t_R _40709_ (.A(_09941_),
    .B(net2804),
    .Y(_11602_));
 NAND3x2_ASAP7_75t_R _40710_ (.B(_11601_),
    .C(_11602_),
    .Y(_11603_),
    .A(net2127));
 NAND2x2_ASAP7_75t_R _40711_ (.A(net1067),
    .B(_09979_),
    .Y(_11604_));
 NOR2x1_ASAP7_75t_R _40712_ (.A(_10005_),
    .B(_11604_),
    .Y(_11605_));
 AO21x1_ASAP7_75t_R _40713_ (.A1(_09946_),
    .A2(net2429),
    .B(_11605_),
    .Y(_11606_));
 OA21x2_ASAP7_75t_R _40714_ (.A1(_09943_),
    .A2(_10255_),
    .B(_10164_),
    .Y(_11607_));
 NOR3x2_ASAP7_75t_R _40715_ (.B(_11606_),
    .C(_11607_),
    .Y(_11609_),
    .A(_11603_));
 NAND2x2_ASAP7_75t_R _40716_ (.A(net2667),
    .B(_09905_),
    .Y(_11610_));
 NOR2x1_ASAP7_75t_R _40717_ (.A(_11610_),
    .B(_10060_),
    .Y(_11611_));
 OA21x2_ASAP7_75t_R _40718_ (.A1(_11212_),
    .A2(_10080_),
    .B(_10133_),
    .Y(_11612_));
 NOR2x1_ASAP7_75t_R _40719_ (.A(_11611_),
    .B(_11612_),
    .Y(_11613_));
 AO21x1_ASAP7_75t_R _40720_ (.A1(net948),
    .A2(net2212),
    .B(net2353),
    .Y(_11614_));
 NAND2x1_ASAP7_75t_R _40721_ (.A(_10157_),
    .B(_10143_),
    .Y(_11615_));
 NOR2x1_ASAP7_75t_R _40722_ (.A(_09925_),
    .B(_10035_),
    .Y(_11616_));
 INVx1_ASAP7_75t_R _40723_ (.A(_11616_),
    .Y(_11617_));
 NAND2x2_ASAP7_75t_R _40724_ (.A(_11615_),
    .B(_11617_),
    .Y(_11618_));
 INVx1_ASAP7_75t_R _40725_ (.A(_11618_),
    .Y(_11620_));
 AND3x1_ASAP7_75t_R _40726_ (.A(_11613_),
    .B(_11614_),
    .C(_11620_),
    .Y(_11621_));
 NOR2x1_ASAP7_75t_R _40727_ (.A(net1799),
    .B(_10040_),
    .Y(_11622_));
 NAND2x1_ASAP7_75t_R _40728_ (.A(net2373),
    .B(_11622_),
    .Y(_11623_));
 AO21x1_ASAP7_75t_R _40729_ (.A1(net948),
    .A2(net2212),
    .B(net2535),
    .Y(_11624_));
 NOR2x2_ASAP7_75t_R _40730_ (.A(_11610_),
    .B(_10246_),
    .Y(_11625_));
 INVx1_ASAP7_75t_R _40731_ (.A(_11625_),
    .Y(_11626_));
 INVx3_ASAP7_75t_R _40732_ (.A(_10207_),
    .Y(_11627_));
 NAND2x2_ASAP7_75t_R _40733_ (.A(_11627_),
    .B(_10140_),
    .Y(_11628_));
 AND4x1_ASAP7_75t_R _40734_ (.A(_11623_),
    .B(_11624_),
    .C(_11626_),
    .D(_11628_),
    .Y(_11629_));
 NAND3x1_ASAP7_75t_R _40735_ (.A(_11609_),
    .B(_11621_),
    .C(_11629_),
    .Y(_11631_));
 OA21x2_ASAP7_75t_R _40736_ (.A1(net2397),
    .A2(net2662),
    .B(_10241_),
    .Y(_11632_));
 AO21x1_ASAP7_75t_R _40737_ (.A1(_09895_),
    .A2(net2235),
    .B(_10035_),
    .Y(_11633_));
 NAND3x1_ASAP7_75t_R _40738_ (.A(_11632_),
    .B(_10230_),
    .C(_11633_),
    .Y(_11634_));
 AO32x1_ASAP7_75t_R _40739_ (.A1(net2591),
    .A2(net2283),
    .A3(_10255_),
    .B1(_10264_),
    .B2(_10099_),
    .Y(_11635_));
 AO21x1_ASAP7_75t_R _40740_ (.A1(_10060_),
    .A2(net2252),
    .B(_10042_),
    .Y(_11636_));
 NOR2x2_ASAP7_75t_R _40741_ (.A(net2374),
    .B(_10011_),
    .Y(_11637_));
 INVx2_ASAP7_75t_R _40742_ (.A(_11637_),
    .Y(_11638_));
 NAND2x2_ASAP7_75t_R _40743_ (.A(_11571_),
    .B(_10255_),
    .Y(_11639_));
 NAND3x1_ASAP7_75t_R _40744_ (.A(_11636_),
    .B(_11638_),
    .C(_11639_),
    .Y(_11640_));
 NOR3x1_ASAP7_75t_R _40745_ (.A(_11634_),
    .B(_11635_),
    .C(_11640_),
    .Y(_11642_));
 AO21x1_ASAP7_75t_R _40746_ (.A1(_09901_),
    .A2(net2660),
    .B(_09895_),
    .Y(_11643_));
 NAND2x1_ASAP7_75t_R _40747_ (.A(_10157_),
    .B(_11558_),
    .Y(_11644_));
 NOR2x1_ASAP7_75t_R _40748_ (.A(net3245),
    .B(net2660),
    .Y(_11645_));
 INVx1_ASAP7_75t_R _40749_ (.A(_11645_),
    .Y(_11646_));
 AND3x1_ASAP7_75t_R _40750_ (.A(_11643_),
    .B(_11644_),
    .C(_11646_),
    .Y(_11647_));
 NAND2x1_ASAP7_75t_R _40751_ (.A(_10161_),
    .B(_10044_),
    .Y(_11648_));
 AND4x1_ASAP7_75t_R _40752_ (.A(_11648_),
    .B(_10170_),
    .C(_10135_),
    .D(_10240_),
    .Y(_11649_));
 NAND2x1_ASAP7_75t_R _40753_ (.A(_11647_),
    .B(_11649_),
    .Y(_11650_));
 NOR2x1_ASAP7_75t_R _40754_ (.A(_09950_),
    .B(_10098_),
    .Y(_11651_));
 INVx1_ASAP7_75t_R _40755_ (.A(_11651_),
    .Y(_11653_));
 NAND2x1_ASAP7_75t_R _40756_ (.A(_09978_),
    .B(_10140_),
    .Y(_11654_));
 AND4x1_ASAP7_75t_R _40757_ (.A(_11653_),
    .B(_11654_),
    .C(_10079_),
    .D(_09944_),
    .Y(_11655_));
 NOR2x2_ASAP7_75t_R _40758_ (.A(net1707),
    .B(net3062),
    .Y(_11656_));
 INVx1_ASAP7_75t_R _40759_ (.A(_11656_),
    .Y(_11657_));
 NAND2x1_ASAP7_75t_R _40760_ (.A(_09978_),
    .B(_10099_),
    .Y(_11658_));
 NAND2x1_ASAP7_75t_R _40761_ (.A(_09876_),
    .B(_09970_),
    .Y(_11659_));
 AND4x1_ASAP7_75t_R _40762_ (.A(_11657_),
    .B(_11658_),
    .C(_11659_),
    .D(_10130_),
    .Y(_11660_));
 NAND2x1_ASAP7_75t_R _40763_ (.A(_11655_),
    .B(_11660_),
    .Y(_11661_));
 NOR2x1_ASAP7_75t_R _40764_ (.A(_11650_),
    .B(_11661_),
    .Y(_11662_));
 NAND2x1_ASAP7_75t_R _40765_ (.A(_11642_),
    .B(_11662_),
    .Y(_11664_));
 NOR2x1_ASAP7_75t_R _40766_ (.A(_11664_),
    .B(_11631_),
    .Y(_11665_));
 NAND2x2_ASAP7_75t_R _40767_ (.A(_11599_),
    .B(_11665_),
    .Y(_11666_));
 AO21x1_ASAP7_75t_R _40768_ (.A1(net1246),
    .A2(net1102),
    .B(net2775),
    .Y(_11667_));
 OAI21x1_ASAP7_75t_R _40769_ (.A1(net3069),
    .A2(net2547),
    .B(_11667_),
    .Y(_11668_));
 NAND2x1_ASAP7_75t_R _40770_ (.A(_09578_),
    .B(_09589_),
    .Y(_11669_));
 NOR2x1_ASAP7_75t_R _40771_ (.A(_11669_),
    .B(_09682_),
    .Y(_11670_));
 INVx1_ASAP7_75t_R _40772_ (.A(_11670_),
    .Y(_11671_));
 OAI22x1_ASAP7_75t_R _40773_ (.A1(_11671_),
    .A2(_09573_),
    .B1(_09779_),
    .B2(_09727_),
    .Y(_11672_));
 NOR2x2_ASAP7_75t_R _40774_ (.A(_11668_),
    .B(_11672_),
    .Y(_11673_));
 NOR2x2_ASAP7_75t_R _40775_ (.A(_09574_),
    .B(_09597_),
    .Y(_11675_));
 AND3x1_ASAP7_75t_R _40776_ (.A(_09701_),
    .B(_09780_),
    .C(net2152),
    .Y(_11676_));
 INVx2_ASAP7_75t_R _40777_ (.A(_09635_),
    .Y(_11677_));
 AND3x2_ASAP7_75t_R _40778_ (.A(_11677_),
    .B(_09701_),
    .C(_09573_),
    .Y(_11678_));
 AOI211x1_ASAP7_75t_R _40779_ (.A1(_11675_),
    .A2(_09696_),
    .B(_11676_),
    .C(_11678_),
    .Y(_11679_));
 NAND3x2_ASAP7_75t_R _40780_ (.B(_11679_),
    .C(_09704_),
    .Y(_11680_),
    .A(_11673_));
 TAPCELL_ASAP7_75t_R PHY_33 ();
 OA21x2_ASAP7_75t_R _40782_ (.A1(_09711_),
    .A2(net2547),
    .B(_09762_),
    .Y(_11682_));
 AO21x1_ASAP7_75t_R _40783_ (.A1(net1387),
    .A2(net1102),
    .B(net2656),
    .Y(_11683_));
 NOR2x1_ASAP7_75t_R _40784_ (.A(_09644_),
    .B(_09770_),
    .Y(_11684_));
 NAND2x1_ASAP7_75t_R _40785_ (.A(net1279),
    .B(_11684_),
    .Y(_11686_));
 AND3x1_ASAP7_75t_R _40786_ (.A(_11682_),
    .B(_11683_),
    .C(_11686_),
    .Y(_11687_));
 NOR2x2_ASAP7_75t_R _40787_ (.A(net1725),
    .B(net1507),
    .Y(_11688_));
 AOI22x1_ASAP7_75t_R _40788_ (.A1(_11688_),
    .A2(net1626),
    .B1(_11675_),
    .B2(_09826_),
    .Y(_11689_));
 INVx3_ASAP7_75t_R _40789_ (.A(_11111_),
    .Y(_11690_));
 AO21x1_ASAP7_75t_R _40790_ (.A1(_09707_),
    .A2(net2085),
    .B(_11690_),
    .Y(_11691_));
 NOR2x1_ASAP7_75t_R _40791_ (.A(_09770_),
    .B(_09858_),
    .Y(_11692_));
 AND2x2_ASAP7_75t_R _40792_ (.A(_09726_),
    .B(_11069_),
    .Y(_11693_));
 NOR2x1_ASAP7_75t_R _40793_ (.A(_11692_),
    .B(_11693_),
    .Y(_11694_));
 AND3x1_ASAP7_75t_R _40794_ (.A(_11689_),
    .B(_11691_),
    .C(_11694_),
    .Y(_11695_));
 NAND2x2_ASAP7_75t_R _40795_ (.A(_11687_),
    .B(_11695_),
    .Y(_11697_));
 AOI22x1_ASAP7_75t_R _40796_ (.A1(_11677_),
    .A2(_09846_),
    .B1(_11168_),
    .B2(_11111_),
    .Y(_11698_));
 AND3x1_ASAP7_75t_R _40797_ (.A(_09726_),
    .B(net2817),
    .C(_09608_),
    .Y(_11699_));
 INVx1_ASAP7_75t_R _40798_ (.A(_11699_),
    .Y(_11700_));
 NAND2x1_ASAP7_75t_R _40799_ (.A(_11698_),
    .B(_11700_),
    .Y(_11701_));
 AO21x1_ASAP7_75t_R _40800_ (.A1(net2553),
    .A2(net2817),
    .B(net1476),
    .Y(_11702_));
 AND3x2_ASAP7_75t_R _40801_ (.A(_09846_),
    .B(net2817),
    .C(_09608_),
    .Y(_11703_));
 INVx1_ASAP7_75t_R _40802_ (.A(_11703_),
    .Y(_11704_));
 OAI21x1_ASAP7_75t_R _40803_ (.A1(net1942),
    .A2(_11702_),
    .B(_11704_),
    .Y(_11705_));
 NOR2x1_ASAP7_75t_R _40804_ (.A(_11701_),
    .B(_11705_),
    .Y(_11706_));
 NOR2x2_ASAP7_75t_R _40805_ (.A(net2861),
    .B(_09597_),
    .Y(_11708_));
 OA21x2_ASAP7_75t_R _40806_ (.A1(_11708_),
    .A2(_11180_),
    .B(net1218),
    .Y(_11709_));
 AO21x2_ASAP7_75t_R _40807_ (.A1(_11161_),
    .A2(_09653_),
    .B(net1871),
    .Y(_11710_));
 AO21x1_ASAP7_75t_R _40808_ (.A1(net1518),
    .A2(_11161_),
    .B(net2692),
    .Y(_11711_));
 NAND2x2_ASAP7_75t_R _40809_ (.A(_11710_),
    .B(_11711_),
    .Y(_11712_));
 AOI211x1_ASAP7_75t_R _40810_ (.A1(net2956),
    .A2(_11090_),
    .B(_11709_),
    .C(_11712_),
    .Y(_11713_));
 NAND2x2_ASAP7_75t_R _40811_ (.A(_11706_),
    .B(_11713_),
    .Y(_11714_));
 NOR3x2_ASAP7_75t_R _40812_ (.B(_11697_),
    .C(_11714_),
    .Y(_11715_),
    .A(_11680_));
 NOR2x1_ASAP7_75t_R _40813_ (.A(net985),
    .B(net1502),
    .Y(_11716_));
 NOR2x1_ASAP7_75t_R _40814_ (.A(_09597_),
    .B(net2501),
    .Y(_11717_));
 OAI21x1_ASAP7_75t_R _40815_ (.A1(_11716_),
    .A2(_11717_),
    .B(_09589_),
    .Y(_11719_));
 NAND2x2_ASAP7_75t_R _40816_ (.A(_11719_),
    .B(_11130_),
    .Y(_11720_));
 AOI21x1_ASAP7_75t_R _40817_ (.A1(_11091_),
    .A2(_11179_),
    .B(net1110),
    .Y(_11721_));
 NOR2x2_ASAP7_75t_R _40818_ (.A(net1481),
    .B(net2291),
    .Y(_11722_));
 OAI21x1_ASAP7_75t_R _40819_ (.A1(_11722_),
    .A2(_11114_),
    .B(net1112),
    .Y(_11723_));
 INVx2_ASAP7_75t_R _40820_ (.A(_11723_),
    .Y(_11724_));
 NOR3x2_ASAP7_75t_R _40821_ (.B(_11721_),
    .C(_11724_),
    .Y(_11725_),
    .A(_11720_));
 NOR2x1_ASAP7_75t_R _40822_ (.A(net2961),
    .B(net2103),
    .Y(_11726_));
 AO22x2_ASAP7_75t_R _40823_ (.A1(_11134_),
    .A2(_09726_),
    .B1(_11726_),
    .B2(net1280),
    .Y(_11727_));
 AO21x1_ASAP7_75t_R _40824_ (.A1(net1544),
    .A2(net2940),
    .B(net1504),
    .Y(_11728_));
 OAI21x1_ASAP7_75t_R _40825_ (.A1(net3069),
    .A2(net1505),
    .B(_11728_),
    .Y(_11730_));
 NOR2x1_ASAP7_75t_R _40826_ (.A(_09739_),
    .B(_09620_),
    .Y(_11731_));
 INVx1_ASAP7_75t_R _40827_ (.A(_11731_),
    .Y(_11732_));
 OAI21x1_ASAP7_75t_R _40828_ (.A1(_09573_),
    .A2(_11067_),
    .B(_11732_),
    .Y(_11733_));
 NOR3x2_ASAP7_75t_R _40829_ (.B(_11730_),
    .C(_11733_),
    .Y(_11734_),
    .A(_11727_));
 NAND2x2_ASAP7_75t_R _40830_ (.A(_11725_),
    .B(_11734_),
    .Y(_11735_));
 INVx1_ASAP7_75t_R _40831_ (.A(_09715_),
    .Y(_11736_));
 NOR2x1_ASAP7_75t_R _40832_ (.A(_09812_),
    .B(net2959),
    .Y(_11737_));
 AOI21x1_ASAP7_75t_R _40833_ (.A1(_11736_),
    .A2(_11056_),
    .B(_11737_),
    .Y(_11738_));
 NAND2x1_ASAP7_75t_R _40834_ (.A(_11168_),
    .B(net3177),
    .Y(_11739_));
 NAND3x1_ASAP7_75t_R _40835_ (.A(_11738_),
    .B(_11185_),
    .C(_11739_),
    .Y(_11741_));
 AOI22x1_ASAP7_75t_R _40836_ (.A1(_11056_),
    .A2(_09832_),
    .B1(_11090_),
    .B2(_09700_),
    .Y(_11742_));
 AO21x1_ASAP7_75t_R _40837_ (.A1(_09674_),
    .A2(_09579_),
    .B(net2942),
    .Y(_11743_));
 NAND2x1_ASAP7_75t_R _40838_ (.A(_09809_),
    .B(_09807_),
    .Y(_11744_));
 NAND3x1_ASAP7_75t_R _40839_ (.A(_11742_),
    .B(_11743_),
    .C(_11744_),
    .Y(_11745_));
 NOR2x1_ASAP7_75t_R _40840_ (.A(_11741_),
    .B(_11745_),
    .Y(_11746_));
 AOI22x1_ASAP7_75t_R _40841_ (.A1(_11096_),
    .A2(_09640_),
    .B1(_09826_),
    .B2(_11111_),
    .Y(_11747_));
 NAND2x1_ASAP7_75t_R _40842_ (.A(_09759_),
    .B(_09754_),
    .Y(_11748_));
 OA21x2_ASAP7_75t_R _40843_ (.A1(net3241),
    .A2(net1246),
    .B(_11748_),
    .Y(_11749_));
 NAND2x1_ASAP7_75t_R _40844_ (.A(_11747_),
    .B(_11749_),
    .Y(_11750_));
 AOI22x1_ASAP7_75t_R _40845_ (.A1(_11090_),
    .A2(_11096_),
    .B1(_09838_),
    .B2(_11677_),
    .Y(_11752_));
 NAND2x1_ASAP7_75t_R _40846_ (.A(net2927),
    .B(_09700_),
    .Y(_11753_));
 NAND3x1_ASAP7_75t_R _40847_ (.A(_11752_),
    .B(_11753_),
    .C(_11097_),
    .Y(_11754_));
 NOR2x1_ASAP7_75t_R _40848_ (.A(_11750_),
    .B(_11754_),
    .Y(_11755_));
 NAND2x2_ASAP7_75t_R _40849_ (.A(_11746_),
    .B(_11755_),
    .Y(_11756_));
 AOI22x1_ASAP7_75t_R _40850_ (.A1(_09807_),
    .A2(_11069_),
    .B1(_09783_),
    .B2(_09759_),
    .Y(_11757_));
 AO21x1_ASAP7_75t_R _40851_ (.A1(net1743),
    .A2(_09801_),
    .B(net2047),
    .Y(_11758_));
 AND3x1_ASAP7_75t_R _40852_ (.A(_11757_),
    .B(_09803_),
    .C(_11758_),
    .Y(_11759_));
 NOR2x1_ASAP7_75t_R _40853_ (.A(net1724),
    .B(_09574_),
    .Y(_11760_));
 AOI22x1_ASAP7_75t_R _40854_ (.A1(net2941),
    .A2(_09838_),
    .B1(_09640_),
    .B2(_11760_),
    .Y(_11761_));
 NAND2x2_ASAP7_75t_R _40855_ (.A(_09726_),
    .B(_11180_),
    .Y(_11763_));
 NAND2x2_ASAP7_75t_R _40856_ (.A(_11708_),
    .B(_09757_),
    .Y(_11764_));
 NAND3x2_ASAP7_75t_R _40857_ (.B(_11763_),
    .C(_11764_),
    .Y(_11765_),
    .A(_11761_));
 CKINVDCx5p33_ASAP7_75t_R _40858_ (.A(_09644_),
    .Y(_11766_));
 AOI22x1_ASAP7_75t_R _40859_ (.A1(_11090_),
    .A2(_11766_),
    .B1(_09612_),
    .B2(_11168_),
    .Y(_11767_));
 NAND2x2_ASAP7_75t_R _40860_ (.A(_11180_),
    .B(_09807_),
    .Y(_11768_));
 NAND2x2_ASAP7_75t_R _40861_ (.A(net2920),
    .B(_11090_),
    .Y(_11769_));
 NAND3x2_ASAP7_75t_R _40862_ (.B(_11768_),
    .C(_11769_),
    .Y(_11770_),
    .A(_11767_));
 NOR2x2_ASAP7_75t_R _40863_ (.A(_11765_),
    .B(_11770_),
    .Y(_11771_));
 NAND2x2_ASAP7_75t_R _40864_ (.A(_11759_),
    .B(_11771_),
    .Y(_11772_));
 NOR3x2_ASAP7_75t_R _40865_ (.B(_11756_),
    .C(_11772_),
    .Y(_11774_),
    .A(_11735_));
 NAND2x2_ASAP7_75t_R _40866_ (.A(_11715_),
    .B(_11774_),
    .Y(_11775_));
 XOR2x2_ASAP7_75t_R _40867_ (.A(_11666_),
    .B(_11775_),
    .Y(_11776_));
 NOR2x1_ASAP7_75t_R _40868_ (.A(_11557_),
    .B(_11776_),
    .Y(_11777_));
 INVx1_ASAP7_75t_R _40869_ (.A(_11557_),
    .Y(_11778_));
 XNOR2x2_ASAP7_75t_R _40870_ (.A(_11775_),
    .B(_11666_),
    .Y(_11779_));
 NOR2x1_ASAP7_75t_R _40871_ (.A(_11778_),
    .B(_11779_),
    .Y(_11780_));
 AO21x1_ASAP7_75t_R _40872_ (.A1(net1446),
    .A2(net1492),
    .B(_10725_),
    .Y(_11781_));
 NAND2x1_ASAP7_75t_R _40873_ (.A(_10968_),
    .B(_11781_),
    .Y(_11782_));
 OR3x2_ASAP7_75t_R _40874_ (.A(_10725_),
    .B(_10623_),
    .C(net1996),
    .Y(_11783_));
 NAND2x1_ASAP7_75t_R _40875_ (.A(_10959_),
    .B(_11783_),
    .Y(_11785_));
 NOR2x1_ASAP7_75t_R _40876_ (.A(_11782_),
    .B(_11785_),
    .Y(_11786_));
 AO21x1_ASAP7_75t_R _40877_ (.A1(_10671_),
    .A2(_10693_),
    .B(_10739_),
    .Y(_11787_));
 AO21x1_ASAP7_75t_R _40878_ (.A1(_10744_),
    .A2(net1446),
    .B(_10739_),
    .Y(_11788_));
 AND3x1_ASAP7_75t_R _40879_ (.A(_10743_),
    .B(_11787_),
    .C(_11788_),
    .Y(_11789_));
 NAND2x1_ASAP7_75t_R _40880_ (.A(_11786_),
    .B(_11789_),
    .Y(_11790_));
 AO21x1_ASAP7_75t_R _40881_ (.A1(_10783_),
    .A2(net2061),
    .B(net3042),
    .Y(_11791_));
 TAPCELL_ASAP7_75t_R PHY_32 ();
 AO21x1_ASAP7_75t_R _40883_ (.A1(_10757_),
    .A2(_10807_),
    .B(net3042),
    .Y(_11793_));
 AO21x1_ASAP7_75t_R _40884_ (.A1(_10624_),
    .A2(_10645_),
    .B(net3042),
    .Y(_11794_));
 AND3x1_ASAP7_75t_R _40885_ (.A(_11791_),
    .B(_11793_),
    .C(_11794_),
    .Y(_11796_));
 AO21x1_ASAP7_75t_R _40886_ (.A1(net3065),
    .A2(net1475),
    .B(_10755_),
    .Y(_11797_));
 NOR2x2_ASAP7_75t_R _40887_ (.A(_10644_),
    .B(_10685_),
    .Y(_11798_));
 NAND2x1_ASAP7_75t_R _40888_ (.A(_10754_),
    .B(_11798_),
    .Y(_11799_));
 AND2x2_ASAP7_75t_R _40889_ (.A(_11797_),
    .B(_11799_),
    .Y(_11800_));
 NAND2x1_ASAP7_75t_R _40890_ (.A(net1346),
    .B(_10754_),
    .Y(_11801_));
 AO21x1_ASAP7_75t_R _40891_ (.A1(net1288),
    .A2(_10660_),
    .B(_10755_),
    .Y(_11802_));
 AND2x2_ASAP7_75t_R _40892_ (.A(_11801_),
    .B(_11802_),
    .Y(_11803_));
 NAND3x1_ASAP7_75t_R _40893_ (.A(_11796_),
    .B(_11800_),
    .C(_11803_),
    .Y(_11804_));
 NOR2x1_ASAP7_75t_R _40894_ (.A(_11790_),
    .B(_11804_),
    .Y(_11805_));
 AO21x1_ASAP7_75t_R _40895_ (.A1(net3022),
    .A2(_10788_),
    .B(_10696_),
    .Y(_11807_));
 NOR2x1_ASAP7_75t_R _40896_ (.A(_10759_),
    .B(_10696_),
    .Y(_11808_));
 INVx1_ASAP7_75t_R _40897_ (.A(_11808_),
    .Y(_11809_));
 AO21x1_ASAP7_75t_R _40898_ (.A1(_10660_),
    .A2(_10656_),
    .B(_10696_),
    .Y(_11810_));
 AND3x1_ASAP7_75t_R _40899_ (.A(_11807_),
    .B(_11809_),
    .C(_11810_),
    .Y(_11811_));
 INVx2_ASAP7_75t_R _40900_ (.A(_10905_),
    .Y(_11812_));
 OA21x2_ASAP7_75t_R _40901_ (.A1(_11812_),
    .A2(_10782_),
    .B(_10713_),
    .Y(_11813_));
 AOI21x1_ASAP7_75t_R _40902_ (.A1(_10713_),
    .A2(_11798_),
    .B(_11813_),
    .Y(_11814_));
 AO21x1_ASAP7_75t_R _40903_ (.A1(_10921_),
    .A2(_10694_),
    .B(_10696_),
    .Y(_11815_));
 NAND3x1_ASAP7_75t_R _40904_ (.A(_11811_),
    .B(_11814_),
    .C(_11815_),
    .Y(_11816_));
 AO21x1_ASAP7_75t_R _40905_ (.A1(net1862),
    .A2(_10671_),
    .B(net3045),
    .Y(_11818_));
 AO21x1_ASAP7_75t_R _40906_ (.A1(_10700_),
    .A2(_10660_),
    .B(net3045),
    .Y(_11819_));
 NAND2x1_ASAP7_75t_R _40907_ (.A(_10681_),
    .B(_10642_),
    .Y(_11820_));
 AND3x1_ASAP7_75t_R _40908_ (.A(_11818_),
    .B(_11819_),
    .C(_11820_),
    .Y(_11821_));
 INVx2_ASAP7_75t_R _40909_ (.A(_10664_),
    .Y(_11822_));
 NAND2x1_ASAP7_75t_R _40910_ (.A(_10711_),
    .B(_11822_),
    .Y(_11823_));
 AO21x1_ASAP7_75t_R _40911_ (.A1(_10767_),
    .A2(_10671_),
    .B(net3021),
    .Y(_11824_));
 NAND2x1_ASAP7_75t_R _40912_ (.A(_11823_),
    .B(_11824_),
    .Y(_11825_));
 NOR2x1_ASAP7_75t_R _40913_ (.A(_10913_),
    .B(_11825_),
    .Y(_11826_));
 AO21x1_ASAP7_75t_R _40914_ (.A1(net1446),
    .A2(net1492),
    .B(net3021),
    .Y(_11827_));
 OA21x2_ASAP7_75t_R _40915_ (.A1(_10740_),
    .A2(net3021),
    .B(_11827_),
    .Y(_11829_));
 NAND3x1_ASAP7_75t_R _40916_ (.A(_11821_),
    .B(_11826_),
    .C(_11829_),
    .Y(_11830_));
 NOR2x1_ASAP7_75t_R _40917_ (.A(_11816_),
    .B(_11830_),
    .Y(_11831_));
 NAND2x2_ASAP7_75t_R _40918_ (.A(_11805_),
    .B(_11831_),
    .Y(_11832_));
 INVx2_ASAP7_75t_R _40919_ (.A(_10796_),
    .Y(_11833_));
 OA21x2_ASAP7_75t_R _40920_ (.A1(_10846_),
    .A2(_11008_),
    .B(_11833_),
    .Y(_11834_));
 NAND2x1_ASAP7_75t_R _40921_ (.A(net1337),
    .B(_11833_),
    .Y(_11835_));
 NOR2x1_ASAP7_75t_R _40922_ (.A(_10807_),
    .B(_10796_),
    .Y(_11836_));
 INVx1_ASAP7_75t_R _40923_ (.A(_11836_),
    .Y(_11837_));
 NAND2x1_ASAP7_75t_R _40924_ (.A(_11835_),
    .B(_11837_),
    .Y(_11838_));
 NOR2x1_ASAP7_75t_R _40925_ (.A(_11834_),
    .B(_11838_),
    .Y(_11840_));
 AO21x1_ASAP7_75t_R _40926_ (.A1(_10678_),
    .A2(_10747_),
    .B(_10785_),
    .Y(_11841_));
 AO31x2_ASAP7_75t_R _40927_ (.A1(net3058),
    .A2(net3057),
    .A3(net1446),
    .B(_10785_),
    .Y(_11842_));
 NAND3x1_ASAP7_75t_R _40928_ (.A(_11840_),
    .B(_11841_),
    .C(_11842_),
    .Y(_11843_));
 TAPCELL_ASAP7_75t_R PHY_31 ();
 AO21x1_ASAP7_75t_R _40930_ (.A1(_10744_),
    .A2(net1492),
    .B(net3056),
    .Y(_11845_));
 AO21x1_ASAP7_75t_R _40931_ (.A1(net1288),
    .A2(_10660_),
    .B(_10816_),
    .Y(_11846_));
 NOR2x1_ASAP7_75t_R _40932_ (.A(_10658_),
    .B(net1997),
    .Y(_11847_));
 OAI21x1_ASAP7_75t_R _40933_ (.A1(net3061),
    .A2(_11847_),
    .B(_10992_),
    .Y(_11848_));
 AND3x1_ASAP7_75t_R _40934_ (.A(_11845_),
    .B(_11846_),
    .C(_11848_),
    .Y(_11849_));
 INVx4_ASAP7_75t_R _40935_ (.A(_10751_),
    .Y(_11851_));
 OA21x2_ASAP7_75t_R _40936_ (.A1(_11851_),
    .A2(_11812_),
    .B(_10809_),
    .Y(_11852_));
 INVx1_ASAP7_75t_R _40937_ (.A(_10807_),
    .Y(_11853_));
 OA21x2_ASAP7_75t_R _40938_ (.A1(_10869_),
    .A2(_11853_),
    .B(_10809_),
    .Y(_11854_));
 AOI211x1_ASAP7_75t_R _40939_ (.A1(_10792_),
    .A2(_10809_),
    .B(_11852_),
    .C(_11854_),
    .Y(_11855_));
 NAND2x1_ASAP7_75t_R _40940_ (.A(_11849_),
    .B(_11855_),
    .Y(_11856_));
 NOR2x1_ASAP7_75t_R _40941_ (.A(_11843_),
    .B(_11856_),
    .Y(_11857_));
 AOI21x1_ASAP7_75t_R _40942_ (.A1(_10807_),
    .A2(_10757_),
    .B(_10851_),
    .Y(_11858_));
 NOR2x1_ASAP7_75t_R _40943_ (.A(_10856_),
    .B(_11858_),
    .Y(_11859_));
 INVx1_ASAP7_75t_R _40944_ (.A(_10851_),
    .Y(_11860_));
 NAND2x1_ASAP7_75t_R _40945_ (.A(_10711_),
    .B(_11860_),
    .Y(_11862_));
 AO21x1_ASAP7_75t_R _40946_ (.A1(net1862),
    .A2(_11039_),
    .B(_10843_),
    .Y(_11863_));
 AOI21x1_ASAP7_75t_R _40947_ (.A1(_10759_),
    .A2(_10832_),
    .B(_10843_),
    .Y(_11864_));
 INVx1_ASAP7_75t_R _40948_ (.A(_11864_),
    .Y(_11865_));
 AND4x1_ASAP7_75t_R _40949_ (.A(_11859_),
    .B(_11862_),
    .C(_11863_),
    .D(_11865_),
    .Y(_11866_));
 AO31x2_ASAP7_75t_R _40950_ (.A1(_10694_),
    .A2(net1475),
    .A3(_10783_),
    .B(_10826_),
    .Y(_11867_));
 NOR2x1_ASAP7_75t_R _40951_ (.A(_10759_),
    .B(_10826_),
    .Y(_11868_));
 NOR2x1_ASAP7_75t_R _40952_ (.A(_10624_),
    .B(net3031),
    .Y(_11869_));
 AOI211x1_ASAP7_75t_R _40953_ (.A1(_10827_),
    .A2(_10831_),
    .B(_11868_),
    .C(_11869_),
    .Y(_11870_));
 NAND2x1_ASAP7_75t_R _40954_ (.A(_11867_),
    .B(_11870_),
    .Y(_11871_));
 TAPCELL_ASAP7_75t_R PHY_30 ();
 AO31x2_ASAP7_75t_R _40956_ (.A1(_10624_),
    .A2(_10645_),
    .A3(net1446),
    .B(_10864_),
    .Y(_11874_));
 AOI211x1_ASAP7_75t_R _40957_ (.A1(net1501),
    .A2(net1420),
    .B(_10864_),
    .C(net2023),
    .Y(_11875_));
 INVx1_ASAP7_75t_R _40958_ (.A(_11875_),
    .Y(_11876_));
 AO21x1_ASAP7_75t_R _40959_ (.A1(net3065),
    .A2(net1475),
    .B(_10864_),
    .Y(_11877_));
 NAND3x1_ASAP7_75t_R _40960_ (.A(_11874_),
    .B(_11876_),
    .C(_11877_),
    .Y(_11878_));
 NOR2x1_ASAP7_75t_R _40961_ (.A(_11871_),
    .B(_11878_),
    .Y(_11879_));
 AND2x2_ASAP7_75t_R _40962_ (.A(_11866_),
    .B(_11879_),
    .Y(_11880_));
 NAND2x2_ASAP7_75t_R _40963_ (.A(_11857_),
    .B(_11880_),
    .Y(_11881_));
 AND3x2_ASAP7_75t_R _40964_ (.A(_10984_),
    .B(_10981_),
    .C(_10982_),
    .Y(_11882_));
 NAND3x2_ASAP7_75t_R _40965_ (.B(net3044),
    .C(_10988_),
    .Y(_11884_),
    .A(_11882_));
 NOR3x2_ASAP7_75t_R _40966_ (.B(_10723_),
    .C(_10734_),
    .Y(_11885_),
    .A(_11884_));
 NOR3x2_ASAP7_75t_R _40967_ (.B(_11881_),
    .C(_11885_),
    .Y(_11886_),
    .A(_11832_));
 XOR2x2_ASAP7_75t_R _40968_ (.A(_11886_),
    .B(_11296_),
    .Y(_11887_));
 OAI21x1_ASAP7_75t_R _40969_ (.A1(_11777_),
    .A2(_11780_),
    .B(_11887_),
    .Y(_11888_));
 NOR2x1_ASAP7_75t_R _40970_ (.A(_11778_),
    .B(_11776_),
    .Y(_11889_));
 NOR2x1_ASAP7_75t_R _40971_ (.A(_11557_),
    .B(_11779_),
    .Y(_11890_));
 INVx1_ASAP7_75t_R _40972_ (.A(_11887_),
    .Y(_11891_));
 OAI21x1_ASAP7_75t_R _40973_ (.A1(_11889_),
    .A2(_11890_),
    .B(_11891_),
    .Y(_11892_));
 AOI21x1_ASAP7_75t_R _40974_ (.A1(_11888_),
    .A2(_11892_),
    .B(net389),
    .Y(_11893_));
 NOR2x1_ASAP7_75t_R _40975_ (.A(_11445_),
    .B(_11893_),
    .Y(_11895_));
 XOR2x2_ASAP7_75t_R _40976_ (.A(_11895_),
    .B(_17438_),
    .Y(_00099_));
 AND2x2_ASAP7_75t_R _40977_ (.A(net389),
    .B(_00816_),
    .Y(_11896_));
 AO21x1_ASAP7_75t_R _40978_ (.A1(_10502_),
    .A2(net3292),
    .B(net2312),
    .Y(_11897_));
 AO21x1_ASAP7_75t_R _40979_ (.A1(net2332),
    .A2(_10410_),
    .B(net2312),
    .Y(_11898_));
 AND3x1_ASAP7_75t_R _40980_ (.A(_11897_),
    .B(_11898_),
    .C(_11550_),
    .Y(_11899_));
 AO21x1_ASAP7_75t_R _40981_ (.A1(_11312_),
    .A2(net2332),
    .B(_10567_),
    .Y(_11900_));
 OAI21x1_ASAP7_75t_R _40982_ (.A1(_10341_),
    .A2(_10567_),
    .B(_11900_),
    .Y(_11901_));
 AO21x1_ASAP7_75t_R _40983_ (.A1(net3157),
    .A2(net1855),
    .B(_10567_),
    .Y(_11902_));
 OAI21x1_ASAP7_75t_R _40984_ (.A1(_10567_),
    .A2(_10502_),
    .B(_11902_),
    .Y(_11903_));
 NOR2x1_ASAP7_75t_R _40985_ (.A(_11901_),
    .B(_11903_),
    .Y(_11905_));
 NAND2x1_ASAP7_75t_R _40986_ (.A(_11899_),
    .B(_11905_),
    .Y(_11906_));
 NAND2x2_ASAP7_75t_R _40987_ (.A(net3018),
    .B(_10589_),
    .Y(_11907_));
 NAND2x1_ASAP7_75t_R _40988_ (.A(_11907_),
    .B(_10587_),
    .Y(_11908_));
 NOR2x1_ASAP7_75t_R _40989_ (.A(_10592_),
    .B(_11908_),
    .Y(_11909_));
 OA21x2_ASAP7_75t_R _40990_ (.A1(_11532_),
    .A2(_10531_),
    .B(_10589_),
    .Y(_11910_));
 OA21x2_ASAP7_75t_R _40991_ (.A1(_10383_),
    .A2(_10385_),
    .B(_10589_),
    .Y(_11911_));
 AOI211x1_ASAP7_75t_R _40992_ (.A1(_10554_),
    .A2(_10589_),
    .B(_11910_),
    .C(_11911_),
    .Y(_11912_));
 NAND2x2_ASAP7_75t_R _40993_ (.A(_11909_),
    .B(_11912_),
    .Y(_11913_));
 AO21x1_ASAP7_75t_R _40994_ (.A1(net2695),
    .A2(_10449_),
    .B(_10600_),
    .Y(_11914_));
 AO21x1_ASAP7_75t_R _40995_ (.A1(net2561),
    .A2(_11306_),
    .B(_10600_),
    .Y(_11916_));
 AND2x2_ASAP7_75t_R _40996_ (.A(_11914_),
    .B(_11916_),
    .Y(_11917_));
 AOI211x1_ASAP7_75t_R _40997_ (.A1(net1373),
    .A2(_10316_),
    .B(_10600_),
    .C(_10341_),
    .Y(_11918_));
 NOR2x2_ASAP7_75t_R _40998_ (.A(net2526),
    .B(net2331),
    .Y(_11919_));
 NOR2x2_ASAP7_75t_R _40999_ (.A(net2526),
    .B(_11312_),
    .Y(_11920_));
 NOR3x2_ASAP7_75t_R _41000_ (.B(_11919_),
    .C(_11920_),
    .Y(_11921_),
    .A(_11918_));
 NAND2x2_ASAP7_75t_R _41001_ (.A(_11917_),
    .B(_11921_),
    .Y(_11922_));
 NOR3x1_ASAP7_75t_R _41002_ (.A(_11906_),
    .B(_11913_),
    .C(_11922_),
    .Y(_11923_));
 AO21x1_ASAP7_75t_R _41003_ (.A1(_10370_),
    .A2(_10471_),
    .B(_10540_),
    .Y(_11924_));
 NAND2x1_ASAP7_75t_R _41004_ (.A(_11499_),
    .B(_11924_),
    .Y(_11925_));
 AO21x2_ASAP7_75t_R _41005_ (.A1(_10485_),
    .A2(_10329_),
    .B(_10540_),
    .Y(_11927_));
 OAI21x1_ASAP7_75t_R _41006_ (.A1(_10341_),
    .A2(_10540_),
    .B(_11927_),
    .Y(_11928_));
 NOR2x1_ASAP7_75t_R _41007_ (.A(_11925_),
    .B(_11928_),
    .Y(_11929_));
 AO21x1_ASAP7_75t_R _41008_ (.A1(_10502_),
    .A2(_10490_),
    .B(net3043),
    .Y(_11930_));
 AO21x1_ASAP7_75t_R _41009_ (.A1(net1077),
    .A2(net2441),
    .B(net3043),
    .Y(_11931_));
 INVx2_ASAP7_75t_R _41010_ (.A(_11364_),
    .Y(_11932_));
 NAND2x2_ASAP7_75t_R _41011_ (.A(_11932_),
    .B(_10547_),
    .Y(_11933_));
 NAND3x1_ASAP7_75t_R _41012_ (.A(_11930_),
    .B(_11931_),
    .C(_11933_),
    .Y(_11934_));
 INVx1_ASAP7_75t_R _41013_ (.A(_11934_),
    .Y(_11935_));
 AND2x2_ASAP7_75t_R _41014_ (.A(_11929_),
    .B(_11935_),
    .Y(_11936_));
 INVx1_ASAP7_75t_R _41015_ (.A(_11936_),
    .Y(_11938_));
 AO21x1_ASAP7_75t_R _41016_ (.A1(net2695),
    .A2(net1855),
    .B(_11355_),
    .Y(_11939_));
 AO21x1_ASAP7_75t_R _41017_ (.A1(_10502_),
    .A2(net3292),
    .B(_11355_),
    .Y(_11940_));
 AO21x1_ASAP7_75t_R _41018_ (.A1(net2841),
    .A2(net1051),
    .B(_11355_),
    .Y(_11941_));
 AND3x1_ASAP7_75t_R _41019_ (.A(_11939_),
    .B(_11940_),
    .C(_11941_),
    .Y(_11942_));
 AO21x1_ASAP7_75t_R _41020_ (.A1(_10449_),
    .A2(net1855),
    .B(_10515_),
    .Y(_11943_));
 AO21x1_ASAP7_75t_R _41021_ (.A1(net2561),
    .A2(net3292),
    .B(_10515_),
    .Y(_11944_));
 NAND2x1_ASAP7_75t_R _41022_ (.A(_10531_),
    .B(_11350_),
    .Y(_11945_));
 AND3x1_ASAP7_75t_R _41023_ (.A(_11943_),
    .B(_11944_),
    .C(_11945_),
    .Y(_11946_));
 AO21x1_ASAP7_75t_R _41024_ (.A1(_10375_),
    .A2(net2332),
    .B(_10515_),
    .Y(_11947_));
 AO21x1_ASAP7_75t_R _41025_ (.A1(net1077),
    .A2(_10410_),
    .B(_10515_),
    .Y(_11949_));
 AND2x2_ASAP7_75t_R _41026_ (.A(_11947_),
    .B(_11949_),
    .Y(_11950_));
 NAND3x1_ASAP7_75t_R _41027_ (.A(_11942_),
    .B(_11946_),
    .C(_11950_),
    .Y(_11951_));
 NOR2x1_ASAP7_75t_R _41028_ (.A(_11938_),
    .B(_11951_),
    .Y(_11952_));
 NAND2x1_ASAP7_75t_R _41029_ (.A(_11923_),
    .B(_11952_),
    .Y(_11953_));
 AO21x2_ASAP7_75t_R _41030_ (.A1(_10382_),
    .A2(_10310_),
    .B(net2187),
    .Y(_11954_));
 AO21x1_ASAP7_75t_R _41031_ (.A1(net3014),
    .A2(net2954),
    .B(net1881),
    .Y(_11955_));
 AO21x1_ASAP7_75t_R _41032_ (.A1(_10370_),
    .A2(net3292),
    .B(net2329),
    .Y(_11956_));
 NAND2x1_ASAP7_75t_R _41033_ (.A(_10350_),
    .B(_10406_),
    .Y(_11957_));
 NAND2x1_ASAP7_75t_R _41034_ (.A(_10406_),
    .B(_10551_),
    .Y(_11958_));
 AND3x1_ASAP7_75t_R _41035_ (.A(_11956_),
    .B(_11957_),
    .C(_11958_),
    .Y(_11960_));
 NAND2x1_ASAP7_75t_R _41036_ (.A(_11955_),
    .B(_11960_),
    .Y(_11961_));
 INVx1_ASAP7_75t_R _41037_ (.A(_11961_),
    .Y(_11962_));
 AO31x2_ASAP7_75t_R _41038_ (.A1(net2955),
    .A2(_10396_),
    .A3(net1114),
    .B(_10336_),
    .Y(_11963_));
 AO21x1_ASAP7_75t_R _41039_ (.A1(net1494),
    .A2(net2851),
    .B(_10336_),
    .Y(_11964_));
 AO21x1_ASAP7_75t_R _41040_ (.A1(net3052),
    .A2(net2354),
    .B(_10336_),
    .Y(_11965_));
 NAND3x1_ASAP7_75t_R _41041_ (.A(_11963_),
    .B(_11964_),
    .C(_11965_),
    .Y(_11966_));
 INVx2_ASAP7_75t_R _41042_ (.A(net2954),
    .Y(_11967_));
 AOI21x1_ASAP7_75t_R _41043_ (.A1(_11967_),
    .A2(_11368_),
    .B(_10376_),
    .Y(_11968_));
 NAND2x1_ASAP7_75t_R _41044_ (.A(_10597_),
    .B(_11368_),
    .Y(_11969_));
 AO21x1_ASAP7_75t_R _41045_ (.A1(_11323_),
    .A2(_10377_),
    .B(_10358_),
    .Y(_11971_));
 NAND3x1_ASAP7_75t_R _41046_ (.A(_11968_),
    .B(_11969_),
    .C(_11971_),
    .Y(_11972_));
 NOR2x1_ASAP7_75t_R _41047_ (.A(_11966_),
    .B(_11972_),
    .Y(_11973_));
 NAND2x2_ASAP7_75t_R _41048_ (.A(_11962_),
    .B(_11973_),
    .Y(_11974_));
 INVx1_ASAP7_75t_R _41049_ (.A(_11974_),
    .Y(_11975_));
 AO21x2_ASAP7_75t_R _41050_ (.A1(_10370_),
    .A2(net3292),
    .B(_10482_),
    .Y(_11976_));
 NAND2x2_ASAP7_75t_R _41051_ (.A(net3319),
    .B(_10483_),
    .Y(_11977_));
 NAND2x2_ASAP7_75t_R _41052_ (.A(net2806),
    .B(_10483_),
    .Y(_11978_));
 NAND3x2_ASAP7_75t_R _41053_ (.B(_11977_),
    .C(_11978_),
    .Y(_11979_),
    .A(_11976_));
 AO31x2_ASAP7_75t_R _41054_ (.A1(net1143),
    .A2(net2442),
    .A3(net2957),
    .B(net2247),
    .Y(_11980_));
 OA21x2_ASAP7_75t_R _41055_ (.A1(_10554_),
    .A2(net3290),
    .B(_11413_),
    .Y(_11982_));
 NOR2x1_ASAP7_75t_R _41056_ (.A(_11412_),
    .B(_11982_),
    .Y(_11983_));
 NAND2x1_ASAP7_75t_R _41057_ (.A(_11980_),
    .B(_11983_),
    .Y(_11984_));
 NOR2x2_ASAP7_75t_R _41058_ (.A(_11979_),
    .B(_11984_),
    .Y(_11985_));
 INVx1_ASAP7_75t_R _41059_ (.A(_11985_),
    .Y(_11986_));
 AO21x1_ASAP7_75t_R _41060_ (.A1(net2562),
    .A2(net2851),
    .B(net1980),
    .Y(_11987_));
 AO21x1_ASAP7_75t_R _41061_ (.A1(_10375_),
    .A2(net2841),
    .B(net1980),
    .Y(_11988_));
 INVx1_ASAP7_75t_R _41062_ (.A(_11467_),
    .Y(_11989_));
 AND4x2_ASAP7_75t_R _41063_ (.A(_11987_),
    .B(_11988_),
    .C(_11464_),
    .D(_11989_),
    .Y(_11990_));
 OAI21x1_ASAP7_75t_R _41064_ (.A1(net1414),
    .A2(net2020),
    .B(_11393_),
    .Y(_11991_));
 AO21x1_ASAP7_75t_R _41065_ (.A1(_10485_),
    .A2(net2333),
    .B(net2464),
    .Y(_11993_));
 INVx1_ASAP7_75t_R _41066_ (.A(_11993_),
    .Y(_11994_));
 AO21x1_ASAP7_75t_R _41067_ (.A1(net2441),
    .A2(net1055),
    .B(_10454_),
    .Y(_11995_));
 OAI21x1_ASAP7_75t_R _41068_ (.A1(net1876),
    .A2(net2020),
    .B(_11995_),
    .Y(_11996_));
 NOR3x2_ASAP7_75t_R _41069_ (.B(_11994_),
    .C(_11996_),
    .Y(_11997_),
    .A(_11991_));
 NAND2x1_ASAP7_75t_R _41070_ (.A(_11990_),
    .B(_11997_),
    .Y(_11998_));
 NOR2x1_ASAP7_75t_R _41071_ (.A(_11986_),
    .B(_11998_),
    .Y(_11999_));
 NAND2x2_ASAP7_75t_R _41072_ (.A(_11975_),
    .B(_11999_),
    .Y(_12000_));
 NOR2x2_ASAP7_75t_R _41073_ (.A(_11953_),
    .B(_12000_),
    .Y(_12001_));
 OAI21x1_ASAP7_75t_R _41074_ (.A1(_11075_),
    .A2(_09825_),
    .B(_09846_),
    .Y(_12002_));
 NOR2x1_ASAP7_75t_R _41075_ (.A(_09649_),
    .B(net1384),
    .Y(_12004_));
 NOR2x1_ASAP7_75t_R _41076_ (.A(_12004_),
    .B(_11703_),
    .Y(_12005_));
 NAND2x1_ASAP7_75t_R _41077_ (.A(_12002_),
    .B(_12005_),
    .Y(_12006_));
 AO21x1_ASAP7_75t_R _41078_ (.A1(_11702_),
    .A2(_09597_),
    .B(_09730_),
    .Y(_12007_));
 NAND2x1_ASAP7_75t_R _41079_ (.A(net2688),
    .B(_11168_),
    .Y(_12008_));
 AO21x1_ASAP7_75t_R _41080_ (.A1(net1562),
    .A2(net1102),
    .B(_09730_),
    .Y(_12009_));
 NAND3x1_ASAP7_75t_R _41081_ (.A(_12007_),
    .B(_12008_),
    .C(_12009_),
    .Y(_12010_));
 NOR2x1_ASAP7_75t_R _41082_ (.A(_12006_),
    .B(_12010_),
    .Y(_12011_));
 AO21x2_ASAP7_75t_R _41083_ (.A1(_09684_),
    .A2(_09798_),
    .B(_09682_),
    .Y(_12012_));
 AO21x2_ASAP7_75t_R _41084_ (.A1(_11161_),
    .A2(_09631_),
    .B(_09682_),
    .Y(_12013_));
 NAND3x2_ASAP7_75t_R _41085_ (.B(_12013_),
    .C(_11151_),
    .Y(_12015_),
    .A(_12012_));
 AO21x1_ASAP7_75t_R _41086_ (.A1(net2503),
    .A2(net2434),
    .B(net2085),
    .Y(_12016_));
 AO21x1_ASAP7_75t_R _41087_ (.A1(net1386),
    .A2(net2939),
    .B(net2085),
    .Y(_12017_));
 NAND2x1_ASAP7_75t_R _41088_ (.A(_12016_),
    .B(_12017_),
    .Y(_12018_));
 AO21x1_ASAP7_75t_R _41089_ (.A1(net2921),
    .A2(_09644_),
    .B(net2085),
    .Y(_12019_));
 AO21x1_ASAP7_75t_R _41090_ (.A1(net3067),
    .A2(_09653_),
    .B(net2085),
    .Y(_12020_));
 NAND2x1_ASAP7_75t_R _41091_ (.A(_12019_),
    .B(_12020_),
    .Y(_12021_));
 NOR3x1_ASAP7_75t_R _41092_ (.A(_12015_),
    .B(_12018_),
    .C(_12021_),
    .Y(_12022_));
 NAND2x1_ASAP7_75t_R _41093_ (.A(_12011_),
    .B(_12022_),
    .Y(_12023_));
 NOR2x1_ASAP7_75t_R _41094_ (.A(net1504),
    .B(net1385),
    .Y(_12024_));
 NOR2x2_ASAP7_75t_R _41095_ (.A(net2103),
    .B(net1504),
    .Y(_12026_));
 AOI211x1_ASAP7_75t_R _41096_ (.A1(_09783_),
    .A2(_09806_),
    .B(_12024_),
    .C(_12026_),
    .Y(_12027_));
 NAND2x2_ASAP7_75t_R _41097_ (.A(_09578_),
    .B(_11688_),
    .Y(_12028_));
 AO21x1_ASAP7_75t_R _41098_ (.A1(_11690_),
    .A2(_09653_),
    .B(net1502),
    .Y(_12029_));
 NAND3x1_ASAP7_75t_R _41099_ (.A(_12027_),
    .B(_12028_),
    .C(_12029_),
    .Y(_12030_));
 NAND2x1_ASAP7_75t_R _41100_ (.A(_11766_),
    .B(_11090_),
    .Y(_12031_));
 NOR2x2_ASAP7_75t_R _41101_ (.A(_09653_),
    .B(net2000),
    .Y(_12032_));
 INVx2_ASAP7_75t_R _41102_ (.A(_12032_),
    .Y(_12033_));
 NAND2x1_ASAP7_75t_R _41103_ (.A(_12031_),
    .B(_12033_),
    .Y(_12034_));
 NOR2x1_ASAP7_75t_R _41104_ (.A(net2001),
    .B(net1924),
    .Y(_12035_));
 OA21x2_ASAP7_75t_R _41105_ (.A1(_11134_),
    .A2(_11167_),
    .B(_11090_),
    .Y(_12037_));
 OR3x1_ASAP7_75t_R _41106_ (.A(_12034_),
    .B(_12035_),
    .C(_12037_),
    .Y(_12038_));
 NOR2x1_ASAP7_75t_R _41107_ (.A(_12030_),
    .B(_12038_),
    .Y(_12039_));
 AO21x1_ASAP7_75t_R _41108_ (.A1(_09817_),
    .A2(_09613_),
    .B(net1871),
    .Y(_12040_));
 AO21x1_ASAP7_75t_R _41109_ (.A1(net1385),
    .A2(net1102),
    .B(net1871),
    .Y(_12041_));
 AND2x2_ASAP7_75t_R _41110_ (.A(_12040_),
    .B(_12041_),
    .Y(_12042_));
 NAND2x1_ASAP7_75t_R _41111_ (.A(_09664_),
    .B(_09759_),
    .Y(_12043_));
 NOR2x1_ASAP7_75t_R _41112_ (.A(net2959),
    .B(net2771),
    .Y(_12044_));
 INVx1_ASAP7_75t_R _41113_ (.A(_12044_),
    .Y(_12045_));
 AND3x1_ASAP7_75t_R _41114_ (.A(_11710_),
    .B(_12043_),
    .C(_12045_),
    .Y(_12046_));
 NAND2x1_ASAP7_75t_R _41115_ (.A(_12042_),
    .B(_12046_),
    .Y(_12048_));
 AO21x2_ASAP7_75t_R _41116_ (.A1(_09714_),
    .A2(net1923),
    .B(net2922),
    .Y(_12049_));
 AO21x1_ASAP7_75t_R _41117_ (.A1(net2828),
    .A2(net1596),
    .B(net1942),
    .Y(_12050_));
 AND2x2_ASAP7_75t_R _41118_ (.A(_12049_),
    .B(_12050_),
    .Y(_12051_));
 AO21x1_ASAP7_75t_R _41119_ (.A1(net1291),
    .A2(_09689_),
    .B(net2922),
    .Y(_12052_));
 NAND2x1_ASAP7_75t_R _41120_ (.A(net3177),
    .B(_09757_),
    .Y(_12053_));
 AO21x1_ASAP7_75t_R _41121_ (.A1(_09658_),
    .A2(_09644_),
    .B(net2924),
    .Y(_12054_));
 AND3x1_ASAP7_75t_R _41122_ (.A(_12052_),
    .B(_12053_),
    .C(_12054_),
    .Y(_12055_));
 NAND2x1_ASAP7_75t_R _41123_ (.A(_12051_),
    .B(_12055_),
    .Y(_12056_));
 NOR2x1_ASAP7_75t_R _41124_ (.A(_12048_),
    .B(_12056_),
    .Y(_12057_));
 NAND2x1_ASAP7_75t_R _41125_ (.A(_12039_),
    .B(_12057_),
    .Y(_12059_));
 NOR2x1_ASAP7_75t_R _41126_ (.A(_12023_),
    .B(_12059_),
    .Y(_12060_));
 AO21x1_ASAP7_75t_R _41127_ (.A1(_11161_),
    .A2(_09689_),
    .B(net2911),
    .Y(_12061_));
 NAND2x1_ASAP7_75t_R _41128_ (.A(_11675_),
    .B(_09826_),
    .Y(_12062_));
 AND2x2_ASAP7_75t_R _41129_ (.A(_12061_),
    .B(_12062_),
    .Y(_12063_));
 AO21x1_ASAP7_75t_R _41130_ (.A1(net1518),
    .A2(net2828),
    .B(net2911),
    .Y(_12064_));
 OA21x2_ASAP7_75t_R _41131_ (.A1(net2046),
    .A2(net2911),
    .B(_12064_),
    .Y(_12065_));
 NAND2x1_ASAP7_75t_R _41132_ (.A(_12063_),
    .B(_12065_),
    .Y(_12066_));
 OA21x2_ASAP7_75t_R _41133_ (.A1(_11675_),
    .A2(_11766_),
    .B(_09701_),
    .Y(_12067_));
 AND3x4_ASAP7_75t_R _41134_ (.A(_09701_),
    .B(_09573_),
    .C(net2152),
    .Y(_12068_));
 NOR2x1_ASAP7_75t_R _41135_ (.A(_12067_),
    .B(_12068_),
    .Y(_12070_));
 NAND2x1_ASAP7_75t_R _41136_ (.A(_09832_),
    .B(_09701_),
    .Y(_12071_));
 NAND3x1_ASAP7_75t_R _41137_ (.A(_12070_),
    .B(_12071_),
    .C(_11144_),
    .Y(_12072_));
 NOR2x1_ASAP7_75t_R _41138_ (.A(_12066_),
    .B(_12072_),
    .Y(_12073_));
 AO21x1_ASAP7_75t_R _41139_ (.A1(_09658_),
    .A2(net2216),
    .B(net2502),
    .Y(_12074_));
 OAI21x1_ASAP7_75t_R _41140_ (.A1(net2502),
    .A2(net1544),
    .B(_12074_),
    .Y(_12075_));
 AO21x1_ASAP7_75t_R _41141_ (.A1(_09714_),
    .A2(_09739_),
    .B(_09655_),
    .Y(_12076_));
 NAND2x1_ASAP7_75t_R _41142_ (.A(_09816_),
    .B(_09661_),
    .Y(_12077_));
 NAND2x2_ASAP7_75t_R _41143_ (.A(_09661_),
    .B(_11069_),
    .Y(_12078_));
 NAND3x1_ASAP7_75t_R _41144_ (.A(_12076_),
    .B(_12077_),
    .C(_12078_),
    .Y(_12079_));
 NOR2x1_ASAP7_75t_R _41145_ (.A(_12075_),
    .B(_12079_),
    .Y(_12081_));
 AO21x1_ASAP7_75t_R _41146_ (.A1(net1518),
    .A2(net1587),
    .B(net2692),
    .Y(_12082_));
 AO21x1_ASAP7_75t_R _41147_ (.A1(net3066),
    .A2(_09597_),
    .B(net2692),
    .Y(_12083_));
 NAND2x1_ASAP7_75t_R _41148_ (.A(_09783_),
    .B(_09696_),
    .Y(_12084_));
 AND3x1_ASAP7_75t_R _41149_ (.A(_12082_),
    .B(_12083_),
    .C(_12084_),
    .Y(_12085_));
 AND2x2_ASAP7_75t_R _41150_ (.A(_12081_),
    .B(_12085_),
    .Y(_12086_));
 NAND2x1_ASAP7_75t_R _41151_ (.A(_12073_),
    .B(_12086_),
    .Y(_12087_));
 AO21x1_ASAP7_75t_R _41152_ (.A1(net1246),
    .A2(net1102),
    .B(_09707_),
    .Y(_12088_));
 NAND2x1_ASAP7_75t_R _41153_ (.A(_09726_),
    .B(_09700_),
    .Y(_12089_));
 NAND2x2_ASAP7_75t_R _41154_ (.A(_09726_),
    .B(_11675_),
    .Y(_12090_));
 AND3x1_ASAP7_75t_R _41155_ (.A(_12088_),
    .B(_12089_),
    .C(_12090_),
    .Y(_12092_));
 NOR2x1_ASAP7_75t_R _41156_ (.A(_09658_),
    .B(net2269),
    .Y(_12093_));
 AND3x2_ASAP7_75t_R _41157_ (.A(_11056_),
    .B(net1930),
    .C(_09780_),
    .Y(_12094_));
 NOR2x1_ASAP7_75t_R _41158_ (.A(_12093_),
    .B(_12094_),
    .Y(_12095_));
 AND2x2_ASAP7_75t_R _41159_ (.A(_12092_),
    .B(_12095_),
    .Y(_12096_));
 AO21x1_ASAP7_75t_R _41160_ (.A1(_09689_),
    .A2(_09653_),
    .B(_09620_),
    .Y(_12097_));
 AO21x1_ASAP7_75t_R _41161_ (.A1(_09858_),
    .A2(_09752_),
    .B(_09620_),
    .Y(_12098_));
 NAND2x1_ASAP7_75t_R _41162_ (.A(_09838_),
    .B(_09809_),
    .Y(_12099_));
 AND3x1_ASAP7_75t_R _41163_ (.A(_12097_),
    .B(_12098_),
    .C(_12099_),
    .Y(_12100_));
 AO21x1_ASAP7_75t_R _41164_ (.A1(net1246),
    .A2(net2828),
    .B(_09594_),
    .Y(_12101_));
 AO21x1_ASAP7_75t_R _41165_ (.A1(net1924),
    .A2(_09739_),
    .B(_09594_),
    .Y(_12103_));
 AND2x2_ASAP7_75t_R _41166_ (.A(_12101_),
    .B(_12103_),
    .Y(_12104_));
 NAND2x2_ASAP7_75t_R _41167_ (.A(net1219),
    .B(net2941),
    .Y(_12105_));
 NAND2x1_ASAP7_75t_R _41168_ (.A(net1219),
    .B(_09809_),
    .Y(_12106_));
 NAND2x1_ASAP7_75t_R _41169_ (.A(net1219),
    .B(_09664_),
    .Y(_12107_));
 AND3x1_ASAP7_75t_R _41170_ (.A(_12105_),
    .B(_12106_),
    .C(_12107_),
    .Y(_12108_));
 AND3x1_ASAP7_75t_R _41171_ (.A(_12100_),
    .B(_12104_),
    .C(_12108_),
    .Y(_12109_));
 NAND2x1_ASAP7_75t_R _41172_ (.A(_12096_),
    .B(_12109_),
    .Y(_12110_));
 NOR2x2_ASAP7_75t_R _41173_ (.A(_12087_),
    .B(_12110_),
    .Y(_12111_));
 NAND2x2_ASAP7_75t_R _41174_ (.A(_12060_),
    .B(_12111_),
    .Y(_12112_));
 NAND2x2_ASAP7_75t_R _41175_ (.A(_12001_),
    .B(_12112_),
    .Y(_12114_));
 NAND3x2_ASAP7_75t_R _41176_ (.B(_11985_),
    .C(_11990_),
    .Y(_12115_),
    .A(_11997_));
 NOR2x2_ASAP7_75t_R _41177_ (.A(_11974_),
    .B(_12115_),
    .Y(_12116_));
 INVx1_ASAP7_75t_R _41178_ (.A(_11906_),
    .Y(_12117_));
 NOR2x1_ASAP7_75t_R _41179_ (.A(_11922_),
    .B(_11913_),
    .Y(_12118_));
 NAND2x1_ASAP7_75t_R _41180_ (.A(_12117_),
    .B(_12118_),
    .Y(_12119_));
 INVx1_ASAP7_75t_R _41181_ (.A(_11942_),
    .Y(_12120_));
 NAND2x1_ASAP7_75t_R _41182_ (.A(_11950_),
    .B(_11946_),
    .Y(_12121_));
 NOR2x1_ASAP7_75t_R _41183_ (.A(_12120_),
    .B(_12121_),
    .Y(_12122_));
 NAND2x1_ASAP7_75t_R _41184_ (.A(_11936_),
    .B(_12122_),
    .Y(_12123_));
 NOR2x1_ASAP7_75t_R _41185_ (.A(_12119_),
    .B(_12123_),
    .Y(_12125_));
 NAND2x2_ASAP7_75t_R _41186_ (.A(_12116_),
    .B(_12125_),
    .Y(_12126_));
 NAND2x1_ASAP7_75t_R _41187_ (.A(_12062_),
    .B(_11710_),
    .Y(_12127_));
 INVx1_ASAP7_75t_R _41188_ (.A(_11144_),
    .Y(_12128_));
 NOR3x1_ASAP7_75t_R _41189_ (.A(_12127_),
    .B(_12128_),
    .C(_11077_),
    .Y(_12129_));
 NAND2x1_ASAP7_75t_R _41190_ (.A(_09624_),
    .B(_09618_),
    .Y(_12130_));
 AO21x1_ASAP7_75t_R _41191_ (.A1(_11161_),
    .A2(_09636_),
    .B(_09730_),
    .Y(_12131_));
 OAI21x1_ASAP7_75t_R _41192_ (.A1(net1102),
    .A2(_12130_),
    .B(_12131_),
    .Y(_12132_));
 NOR3x1_ASAP7_75t_R _41193_ (.A(_12132_),
    .B(_11678_),
    .C(_11703_),
    .Y(_12133_));
 NAND2x1_ASAP7_75t_R _41194_ (.A(_12129_),
    .B(_12133_),
    .Y(_12134_));
 OAI22x1_ASAP7_75t_R _41195_ (.A1(_11097_),
    .A2(_09573_),
    .B1(_11136_),
    .B2(_09589_),
    .Y(_12136_));
 NAND3x1_ASAP7_75t_R _41196_ (.A(_09719_),
    .B(_09758_),
    .C(_09760_),
    .Y(_12137_));
 NOR2x1_ASAP7_75t_R _41197_ (.A(_12136_),
    .B(_12137_),
    .Y(_12138_));
 AO21x1_ASAP7_75t_R _41198_ (.A1(net1544),
    .A2(net2453),
    .B(net3241),
    .Y(_12139_));
 AND4x1_ASAP7_75t_R _41199_ (.A(_09750_),
    .B(_12097_),
    .C(_09740_),
    .D(_12139_),
    .Y(_12140_));
 NAND2x1_ASAP7_75t_R _41200_ (.A(_12138_),
    .B(_12140_),
    .Y(_12141_));
 NOR2x1_ASAP7_75t_R _41201_ (.A(_12134_),
    .B(_12141_),
    .Y(_12142_));
 AO21x1_ASAP7_75t_R _41202_ (.A1(_11766_),
    .A2(_11090_),
    .B(_12026_),
    .Y(_12143_));
 AOI211x1_ASAP7_75t_R _41203_ (.A1(_09838_),
    .A2(_09754_),
    .B(_12143_),
    .C(_12094_),
    .Y(_12144_));
 OR3x1_ASAP7_75t_R _41204_ (.A(net3016),
    .B(_09573_),
    .C(_09635_),
    .Y(_12145_));
 NAND2x1_ASAP7_75t_R _41205_ (.A(_12028_),
    .B(_12145_),
    .Y(_12147_));
 AO21x1_ASAP7_75t_R _41206_ (.A1(_09846_),
    .A2(_09825_),
    .B(_12068_),
    .Y(_12148_));
 NOR2x1_ASAP7_75t_R _41207_ (.A(_12147_),
    .B(_12148_),
    .Y(_12149_));
 NAND2x1_ASAP7_75t_R _41208_ (.A(_12144_),
    .B(_12149_),
    .Y(_12150_));
 NAND2x1_ASAP7_75t_R _41209_ (.A(_12106_),
    .B(_12013_),
    .Y(_12151_));
 AND3x1_ASAP7_75t_R _41210_ (.A(_09759_),
    .B(_09573_),
    .C(_11096_),
    .Y(_12152_));
 OA21x2_ASAP7_75t_R _41211_ (.A1(_09757_),
    .A2(_09661_),
    .B(net2956),
    .Y(_12153_));
 NOR3x1_ASAP7_75t_R _41212_ (.A(_12151_),
    .B(_12152_),
    .C(_12153_),
    .Y(_12154_));
 NOR2x1_ASAP7_75t_R _41213_ (.A(_12044_),
    .B(_12093_),
    .Y(_12155_));
 NAND2x1_ASAP7_75t_R _41214_ (.A(net1220),
    .B(_11128_),
    .Y(_12156_));
 AND4x1_ASAP7_75t_R _41215_ (.A(_12155_),
    .B(_12077_),
    .C(_12156_),
    .D(_12090_),
    .Y(_12158_));
 NAND2x1_ASAP7_75t_R _41216_ (.A(_12154_),
    .B(_12158_),
    .Y(_12159_));
 NOR2x1_ASAP7_75t_R _41217_ (.A(_12150_),
    .B(_12159_),
    .Y(_12160_));
 NAND2x1_ASAP7_75t_R _41218_ (.A(_12142_),
    .B(_12160_),
    .Y(_12161_));
 OA21x2_ASAP7_75t_R _41219_ (.A1(net3016),
    .A2(_09858_),
    .B(_12053_),
    .Y(_12162_));
 AO21x1_ASAP7_75t_R _41220_ (.A1(net1387),
    .A2(_11177_),
    .B(net2607),
    .Y(_12163_));
 NAND3x2_ASAP7_75t_R _41221_ (.B(_12163_),
    .C(_12012_),
    .Y(_12164_),
    .A(_12162_));
 AOI22x1_ASAP7_75t_R _41222_ (.A1(_09701_),
    .A2(net1931),
    .B1(_09726_),
    .B2(_09608_),
    .Y(_12165_));
 OA21x2_ASAP7_75t_R _41223_ (.A1(_12165_),
    .A2(net2554),
    .B(_12082_),
    .Y(_12166_));
 NAND2x1_ASAP7_75t_R _41224_ (.A(net3067),
    .B(net1384),
    .Y(_12167_));
 OA21x2_ASAP7_75t_R _41225_ (.A1(_12167_),
    .A2(_09741_),
    .B(_09807_),
    .Y(_12169_));
 NOR2x1_ASAP7_75t_R _41226_ (.A(_12169_),
    .B(_11727_),
    .Y(_12170_));
 NAND2x1_ASAP7_75t_R _41227_ (.A(_12166_),
    .B(_12170_),
    .Y(_12171_));
 NOR2x2_ASAP7_75t_R _41228_ (.A(_12164_),
    .B(_12171_),
    .Y(_12172_));
 NOR2x1_ASAP7_75t_R _41229_ (.A(net1246),
    .B(net2913),
    .Y(_12173_));
 OR4x2_ASAP7_75t_R _41230_ (.A(_12004_),
    .B(_12173_),
    .C(_12024_),
    .D(_12032_),
    .Y(_12174_));
 NAND2x2_ASAP7_75t_R _41231_ (.A(_11766_),
    .B(_09757_),
    .Y(_12175_));
 NAND3x2_ASAP7_75t_R _41232_ (.B(_12105_),
    .C(_12175_),
    .Y(_12176_),
    .A(_12049_));
 NAND2x2_ASAP7_75t_R _41233_ (.A(_12083_),
    .B(net2926),
    .Y(_12177_));
 NOR3x2_ASAP7_75t_R _41234_ (.B(_12176_),
    .C(_12177_),
    .Y(_12178_),
    .A(_12174_));
 NAND2x1_ASAP7_75t_R _41235_ (.A(_11124_),
    .B(_12078_),
    .Y(_12180_));
 NAND2x1_ASAP7_75t_R _41236_ (.A(_12008_),
    .B(_11758_),
    .Y(_12181_));
 NOR2x1_ASAP7_75t_R _41237_ (.A(_12180_),
    .B(_12181_),
    .Y(_12182_));
 AO21x1_ASAP7_75t_R _41238_ (.A1(_09707_),
    .A2(net2911),
    .B(net1246),
    .Y(_12183_));
 NAND2x1_ASAP7_75t_R _41239_ (.A(_09701_),
    .B(_11766_),
    .Y(_12184_));
 AND3x1_ASAP7_75t_R _41240_ (.A(_12183_),
    .B(_12184_),
    .C(_12107_),
    .Y(_12185_));
 NAND2x1_ASAP7_75t_R _41241_ (.A(_12182_),
    .B(_12185_),
    .Y(_12186_));
 AO21x1_ASAP7_75t_R _41242_ (.A1(_09640_),
    .A2(net2686),
    .B(_11114_),
    .Y(_12187_));
 AO22x1_ASAP7_75t_R _41243_ (.A1(_11090_),
    .A2(_11167_),
    .B1(_11096_),
    .B2(_09807_),
    .Y(_12188_));
 NOR2x1_ASAP7_75t_R _41244_ (.A(_12187_),
    .B(_12188_),
    .Y(_12189_));
 NAND2x1_ASAP7_75t_R _41245_ (.A(_11753_),
    .B(_11067_),
    .Y(_12191_));
 AOI211x1_ASAP7_75t_R _41246_ (.A1(_11111_),
    .A2(_09806_),
    .B(_12191_),
    .C(_11684_),
    .Y(_12192_));
 NAND2x2_ASAP7_75t_R _41247_ (.A(_12189_),
    .B(_12192_),
    .Y(_12193_));
 NOR2x2_ASAP7_75t_R _41248_ (.A(_12186_),
    .B(_12193_),
    .Y(_12194_));
 NAND3x2_ASAP7_75t_R _41249_ (.B(_12178_),
    .C(_12194_),
    .Y(_12195_),
    .A(_12172_));
 NOR2x2_ASAP7_75t_R _41250_ (.A(_12161_),
    .B(_12195_),
    .Y(_12196_));
 NAND2x2_ASAP7_75t_R _41251_ (.A(_12126_),
    .B(_12196_),
    .Y(_12197_));
 NAND2x2_ASAP7_75t_R _41252_ (.A(_12114_),
    .B(_12197_),
    .Y(_12198_));
 AO21x1_ASAP7_75t_R _41253_ (.A1(_10678_),
    .A2(_10767_),
    .B(_10755_),
    .Y(_12199_));
 AO21x1_ASAP7_75t_R _41254_ (.A1(net3049),
    .A2(net3058),
    .B(_10755_),
    .Y(_12200_));
 NOR2x2_ASAP7_75t_R _41255_ (.A(_10710_),
    .B(_10732_),
    .Y(_12202_));
 NAND2x1_ASAP7_75t_R _41256_ (.A(_10754_),
    .B(_12202_),
    .Y(_12203_));
 AND3x1_ASAP7_75t_R _41257_ (.A(_12199_),
    .B(_12200_),
    .C(_12203_),
    .Y(_12204_));
 AO21x1_ASAP7_75t_R _41258_ (.A1(net3048),
    .A2(net3058),
    .B(net3040),
    .Y(_12205_));
 NAND2x1_ASAP7_75t_R _41259_ (.A(_10792_),
    .B(_10774_),
    .Y(_12206_));
 NOR2x1_ASAP7_75t_R _41260_ (.A(_10771_),
    .B(net3040),
    .Y(_12207_));
 INVx1_ASAP7_75t_R _41261_ (.A(_12207_),
    .Y(_12208_));
 INVx1_ASAP7_75t_R _41262_ (.A(_10776_),
    .Y(_12209_));
 AND4x1_ASAP7_75t_R _41263_ (.A(_12205_),
    .B(_12206_),
    .C(_12208_),
    .D(_12209_),
    .Y(_12210_));
 NAND2x1_ASAP7_75t_R _41264_ (.A(_12204_),
    .B(_12210_),
    .Y(_12211_));
 AO21x1_ASAP7_75t_R _41265_ (.A1(_10788_),
    .A2(_10759_),
    .B(_10725_),
    .Y(_12213_));
 NAND2x1_ASAP7_75t_R _41266_ (.A(_10736_),
    .B(_11012_),
    .Y(_12214_));
 AND3x1_ASAP7_75t_R _41267_ (.A(_12213_),
    .B(_10968_),
    .C(_12214_),
    .Y(_12215_));
 OA21x2_ASAP7_75t_R _41268_ (.A1(net3053),
    .A2(_10725_),
    .B(_10962_),
    .Y(_12216_));
 AO21x1_ASAP7_75t_R _41269_ (.A1(_10807_),
    .A2(net3048),
    .B(_10739_),
    .Y(_12217_));
 AO21x1_ASAP7_75t_R _41270_ (.A1(_10771_),
    .A2(_10694_),
    .B(_10739_),
    .Y(_12218_));
 AND2x2_ASAP7_75t_R _41271_ (.A(_12217_),
    .B(_12218_),
    .Y(_12219_));
 NAND3x1_ASAP7_75t_R _41272_ (.A(_12215_),
    .B(_12216_),
    .C(_12219_),
    .Y(_12220_));
 NOR2x1_ASAP7_75t_R _41273_ (.A(_12211_),
    .B(_12220_),
    .Y(_12221_));
 AO21x1_ASAP7_75t_R _41274_ (.A1(_10768_),
    .A2(_10672_),
    .B(net3021),
    .Y(_12222_));
 AO21x1_ASAP7_75t_R _41275_ (.A1(net3053),
    .A2(_10678_),
    .B(net3021),
    .Y(_12224_));
 NAND2x1_ASAP7_75t_R _41276_ (.A(_12222_),
    .B(_12224_),
    .Y(_12225_));
 AO21x1_ASAP7_75t_R _41277_ (.A1(_10656_),
    .A2(net3058),
    .B(_10664_),
    .Y(_12226_));
 OAI21x1_ASAP7_75t_R _41278_ (.A1(_10757_),
    .A2(net3021),
    .B(_12226_),
    .Y(_12227_));
 NOR2x1_ASAP7_75t_R _41279_ (.A(_12225_),
    .B(_12227_),
    .Y(_12228_));
 AO21x1_ASAP7_75t_R _41280_ (.A1(net3023),
    .A2(_10788_),
    .B(_10637_),
    .Y(_12229_));
 AO21x1_ASAP7_75t_R _41281_ (.A1(net2053),
    .A2(_10771_),
    .B(_10637_),
    .Y(_12230_));
 NAND2x1_ASAP7_75t_R _41282_ (.A(_10642_),
    .B(_10869_),
    .Y(_12231_));
 AND4x1_ASAP7_75t_R _41283_ (.A(_12229_),
    .B(_12230_),
    .C(_10638_),
    .D(_12231_),
    .Y(_12232_));
 NAND2x1_ASAP7_75t_R _41284_ (.A(_12228_),
    .B(_12232_),
    .Y(_12233_));
 AO21x1_ASAP7_75t_R _41285_ (.A1(_10783_),
    .A2(net3053),
    .B(_10696_),
    .Y(_12235_));
 AO21x1_ASAP7_75t_R _41286_ (.A1(_10767_),
    .A2(net2053),
    .B(_10696_),
    .Y(_12236_));
 AO21x1_ASAP7_75t_R _41287_ (.A1(_10788_),
    .A2(_11036_),
    .B(_10696_),
    .Y(_12237_));
 AND3x1_ASAP7_75t_R _41288_ (.A(_12235_),
    .B(_12236_),
    .C(_12237_),
    .Y(_12238_));
 AO21x1_ASAP7_75t_R _41289_ (.A1(_10757_),
    .A2(_10807_),
    .B(_10705_),
    .Y(_12239_));
 AO21x1_ASAP7_75t_R _41290_ (.A1(_10938_),
    .A2(_10685_),
    .B(_10705_),
    .Y(_12240_));
 OA211x2_ASAP7_75t_R _41291_ (.A1(net3058),
    .A2(_10705_),
    .B(_12239_),
    .C(_12240_),
    .Y(_12241_));
 NAND2x1_ASAP7_75t_R _41292_ (.A(_12238_),
    .B(_12241_),
    .Y(_12242_));
 NOR2x1_ASAP7_75t_R _41293_ (.A(_12233_),
    .B(_12242_),
    .Y(_12243_));
 NAND2x1_ASAP7_75t_R _41294_ (.A(_12221_),
    .B(_12243_),
    .Y(_12244_));
 AO21x1_ASAP7_75t_R _41295_ (.A1(_10783_),
    .A2(_10771_),
    .B(_10843_),
    .Y(_12246_));
 AO21x1_ASAP7_75t_R _41296_ (.A1(_10700_),
    .A2(_11036_),
    .B(_10843_),
    .Y(_12247_));
 AND3x1_ASAP7_75t_R _41297_ (.A(_12246_),
    .B(_10848_),
    .C(_12247_),
    .Y(_12248_));
 OR3x1_ASAP7_75t_R _41298_ (.A(net3033),
    .B(_10740_),
    .C(_10659_),
    .Y(_12249_));
 AO21x1_ASAP7_75t_R _41299_ (.A1(net2053),
    .A2(_10672_),
    .B(net3033),
    .Y(_12250_));
 AO21x1_ASAP7_75t_R _41300_ (.A1(net3057),
    .A2(_10757_),
    .B(net3033),
    .Y(_12251_));
 AND3x1_ASAP7_75t_R _41301_ (.A(_12249_),
    .B(_12250_),
    .C(_12251_),
    .Y(_12252_));
 NAND2x1_ASAP7_75t_R _41302_ (.A(_12248_),
    .B(_12252_),
    .Y(_12253_));
 AO21x1_ASAP7_75t_R _41303_ (.A1(net2053),
    .A2(net1982),
    .B(net3054),
    .Y(_12254_));
 AO21x1_ASAP7_75t_R _41304_ (.A1(_10678_),
    .A2(_10771_),
    .B(net3054),
    .Y(_12255_));
 NAND2x1_ASAP7_75t_R _41305_ (.A(_10870_),
    .B(_11851_),
    .Y(_12257_));
 AND3x2_ASAP7_75t_R _41306_ (.A(_12254_),
    .B(_12255_),
    .C(_12257_),
    .Y(_12258_));
 AO21x1_ASAP7_75t_R _41307_ (.A1(_10678_),
    .A2(_10771_),
    .B(net3029),
    .Y(_12259_));
 NAND2x1_ASAP7_75t_R _41308_ (.A(_10668_),
    .B(_10627_),
    .Y(_12260_));
 AO21x1_ASAP7_75t_R _41309_ (.A1(_10700_),
    .A2(_12260_),
    .B(net3029),
    .Y(_12261_));
 NAND2x1_ASAP7_75t_R _41310_ (.A(_10669_),
    .B(_10827_),
    .Y(_12262_));
 AND3x2_ASAP7_75t_R _41311_ (.A(_12259_),
    .B(_12261_),
    .C(_12262_),
    .Y(_12263_));
 AO21x1_ASAP7_75t_R _41312_ (.A1(_10832_),
    .A2(net3020),
    .B(net3054),
    .Y(_12264_));
 AO21x1_ASAP7_75t_R _41313_ (.A1(net3057),
    .A2(_10757_),
    .B(net3054),
    .Y(_12265_));
 AND2x2_ASAP7_75t_R _41314_ (.A(_12264_),
    .B(_12265_),
    .Y(_12266_));
 NAND3x2_ASAP7_75t_R _41315_ (.B(_12263_),
    .C(_12266_),
    .Y(_12268_),
    .A(_12258_));
 NOR2x2_ASAP7_75t_R _41316_ (.A(_12253_),
    .B(_12268_),
    .Y(_12269_));
 AO21x1_ASAP7_75t_R _41317_ (.A1(net2053),
    .A2(_11039_),
    .B(net3056),
    .Y(_12270_));
 AO21x1_ASAP7_75t_R _41318_ (.A1(_10757_),
    .A2(_10807_),
    .B(net3056),
    .Y(_12271_));
 AO21x1_ASAP7_75t_R _41319_ (.A1(net3020),
    .A2(net3049),
    .B(net3056),
    .Y(_12272_));
 NAND2x1_ASAP7_75t_R _41320_ (.A(_10996_),
    .B(_10992_),
    .Y(_12273_));
 AND4x1_ASAP7_75t_R _41321_ (.A(_12270_),
    .B(_12271_),
    .C(_12272_),
    .D(_12273_),
    .Y(_12274_));
 OA211x2_ASAP7_75t_R _41322_ (.A1(_10626_),
    .A2(_10658_),
    .B(_10809_),
    .C(net2118),
    .Y(_12275_));
 OA21x2_ASAP7_75t_R _41323_ (.A1(_10967_),
    .A2(_11012_),
    .B(_10809_),
    .Y(_12276_));
 AO21x1_ASAP7_75t_R _41324_ (.A1(_12202_),
    .A2(_10809_),
    .B(_12276_),
    .Y(_12277_));
 NOR2x1_ASAP7_75t_R _41325_ (.A(_12275_),
    .B(_12277_),
    .Y(_12279_));
 NAND2x1_ASAP7_75t_R _41326_ (.A(_12274_),
    .B(_12279_),
    .Y(_12280_));
 AO21x1_ASAP7_75t_R _41327_ (.A1(_10732_),
    .A2(_10656_),
    .B(_10785_),
    .Y(_12281_));
 OA211x2_ASAP7_75t_R _41328_ (.A1(_10785_),
    .A2(_10938_),
    .B(_12281_),
    .C(_11007_),
    .Y(_12282_));
 AO21x1_ASAP7_75t_R _41329_ (.A1(_10807_),
    .A2(_10759_),
    .B(_10796_),
    .Y(_12283_));
 NAND2x1_ASAP7_75t_R _41330_ (.A(_11812_),
    .B(_11833_),
    .Y(_12284_));
 OA211x2_ASAP7_75t_R _41331_ (.A1(_10796_),
    .A2(_10656_),
    .B(_12283_),
    .C(_12284_),
    .Y(_12285_));
 NAND2x1_ASAP7_75t_R _41332_ (.A(_12282_),
    .B(_12285_),
    .Y(_12286_));
 NOR2x1_ASAP7_75t_R _41333_ (.A(_12280_),
    .B(_12286_),
    .Y(_12287_));
 NAND2x2_ASAP7_75t_R _41334_ (.A(_12269_),
    .B(_12287_),
    .Y(_12288_));
 NOR2x2_ASAP7_75t_R _41335_ (.A(_12244_),
    .B(_12288_),
    .Y(_12290_));
 XOR2x2_ASAP7_75t_R _41336_ (.A(_12290_),
    .B(net2515),
    .Y(_12291_));
 XOR2x1_ASAP7_75t_R _41337_ (.A(_12198_),
    .Y(_12292_),
    .B(_12291_));
 XOR2x2_ASAP7_75t_R _41338_ (.A(_11666_),
    .B(net1882),
    .Y(_12293_));
 AO21x1_ASAP7_75t_R _41339_ (.A1(_10008_),
    .A2(net1757),
    .B(net2535),
    .Y(_12294_));
 AO21x1_ASAP7_75t_R _41340_ (.A1(net1660),
    .A2(_09950_),
    .B(net2535),
    .Y(_12295_));
 NAND3x1_ASAP7_75t_R _41341_ (.A(_12294_),
    .B(_12295_),
    .C(_11562_),
    .Y(_12296_));
 NOR3x1_ASAP7_75t_R _41342_ (.A(_10112_),
    .B(_10180_),
    .C(_10261_),
    .Y(_12297_));
 NAND2x1_ASAP7_75t_R _41343_ (.A(_10126_),
    .B(_10114_),
    .Y(_12298_));
 AO21x1_ASAP7_75t_R _41344_ (.A1(_10015_),
    .A2(net2445),
    .B(net2925),
    .Y(_12299_));
 NAND3x1_ASAP7_75t_R _41345_ (.A(_12297_),
    .B(_12298_),
    .C(_12299_),
    .Y(_12300_));
 NOR2x1_ASAP7_75t_R _41346_ (.A(_12296_),
    .B(_12300_),
    .Y(_12301_));
 AO31x2_ASAP7_75t_R _41347_ (.A1(net944),
    .A2(net2235),
    .A3(_10042_),
    .B(net2253),
    .Y(_12302_));
 AO21x1_ASAP7_75t_R _41348_ (.A1(_10008_),
    .A2(net1757),
    .B(net2253),
    .Y(_12303_));
 AO21x1_ASAP7_75t_R _41349_ (.A1(_10107_),
    .A2(_10153_),
    .B(net2253),
    .Y(_12304_));
 NAND3x1_ASAP7_75t_R _41350_ (.A(_12302_),
    .B(_12303_),
    .C(_12304_),
    .Y(_12305_));
 AO21x1_ASAP7_75t_R _41351_ (.A1(_09906_),
    .A2(net2160),
    .B(net2353),
    .Y(_12306_));
 AO21x1_ASAP7_75t_R _41352_ (.A1(_09913_),
    .A2(_10038_),
    .B(net2353),
    .Y(_12307_));
 AND2x2_ASAP7_75t_R _41353_ (.A(_12306_),
    .B(_12307_),
    .Y(_12308_));
 AO21x1_ASAP7_75t_R _41354_ (.A1(_10111_),
    .A2(net1661),
    .B(net3244),
    .Y(_12309_));
 AO21x1_ASAP7_75t_R _41355_ (.A1(net2235),
    .A2(_09882_),
    .B(_10086_),
    .Y(_12311_));
 NAND2x1_ASAP7_75t_R _41356_ (.A(_10140_),
    .B(_10264_),
    .Y(_12312_));
 AND3x1_ASAP7_75t_R _41357_ (.A(_12309_),
    .B(_12311_),
    .C(_12312_),
    .Y(_12313_));
 NAND2x1_ASAP7_75t_R _41358_ (.A(_12308_),
    .B(_12313_),
    .Y(_12314_));
 NOR2x1_ASAP7_75t_R _41359_ (.A(_12305_),
    .B(_12314_),
    .Y(_12315_));
 NAND2x1_ASAP7_75t_R _41360_ (.A(_12301_),
    .B(_12315_),
    .Y(_12316_));
 AO21x1_ASAP7_75t_R _41361_ (.A1(_10008_),
    .A2(_11610_),
    .B(_10060_),
    .Y(_12317_));
 NAND2x2_ASAP7_75t_R _41362_ (.A(_09982_),
    .B(net2805),
    .Y(_12318_));
 NAND3x1_ASAP7_75t_R _41363_ (.A(_12317_),
    .B(_10210_),
    .C(_12318_),
    .Y(_12319_));
 NAND2x1_ASAP7_75t_R _41364_ (.A(_10152_),
    .B(_10157_),
    .Y(_12320_));
 AO21x1_ASAP7_75t_R _41365_ (.A1(net2356),
    .A2(net1757),
    .B(_10048_),
    .Y(_12322_));
 NAND2x1_ASAP7_75t_R _41366_ (.A(_12320_),
    .B(_12322_),
    .Y(_12323_));
 NAND2x1_ASAP7_75t_R _41367_ (.A(net1250),
    .B(_10157_),
    .Y(_12324_));
 NAND2x1_ASAP7_75t_R _41368_ (.A(_12324_),
    .B(_10052_),
    .Y(_12325_));
 NOR3x1_ASAP7_75t_R _41369_ (.A(_12319_),
    .B(_12323_),
    .C(_12325_),
    .Y(_12326_));
 AO21x1_ASAP7_75t_R _41370_ (.A1(_09895_),
    .A2(_09882_),
    .B(_10035_),
    .Y(_12327_));
 AO21x1_ASAP7_75t_R _41371_ (.A1(_10289_),
    .A2(_10153_),
    .B(_10035_),
    .Y(_12328_));
 NAND2x1_ASAP7_75t_R _41372_ (.A(_12327_),
    .B(_12328_),
    .Y(_12329_));
 AOI211x1_ASAP7_75t_R _41373_ (.A1(net1024),
    .A2(_09892_),
    .B(_10040_),
    .C(net1703),
    .Y(_12330_));
 NOR2x1_ASAP7_75t_R _41374_ (.A(_10040_),
    .B(net2445),
    .Y(_12331_));
 AOI211x1_ASAP7_75t_R _41375_ (.A1(_10077_),
    .A2(_10044_),
    .B(_12330_),
    .C(_12331_),
    .Y(_12333_));
 AO21x1_ASAP7_75t_R _41376_ (.A1(_10063_),
    .A2(net1661),
    .B(_10040_),
    .Y(_12334_));
 AO21x1_ASAP7_75t_R _41377_ (.A1(net2235),
    .A2(_09882_),
    .B(_10040_),
    .Y(_12335_));
 NAND2x1_ASAP7_75t_R _41378_ (.A(_10044_),
    .B(_09970_),
    .Y(_12336_));
 AND3x1_ASAP7_75t_R _41379_ (.A(_12334_),
    .B(_12335_),
    .C(_12336_),
    .Y(_12337_));
 NAND2x1_ASAP7_75t_R _41380_ (.A(_12333_),
    .B(_12337_),
    .Y(_12338_));
 NOR2x1_ASAP7_75t_R _41381_ (.A(_12329_),
    .B(_12338_),
    .Y(_12339_));
 NAND2x1_ASAP7_75t_R _41382_ (.A(_12326_),
    .B(_12339_),
    .Y(_12340_));
 NOR2x1_ASAP7_75t_R _41383_ (.A(_12340_),
    .B(_12316_),
    .Y(_12341_));
 AO21x1_ASAP7_75t_R _41384_ (.A1(_10063_),
    .A2(_09895_),
    .B(_09937_),
    .Y(_12342_));
 AND2x2_ASAP7_75t_R _41385_ (.A(_12342_),
    .B(_11573_),
    .Y(_12344_));
 AO21x1_ASAP7_75t_R _41386_ (.A1(_09913_),
    .A2(net2356),
    .B(_09937_),
    .Y(_12345_));
 OA21x2_ASAP7_75t_R _41387_ (.A1(net2444),
    .A2(_09937_),
    .B(_12345_),
    .Y(_12346_));
 NAND2x1_ASAP7_75t_R _41388_ (.A(_12344_),
    .B(_12346_),
    .Y(_12347_));
 NAND2x1_ASAP7_75t_R _41389_ (.A(net2382),
    .B(_11212_),
    .Y(_12348_));
 AND2x2_ASAP7_75t_R _41390_ (.A(_11231_),
    .B(_12348_),
    .Y(_12349_));
 AO21x2_ASAP7_75t_R _41391_ (.A1(net945),
    .A2(_09919_),
    .B(_09953_),
    .Y(_12350_));
 AO21x1_ASAP7_75t_R _41392_ (.A1(_09928_),
    .A2(_09950_),
    .B(_09953_),
    .Y(_12351_));
 NAND3x1_ASAP7_75t_R _41393_ (.A(_12349_),
    .B(_12350_),
    .C(_12351_),
    .Y(_12352_));
 NOR2x1_ASAP7_75t_R _41394_ (.A(_12347_),
    .B(_12352_),
    .Y(_12353_));
 AO21x1_ASAP7_75t_R _41395_ (.A1(_09998_),
    .A2(net2734),
    .B(_09901_),
    .Y(_12355_));
 AND2x2_ASAP7_75t_R _41396_ (.A(_12355_),
    .B(_11242_),
    .Y(_12356_));
 AO21x1_ASAP7_75t_R _41397_ (.A1(_09988_),
    .A2(net2444),
    .B(_09901_),
    .Y(_12357_));
 NAND3x1_ASAP7_75t_R _41398_ (.A(_12356_),
    .B(_10225_),
    .C(_12357_),
    .Y(_12358_));
 AO21x1_ASAP7_75t_R _41399_ (.A1(net2397),
    .A2(net2235),
    .B(net2660),
    .Y(_12359_));
 OA21x2_ASAP7_75t_R _41400_ (.A1(net943),
    .A2(net2660),
    .B(_12359_),
    .Y(_12360_));
 AO21x1_ASAP7_75t_R _41401_ (.A1(net2160),
    .A2(net2444),
    .B(net2660),
    .Y(_12361_));
 NAND2x1_ASAP7_75t_R _41402_ (.A(_10027_),
    .B(_10133_),
    .Y(_12362_));
 AND3x1_ASAP7_75t_R _41403_ (.A(_12361_),
    .B(_12362_),
    .C(_11224_),
    .Y(_12363_));
 NAND2x1_ASAP7_75t_R _41404_ (.A(_12360_),
    .B(_12363_),
    .Y(_12364_));
 NOR2x1_ASAP7_75t_R _41405_ (.A(_12358_),
    .B(_12364_),
    .Y(_12366_));
 NAND2x1_ASAP7_75t_R _41406_ (.A(_12353_),
    .B(_12366_),
    .Y(_12367_));
 NAND2x2_ASAP7_75t_R _41407_ (.A(_10255_),
    .B(_10264_),
    .Y(_12368_));
 INVx2_ASAP7_75t_R _41408_ (.A(_12368_),
    .Y(_12369_));
 NOR2x1_ASAP7_75t_R _41409_ (.A(_12369_),
    .B(_10257_),
    .Y(_12370_));
 AO21x1_ASAP7_75t_R _41410_ (.A1(net2358),
    .A2(_10008_),
    .B(_10011_),
    .Y(_12371_));
 NAND2x2_ASAP7_75t_R _41411_ (.A(_10255_),
    .B(net2772),
    .Y(_12372_));
 AND3x1_ASAP7_75t_R _41412_ (.A(_12370_),
    .B(_12371_),
    .C(_12372_),
    .Y(_12373_));
 OA21x2_ASAP7_75t_R _41413_ (.A1(_10264_),
    .A2(net2627),
    .B(net1890),
    .Y(_12374_));
 AOI211x1_ASAP7_75t_R _41414_ (.A1(_10143_),
    .A2(net1890),
    .B(_12374_),
    .C(_10292_),
    .Y(_12375_));
 AO21x1_ASAP7_75t_R _41415_ (.A1(_10008_),
    .A2(net1757),
    .B(_09990_),
    .Y(_12377_));
 NAND2x1_ASAP7_75t_R _41416_ (.A(net1800),
    .B(net1029),
    .Y(_12378_));
 AO21x1_ASAP7_75t_R _41417_ (.A1(_12378_),
    .A2(net1757),
    .B(_10246_),
    .Y(_12379_));
 NAND2x1_ASAP7_75t_R _41418_ (.A(_09992_),
    .B(_10264_),
    .Y(_12380_));
 AND3x1_ASAP7_75t_R _41419_ (.A(_12377_),
    .B(_12379_),
    .C(_12380_),
    .Y(_12381_));
 NAND3x1_ASAP7_75t_R _41420_ (.A(_12373_),
    .B(_12375_),
    .C(_12381_),
    .Y(_12382_));
 NOR2x1_ASAP7_75t_R _41421_ (.A(_12367_),
    .B(_12382_),
    .Y(_12383_));
 NAND2x2_ASAP7_75t_R _41422_ (.A(_12341_),
    .B(_12383_),
    .Y(_12384_));
 XOR2x1_ASAP7_75t_R _41423_ (.A(_12293_),
    .Y(_12385_),
    .B(_12384_));
 NAND2x1_ASAP7_75t_R _41424_ (.A(_12292_),
    .B(_12385_),
    .Y(_12386_));
 XNOR2x2_ASAP7_75t_R _41425_ (.A(_10877_),
    .B(_12290_),
    .Y(_12388_));
 XOR2x1_ASAP7_75t_R _41426_ (.A(_12198_),
    .Y(_12389_),
    .B(_12388_));
 XOR2x2_ASAP7_75t_R _41427_ (.A(_11666_),
    .B(_10883_),
    .Y(_12390_));
 XOR2x1_ASAP7_75t_R _41428_ (.A(_12390_),
    .Y(_12391_),
    .B(_12384_));
 NAND2x1_ASAP7_75t_R _41429_ (.A(_12389_),
    .B(_12391_),
    .Y(_12392_));
 AOI21x1_ASAP7_75t_R _41430_ (.A1(_12386_),
    .A2(_12392_),
    .B(net389),
    .Y(_12393_));
 INVx1_ASAP7_75t_R _41431_ (.A(_00523_),
    .Y(_12394_));
 OAI21x1_ASAP7_75t_R _41432_ (.A1(_11896_),
    .A2(_12393_),
    .B(_12394_),
    .Y(_12395_));
 NOR2x1_ASAP7_75t_R _41433_ (.A(net393),
    .B(_00816_),
    .Y(_12396_));
 NAND2x1_ASAP7_75t_R _41434_ (.A(_12292_),
    .B(_12391_),
    .Y(_12397_));
 NAND2x1_ASAP7_75t_R _41435_ (.A(_12389_),
    .B(_12385_),
    .Y(_12399_));
 AOI21x1_ASAP7_75t_R _41436_ (.A1(_12397_),
    .A2(_12399_),
    .B(net389),
    .Y(_12400_));
 OAI21x1_ASAP7_75t_R _41437_ (.A1(_12396_),
    .A2(_12400_),
    .B(_00523_),
    .Y(_12401_));
 NAND2x1_ASAP7_75t_R _41438_ (.A(_12401_),
    .B(_12395_),
    .Y(_00100_));
 OR2x2_ASAP7_75t_R _41439_ (.A(net392),
    .B(_00815_),
    .Y(_12402_));
 XOR2x1_ASAP7_75t_R _41440_ (.A(_12384_),
    .Y(_12403_),
    .B(_10883_));
 AO21x1_ASAP7_75t_R _41441_ (.A1(net2356),
    .A2(_10085_),
    .B(_09901_),
    .Y(_12404_));
 AO21x1_ASAP7_75t_R _41442_ (.A1(net2235),
    .A2(_10042_),
    .B(_09901_),
    .Y(_12405_));
 NAND2x1_ASAP7_75t_R _41443_ (.A(_10014_),
    .B(_09876_),
    .Y(_12406_));
 AND3x1_ASAP7_75t_R _41444_ (.A(_12404_),
    .B(_12405_),
    .C(_12406_),
    .Y(_12407_));
 NOR2x1_ASAP7_75t_R _41445_ (.A(_10008_),
    .B(_09922_),
    .Y(_12409_));
 NOR2x1_ASAP7_75t_R _41446_ (.A(_09913_),
    .B(net2559),
    .Y(_12410_));
 NOR2x1_ASAP7_75t_R _41447_ (.A(_09908_),
    .B(net2559),
    .Y(_12411_));
 OR3x1_ASAP7_75t_R _41448_ (.A(_12409_),
    .B(_12410_),
    .C(_12411_),
    .Y(_12412_));
 NOR2x1_ASAP7_75t_R _41449_ (.A(_12412_),
    .B(_11223_),
    .Y(_12413_));
 NAND2x1_ASAP7_75t_R _41450_ (.A(_12407_),
    .B(_12413_),
    .Y(_12414_));
 AO21x1_ASAP7_75t_R _41451_ (.A1(_10038_),
    .A2(_10085_),
    .B(_09937_),
    .Y(_12415_));
 NAND2x1_ASAP7_75t_R _41452_ (.A(_10278_),
    .B(_12415_),
    .Y(_12416_));
 NOR3x1_ASAP7_75t_R _41453_ (.A(_12416_),
    .B(_09948_),
    .C(_09938_),
    .Y(_12417_));
 AO21x1_ASAP7_75t_R _41454_ (.A1(_10059_),
    .A2(_09913_),
    .B(_09953_),
    .Y(_12418_));
 AO21x1_ASAP7_75t_R _41455_ (.A1(net2235),
    .A2(_10003_),
    .B(_09953_),
    .Y(_12420_));
 AND3x1_ASAP7_75t_R _41456_ (.A(_12418_),
    .B(_12350_),
    .C(_12420_),
    .Y(_12421_));
 NAND2x1_ASAP7_75t_R _41457_ (.A(_12417_),
    .B(_12421_),
    .Y(_12422_));
 NOR2x1_ASAP7_75t_R _41458_ (.A(_12414_),
    .B(_12422_),
    .Y(_12423_));
 AOI211x1_ASAP7_75t_R _41459_ (.A1(net3015),
    .A2(net1159),
    .B(_09990_),
    .C(net1703),
    .Y(_12424_));
 INVx1_ASAP7_75t_R _41460_ (.A(_12424_),
    .Y(_12425_));
 NAND2x1_ASAP7_75t_R _41461_ (.A(_09981_),
    .B(_09992_),
    .Y(_12426_));
 AO21x1_ASAP7_75t_R _41462_ (.A1(net2235),
    .A2(net3245),
    .B(_09990_),
    .Y(_12427_));
 AND3x1_ASAP7_75t_R _41463_ (.A(_12425_),
    .B(_12426_),
    .C(_12427_),
    .Y(_12428_));
 AO21x1_ASAP7_75t_R _41464_ (.A1(_10063_),
    .A2(net1661),
    .B(_10246_),
    .Y(_12429_));
 INVx1_ASAP7_75t_R _41465_ (.A(_11593_),
    .Y(_12431_));
 NAND2x1_ASAP7_75t_R _41466_ (.A(_09979_),
    .B(_09974_),
    .Y(_12432_));
 AND4x1_ASAP7_75t_R _41467_ (.A(_12429_),
    .B(_11201_),
    .C(_12431_),
    .D(_12432_),
    .Y(_12433_));
 NAND2x1_ASAP7_75t_R _41468_ (.A(_12428_),
    .B(_12433_),
    .Y(_12434_));
 AO21x1_ASAP7_75t_R _41469_ (.A1(net1961),
    .A2(_09963_),
    .B(_10005_),
    .Y(_12435_));
 AO21x1_ASAP7_75t_R _41470_ (.A1(_10063_),
    .A2(_10207_),
    .B(_10005_),
    .Y(_12436_));
 NAND2x1_ASAP7_75t_R _41471_ (.A(net1890),
    .B(_10126_),
    .Y(_12437_));
 AND3x1_ASAP7_75t_R _41472_ (.A(_12435_),
    .B(_12436_),
    .C(_12437_),
    .Y(_12438_));
 NAND2x1_ASAP7_75t_R _41473_ (.A(_10255_),
    .B(net2575),
    .Y(_12439_));
 NOR2x1_ASAP7_75t_R _41474_ (.A(_09908_),
    .B(_10011_),
    .Y(_12440_));
 INVx1_ASAP7_75t_R _41475_ (.A(_12440_),
    .Y(_12442_));
 AND3x1_ASAP7_75t_R _41476_ (.A(_12371_),
    .B(_12439_),
    .C(_12442_),
    .Y(_12443_));
 NAND2x1_ASAP7_75t_R _41477_ (.A(_10255_),
    .B(_10161_),
    .Y(_12444_));
 AND3x1_ASAP7_75t_R _41478_ (.A(_11638_),
    .B(_12368_),
    .C(_12444_),
    .Y(_12445_));
 NAND3x1_ASAP7_75t_R _41479_ (.A(_12438_),
    .B(_12443_),
    .C(_12445_),
    .Y(_12446_));
 NOR2x1_ASAP7_75t_R _41480_ (.A(_12434_),
    .B(_12446_),
    .Y(_12447_));
 NAND2x1_ASAP7_75t_R _41481_ (.A(_12423_),
    .B(_12447_),
    .Y(_12448_));
 AO21x1_ASAP7_75t_R _41482_ (.A1(_09913_),
    .A2(net2444),
    .B(_10048_),
    .Y(_12449_));
 AO21x1_ASAP7_75t_R _41483_ (.A1(net2213),
    .A2(net1661),
    .B(_10048_),
    .Y(_12450_));
 NAND2x1_ASAP7_75t_R _41484_ (.A(_10157_),
    .B(_11627_),
    .Y(_12451_));
 AND3x1_ASAP7_75t_R _41485_ (.A(_12449_),
    .B(_12450_),
    .C(_12451_),
    .Y(_12453_));
 INVx1_ASAP7_75t_R _41486_ (.A(_11266_),
    .Y(_12454_));
 AND3x1_ASAP7_75t_R _41487_ (.A(_10210_),
    .B(_10211_),
    .C(_12318_),
    .Y(_12455_));
 NAND3x1_ASAP7_75t_R _41488_ (.A(_12453_),
    .B(_12454_),
    .C(_12455_),
    .Y(_12456_));
 AO21x1_ASAP7_75t_R _41489_ (.A1(net946),
    .A2(_09895_),
    .B(_10040_),
    .Y(_12457_));
 AO21x1_ASAP7_75t_R _41490_ (.A1(net2160),
    .A2(net2357),
    .B(net2662),
    .Y(_12458_));
 AND3x1_ASAP7_75t_R _41491_ (.A(_12457_),
    .B(_12458_),
    .C(_12336_),
    .Y(_12459_));
 OA211x2_ASAP7_75t_R _41492_ (.A1(_10035_),
    .A2(_11604_),
    .B(_10209_),
    .C(_11617_),
    .Y(_12460_));
 NAND2x1_ASAP7_75t_R _41493_ (.A(_12459_),
    .B(_12460_),
    .Y(_12461_));
 NOR2x1_ASAP7_75t_R _41494_ (.A(_12456_),
    .B(_12461_),
    .Y(_12462_));
 AO21x1_ASAP7_75t_R _41495_ (.A1(_09895_),
    .A2(net1660),
    .B(net2535),
    .Y(_12464_));
 NAND2x1_ASAP7_75t_R _41496_ (.A(_09981_),
    .B(_10099_),
    .Y(_12465_));
 AND3x1_ASAP7_75t_R _41497_ (.A(_12464_),
    .B(_11653_),
    .C(_12465_),
    .Y(_12466_));
 AO21x1_ASAP7_75t_R _41498_ (.A1(_10107_),
    .A2(net2808),
    .B(net2535),
    .Y(_12467_));
 NAND2x2_ASAP7_75t_R _41499_ (.A(net2583),
    .B(_10099_),
    .Y(_12468_));
 AND3x2_ASAP7_75t_R _41500_ (.A(_12467_),
    .B(_10277_),
    .C(_12468_),
    .Y(_12469_));
 NAND2x2_ASAP7_75t_R _41501_ (.A(_12466_),
    .B(_12469_),
    .Y(_12470_));
 NAND2x1_ASAP7_75t_R _41502_ (.A(_10126_),
    .B(_10071_),
    .Y(_12471_));
 AND3x1_ASAP7_75t_R _41503_ (.A(_10075_),
    .B(_12471_),
    .C(_10073_),
    .Y(_12472_));
 AO21x1_ASAP7_75t_R _41504_ (.A1(net2808),
    .A2(_10153_),
    .B(net2353),
    .Y(_12473_));
 AO21x1_ASAP7_75t_R _41505_ (.A1(net2358),
    .A2(net1757),
    .B(net3244),
    .Y(_12475_));
 AO21x1_ASAP7_75t_R _41506_ (.A1(_10111_),
    .A2(_10137_),
    .B(net3244),
    .Y(_12476_));
 AND3x1_ASAP7_75t_R _41507_ (.A(_12473_),
    .B(_12475_),
    .C(_12476_),
    .Y(_12477_));
 NAND2x2_ASAP7_75t_R _41508_ (.A(_12472_),
    .B(_12477_),
    .Y(_12478_));
 NAND2x1_ASAP7_75t_R _41509_ (.A(_10014_),
    .B(_10114_),
    .Y(_12479_));
 NAND2x2_ASAP7_75t_R _41510_ (.A(net2583),
    .B(_10114_),
    .Y(_12480_));
 AND3x1_ASAP7_75t_R _41511_ (.A(_12479_),
    .B(_12480_),
    .C(_12298_),
    .Y(_12481_));
 NAND2x2_ASAP7_75t_R _41512_ (.A(_11588_),
    .B(_12481_),
    .Y(_12482_));
 NOR3x2_ASAP7_75t_R _41513_ (.B(_12478_),
    .C(_12482_),
    .Y(_12483_),
    .A(_12470_));
 NAND2x2_ASAP7_75t_R _41514_ (.A(_12462_),
    .B(_12483_),
    .Y(_12484_));
 NOR2x2_ASAP7_75t_R _41515_ (.A(_12448_),
    .B(_12484_),
    .Y(_12486_));
 AO21x1_ASAP7_75t_R _41516_ (.A1(net1387),
    .A2(net2434),
    .B(net2912),
    .Y(_12487_));
 OA21x2_ASAP7_75t_R _41517_ (.A1(_11708_),
    .A2(_11075_),
    .B(_11168_),
    .Y(_12488_));
 INVx1_ASAP7_75t_R _41518_ (.A(_12488_),
    .Y(_12489_));
 NAND2x1_ASAP7_75t_R _41519_ (.A(_12487_),
    .B(_12489_),
    .Y(_12490_));
 NAND3x2_ASAP7_75t_R _41520_ (.B(_09650_),
    .C(_11124_),
    .Y(_12491_),
    .A(_11087_));
 NOR2x2_ASAP7_75t_R _41521_ (.A(_12490_),
    .B(_12491_),
    .Y(_12492_));
 AO21x1_ASAP7_75t_R _41522_ (.A1(net1246),
    .A2(net2732),
    .B(net2085),
    .Y(_12493_));
 AO21x1_ASAP7_75t_R _41523_ (.A1(_11161_),
    .A2(net1292),
    .B(net2085),
    .Y(_12494_));
 NOR2x1_ASAP7_75t_R _41524_ (.A(net2340),
    .B(net2921),
    .Y(_12495_));
 INVx1_ASAP7_75t_R _41525_ (.A(_12495_),
    .Y(_12497_));
 NAND3x1_ASAP7_75t_R _41526_ (.A(_12493_),
    .B(_12494_),
    .C(_12497_),
    .Y(_12498_));
 NAND2x1_ASAP7_75t_R _41527_ (.A(_09640_),
    .B(_11134_),
    .Y(_12499_));
 AO21x1_ASAP7_75t_R _41528_ (.A1(net2732),
    .A2(net2503),
    .B(_09682_),
    .Y(_12500_));
 NAND3x1_ASAP7_75t_R _41529_ (.A(_09641_),
    .B(_12499_),
    .C(_12500_),
    .Y(_12501_));
 NOR2x1_ASAP7_75t_R _41530_ (.A(_12498_),
    .B(_12501_),
    .Y(_12502_));
 NAND2x2_ASAP7_75t_R _41531_ (.A(_12492_),
    .B(_12502_),
    .Y(_12503_));
 AO21x1_ASAP7_75t_R _41532_ (.A1(_11128_),
    .A2(_09806_),
    .B(_12024_),
    .Y(_12504_));
 NOR3x2_ASAP7_75t_R _41533_ (.B(_12504_),
    .C(_12026_),
    .Y(_12505_),
    .A(net3242));
 AO21x1_ASAP7_75t_R _41534_ (.A1(net2732),
    .A2(net2103),
    .B(net2001),
    .Y(_12506_));
 AO21x1_ASAP7_75t_R _41535_ (.A1(net1544),
    .A2(net1577),
    .B(net2001),
    .Y(_12508_));
 NAND2x1_ASAP7_75t_R _41536_ (.A(_11128_),
    .B(_11090_),
    .Y(_12509_));
 AND4x1_ASAP7_75t_R _41537_ (.A(_12506_),
    .B(_12508_),
    .C(_12509_),
    .D(_12031_),
    .Y(_12510_));
 NAND2x2_ASAP7_75t_R _41538_ (.A(_12505_),
    .B(_12510_),
    .Y(_12511_));
 OAI21x1_ASAP7_75t_R _41539_ (.A1(net1942),
    .A2(_09812_),
    .B(_12052_),
    .Y(_12512_));
 AO21x1_ASAP7_75t_R _41540_ (.A1(net1291),
    .A2(_09597_),
    .B(net1871),
    .Y(_12513_));
 OAI21x1_ASAP7_75t_R _41541_ (.A1(net1872),
    .A2(net1385),
    .B(_12513_),
    .Y(_12514_));
 AO21x1_ASAP7_75t_R _41542_ (.A1(net1246),
    .A2(net3243),
    .B(net2922),
    .Y(_12515_));
 AO21x1_ASAP7_75t_R _41543_ (.A1(net2503),
    .A2(_09613_),
    .B(net2923),
    .Y(_12516_));
 NAND2x1_ASAP7_75t_R _41544_ (.A(_12515_),
    .B(_12516_),
    .Y(_12517_));
 OR3x4_ASAP7_75t_R _41545_ (.A(_12512_),
    .B(_12514_),
    .C(_12517_),
    .Y(_12519_));
 NOR3x2_ASAP7_75t_R _41546_ (.B(_12511_),
    .C(_12519_),
    .Y(_12520_),
    .A(_12503_));
 INVx2_ASAP7_75t_R _41547_ (.A(_11708_),
    .Y(_12521_));
 AO21x1_ASAP7_75t_R _41548_ (.A1(_12521_),
    .A2(_09689_),
    .B(net2917),
    .Y(_12522_));
 NOR2x1_ASAP7_75t_R _41549_ (.A(net1385),
    .B(net2917),
    .Y(_12523_));
 INVx1_ASAP7_75t_R _41550_ (.A(_12523_),
    .Y(_12524_));
 NAND3x1_ASAP7_75t_R _41551_ (.A(_12522_),
    .B(_09614_),
    .C(_12524_),
    .Y(_12525_));
 AO21x1_ASAP7_75t_R _41552_ (.A1(_09752_),
    .A2(net1587),
    .B(net2290),
    .Y(_12526_));
 AND2x2_ASAP7_75t_R _41553_ (.A(_12526_),
    .B(_11732_),
    .Y(_12527_));
 AO21x1_ASAP7_75t_R _41554_ (.A1(_09658_),
    .A2(net2217),
    .B(net2290),
    .Y(_12528_));
 OA21x2_ASAP7_75t_R _41555_ (.A1(net2290),
    .A2(net1544),
    .B(_12528_),
    .Y(_12530_));
 NAND2x1_ASAP7_75t_R _41556_ (.A(_12527_),
    .B(_12530_),
    .Y(_12531_));
 NOR2x1_ASAP7_75t_R _41557_ (.A(_12525_),
    .B(_12531_),
    .Y(_12532_));
 NAND2x1_ASAP7_75t_R _41558_ (.A(net2152),
    .B(_09726_),
    .Y(_12533_));
 OAI21x1_ASAP7_75t_R _41559_ (.A1(_09781_),
    .A2(_12533_),
    .B(_09727_),
    .Y(_12534_));
 INVx1_ASAP7_75t_R _41560_ (.A(_09716_),
    .Y(_12535_));
 NOR3x1_ASAP7_75t_R _41561_ (.A(_12534_),
    .B(_12535_),
    .C(_11693_),
    .Y(_12536_));
 OA21x2_ASAP7_75t_R _41562_ (.A1(_11766_),
    .A2(net2919),
    .B(_11056_),
    .Y(_12537_));
 OA21x2_ASAP7_75t_R _41563_ (.A1(_09832_),
    .A2(_11167_),
    .B(_11056_),
    .Y(_12538_));
 AOI211x1_ASAP7_75t_R _41564_ (.A1(_11134_),
    .A2(_11056_),
    .B(_12537_),
    .C(_12538_),
    .Y(_12539_));
 AND2x2_ASAP7_75t_R _41565_ (.A(_12536_),
    .B(_12539_),
    .Y(_12541_));
 NAND2x1_ASAP7_75t_R _41566_ (.A(_12532_),
    .B(_12541_),
    .Y(_12542_));
 AO21x1_ASAP7_75t_R _41567_ (.A1(net1246),
    .A2(net2937),
    .B(net1743),
    .Y(_12543_));
 AO21x1_ASAP7_75t_R _41568_ (.A1(net1577),
    .A2(net2453),
    .B(net1743),
    .Y(_12544_));
 NAND3x2_ASAP7_75t_R _41569_ (.B(_12544_),
    .C(_11123_),
    .Y(_12545_),
    .A(_12543_));
 NAND2x2_ASAP7_75t_R _41570_ (.A(_11179_),
    .B(_09656_),
    .Y(_12546_));
 AO21x1_ASAP7_75t_R _41571_ (.A1(net2434),
    .A2(_11165_),
    .B(net2501),
    .Y(_12547_));
 INVx1_ASAP7_75t_R _41572_ (.A(_12547_),
    .Y(_12548_));
 NOR3x2_ASAP7_75t_R _41573_ (.B(_12546_),
    .C(_12548_),
    .Y(_12549_),
    .A(_12545_));
 AO21x1_ASAP7_75t_R _41574_ (.A1(_09752_),
    .A2(net2937),
    .B(net2605),
    .Y(_12550_));
 OAI21x1_ASAP7_75t_R _41575_ (.A1(_09817_),
    .A2(net2606),
    .B(_12550_),
    .Y(_12552_));
 AO21x1_ASAP7_75t_R _41576_ (.A1(_11690_),
    .A2(_11161_),
    .B(net2605),
    .Y(_12553_));
 OAI21x1_ASAP7_75t_R _41577_ (.A1(_09597_),
    .A2(net2605),
    .B(_12553_),
    .Y(_12554_));
 NOR2x1_ASAP7_75t_R _41578_ (.A(_12552_),
    .B(_12554_),
    .Y(_12555_));
 INVx1_ASAP7_75t_R _41579_ (.A(_12555_),
    .Y(_12556_));
 AO21x1_ASAP7_75t_R _41580_ (.A1(_09817_),
    .A2(_09739_),
    .B(_09672_),
    .Y(_12557_));
 OA21x2_ASAP7_75t_R _41581_ (.A1(net1387),
    .A2(_09672_),
    .B(_12557_),
    .Y(_12558_));
 OA21x2_ASAP7_75t_R _41582_ (.A1(_09809_),
    .A2(_11675_),
    .B(_09701_),
    .Y(_12559_));
 NOR3x2_ASAP7_75t_R _41583_ (.B(_12559_),
    .C(_11129_),
    .Y(_12560_),
    .A(_12068_));
 NAND2x1_ASAP7_75t_R _41584_ (.A(_12558_),
    .B(_12560_),
    .Y(_12561_));
 NOR2x1_ASAP7_75t_R _41585_ (.A(_12556_),
    .B(_12561_),
    .Y(_12563_));
 NAND2x1_ASAP7_75t_R _41586_ (.A(_12549_),
    .B(_12563_),
    .Y(_12564_));
 NOR2x1_ASAP7_75t_R _41587_ (.A(_12542_),
    .B(_12564_),
    .Y(_12565_));
 NAND2x2_ASAP7_75t_R _41588_ (.A(_12520_),
    .B(_12565_),
    .Y(_12566_));
 XOR2x2_ASAP7_75t_R _41589_ (.A(_12486_),
    .B(_12566_),
    .Y(_12567_));
 XOR2x1_ASAP7_75t_R _41590_ (.A(_12403_),
    .Y(_12568_),
    .B(_12567_));
 AO21x1_ASAP7_75t_R _41591_ (.A1(_10832_),
    .A2(net1492),
    .B(_10864_),
    .Y(_12569_));
 AO21x1_ASAP7_75t_R _41592_ (.A1(_10671_),
    .A2(net1982),
    .B(_10864_),
    .Y(_12570_));
 AND3x1_ASAP7_75t_R _41593_ (.A(_12569_),
    .B(_12257_),
    .C(_12570_),
    .Y(_12571_));
 AO21x1_ASAP7_75t_R _41594_ (.A1(_10682_),
    .A2(net1475),
    .B(net3031),
    .Y(_12572_));
 OAI21x1_ASAP7_75t_R _41595_ (.A1(_10671_),
    .A2(net3031),
    .B(_12572_),
    .Y(_12574_));
 NOR2x1_ASAP7_75t_R _41596_ (.A(_10740_),
    .B(_10826_),
    .Y(_12575_));
 OR3x1_ASAP7_75t_R _41597_ (.A(_10828_),
    .B(_11868_),
    .C(_12575_),
    .Y(_12576_));
 NOR2x1_ASAP7_75t_R _41598_ (.A(_12574_),
    .B(_12576_),
    .Y(_12577_));
 NAND2x1_ASAP7_75t_R _41599_ (.A(_12571_),
    .B(_12577_),
    .Y(_12578_));
 AO21x1_ASAP7_75t_R _41600_ (.A1(_10783_),
    .A2(_10905_),
    .B(_10843_),
    .Y(_12579_));
 AO21x1_ASAP7_75t_R _41601_ (.A1(_10671_),
    .A2(net1982),
    .B(_10843_),
    .Y(_12580_));
 AO21x1_ASAP7_75t_R _41602_ (.A1(_10717_),
    .A2(net3049),
    .B(_10843_),
    .Y(_12581_));
 AND3x2_ASAP7_75t_R _41603_ (.A(_12579_),
    .B(_12580_),
    .C(_12581_),
    .Y(_12582_));
 AO21x1_ASAP7_75t_R _41604_ (.A1(_10730_),
    .A2(_10710_),
    .B(net1994),
    .Y(_12583_));
 NOR2x1_ASAP7_75t_R _41605_ (.A(net3033),
    .B(_12583_),
    .Y(_12585_));
 INVx1_ASAP7_75t_R _41606_ (.A(_11040_),
    .Y(_12586_));
 NAND2x1_ASAP7_75t_R _41607_ (.A(_11862_),
    .B(_12586_),
    .Y(_12587_));
 NOR2x2_ASAP7_75t_R _41608_ (.A(_12585_),
    .B(_12587_),
    .Y(_12588_));
 AO21x1_ASAP7_75t_R _41609_ (.A1(_10832_),
    .A2(net3020),
    .B(_10851_),
    .Y(_12589_));
 AO21x1_ASAP7_75t_R _41610_ (.A1(_10807_),
    .A2(net1492),
    .B(net3033),
    .Y(_12590_));
 AND2x2_ASAP7_75t_R _41611_ (.A(_12589_),
    .B(_12590_),
    .Y(_12591_));
 NAND3x2_ASAP7_75t_R _41612_ (.B(_12588_),
    .C(_12591_),
    .Y(_12592_),
    .A(_12582_));
 NOR2x2_ASAP7_75t_R _41613_ (.A(_12578_),
    .B(_12592_),
    .Y(_12593_));
 AND3x1_ASAP7_75t_R _41614_ (.A(_10791_),
    .B(_10626_),
    .C(net1344),
    .Y(_12594_));
 INVx1_ASAP7_75t_R _41615_ (.A(_12594_),
    .Y(_12596_));
 AO21x1_ASAP7_75t_R _41616_ (.A1(_10671_),
    .A2(_10938_),
    .B(_10785_),
    .Y(_12597_));
 AO21x1_ASAP7_75t_R _41617_ (.A1(net1288),
    .A2(net3049),
    .B(_10785_),
    .Y(_12598_));
 AND3x1_ASAP7_75t_R _41618_ (.A(_12596_),
    .B(_12597_),
    .C(_12598_),
    .Y(_12599_));
 AO21x1_ASAP7_75t_R _41619_ (.A1(_10767_),
    .A2(net1982),
    .B(_10796_),
    .Y(_12600_));
 AND4x1_ASAP7_75t_R _41620_ (.A(_10804_),
    .B(_12600_),
    .C(_12284_),
    .D(_11835_),
    .Y(_12601_));
 NAND2x1_ASAP7_75t_R _41621_ (.A(_12599_),
    .B(_12601_),
    .Y(_12602_));
 AO21x1_ASAP7_75t_R _41622_ (.A1(_10788_),
    .A2(_10759_),
    .B(_10816_),
    .Y(_12603_));
 AO21x1_ASAP7_75t_R _41623_ (.A1(net3049),
    .A2(_10645_),
    .B(_10816_),
    .Y(_12604_));
 NOR2x1_ASAP7_75t_R _41624_ (.A(net3046),
    .B(_10816_),
    .Y(_12605_));
 INVx1_ASAP7_75t_R _41625_ (.A(_12605_),
    .Y(_12607_));
 AND3x1_ASAP7_75t_R _41626_ (.A(_12603_),
    .B(_12604_),
    .C(_12607_),
    .Y(_12608_));
 OA21x2_ASAP7_75t_R _41627_ (.A1(_10647_),
    .A2(_12202_),
    .B(_10809_),
    .Y(_12609_));
 OA21x2_ASAP7_75t_R _41628_ (.A1(_10708_),
    .A2(_11043_),
    .B(_10809_),
    .Y(_12610_));
 AOI211x1_ASAP7_75t_R _41629_ (.A1(_10809_),
    .A2(_11812_),
    .B(_12609_),
    .C(_12610_),
    .Y(_12611_));
 AOI211x1_ASAP7_75t_R _41630_ (.A1(net1501),
    .A2(_10658_),
    .B(net3056),
    .C(net2024),
    .Y(_12612_));
 NOR2x1_ASAP7_75t_R _41631_ (.A(_10816_),
    .B(net1475),
    .Y(_12613_));
 AOI211x1_ASAP7_75t_R _41632_ (.A1(_11851_),
    .A2(_10992_),
    .B(_12612_),
    .C(_12613_),
    .Y(_12614_));
 NAND3x1_ASAP7_75t_R _41633_ (.A(_12608_),
    .B(_12611_),
    .C(_12614_),
    .Y(_12615_));
 NOR2x1_ASAP7_75t_R _41634_ (.A(_12602_),
    .B(_12615_),
    .Y(_12616_));
 NAND2x2_ASAP7_75t_R _41635_ (.A(_12593_),
    .B(_12616_),
    .Y(_12618_));
 AO21x1_ASAP7_75t_R _41636_ (.A1(_10767_),
    .A2(_10672_),
    .B(_10705_),
    .Y(_12619_));
 NOR2x1_ASAP7_75t_R _41637_ (.A(_10705_),
    .B(_10751_),
    .Y(_12620_));
 INVx1_ASAP7_75t_R _41638_ (.A(_12620_),
    .Y(_12621_));
 AND2x2_ASAP7_75t_R _41639_ (.A(_12619_),
    .B(_12621_),
    .Y(_12622_));
 NAND2x1_ASAP7_75t_R _41640_ (.A(_10713_),
    .B(_11012_),
    .Y(_12623_));
 AO21x1_ASAP7_75t_R _41641_ (.A1(_10686_),
    .A2(_10624_),
    .B(_10696_),
    .Y(_12624_));
 AND3x2_ASAP7_75t_R _41642_ (.A(_12622_),
    .B(_12623_),
    .C(_12624_),
    .Y(_12625_));
 NOR2x1_ASAP7_75t_R _41643_ (.A(_10624_),
    .B(_10637_),
    .Y(_12626_));
 NOR2x1_ASAP7_75t_R _41644_ (.A(_12626_),
    .B(_10903_),
    .Y(_12627_));
 AND2x2_ASAP7_75t_R _41645_ (.A(_10996_),
    .B(_10642_),
    .Y(_12629_));
 NOR2x1_ASAP7_75t_R _41646_ (.A(_10767_),
    .B(_10637_),
    .Y(_12630_));
 AOI211x1_ASAP7_75t_R _41647_ (.A1(_10642_),
    .A2(_11043_),
    .B(_12629_),
    .C(_12630_),
    .Y(_12631_));
 NAND2x1_ASAP7_75t_R _41648_ (.A(_12627_),
    .B(_12631_),
    .Y(_12632_));
 AO21x1_ASAP7_75t_R _41649_ (.A1(_10767_),
    .A2(_10768_),
    .B(_10664_),
    .Y(_12633_));
 AO21x1_ASAP7_75t_R _41650_ (.A1(_10751_),
    .A2(_10771_),
    .B(_10664_),
    .Y(_12634_));
 AND2x2_ASAP7_75t_R _41651_ (.A(_12633_),
    .B(_12634_),
    .Y(_12635_));
 AO21x1_ASAP7_75t_R _41652_ (.A1(_10624_),
    .A2(_10660_),
    .B(_10664_),
    .Y(_12636_));
 OA21x2_ASAP7_75t_R _41653_ (.A1(_10759_),
    .A2(_10664_),
    .B(_12636_),
    .Y(_12637_));
 NAND2x1_ASAP7_75t_R _41654_ (.A(_12635_),
    .B(_12637_),
    .Y(_12638_));
 NOR2x2_ASAP7_75t_R _41655_ (.A(_12632_),
    .B(_12638_),
    .Y(_12640_));
 NAND2x2_ASAP7_75t_R _41656_ (.A(_12625_),
    .B(_12640_),
    .Y(_12641_));
 INVx1_ASAP7_75t_R _41657_ (.A(_12641_),
    .Y(_12642_));
 INVx3_ASAP7_75t_R _41658_ (.A(_10771_),
    .Y(_12643_));
 NAND2x1_ASAP7_75t_R _41659_ (.A(_10754_),
    .B(_12643_),
    .Y(_12644_));
 NAND2x1_ASAP7_75t_R _41660_ (.A(_10782_),
    .B(_10754_),
    .Y(_12645_));
 NAND2x1_ASAP7_75t_R _41661_ (.A(_10754_),
    .B(_11008_),
    .Y(_12646_));
 AND4x2_ASAP7_75t_R _41662_ (.A(_12644_),
    .B(_12645_),
    .C(_11799_),
    .D(_12646_),
    .Y(_12647_));
 AO21x1_ASAP7_75t_R _41663_ (.A1(net1475),
    .A2(_10694_),
    .B(net3040),
    .Y(_12648_));
 AO21x1_ASAP7_75t_R _41664_ (.A1(_10807_),
    .A2(_10740_),
    .B(net3040),
    .Y(_12649_));
 INVx1_ASAP7_75t_R _41665_ (.A(_10700_),
    .Y(_12651_));
 NAND2x1_ASAP7_75t_R _41666_ (.A(_12651_),
    .B(_10774_),
    .Y(_12652_));
 AND3x2_ASAP7_75t_R _41667_ (.A(_12648_),
    .B(_12649_),
    .C(_12652_),
    .Y(_12653_));
 AO21x1_ASAP7_75t_R _41668_ (.A1(net3020),
    .A2(net3049),
    .B(_10755_),
    .Y(_12654_));
 OA21x2_ASAP7_75t_R _41669_ (.A1(_10755_),
    .A2(net3057),
    .B(_12654_),
    .Y(_12655_));
 NAND3x2_ASAP7_75t_R _41670_ (.B(_12653_),
    .C(_12655_),
    .Y(_12656_),
    .A(_12647_));
 NAND2x1_ASAP7_75t_R _41671_ (.A(_12214_),
    .B(_10726_),
    .Y(_12657_));
 NOR2x2_ASAP7_75t_R _41672_ (.A(net1423),
    .B(_10966_),
    .Y(_12658_));
 NOR2x2_ASAP7_75t_R _41673_ (.A(_12657_),
    .B(_12658_),
    .Y(_12659_));
 OA21x2_ASAP7_75t_R _41674_ (.A1(_10767_),
    .A2(_10725_),
    .B(_11783_),
    .Y(_12660_));
 AO21x1_ASAP7_75t_R _41675_ (.A1(_10767_),
    .A2(net2053),
    .B(_10739_),
    .Y(_12662_));
 AO21x1_ASAP7_75t_R _41676_ (.A1(_10745_),
    .A2(net3048),
    .B(_10739_),
    .Y(_12663_));
 INVx2_ASAP7_75t_R _41677_ (.A(_10739_),
    .Y(_12664_));
 NAND2x1_ASAP7_75t_R _41678_ (.A(_12664_),
    .B(_12643_),
    .Y(_12665_));
 AND3x2_ASAP7_75t_R _41679_ (.A(_12662_),
    .B(_12663_),
    .C(_12665_),
    .Y(_12666_));
 NAND3x2_ASAP7_75t_R _41680_ (.B(_12660_),
    .C(_12666_),
    .Y(_12667_),
    .A(_12659_));
 NOR2x1_ASAP7_75t_R _41681_ (.A(_12656_),
    .B(_12667_),
    .Y(_12668_));
 NAND2x1_ASAP7_75t_R _41682_ (.A(_12642_),
    .B(_12668_),
    .Y(_12669_));
 NOR2x2_ASAP7_75t_R _41683_ (.A(_12618_),
    .B(_12669_),
    .Y(_12670_));
 XOR2x2_ASAP7_75t_R _41684_ (.A(_12670_),
    .B(_10877_),
    .Y(_12671_));
 INVx1_ASAP7_75t_R _41685_ (.A(_11347_),
    .Y(_12673_));
 NAND3x1_ASAP7_75t_R _41686_ (.A(_12673_),
    .B(_11933_),
    .C(_10552_),
    .Y(_12674_));
 AND3x1_ASAP7_75t_R _41687_ (.A(_10537_),
    .B(net2962),
    .C(net1271),
    .Y(_12675_));
 NOR2x1_ASAP7_75t_R _41688_ (.A(net2953),
    .B(_10540_),
    .Y(_12676_));
 OA21x2_ASAP7_75t_R _41689_ (.A1(net2807),
    .A2(_11317_),
    .B(_10537_),
    .Y(_12677_));
 OR3x1_ASAP7_75t_R _41690_ (.A(_12675_),
    .B(_12676_),
    .C(_12677_),
    .Y(_12678_));
 NOR2x1_ASAP7_75t_R _41691_ (.A(_12674_),
    .B(_12678_),
    .Y(_12679_));
 OA21x2_ASAP7_75t_R _41692_ (.A1(net2456),
    .A2(_10576_),
    .B(_11350_),
    .Y(_12680_));
 OA21x2_ASAP7_75t_R _41693_ (.A1(net1264),
    .A2(_11338_),
    .B(_11350_),
    .Y(_12681_));
 NOR2x1_ASAP7_75t_R _41694_ (.A(net1876),
    .B(net2228),
    .Y(_12682_));
 OR3x1_ASAP7_75t_R _41695_ (.A(_12680_),
    .B(_12681_),
    .C(_12682_),
    .Y(_12684_));
 NAND2x1_ASAP7_75t_R _41696_ (.A(_10530_),
    .B(_10529_),
    .Y(_12685_));
 NOR2x1_ASAP7_75t_R _41697_ (.A(net1306),
    .B(_11355_),
    .Y(_12686_));
 OA21x2_ASAP7_75t_R _41698_ (.A1(_10385_),
    .A2(net2714),
    .B(_10528_),
    .Y(_12687_));
 OR3x1_ASAP7_75t_R _41699_ (.A(_12685_),
    .B(_12686_),
    .C(_12687_),
    .Y(_12688_));
 NOR2x1_ASAP7_75t_R _41700_ (.A(_12684_),
    .B(_12688_),
    .Y(_12689_));
 NAND2x1_ASAP7_75t_R _41701_ (.A(_12679_),
    .B(_12689_),
    .Y(_12690_));
 AOI211x1_ASAP7_75t_R _41702_ (.A1(net975),
    .A2(net1318),
    .B(net966),
    .C(net2180),
    .Y(_12691_));
 INVx1_ASAP7_75t_R _41703_ (.A(_12691_),
    .Y(_12692_));
 AO21x1_ASAP7_75t_R _41704_ (.A1(net3318),
    .A2(net1306),
    .B(net2180),
    .Y(_12693_));
 AND2x2_ASAP7_75t_R _41705_ (.A(_12692_),
    .B(_12693_),
    .Y(_12695_));
 NAND2x1_ASAP7_75t_R _41706_ (.A(_10531_),
    .B(_10589_),
    .Y(_12696_));
 AND3x1_ASAP7_75t_R _41707_ (.A(_12696_),
    .B(_11907_),
    .C(_11525_),
    .Y(_12697_));
 NOR2x1_ASAP7_75t_R _41708_ (.A(_11920_),
    .B(_10607_),
    .Y(_12698_));
 AND3x1_ASAP7_75t_R _41709_ (.A(_12695_),
    .B(_12697_),
    .C(_12698_),
    .Y(_12699_));
 AO21x1_ASAP7_75t_R _41710_ (.A1(net1115),
    .A2(_10502_),
    .B(net2211),
    .Y(_12700_));
 OA21x2_ASAP7_75t_R _41711_ (.A1(net3158),
    .A2(net2211),
    .B(_12700_),
    .Y(_12701_));
 NAND2x1_ASAP7_75t_R _41712_ (.A(_11539_),
    .B(_12701_),
    .Y(_12702_));
 AOI211x1_ASAP7_75t_R _41713_ (.A1(net975),
    .A2(net1318),
    .B(net1515),
    .C(net1840),
    .Y(_12703_));
 AOI21x1_ASAP7_75t_R _41714_ (.A1(_10550_),
    .A2(_10579_),
    .B(_12703_),
    .Y(_12704_));
 OA21x2_ASAP7_75t_R _41715_ (.A1(_10554_),
    .A2(net2715),
    .B(_10579_),
    .Y(_12706_));
 NOR2x1_ASAP7_75t_R _41716_ (.A(net1840),
    .B(net1115),
    .Y(_12707_));
 AOI211x1_ASAP7_75t_R _41717_ (.A1(_10579_),
    .A2(net2455),
    .B(_12706_),
    .C(_12707_),
    .Y(_12708_));
 NAND2x1_ASAP7_75t_R _41718_ (.A(_12704_),
    .B(_12708_),
    .Y(_12709_));
 NOR2x1_ASAP7_75t_R _41719_ (.A(_12702_),
    .B(_12709_),
    .Y(_12710_));
 NAND2x1_ASAP7_75t_R _41720_ (.A(_12699_),
    .B(_12710_),
    .Y(_12711_));
 NOR2x1_ASAP7_75t_R _41721_ (.A(_12690_),
    .B(_12711_),
    .Y(_12712_));
 AND2x2_ASAP7_75t_R _41722_ (.A(_10439_),
    .B(_10367_),
    .Y(_12713_));
 NOR2x1_ASAP7_75t_R _41723_ (.A(net1881),
    .B(net2957),
    .Y(_12714_));
 AOI21x1_ASAP7_75t_R _41724_ (.A1(net3318),
    .A2(net3014),
    .B(net1881),
    .Y(_12715_));
 OR3x1_ASAP7_75t_R _41725_ (.A(_12713_),
    .B(_12714_),
    .C(_12715_),
    .Y(_12717_));
 AO21x1_ASAP7_75t_R _41726_ (.A1(_10375_),
    .A2(net1114),
    .B(net2536),
    .Y(_12718_));
 AO21x1_ASAP7_75t_R _41727_ (.A1(net3297),
    .A2(_10410_),
    .B(net2536),
    .Y(_12719_));
 AND2x2_ASAP7_75t_R _41728_ (.A(_12718_),
    .B(_12719_),
    .Y(_12720_));
 NAND3x1_ASAP7_75t_R _41729_ (.A(_12720_),
    .B(_11380_),
    .C(_10422_),
    .Y(_12721_));
 NOR2x1_ASAP7_75t_R _41730_ (.A(_12717_),
    .B(_12721_),
    .Y(_12722_));
 OA21x2_ASAP7_75t_R _41731_ (.A1(_10557_),
    .A2(net2806),
    .B(_11368_),
    .Y(_12723_));
 NAND2x1_ASAP7_75t_R _41732_ (.A(_11368_),
    .B(net3019),
    .Y(_12724_));
 INVx1_ASAP7_75t_R _41733_ (.A(_12724_),
    .Y(_12725_));
 OA21x2_ASAP7_75t_R _41734_ (.A1(_11967_),
    .A2(_11349_),
    .B(_11368_),
    .Y(_12726_));
 OR3x1_ASAP7_75t_R _41735_ (.A(_12723_),
    .B(_12725_),
    .C(_12726_),
    .Y(_12728_));
 AND3x1_ASAP7_75t_R _41736_ (.A(_10323_),
    .B(net2962),
    .C(net2566),
    .Y(_12729_));
 NOR2x1_ASAP7_75t_R _41737_ (.A(_10375_),
    .B(_10336_),
    .Y(_12730_));
 INVx1_ASAP7_75t_R _41738_ (.A(_10351_),
    .Y(_12731_));
 NOR2x1_ASAP7_75t_R _41739_ (.A(_10502_),
    .B(_10336_),
    .Y(_12732_));
 OR4x1_ASAP7_75t_R _41740_ (.A(_12729_),
    .B(_12730_),
    .C(_12731_),
    .D(_12732_),
    .Y(_12733_));
 NOR2x1_ASAP7_75t_R _41741_ (.A(_12728_),
    .B(_12733_),
    .Y(_12734_));
 NAND2x1_ASAP7_75t_R _41742_ (.A(_12722_),
    .B(_12734_),
    .Y(_12735_));
 AO21x1_ASAP7_75t_R _41743_ (.A1(net1090),
    .A2(_10505_),
    .B(net2020),
    .Y(_12736_));
 AND2x2_ASAP7_75t_R _41744_ (.A(_12736_),
    .B(_11993_),
    .Y(_12737_));
 NAND2x1_ASAP7_75t_R _41745_ (.A(_11317_),
    .B(_10462_),
    .Y(_12739_));
 AO21x1_ASAP7_75t_R _41746_ (.A1(_11323_),
    .A2(net1125),
    .B(net2020),
    .Y(_12740_));
 NAND3x1_ASAP7_75t_R _41747_ (.A(_12737_),
    .B(_12739_),
    .C(_12740_),
    .Y(_12741_));
 AO21x1_ASAP7_75t_R _41748_ (.A1(_11323_),
    .A2(net2189),
    .B(net2233),
    .Y(_12742_));
 NAND2x1_ASAP7_75t_R _41749_ (.A(net958),
    .B(net2566),
    .Y(_12743_));
 AO21x1_ASAP7_75t_R _41750_ (.A1(_10329_),
    .A2(_12743_),
    .B(_10468_),
    .Y(_12744_));
 NAND2x2_ASAP7_75t_R _41751_ (.A(_11463_),
    .B(_12744_),
    .Y(_12745_));
 AOI21x1_ASAP7_75t_R _41752_ (.A1(_11967_),
    .A2(_11397_),
    .B(_12745_),
    .Y(_12746_));
 NAND2x1_ASAP7_75t_R _41753_ (.A(_12742_),
    .B(_12746_),
    .Y(_12747_));
 NOR2x1_ASAP7_75t_R _41754_ (.A(_12747_),
    .B(_12741_),
    .Y(_12748_));
 AO21x1_ASAP7_75t_R _41755_ (.A1(_11323_),
    .A2(net3052),
    .B(net2069),
    .Y(_12750_));
 NAND2x1_ASAP7_75t_R _41756_ (.A(_10576_),
    .B(_10483_),
    .Y(_12751_));
 AND3x1_ASAP7_75t_R _41757_ (.A(_12750_),
    .B(_10494_),
    .C(_12751_),
    .Y(_12752_));
 AO21x1_ASAP7_75t_R _41758_ (.A1(net1494),
    .A2(_10502_),
    .B(net2247),
    .Y(_12753_));
 NAND2x1_ASAP7_75t_R _41759_ (.A(net2806),
    .B(_11413_),
    .Y(_12754_));
 AND3x1_ASAP7_75t_R _41760_ (.A(_12753_),
    .B(_11418_),
    .C(_12754_),
    .Y(_12755_));
 AO21x1_ASAP7_75t_R _41761_ (.A1(net2952),
    .A2(net1090),
    .B(net2069),
    .Y(_12756_));
 AND3x1_ASAP7_75t_R _41762_ (.A(_12752_),
    .B(_12755_),
    .C(_12756_),
    .Y(_12757_));
 NAND2x1_ASAP7_75t_R _41763_ (.A(_12748_),
    .B(_12757_),
    .Y(_12758_));
 NOR2x2_ASAP7_75t_R _41764_ (.A(_12758_),
    .B(_12735_),
    .Y(_12759_));
 NAND2x2_ASAP7_75t_R _41765_ (.A(_12712_),
    .B(_12759_),
    .Y(_12761_));
 INVx2_ASAP7_75t_R _41766_ (.A(_12761_),
    .Y(_12762_));
 XOR2x1_ASAP7_75t_R _41767_ (.A(_12671_),
    .Y(_12763_),
    .B(_12762_));
 NOR2x1_ASAP7_75t_R _41768_ (.A(_12568_),
    .B(_12763_),
    .Y(_12764_));
 XOR2x1_ASAP7_75t_R _41769_ (.A(_12671_),
    .Y(_12765_),
    .B(_12761_));
 INVx1_ASAP7_75t_R _41770_ (.A(_12568_),
    .Y(_12766_));
 NOR2x1_ASAP7_75t_R _41771_ (.A(_12765_),
    .B(_12766_),
    .Y(_12767_));
 OAI21x1_ASAP7_75t_R _41772_ (.A1(_12764_),
    .A2(_12767_),
    .B(net392),
    .Y(_12768_));
 AOI21x1_ASAP7_75t_R _41773_ (.A1(_12402_),
    .A2(_12768_),
    .B(_00522_),
    .Y(_12769_));
 NAND2x1_ASAP7_75t_R _41774_ (.A(_00815_),
    .B(net389),
    .Y(_12770_));
 NOR2x1_ASAP7_75t_R _41775_ (.A(_12566_),
    .B(_12486_),
    .Y(_12772_));
 INVx1_ASAP7_75t_R _41776_ (.A(_12503_),
    .Y(_12773_));
 NOR2x1_ASAP7_75t_R _41777_ (.A(_12519_),
    .B(_12511_),
    .Y(_12774_));
 NAND2x1_ASAP7_75t_R _41778_ (.A(_12773_),
    .B(_12774_),
    .Y(_12775_));
 INVx1_ASAP7_75t_R _41779_ (.A(_12542_),
    .Y(_12776_));
 INVx1_ASAP7_75t_R _41780_ (.A(_12549_),
    .Y(_12777_));
 NAND3x1_ASAP7_75t_R _41781_ (.A(_12555_),
    .B(_12560_),
    .C(_12558_),
    .Y(_12778_));
 NOR2x1_ASAP7_75t_R _41782_ (.A(_12777_),
    .B(_12778_),
    .Y(_12779_));
 NAND2x1_ASAP7_75t_R _41783_ (.A(_12776_),
    .B(_12779_),
    .Y(_12780_));
 NOR2x2_ASAP7_75t_R _41784_ (.A(_12775_),
    .B(_12780_),
    .Y(_12781_));
 AND4x1_ASAP7_75t_R _41785_ (.A(_12427_),
    .B(_12439_),
    .C(_12426_),
    .D(_12465_),
    .Y(_12783_));
 NAND3x1_ASAP7_75t_R _41786_ (.A(_12435_),
    .B(_12350_),
    .C(_12318_),
    .Y(_12784_));
 INVx1_ASAP7_75t_R _41787_ (.A(_12784_),
    .Y(_12785_));
 NAND3x1_ASAP7_75t_R _41788_ (.A(_12783_),
    .B(_10212_),
    .C(_12785_),
    .Y(_12786_));
 AOI21x1_ASAP7_75t_R _41789_ (.A1(_09876_),
    .A2(_11212_),
    .B(_12409_),
    .Y(_12787_));
 NOR2x1_ASAP7_75t_R _41790_ (.A(net3309),
    .B(_10079_),
    .Y(_12788_));
 NOR2x1_ASAP7_75t_R _41791_ (.A(_09948_),
    .B(_12788_),
    .Y(_12789_));
 NAND2x1_ASAP7_75t_R _41792_ (.A(_12787_),
    .B(_12789_),
    .Y(_12790_));
 NAND2x1_ASAP7_75t_R _41793_ (.A(_11653_),
    .B(_12479_),
    .Y(_12791_));
 NOR2x1_ASAP7_75t_R _41794_ (.A(_11618_),
    .B(_12791_),
    .Y(_12792_));
 AOI221x1_ASAP7_75t_R _41795_ (.A1(net2382),
    .A2(net2627),
    .B1(_09959_),
    .B2(net1950),
    .C(_10074_),
    .Y(_12794_));
 NAND2x1_ASAP7_75t_R _41796_ (.A(_12792_),
    .B(_12794_),
    .Y(_12795_));
 NOR2x1_ASAP7_75t_R _41797_ (.A(_12790_),
    .B(_12795_),
    .Y(_12796_));
 AND2x2_ASAP7_75t_R _41798_ (.A(_12457_),
    .B(_11638_),
    .Y(_12797_));
 AO21x1_ASAP7_75t_R _41799_ (.A1(net1963),
    .A2(_09928_),
    .B(net2662),
    .Y(_12798_));
 AO21x1_ASAP7_75t_R _41800_ (.A1(_10015_),
    .A2(_10042_),
    .B(net2535),
    .Y(_12799_));
 AND2x2_ASAP7_75t_R _41801_ (.A(_12798_),
    .B(_12799_),
    .Y(_12800_));
 AND3x1_ASAP7_75t_R _41802_ (.A(_10255_),
    .B(net1022),
    .C(net2283),
    .Y(_12801_));
 NOR2x1_ASAP7_75t_R _41803_ (.A(_12369_),
    .B(_12801_),
    .Y(_12802_));
 OA21x2_ASAP7_75t_R _41804_ (.A1(_10289_),
    .A2(_09990_),
    .B(_12480_),
    .Y(_12803_));
 AND4x1_ASAP7_75t_R _41805_ (.A(_12797_),
    .B(_12800_),
    .C(_12802_),
    .D(_12803_),
    .Y(_12805_));
 NAND2x1_ASAP7_75t_R _41806_ (.A(_12796_),
    .B(_12805_),
    .Y(_12806_));
 NOR2x1_ASAP7_75t_R _41807_ (.A(_12786_),
    .B(_12806_),
    .Y(_12807_));
 NAND2x1_ASAP7_75t_R _41808_ (.A(_12437_),
    .B(_12444_),
    .Y(_12808_));
 NOR2x1_ASAP7_75t_R _41809_ (.A(_12808_),
    .B(_11266_),
    .Y(_12809_));
 AOI22x1_ASAP7_75t_R _41810_ (.A1(_11656_),
    .A2(_09994_),
    .B1(_10140_),
    .B2(_10077_),
    .Y(_12810_));
 AND3x1_ASAP7_75t_R _41811_ (.A(_12809_),
    .B(_11588_),
    .C(_12810_),
    .Y(_12811_));
 NAND2x2_ASAP7_75t_R _41812_ (.A(net1700),
    .B(_09974_),
    .Y(_12812_));
 OAI21x1_ASAP7_75t_R _41813_ (.A1(_09953_),
    .A2(net1353),
    .B(_12812_),
    .Y(_12813_));
 OAI22x1_ASAP7_75t_R _41814_ (.A1(_11604_),
    .A2(_10035_),
    .B1(_10085_),
    .B2(_09937_),
    .Y(_12814_));
 AO21x1_ASAP7_75t_R _41815_ (.A1(_10254_),
    .A2(_12813_),
    .B(_12814_),
    .Y(_12816_));
 AO21x2_ASAP7_75t_R _41816_ (.A1(net2382),
    .A2(net2583),
    .B(_12440_),
    .Y(_12817_));
 AO21x1_ASAP7_75t_R _41817_ (.A1(_11627_),
    .A2(_10157_),
    .B(_12410_),
    .Y(_12818_));
 NOR3x1_ASAP7_75t_R _41818_ (.A(_12816_),
    .B(_12817_),
    .C(_12818_),
    .Y(_12819_));
 NAND2x1_ASAP7_75t_R _41819_ (.A(_12811_),
    .B(_12819_),
    .Y(_12820_));
 AOI21x1_ASAP7_75t_R _41820_ (.A1(net1890),
    .A2(_11627_),
    .B(_12411_),
    .Y(_12821_));
 AOI22x1_ASAP7_75t_R _41821_ (.A1(_10140_),
    .A2(net2576),
    .B1(_09946_),
    .B2(_10157_),
    .Y(_12822_));
 AND2x2_ASAP7_75t_R _41822_ (.A(_12821_),
    .B(_12822_),
    .Y(_12823_));
 NOR2x1_ASAP7_75t_R _41823_ (.A(_10100_),
    .B(_11223_),
    .Y(_12824_));
 NOR2x1_ASAP7_75t_R _41824_ (.A(_09870_),
    .B(_09942_),
    .Y(_12825_));
 NOR2x1_ASAP7_75t_R _41825_ (.A(_10063_),
    .B(_10005_),
    .Y(_12827_));
 NOR2x1_ASAP7_75t_R _41826_ (.A(_10042_),
    .B(_09901_),
    .Y(_12828_));
 AOI211x1_ASAP7_75t_R _41827_ (.A1(_11212_),
    .A2(_12825_),
    .B(_12827_),
    .C(_12828_),
    .Y(_12829_));
 AND3x1_ASAP7_75t_R _41828_ (.A(_12823_),
    .B(_12824_),
    .C(_12829_),
    .Y(_12830_));
 OAI21x1_ASAP7_75t_R _41829_ (.A1(net2353),
    .A2(net2358),
    .B(_10073_),
    .Y(_12831_));
 AO21x1_ASAP7_75t_R _41830_ (.A1(_10164_),
    .A2(_10157_),
    .B(_11593_),
    .Y(_12832_));
 NOR2x1_ASAP7_75t_R _41831_ (.A(_12831_),
    .B(_12832_),
    .Y(_12833_));
 OAI21x1_ASAP7_75t_R _41832_ (.A1(_10111_),
    .A2(net2353),
    .B(_11201_),
    .Y(_12834_));
 AOI211x1_ASAP7_75t_R _41833_ (.A1(net2222),
    .A2(_10157_),
    .B(_12834_),
    .C(_09938_),
    .Y(_12835_));
 NAND2x1_ASAP7_75t_R _41834_ (.A(_12833_),
    .B(_12835_),
    .Y(_12836_));
 AND4x1_ASAP7_75t_R _41835_ (.A(_10141_),
    .B(_12406_),
    .C(_10132_),
    .D(_12432_),
    .Y(_12838_));
 AOI22x1_ASAP7_75t_R _41836_ (.A1(net2382),
    .A2(_11558_),
    .B1(net2627),
    .B2(_09876_),
    .Y(_12839_));
 NAND2x1_ASAP7_75t_R _41837_ (.A(_10152_),
    .B(_10140_),
    .Y(_12840_));
 AND3x1_ASAP7_75t_R _41838_ (.A(_12839_),
    .B(_12840_),
    .C(_10278_),
    .Y(_12841_));
 NAND2x1_ASAP7_75t_R _41839_ (.A(_12838_),
    .B(_12841_),
    .Y(_12842_));
 NOR2x1_ASAP7_75t_R _41840_ (.A(_12836_),
    .B(_12842_),
    .Y(_12843_));
 NAND2x1_ASAP7_75t_R _41841_ (.A(_12830_),
    .B(_12843_),
    .Y(_12844_));
 NOR2x2_ASAP7_75t_R _41842_ (.A(_12820_),
    .B(_12844_),
    .Y(_12845_));
 NAND2x2_ASAP7_75t_R _41843_ (.A(_12807_),
    .B(_12845_),
    .Y(_12846_));
 NOR2x1_ASAP7_75t_R _41844_ (.A(_12781_),
    .B(_12846_),
    .Y(_12847_));
 OAI21x1_ASAP7_75t_R _41845_ (.A1(_12772_),
    .A2(_12847_),
    .B(_12762_),
    .Y(_12849_));
 NOR2x1_ASAP7_75t_R _41846_ (.A(_12486_),
    .B(_12781_),
    .Y(_12850_));
 NOR2x1_ASAP7_75t_R _41847_ (.A(_12566_),
    .B(_12846_),
    .Y(_12851_));
 OAI21x1_ASAP7_75t_R _41848_ (.A1(_12850_),
    .A2(_12851_),
    .B(_12761_),
    .Y(_12852_));
 NAND2x1_ASAP7_75t_R _41849_ (.A(_12849_),
    .B(_12852_),
    .Y(_12853_));
 INVx1_ASAP7_75t_R _41850_ (.A(_12853_),
    .Y(_12854_));
 XOR2x2_ASAP7_75t_R _41851_ (.A(_12384_),
    .B(net1882),
    .Y(_12855_));
 XOR2x1_ASAP7_75t_R _41852_ (.A(_12671_),
    .Y(_12856_),
    .B(_12855_));
 NAND2x1_ASAP7_75t_R _41853_ (.A(_12856_),
    .B(_12854_),
    .Y(_12857_));
 NOR2x1_ASAP7_75t_R _41854_ (.A(_12855_),
    .B(_12671_),
    .Y(_12858_));
 AND2x2_ASAP7_75t_R _41855_ (.A(_12671_),
    .B(_12855_),
    .Y(_12860_));
 OAI21x1_ASAP7_75t_R _41856_ (.A1(_12858_),
    .A2(_12860_),
    .B(_12853_),
    .Y(_12861_));
 NAND3x1_ASAP7_75t_R _41857_ (.A(_12857_),
    .B(_12861_),
    .C(net392),
    .Y(_12862_));
 INVx1_ASAP7_75t_R _41858_ (.A(_00522_),
    .Y(_12863_));
 AOI21x1_ASAP7_75t_R _41859_ (.A1(_12770_),
    .A2(_12862_),
    .B(_12863_),
    .Y(_12864_));
 NOR2x2_ASAP7_75t_R _41860_ (.A(_12864_),
    .B(_12769_),
    .Y(_00101_));
 OR2x2_ASAP7_75t_R _41861_ (.A(net393),
    .B(_00814_),
    .Y(_12865_));
 AO21x1_ASAP7_75t_R _41862_ (.A1(_10678_),
    .A2(_10767_),
    .B(_10816_),
    .Y(_12866_));
 AO21x1_ASAP7_75t_R _41863_ (.A1(net3057),
    .A2(_10757_),
    .B(_10816_),
    .Y(_12867_));
 AND3x2_ASAP7_75t_R _41864_ (.A(_12866_),
    .B(_12867_),
    .C(_12607_),
    .Y(_12868_));
 AO21x1_ASAP7_75t_R _41865_ (.A1(_12583_),
    .A2(net1982),
    .B(_10810_),
    .Y(_12870_));
 NAND3x2_ASAP7_75t_R _41866_ (.B(_11003_),
    .C(_12870_),
    .Y(_12871_),
    .A(_12868_));
 AND3x1_ASAP7_75t_R _41867_ (.A(_12596_),
    .B(_11841_),
    .C(_11013_),
    .Y(_12872_));
 AO21x1_ASAP7_75t_R _41868_ (.A1(net1862),
    .A2(net1475),
    .B(_10796_),
    .Y(_12873_));
 AO21x1_ASAP7_75t_R _41869_ (.A1(_10645_),
    .A2(_10656_),
    .B(_10796_),
    .Y(_12874_));
 OA211x2_ASAP7_75t_R _41870_ (.A1(_10700_),
    .A2(_10796_),
    .B(_12873_),
    .C(_12874_),
    .Y(_12875_));
 NAND2x1_ASAP7_75t_R _41871_ (.A(_12872_),
    .B(_12875_),
    .Y(_12876_));
 NOR2x2_ASAP7_75t_R _41872_ (.A(_12871_),
    .B(_12876_),
    .Y(_12877_));
 AO21x1_ASAP7_75t_R _41873_ (.A1(net3057),
    .A2(_10740_),
    .B(_10843_),
    .Y(_12878_));
 NAND2x1_ASAP7_75t_R _41874_ (.A(_11044_),
    .B(_12878_),
    .Y(_12879_));
 OA21x2_ASAP7_75t_R _41875_ (.A1(_10792_),
    .A2(_10708_),
    .B(_11860_),
    .Y(_12881_));
 AOI211x1_ASAP7_75t_R _41876_ (.A1(net1501),
    .A2(net1419),
    .B(net1990),
    .C(net3033),
    .Y(_12882_));
 AOI21x1_ASAP7_75t_R _41877_ (.A1(_11036_),
    .A2(_10807_),
    .B(net3033),
    .Y(_12883_));
 OR4x2_ASAP7_75t_R _41878_ (.A(_12879_),
    .B(_12881_),
    .C(_12882_),
    .D(_12883_),
    .Y(_12884_));
 NOR2x1_ASAP7_75t_R _41879_ (.A(net3054),
    .B(net1862),
    .Y(_12885_));
 OA211x2_ASAP7_75t_R _41880_ (.A1(net1501),
    .A2(net1418),
    .B(_10870_),
    .C(_10677_),
    .Y(_12886_));
 NOR2x2_ASAP7_75t_R _41881_ (.A(_12885_),
    .B(_12886_),
    .Y(_12887_));
 NOR2x1_ASAP7_75t_R _41882_ (.A(net3054),
    .B(_10832_),
    .Y(_12888_));
 OA211x2_ASAP7_75t_R _41883_ (.A1(_10626_),
    .A2(_10658_),
    .B(_10870_),
    .C(net2148),
    .Y(_12889_));
 NOR2x2_ASAP7_75t_R _41884_ (.A(_12888_),
    .B(_12889_),
    .Y(_12890_));
 AO21x1_ASAP7_75t_R _41885_ (.A1(net1862),
    .A2(_10671_),
    .B(net3029),
    .Y(_12892_));
 NAND2x1_ASAP7_75t_R _41886_ (.A(_10681_),
    .B(_10827_),
    .Y(_12893_));
 AND3x2_ASAP7_75t_R _41887_ (.A(_12892_),
    .B(_12261_),
    .C(_12893_),
    .Y(_12894_));
 NAND3x2_ASAP7_75t_R _41888_ (.B(_12890_),
    .C(_12894_),
    .Y(_12895_),
    .A(_12887_));
 NOR2x2_ASAP7_75t_R _41889_ (.A(_12884_),
    .B(_12895_),
    .Y(_12896_));
 NAND2x2_ASAP7_75t_R _41890_ (.A(_12877_),
    .B(_12896_),
    .Y(_12897_));
 AO21x1_ASAP7_75t_R _41891_ (.A1(net1862),
    .A2(_10671_),
    .B(_10755_),
    .Y(_12898_));
 AND3x1_ASAP7_75t_R _41892_ (.A(_12898_),
    .B(_11801_),
    .C(_12644_),
    .Y(_12899_));
 INVx1_ASAP7_75t_R _41893_ (.A(_10942_),
    .Y(_12900_));
 AO21x1_ASAP7_75t_R _41894_ (.A1(_10700_),
    .A2(net3049),
    .B(net3040),
    .Y(_12901_));
 NAND2x1_ASAP7_75t_R _41895_ (.A(_10681_),
    .B(_10774_),
    .Y(_12903_));
 AND4x1_ASAP7_75t_R _41896_ (.A(_12900_),
    .B(_12901_),
    .C(_12206_),
    .D(_12903_),
    .Y(_12904_));
 NAND2x1_ASAP7_75t_R _41897_ (.A(_12899_),
    .B(_12904_),
    .Y(_12905_));
 NAND2x1_ASAP7_75t_R _41898_ (.A(_10782_),
    .B(_12664_),
    .Y(_12906_));
 AO21x1_ASAP7_75t_R _41899_ (.A1(net1862),
    .A2(_10747_),
    .B(_10739_),
    .Y(_12907_));
 NAND2x1_ASAP7_75t_R _41900_ (.A(_12906_),
    .B(_12907_),
    .Y(_12908_));
 INVx1_ASAP7_75t_R _41901_ (.A(_10746_),
    .Y(_12909_));
 NOR2x1_ASAP7_75t_R _41902_ (.A(_10740_),
    .B(_10739_),
    .Y(_12910_));
 NOR3x1_ASAP7_75t_R _41903_ (.A(_12908_),
    .B(_12909_),
    .C(_12910_),
    .Y(_12911_));
 OA211x2_ASAP7_75t_R _41904_ (.A1(net1501),
    .A2(net1422),
    .B(_10736_),
    .C(net1336),
    .Y(_12912_));
 NOR2x1_ASAP7_75t_R _41905_ (.A(_12912_),
    .B(_12658_),
    .Y(_12914_));
 NAND2x1_ASAP7_75t_R _41906_ (.A(net3061),
    .B(_10736_),
    .Y(_12915_));
 AO21x1_ASAP7_75t_R _41907_ (.A1(_10783_),
    .A2(net1475),
    .B(_10725_),
    .Y(_12916_));
 NAND2x1_ASAP7_75t_R _41908_ (.A(_12915_),
    .B(_12916_),
    .Y(_12917_));
 INVx1_ASAP7_75t_R _41909_ (.A(_12917_),
    .Y(_12918_));
 NAND3x1_ASAP7_75t_R _41910_ (.A(_12911_),
    .B(_12914_),
    .C(_12918_),
    .Y(_12919_));
 NOR2x1_ASAP7_75t_R _41911_ (.A(_12905_),
    .B(_12919_),
    .Y(_12920_));
 AO21x1_ASAP7_75t_R _41912_ (.A1(net3020),
    .A2(net3049),
    .B(_10637_),
    .Y(_12921_));
 OAI21x1_ASAP7_75t_R _41913_ (.A1(_10637_),
    .A2(net3023),
    .B(_12921_),
    .Y(_12922_));
 NOR2x1_ASAP7_75t_R _41914_ (.A(_10771_),
    .B(_10637_),
    .Y(_12923_));
 OR3x1_ASAP7_75t_R _41915_ (.A(_10688_),
    .B(_12630_),
    .C(_12923_),
    .Y(_12925_));
 NOR2x1_ASAP7_75t_R _41916_ (.A(_12922_),
    .B(_12925_),
    .Y(_12926_));
 AO21x1_ASAP7_75t_R _41917_ (.A1(_10832_),
    .A2(net3022),
    .B(_10696_),
    .Y(_12927_));
 NOR2x1_ASAP7_75t_R _41918_ (.A(net1982),
    .B(_10696_),
    .Y(_12928_));
 INVx1_ASAP7_75t_R _41919_ (.A(_12928_),
    .Y(_12929_));
 AO21x1_ASAP7_75t_R _41920_ (.A1(_10767_),
    .A2(_10671_),
    .B(_10696_),
    .Y(_12930_));
 NAND3x1_ASAP7_75t_R _41921_ (.A(_12927_),
    .B(_12929_),
    .C(_12930_),
    .Y(_12931_));
 AOI21x1_ASAP7_75t_R _41922_ (.A1(_10713_),
    .A2(_11798_),
    .B(_10707_),
    .Y(_12932_));
 AO21x1_ASAP7_75t_R _41923_ (.A1(_10788_),
    .A2(net1492),
    .B(_10705_),
    .Y(_12933_));
 AO21x1_ASAP7_75t_R _41924_ (.A1(_10832_),
    .A2(_10656_),
    .B(_10705_),
    .Y(_12934_));
 NAND3x1_ASAP7_75t_R _41925_ (.A(_12932_),
    .B(_12933_),
    .C(_12934_),
    .Y(_12936_));
 NOR2x1_ASAP7_75t_R _41926_ (.A(_12931_),
    .B(_12936_),
    .Y(_12937_));
 OAI21x1_ASAP7_75t_R _41927_ (.A1(net3021),
    .A2(_10788_),
    .B(_12226_),
    .Y(_12938_));
 NAND2x1_ASAP7_75t_R _41928_ (.A(_11851_),
    .B(_11822_),
    .Y(_12939_));
 NAND2x1_ASAP7_75t_R _41929_ (.A(_12939_),
    .B(_10912_),
    .Y(_12940_));
 AOI211x1_ASAP7_75t_R _41930_ (.A1(_11043_),
    .A2(_11822_),
    .B(_12938_),
    .C(_12940_),
    .Y(_12941_));
 AND3x2_ASAP7_75t_R _41931_ (.A(_12926_),
    .B(_12937_),
    .C(_12941_),
    .Y(_12942_));
 NAND2x2_ASAP7_75t_R _41932_ (.A(_12920_),
    .B(_12942_),
    .Y(_12943_));
 NOR2x2_ASAP7_75t_R _41933_ (.A(_12897_),
    .B(_12943_),
    .Y(_12944_));
 NAND2x2_ASAP7_75t_R _41934_ (.A(_12486_),
    .B(_12944_),
    .Y(_12945_));
 OAI21x1_ASAP7_75t_R _41935_ (.A1(_12897_),
    .A2(_12943_),
    .B(_12846_),
    .Y(_12947_));
 AO21x1_ASAP7_75t_R _41936_ (.A1(net1876),
    .A2(net1055),
    .B(net2464),
    .Y(_12948_));
 AND4x2_ASAP7_75t_R _41937_ (.A(_11393_),
    .B(_11993_),
    .C(_12739_),
    .D(_12948_),
    .Y(_12949_));
 AO21x1_ASAP7_75t_R _41938_ (.A1(net1876),
    .A2(net1090),
    .B(net1981),
    .Y(_12950_));
 AO21x1_ASAP7_75t_R _41939_ (.A1(net1115),
    .A2(net1306),
    .B(net1981),
    .Y(_12951_));
 AO21x1_ASAP7_75t_R _41940_ (.A1(_11312_),
    .A2(net3161),
    .B(net1981),
    .Y(_12952_));
 NAND2x1_ASAP7_75t_R _41941_ (.A(net2716),
    .B(_11397_),
    .Y(_12953_));
 AND4x2_ASAP7_75t_R _41942_ (.A(_12950_),
    .B(_12951_),
    .C(_12952_),
    .D(_12953_),
    .Y(_12954_));
 AO21x1_ASAP7_75t_R _41943_ (.A1(net3051),
    .A2(net2952),
    .B(net2070),
    .Y(_12955_));
 AO21x1_ASAP7_75t_R _41944_ (.A1(_11379_),
    .A2(net1125),
    .B(net2070),
    .Y(_12956_));
 NAND2x2_ASAP7_75t_R _41945_ (.A(_12955_),
    .B(_12956_),
    .Y(_12958_));
 NAND2x2_ASAP7_75t_R _41946_ (.A(_10507_),
    .B(_10501_),
    .Y(_12959_));
 AO21x1_ASAP7_75t_R _41947_ (.A1(net1414),
    .A2(net1306),
    .B(net2249),
    .Y(_12960_));
 NAND2x2_ASAP7_75t_R _41948_ (.A(_11448_),
    .B(_12960_),
    .Y(_12961_));
 NOR3x2_ASAP7_75t_R _41949_ (.B(_12959_),
    .C(_12961_),
    .Y(_12962_),
    .A(_12958_));
 NAND3x2_ASAP7_75t_R _41950_ (.B(_12954_),
    .C(_12962_),
    .Y(_12963_),
    .A(_12949_));
 NOR2x1_ASAP7_75t_R _41951_ (.A(net2449),
    .B(_10420_),
    .Y(_12964_));
 NOR2x1_ASAP7_75t_R _41952_ (.A(net2333),
    .B(net2449),
    .Y(_12965_));
 OR3x2_ASAP7_75t_R _41953_ (.A(_12964_),
    .B(_12965_),
    .C(_10439_),
    .Y(_12966_));
 OAI21x1_ASAP7_75t_R _41954_ (.A1(net2868),
    .A2(_11486_),
    .B(_11380_),
    .Y(_12967_));
 AO21x1_ASAP7_75t_R _41955_ (.A1(_11312_),
    .A2(_11364_),
    .B(net2329),
    .Y(_12969_));
 AO21x1_ASAP7_75t_R _41956_ (.A1(net2954),
    .A2(net1090),
    .B(net2329),
    .Y(_12970_));
 NAND2x2_ASAP7_75t_R _41957_ (.A(_12969_),
    .B(_12970_),
    .Y(_12971_));
 NOR3x2_ASAP7_75t_R _41958_ (.B(_12967_),
    .C(_12971_),
    .Y(_12972_),
    .A(_12966_));
 AO221x1_ASAP7_75t_R _41959_ (.A1(net975),
    .A2(net3338),
    .B1(_10341_),
    .B2(net1510),
    .C(_10336_),
    .Y(_12973_));
 NOR2x1_ASAP7_75t_R _41960_ (.A(_12731_),
    .B(_11373_),
    .Y(_12974_));
 AND2x2_ASAP7_75t_R _41961_ (.A(_12973_),
    .B(_12974_),
    .Y(_12975_));
 AO21x1_ASAP7_75t_R _41962_ (.A1(net3014),
    .A2(net1125),
    .B(net2240),
    .Y(_12976_));
 AO21x1_ASAP7_75t_R _41963_ (.A1(net3051),
    .A2(_11364_),
    .B(net2240),
    .Y(_12977_));
 AO21x1_ASAP7_75t_R _41964_ (.A1(net1080),
    .A2(net1090),
    .B(net2240),
    .Y(_12978_));
 AND3x2_ASAP7_75t_R _41965_ (.A(_12976_),
    .B(_12977_),
    .C(_12978_),
    .Y(_12980_));
 NAND3x2_ASAP7_75t_R _41966_ (.B(_12975_),
    .C(_12980_),
    .Y(_12981_),
    .A(_12972_));
 NOR2x2_ASAP7_75t_R _41967_ (.A(_12963_),
    .B(_12981_),
    .Y(_12982_));
 OA211x2_ASAP7_75t_R _41968_ (.A1(net1270),
    .A2(_11932_),
    .B(_10589_),
    .C(net1318),
    .Y(_12983_));
 AO21x1_ASAP7_75t_R _41969_ (.A1(net1090),
    .A2(net1114),
    .B(net2180),
    .Y(_12984_));
 AO21x1_ASAP7_75t_R _41970_ (.A1(_10502_),
    .A2(net3157),
    .B(net2180),
    .Y(_12985_));
 NAND2x2_ASAP7_75t_R _41971_ (.A(_12984_),
    .B(_12985_),
    .Y(_12986_));
 OA31x2_ASAP7_75t_R _41972_ (.A1(_11532_),
    .A2(_10597_),
    .A3(net2714),
    .B1(_10589_),
    .Y(_12987_));
 NOR3x2_ASAP7_75t_R _41973_ (.B(_12986_),
    .C(_12987_),
    .Y(_12988_),
    .A(_12983_));
 AO21x1_ASAP7_75t_R _41974_ (.A1(net1115),
    .A2(net3318),
    .B(net2211),
    .Y(_12989_));
 AO21x1_ASAP7_75t_R _41975_ (.A1(_10375_),
    .A2(net1659),
    .B(net2211),
    .Y(_12991_));
 NAND2x1_ASAP7_75t_R _41976_ (.A(net2951),
    .B(_10572_),
    .Y(_12992_));
 AND4x1_ASAP7_75t_R _41977_ (.A(_12989_),
    .B(_12991_),
    .C(_11538_),
    .D(_12992_),
    .Y(_12993_));
 AO21x1_ASAP7_75t_R _41978_ (.A1(net2854),
    .A2(net3051),
    .B(net1840),
    .Y(_12994_));
 AO21x1_ASAP7_75t_R _41979_ (.A1(net1115),
    .A2(net967),
    .B(net1840),
    .Y(_12995_));
 NOR2x1_ASAP7_75t_R _41980_ (.A(net3333),
    .B(_10333_),
    .Y(_12996_));
 INVx1_ASAP7_75t_R _41981_ (.A(_12996_),
    .Y(_12997_));
 NAND3x1_ASAP7_75t_R _41982_ (.A(_12994_),
    .B(_12995_),
    .C(_12997_),
    .Y(_12998_));
 INVx1_ASAP7_75t_R _41983_ (.A(_12998_),
    .Y(_12999_));
 NAND3x1_ASAP7_75t_R _41984_ (.A(_12988_),
    .B(_12993_),
    .C(_12999_),
    .Y(_13000_));
 OA21x2_ASAP7_75t_R _41985_ (.A1(net1306),
    .A2(net2228),
    .B(_11515_),
    .Y(_13002_));
 AOI211x1_ASAP7_75t_R _41986_ (.A1(net975),
    .A2(net3338),
    .B(net2228),
    .C(net1516),
    .Y(_13003_));
 INVx1_ASAP7_75t_R _41987_ (.A(_13003_),
    .Y(_13004_));
 AO21x1_ASAP7_75t_R _41988_ (.A1(net1090),
    .A2(_10505_),
    .B(net2228),
    .Y(_13005_));
 AND3x1_ASAP7_75t_R _41989_ (.A(_13002_),
    .B(_13004_),
    .C(_13005_),
    .Y(_13006_));
 AO21x1_ASAP7_75t_R _41990_ (.A1(_11323_),
    .A2(_11306_),
    .B(_10540_),
    .Y(_13007_));
 NAND2x1_ASAP7_75t_R _41991_ (.A(_11927_),
    .B(_13007_),
    .Y(_13008_));
 AO21x1_ASAP7_75t_R _41992_ (.A1(net2957),
    .A2(net2952),
    .B(net3043),
    .Y(_13009_));
 AO21x1_ASAP7_75t_R _41993_ (.A1(net1143),
    .A2(net1054),
    .B(net3043),
    .Y(_13010_));
 NAND2x1_ASAP7_75t_R _41994_ (.A(net2807),
    .B(_10547_),
    .Y(_13011_));
 NAND3x1_ASAP7_75t_R _41995_ (.A(_13009_),
    .B(_13010_),
    .C(_13011_),
    .Y(_13013_));
 NOR2x1_ASAP7_75t_R _41996_ (.A(_13008_),
    .B(_13013_),
    .Y(_13014_));
 OA211x2_ASAP7_75t_R _41997_ (.A1(net975),
    .A2(net1318),
    .B(_10528_),
    .C(net2951),
    .Y(_13015_));
 AND3x1_ASAP7_75t_R _41998_ (.A(_10528_),
    .B(net3319),
    .C(_10367_),
    .Y(_13016_));
 AOI211x1_ASAP7_75t_R _41999_ (.A1(_11317_),
    .A2(_10528_),
    .B(_13015_),
    .C(_13016_),
    .Y(_13017_));
 NAND3x1_ASAP7_75t_R _42000_ (.A(_13006_),
    .B(_13014_),
    .C(_13017_),
    .Y(_13018_));
 NOR2x1_ASAP7_75t_R _42001_ (.A(_13000_),
    .B(_13018_),
    .Y(_13019_));
 NAND2x2_ASAP7_75t_R _42002_ (.A(_12982_),
    .B(_13019_),
    .Y(_13020_));
 NOR2x2_ASAP7_75t_R _42003_ (.A(_10364_),
    .B(_13020_),
    .Y(_13021_));
 AOI21x1_ASAP7_75t_R _42004_ (.A1(_12945_),
    .A2(_12947_),
    .B(net3294),
    .Y(_13022_));
 INVx1_ASAP7_75t_R _42005_ (.A(_12945_),
    .Y(_13024_));
 NOR2x1_ASAP7_75t_R _42006_ (.A(_12486_),
    .B(_12944_),
    .Y(_13025_));
 INVx1_ASAP7_75t_R _42007_ (.A(net3294),
    .Y(_13026_));
 NOR3x1_ASAP7_75t_R _42008_ (.A(_13024_),
    .B(_13025_),
    .C(_13026_),
    .Y(_13027_));
 OAI22x1_ASAP7_75t_R _42009_ (.A1(_10247_),
    .A2(_10005_),
    .B1(_10042_),
    .B2(_10011_),
    .Y(_13028_));
 NOR2x1_ASAP7_75t_R _42010_ (.A(_12808_),
    .B(_13028_),
    .Y(_13029_));
 AND3x4_ASAP7_75t_R _42011_ (.A(_12785_),
    .B(_10219_),
    .C(_13029_),
    .Y(_13030_));
 NOR2x1_ASAP7_75t_R _42012_ (.A(_09934_),
    .B(_10011_),
    .Y(_13031_));
 AOI22x1_ASAP7_75t_R _42013_ (.A1(_13031_),
    .A2(net2049),
    .B1(net2627),
    .B2(net2431),
    .Y(_13032_));
 OA22x2_ASAP7_75t_R _42014_ (.A1(net2808),
    .A2(_09937_),
    .B1(_10123_),
    .B2(net1161),
    .Y(_13033_));
 NAND2x1_ASAP7_75t_R _42015_ (.A(_13032_),
    .B(_13033_),
    .Y(_13035_));
 AO21x1_ASAP7_75t_R _42016_ (.A1(net2391),
    .A2(net3245),
    .B(_10060_),
    .Y(_13036_));
 OAI21x1_ASAP7_75t_R _42017_ (.A1(net3309),
    .A2(_10132_),
    .B(_13036_),
    .Y(_13037_));
 AO21x1_ASAP7_75t_R _42018_ (.A1(net3015),
    .A2(_10294_),
    .B(_13037_),
    .Y(_13038_));
 NOR2x2_ASAP7_75t_R _42019_ (.A(_13035_),
    .B(_13038_),
    .Y(_13039_));
 NOR2x2_ASAP7_75t_R _42020_ (.A(_11625_),
    .B(_11612_),
    .Y(_13040_));
 NOR2x2_ASAP7_75t_R _42021_ (.A(_09990_),
    .B(net2936),
    .Y(_13041_));
 AOI21x1_ASAP7_75t_R _42022_ (.A1(_10157_),
    .A2(_09959_),
    .B(_13041_),
    .Y(_13042_));
 NAND3x2_ASAP7_75t_R _42023_ (.B(_10012_),
    .C(_13042_),
    .Y(_13043_),
    .A(_13040_));
 NOR2x1_ASAP7_75t_R _42024_ (.A(_10003_),
    .B(_10005_),
    .Y(_13044_));
 AOI22x1_ASAP7_75t_R _42025_ (.A1(_13044_),
    .A2(net1161),
    .B1(net2575),
    .B2(_10071_),
    .Y(_13046_));
 AO21x1_ASAP7_75t_R _42026_ (.A1(_10063_),
    .A2(_10008_),
    .B(_09901_),
    .Y(_13047_));
 NAND3x2_ASAP7_75t_R _42027_ (.B(_12480_),
    .C(_13047_),
    .Y(_13048_),
    .A(_13046_));
 NOR2x2_ASAP7_75t_R _42028_ (.A(_13048_),
    .B(_13043_),
    .Y(_13049_));
 NAND3x2_ASAP7_75t_R _42029_ (.B(_13039_),
    .C(_13049_),
    .Y(_13050_),
    .A(_13030_));
 OAI21x1_ASAP7_75t_R _42030_ (.A1(net2353),
    .A2(_10015_),
    .B(_12468_),
    .Y(_13051_));
 NOR2x2_ASAP7_75t_R _42031_ (.A(net3309),
    .B(_10073_),
    .Y(_13052_));
 NOR3x2_ASAP7_75t_R _42032_ (.B(_10252_),
    .C(_13052_),
    .Y(_13053_),
    .A(_13051_));
 AND4x2_ASAP7_75t_R _42033_ (.A(_10052_),
    .B(_10043_),
    .C(_11231_),
    .D(_10031_),
    .Y(_13054_));
 NAND2x2_ASAP7_75t_R _42034_ (.A(_13054_),
    .B(_13053_),
    .Y(_13055_));
 OA22x2_ASAP7_75t_R _42035_ (.A1(_10098_),
    .A2(_09919_),
    .B1(net3062),
    .B2(_11561_),
    .Y(_13057_));
 OA21x2_ASAP7_75t_R _42036_ (.A1(_09925_),
    .A2(_09922_),
    .B(_11201_),
    .Y(_13058_));
 NAND2x1_ASAP7_75t_R _42037_ (.A(_13057_),
    .B(_13058_),
    .Y(_13059_));
 AOI22x1_ASAP7_75t_R _42038_ (.A1(_11566_),
    .A2(_10044_),
    .B1(_09992_),
    .B2(_10080_),
    .Y(_13060_));
 NAND3x1_ASAP7_75t_R _42039_ (.A(_13060_),
    .B(_10168_),
    .C(_10173_),
    .Y(_13061_));
 NOR2x1_ASAP7_75t_R _42040_ (.A(_13059_),
    .B(_13061_),
    .Y(_13062_));
 AND2x2_ASAP7_75t_R _42041_ (.A(_09944_),
    .B(_10272_),
    .Y(_13063_));
 OA21x2_ASAP7_75t_R _42042_ (.A1(_09934_),
    .A2(_09990_),
    .B(_10170_),
    .Y(_13064_));
 NAND2x1_ASAP7_75t_R _42043_ (.A(_13063_),
    .B(_13064_),
    .Y(_13065_));
 NAND2x1_ASAP7_75t_R _42044_ (.A(_09910_),
    .B(_09888_),
    .Y(_13066_));
 OA21x2_ASAP7_75t_R _42045_ (.A1(_10035_),
    .A2(_13066_),
    .B(_10079_),
    .Y(_13068_));
 NAND2x1_ASAP7_75t_R _42046_ (.A(_11590_),
    .B(_13068_),
    .Y(_13069_));
 NOR2x1_ASAP7_75t_R _42047_ (.A(_13065_),
    .B(_13069_),
    .Y(_13070_));
 NAND2x1_ASAP7_75t_R _42048_ (.A(_13062_),
    .B(_13070_),
    .Y(_13071_));
 NOR2x2_ASAP7_75t_R _42049_ (.A(_13071_),
    .B(_13055_),
    .Y(_13072_));
 AO22x1_ASAP7_75t_R _42050_ (.A1(_10164_),
    .A2(net2804),
    .B1(_10044_),
    .B2(_11558_),
    .Y(_13073_));
 NAND2x2_ASAP7_75t_R _42051_ (.A(net1165),
    .B(net1699),
    .Y(_13074_));
 NOR2x2_ASAP7_75t_R _42052_ (.A(_13074_),
    .B(net3062),
    .Y(_13075_));
 AO21x1_ASAP7_75t_R _42053_ (.A1(_09941_),
    .A2(_10099_),
    .B(_13075_),
    .Y(_13076_));
 NOR2x1_ASAP7_75t_R _42054_ (.A(_13073_),
    .B(_13076_),
    .Y(_13077_));
 AO21x1_ASAP7_75t_R _42055_ (.A1(_10008_),
    .A2(net2958),
    .B(_10086_),
    .Y(_13079_));
 NAND2x1_ASAP7_75t_R _42056_ (.A(_09946_),
    .B(_10071_),
    .Y(_13080_));
 AND3x1_ASAP7_75t_R _42057_ (.A(_13079_),
    .B(_11639_),
    .C(_13080_),
    .Y(_13081_));
 NAND2x2_ASAP7_75t_R _42058_ (.A(_13077_),
    .B(_13081_),
    .Y(_13082_));
 NOR2x2_ASAP7_75t_R _42059_ (.A(_12817_),
    .B(_12814_),
    .Y(_13083_));
 AND2x2_ASAP7_75t_R _42060_ (.A(_10187_),
    .B(_11600_),
    .Y(_13084_));
 NAND2x2_ASAP7_75t_R _42061_ (.A(_13083_),
    .B(_13084_),
    .Y(_13085_));
 OAI21x1_ASAP7_75t_R _42062_ (.A1(net2353),
    .A2(net1661),
    .B(_12812_),
    .Y(_13086_));
 NOR2x1_ASAP7_75t_R _42063_ (.A(_13086_),
    .B(_11568_),
    .Y(_13087_));
 AO21x1_ASAP7_75t_R _42064_ (.A1(_11571_),
    .A2(_10044_),
    .B(_12828_),
    .Y(_13088_));
 AO21x1_ASAP7_75t_R _42065_ (.A1(_10027_),
    .A2(_10157_),
    .B(_12827_),
    .Y(_13090_));
 NOR2x1_ASAP7_75t_R _42066_ (.A(_13088_),
    .B(_13090_),
    .Y(_13091_));
 NAND2x2_ASAP7_75t_R _42067_ (.A(_13087_),
    .B(_13091_),
    .Y(_13092_));
 NOR3x2_ASAP7_75t_R _42068_ (.B(_13085_),
    .C(_13092_),
    .Y(_13093_),
    .A(_13082_));
 NAND2x2_ASAP7_75t_R _42069_ (.A(_13072_),
    .B(_13093_),
    .Y(_13094_));
 NOR2x2_ASAP7_75t_R _42070_ (.A(_13050_),
    .B(_13094_),
    .Y(_13095_));
 NAND2x2_ASAP7_75t_R _42071_ (.A(net2681),
    .B(_13095_),
    .Y(_13096_));
 INVx2_ASAP7_75t_R _42072_ (.A(_09628_),
    .Y(_13097_));
 AO21x1_ASAP7_75t_R _42073_ (.A1(_09817_),
    .A2(_09752_),
    .B(net2912),
    .Y(_13098_));
 NAND2x1_ASAP7_75t_R _42074_ (.A(_12131_),
    .B(_13098_),
    .Y(_13099_));
 NOR2x1_ASAP7_75t_R _42075_ (.A(net2434),
    .B(_09649_),
    .Y(_13100_));
 OA21x2_ASAP7_75t_R _42076_ (.A1(_09633_),
    .A2(_09809_),
    .B(_09846_),
    .Y(_13101_));
 NAND2x1_ASAP7_75t_R _42077_ (.A(_11187_),
    .B(_11124_),
    .Y(_13102_));
 OR4x2_ASAP7_75t_R _42078_ (.A(_13099_),
    .B(_13100_),
    .C(_13101_),
    .D(_13102_),
    .Y(_13103_));
 AOI211x1_ASAP7_75t_R _42079_ (.A1(net1105),
    .A2(_09573_),
    .B(_09770_),
    .C(_09579_),
    .Y(_13104_));
 OA21x2_ASAP7_75t_R _42080_ (.A1(_11677_),
    .A2(_09664_),
    .B(_09807_),
    .Y(_13105_));
 OR2x2_ASAP7_75t_R _42081_ (.A(_13104_),
    .B(_13105_),
    .Y(_13106_));
 AO21x1_ASAP7_75t_R _42082_ (.A1(net2732),
    .A2(_09715_),
    .B(_09682_),
    .Y(_13107_));
 NOR2x1_ASAP7_75t_R _42083_ (.A(_09682_),
    .B(_09711_),
    .Y(_13108_));
 INVx1_ASAP7_75t_R _42084_ (.A(_13108_),
    .Y(_13109_));
 NAND3x1_ASAP7_75t_R _42085_ (.A(_13107_),
    .B(_13109_),
    .C(_11671_),
    .Y(_13111_));
 AO21x1_ASAP7_75t_R _42086_ (.A1(_09858_),
    .A2(_09798_),
    .B(net2339),
    .Y(_13112_));
 INVx1_ASAP7_75t_R _42087_ (.A(_13112_),
    .Y(_13113_));
 OR3x4_ASAP7_75t_R _42088_ (.A(_13106_),
    .B(_13111_),
    .C(_13113_),
    .Y(_13114_));
 AO21x1_ASAP7_75t_R _42089_ (.A1(net1246),
    .A2(net1387),
    .B(net1503),
    .Y(_13115_));
 AOI21x1_ASAP7_75t_R _42090_ (.A1(_11177_),
    .A2(net2921),
    .B(net1503),
    .Y(_13116_));
 INVx1_ASAP7_75t_R _42091_ (.A(_13116_),
    .Y(_13117_));
 INVx1_ASAP7_75t_R _42092_ (.A(_11716_),
    .Y(_13118_));
 NAND3x1_ASAP7_75t_R _42093_ (.A(_13115_),
    .B(_13117_),
    .C(_13118_),
    .Y(_13119_));
 AO21x1_ASAP7_75t_R _42094_ (.A1(net1290),
    .A2(net3067),
    .B(net1999),
    .Y(_13120_));
 AO21x1_ASAP7_75t_R _42095_ (.A1(net1387),
    .A2(net986),
    .B(net1999),
    .Y(_13122_));
 NAND3x1_ASAP7_75t_R _42096_ (.A(_13120_),
    .B(_13122_),
    .C(_12033_),
    .Y(_13123_));
 NOR2x1_ASAP7_75t_R _42097_ (.A(_13119_),
    .B(_13123_),
    .Y(_13124_));
 AO21x1_ASAP7_75t_R _42098_ (.A1(_09658_),
    .A2(net2327),
    .B(net1868),
    .Y(_13125_));
 OAI21x1_ASAP7_75t_R _42099_ (.A1(_11161_),
    .A2(net1870),
    .B(_13125_),
    .Y(_13126_));
 AO21x1_ASAP7_75t_R _42100_ (.A1(_09653_),
    .A2(net2328),
    .B(net1942),
    .Y(_13127_));
 AO21x1_ASAP7_75t_R _42101_ (.A1(_09684_),
    .A2(net2105),
    .B(net1942),
    .Y(_13128_));
 NAND2x1_ASAP7_75t_R _42102_ (.A(_13127_),
    .B(_13128_),
    .Y(_13129_));
 AO21x1_ASAP7_75t_R _42103_ (.A1(net1596),
    .A2(net1102),
    .B(net1868),
    .Y(_13130_));
 NAND2x1_ASAP7_75t_R _42104_ (.A(_09859_),
    .B(_13130_),
    .Y(_13131_));
 NOR3x1_ASAP7_75t_R _42105_ (.A(_13126_),
    .B(_13129_),
    .C(_13131_),
    .Y(_13133_));
 NAND2x1_ASAP7_75t_R _42106_ (.A(_13124_),
    .B(_13133_),
    .Y(_13134_));
 NOR3x1_ASAP7_75t_R _42107_ (.A(_13103_),
    .B(_13114_),
    .C(_13134_),
    .Y(_13135_));
 OA211x2_ASAP7_75t_R _42108_ (.A1(net2152),
    .A2(net1101),
    .B(_09701_),
    .C(_09573_),
    .Y(_13136_));
 INVx1_ASAP7_75t_R _42109_ (.A(_13136_),
    .Y(_13137_));
 OA21x2_ASAP7_75t_R _42110_ (.A1(net1387),
    .A2(_09672_),
    .B(_11144_),
    .Y(_13138_));
 NAND2x1_ASAP7_75t_R _42111_ (.A(_13137_),
    .B(_13138_),
    .Y(_13139_));
 OA21x2_ASAP7_75t_R _42112_ (.A1(_11096_),
    .A2(_09700_),
    .B(_09826_),
    .Y(_13140_));
 OA21x2_ASAP7_75t_R _42113_ (.A1(_11675_),
    .A2(_09664_),
    .B(_09826_),
    .Y(_13141_));
 OA21x2_ASAP7_75t_R _42114_ (.A1(net2941),
    .A2(_11111_),
    .B(_09826_),
    .Y(_13142_));
 OR3x1_ASAP7_75t_R _42115_ (.A(_13140_),
    .B(_13141_),
    .C(_13142_),
    .Y(_13144_));
 NOR2x1_ASAP7_75t_R _42116_ (.A(_13139_),
    .B(_13144_),
    .Y(_13145_));
 AO21x1_ASAP7_75t_R _42117_ (.A1(net1387),
    .A2(net1596),
    .B(net1743),
    .Y(_13146_));
 AO21x1_ASAP7_75t_R _42118_ (.A1(net3067),
    .A2(net1577),
    .B(net1743),
    .Y(_13147_));
 NAND3x1_ASAP7_75t_R _42119_ (.A(_13146_),
    .B(_13147_),
    .C(_12084_),
    .Y(_13148_));
 AO21x1_ASAP7_75t_R _42120_ (.A1(net1246),
    .A2(net1102),
    .B(net2501),
    .Y(_13149_));
 OA21x2_ASAP7_75t_R _42121_ (.A1(net2501),
    .A2(net2732),
    .B(_13149_),
    .Y(_13150_));
 NAND2x1_ASAP7_75t_R _42122_ (.A(_13150_),
    .B(_09667_),
    .Y(_13151_));
 NOR2x1_ASAP7_75t_R _42123_ (.A(_13148_),
    .B(_13151_),
    .Y(_13152_));
 NAND2x1_ASAP7_75t_R _42124_ (.A(_13145_),
    .B(_13152_),
    .Y(_13153_));
 NAND2x1_ASAP7_75t_R _42125_ (.A(_09761_),
    .B(_11056_),
    .Y(_13155_));
 AND3x1_ASAP7_75t_R _42126_ (.A(_13155_),
    .B(_11106_),
    .C(_11057_),
    .Y(_13156_));
 INVx1_ASAP7_75t_R _42127_ (.A(_13156_),
    .Y(_13157_));
 NOR2x1_ASAP7_75t_R _42128_ (.A(_11693_),
    .B(_11699_),
    .Y(_13158_));
 AO21x1_ASAP7_75t_R _42129_ (.A1(_09658_),
    .A2(net2558),
    .B(_09707_),
    .Y(_13159_));
 AND2x2_ASAP7_75t_R _42130_ (.A(_13159_),
    .B(_12533_),
    .Y(_13160_));
 NAND2x1_ASAP7_75t_R _42131_ (.A(_13158_),
    .B(_13160_),
    .Y(_13161_));
 NOR2x2_ASAP7_75t_R _42132_ (.A(_13157_),
    .B(_13161_),
    .Y(_13162_));
 OA21x2_ASAP7_75t_R _42133_ (.A1(_11134_),
    .A2(_11167_),
    .B(_09838_),
    .Y(_13163_));
 NOR2x1_ASAP7_75t_R _42134_ (.A(_11731_),
    .B(_13163_),
    .Y(_13164_));
 AO21x1_ASAP7_75t_R _42135_ (.A1(net3067),
    .A2(net1577),
    .B(net2290),
    .Y(_13166_));
 AO21x1_ASAP7_75t_R _42136_ (.A1(net3069),
    .A2(net2217),
    .B(net2290),
    .Y(_13167_));
 AND3x2_ASAP7_75t_R _42137_ (.A(_13164_),
    .B(_13166_),
    .C(_13167_),
    .Y(_13168_));
 AO21x1_ASAP7_75t_R _42138_ (.A1(_09689_),
    .A2(net1577),
    .B(net2917),
    .Y(_13169_));
 AO21x1_ASAP7_75t_R _42139_ (.A1(_09658_),
    .A2(_09644_),
    .B(net2917),
    .Y(_13170_));
 AND4x2_ASAP7_75t_R _42140_ (.A(_11072_),
    .B(_09614_),
    .C(_13169_),
    .D(_13170_),
    .Y(_13171_));
 NAND3x1_ASAP7_75t_R _42141_ (.A(_13162_),
    .B(_13168_),
    .C(_13171_),
    .Y(_13172_));
 NOR2x1_ASAP7_75t_R _42142_ (.A(_13153_),
    .B(_13172_),
    .Y(_13173_));
 NAND2x1_ASAP7_75t_R _42143_ (.A(_13135_),
    .B(_13173_),
    .Y(_13174_));
 NOR2x2_ASAP7_75t_R _42144_ (.A(_13097_),
    .B(_13174_),
    .Y(_13175_));
 XNOR2x2_ASAP7_75t_R _42145_ (.A(_13096_),
    .B(_13175_),
    .Y(_13177_));
 INVx2_ASAP7_75t_R _42146_ (.A(_13177_),
    .Y(_13178_));
 OAI21x1_ASAP7_75t_R _42147_ (.A1(_13022_),
    .A2(_13027_),
    .B(_13178_),
    .Y(_13179_));
 INVx1_ASAP7_75t_R _42148_ (.A(_13179_),
    .Y(_13180_));
 NAND3x2_ASAP7_75t_R _42149_ (.B(_12945_),
    .C(net3294),
    .Y(_13181_),
    .A(_12947_));
 INVx1_ASAP7_75t_R _42150_ (.A(_13022_),
    .Y(_13182_));
 NAND3x2_ASAP7_75t_R _42151_ (.B(_13182_),
    .C(_13177_),
    .Y(_13183_),
    .A(_13181_));
 INVx1_ASAP7_75t_R _42152_ (.A(_13183_),
    .Y(_13184_));
 OAI21x1_ASAP7_75t_R _42153_ (.A1(_13180_),
    .A2(_13184_),
    .B(net393),
    .Y(_13185_));
 AOI21x1_ASAP7_75t_R _42154_ (.A1(_12865_),
    .A2(_13185_),
    .B(_00521_),
    .Y(_13186_));
 NAND2x1_ASAP7_75t_R _42155_ (.A(_00814_),
    .B(net389),
    .Y(_13188_));
 NAND3x1_ASAP7_75t_R _42156_ (.A(_13183_),
    .B(_13179_),
    .C(net393),
    .Y(_13189_));
 AOI21x1_ASAP7_75t_R _42157_ (.A1(_13188_),
    .A2(_13189_),
    .B(_17446_),
    .Y(_13190_));
 NOR2x1_ASAP7_75t_R _42158_ (.A(_13190_),
    .B(_13186_),
    .Y(_00102_));
 NOR2x2_ASAP7_75t_R _42159_ (.A(net393),
    .B(_00813_),
    .Y(_13191_));
 AO21x1_ASAP7_75t_R _42160_ (.A1(net1519),
    .A2(net2938),
    .B(net1868),
    .Y(_13192_));
 AO21x1_ASAP7_75t_R _42161_ (.A1(net3067),
    .A2(net2921),
    .B(net1869),
    .Y(_13193_));
 AND2x2_ASAP7_75t_R _42162_ (.A(_13192_),
    .B(_13193_),
    .Y(_13194_));
 AO21x1_ASAP7_75t_R _42163_ (.A1(_12521_),
    .A2(_09653_),
    .B(net1942),
    .Y(_13195_));
 AO21x1_ASAP7_75t_R _42164_ (.A1(net2105),
    .A2(net1596),
    .B(net1942),
    .Y(_13196_));
 AND2x2_ASAP7_75t_R _42165_ (.A(_13195_),
    .B(_13196_),
    .Y(_13198_));
 NAND2x1_ASAP7_75t_R _42166_ (.A(_13194_),
    .B(_13198_),
    .Y(_13199_));
 AO21x1_ASAP7_75t_R _42167_ (.A1(_11690_),
    .A2(_11161_),
    .B(net1503),
    .Y(_13200_));
 NAND2x1_ASAP7_75t_R _42168_ (.A(net2956),
    .B(_09806_),
    .Y(_13201_));
 AO21x1_ASAP7_75t_R _42169_ (.A1(net2503),
    .A2(net1102),
    .B(net1503),
    .Y(_13202_));
 NAND3x1_ASAP7_75t_R _42170_ (.A(_13200_),
    .B(_13201_),
    .C(_13202_),
    .Y(_13203_));
 AO21x1_ASAP7_75t_R _42171_ (.A1(net2921),
    .A2(_11177_),
    .B(net1999),
    .Y(_13204_));
 AO21x2_ASAP7_75t_R _42172_ (.A1(_09779_),
    .A2(_09581_),
    .B(net987),
    .Y(_13205_));
 AO21x1_ASAP7_75t_R _42173_ (.A1(_13205_),
    .A2(_11165_),
    .B(net1999),
    .Y(_13206_));
 NAND2x1_ASAP7_75t_R _42174_ (.A(_13204_),
    .B(_13206_),
    .Y(_13207_));
 NOR3x1_ASAP7_75t_R _42175_ (.A(_13199_),
    .B(_13203_),
    .C(_13207_),
    .Y(_13209_));
 AO21x1_ASAP7_75t_R _42176_ (.A1(_11160_),
    .A2(_09644_),
    .B(_09682_),
    .Y(_13210_));
 NAND2x1_ASAP7_75t_R _42177_ (.A(_09816_),
    .B(_09640_),
    .Y(_13211_));
 AND3x1_ASAP7_75t_R _42178_ (.A(_12012_),
    .B(_13210_),
    .C(_13211_),
    .Y(_13212_));
 AO21x1_ASAP7_75t_R _42179_ (.A1(net1562),
    .A2(_09711_),
    .B(net2085),
    .Y(_13213_));
 AO21x1_ASAP7_75t_R _42180_ (.A1(net2434),
    .A2(net2104),
    .B(net2085),
    .Y(_13214_));
 AO21x1_ASAP7_75t_R _42181_ (.A1(_09635_),
    .A2(net1479),
    .B(net2085),
    .Y(_13215_));
 AND3x1_ASAP7_75t_R _42182_ (.A(_13213_),
    .B(_13214_),
    .C(_13215_),
    .Y(_13216_));
 NAND2x1_ASAP7_75t_R _42183_ (.A(_13212_),
    .B(_13216_),
    .Y(_13217_));
 AO21x1_ASAP7_75t_R _42184_ (.A1(_09817_),
    .A2(_09613_),
    .B(net2912),
    .Y(_13218_));
 AO21x1_ASAP7_75t_R _42185_ (.A1(_12521_),
    .A2(_11690_),
    .B(net2912),
    .Y(_13220_));
 NAND2x1_ASAP7_75t_R _42186_ (.A(_13218_),
    .B(_13220_),
    .Y(_13221_));
 AO21x1_ASAP7_75t_R _42187_ (.A1(_09711_),
    .A2(_09684_),
    .B(net2943),
    .Y(_13222_));
 OAI21x1_ASAP7_75t_R _42188_ (.A1(net2943),
    .A2(_13205_),
    .B(_13222_),
    .Y(_13223_));
 AO21x1_ASAP7_75t_R _42189_ (.A1(_09635_),
    .A2(_09631_),
    .B(net2943),
    .Y(_13224_));
 AO21x1_ASAP7_75t_R _42190_ (.A1(_11161_),
    .A2(net3067),
    .B(net2943),
    .Y(_13225_));
 NAND2x1_ASAP7_75t_R _42191_ (.A(_13224_),
    .B(_13225_),
    .Y(_13226_));
 OR3x1_ASAP7_75t_R _42192_ (.A(_13221_),
    .B(_13223_),
    .C(_13226_),
    .Y(_13227_));
 NOR2x1_ASAP7_75t_R _42193_ (.A(_13217_),
    .B(_13227_),
    .Y(_13228_));
 NAND2x1_ASAP7_75t_R _42194_ (.A(_13209_),
    .B(_13228_),
    .Y(_13229_));
 AO21x1_ASAP7_75t_R _42195_ (.A1(_09658_),
    .A2(_09631_),
    .B(net2547),
    .Y(_13231_));
 NAND2x1_ASAP7_75t_R _42196_ (.A(_09741_),
    .B(_11056_),
    .Y(_13232_));
 NAND3x1_ASAP7_75t_R _42197_ (.A(_13231_),
    .B(_11057_),
    .C(_13232_),
    .Y(_13233_));
 AO21x1_ASAP7_75t_R _42198_ (.A1(_09711_),
    .A2(_09798_),
    .B(_09707_),
    .Y(_13234_));
 AO21x1_ASAP7_75t_R _42199_ (.A1(net1577),
    .A2(_09635_),
    .B(_09707_),
    .Y(_13235_));
 NAND3x1_ASAP7_75t_R _42200_ (.A(_13234_),
    .B(_13235_),
    .C(_12089_),
    .Y(_13236_));
 OR2x2_ASAP7_75t_R _42201_ (.A(_13233_),
    .B(_13236_),
    .Y(_13237_));
 AO21x1_ASAP7_75t_R _42202_ (.A1(_09858_),
    .A2(_09674_),
    .B(net3016),
    .Y(_13238_));
 AO21x1_ASAP7_75t_R _42203_ (.A1(net1544),
    .A2(_09644_),
    .B(net3016),
    .Y(_13239_));
 NAND2x1_ASAP7_75t_R _42204_ (.A(_13238_),
    .B(_13239_),
    .Y(_13240_));
 OR3x1_ASAP7_75t_R _42205_ (.A(_13240_),
    .B(_09615_),
    .C(_11709_),
    .Y(_13242_));
 NOR2x2_ASAP7_75t_R _42206_ (.A(_13237_),
    .B(_13242_),
    .Y(_13243_));
 OA21x2_ASAP7_75t_R _42207_ (.A1(_09832_),
    .A2(_11128_),
    .B(_09661_),
    .Y(_13244_));
 NOR3x1_ASAP7_75t_R _42208_ (.A(_13244_),
    .B(_11178_),
    .C(_11103_),
    .Y(_13245_));
 OA21x2_ASAP7_75t_R _42209_ (.A1(_09597_),
    .A2(net1743),
    .B(_11094_),
    .Y(_13246_));
 AO21x1_ASAP7_75t_R _42210_ (.A1(net2434),
    .A2(net2103),
    .B(net1743),
    .Y(_13247_));
 AND2x2_ASAP7_75t_R _42211_ (.A(_12082_),
    .B(_13247_),
    .Y(_13248_));
 NAND3x1_ASAP7_75t_R _42212_ (.A(_13245_),
    .B(_13246_),
    .C(_13248_),
    .Y(_13249_));
 NOR2x1_ASAP7_75t_R _42213_ (.A(net984),
    .B(_09801_),
    .Y(_13250_));
 INVx1_ASAP7_75t_R _42214_ (.A(_11183_),
    .Y(_13251_));
 NOR2x1_ASAP7_75t_R _42215_ (.A(_09798_),
    .B(_09801_),
    .Y(_13253_));
 AOI211x1_ASAP7_75t_R _42216_ (.A1(net1287),
    .A2(_13250_),
    .B(_13251_),
    .C(_13253_),
    .Y(_13254_));
 AO21x1_ASAP7_75t_R _42217_ (.A1(net1562),
    .A2(net2724),
    .B(net2916),
    .Y(_13255_));
 AO21x1_ASAP7_75t_R _42218_ (.A1(net2434),
    .A2(_09715_),
    .B(net2916),
    .Y(_13256_));
 AND2x2_ASAP7_75t_R _42219_ (.A(_13255_),
    .B(_13256_),
    .Y(_13257_));
 AOI211x1_ASAP7_75t_R _42220_ (.A1(_09589_),
    .A2(net1282),
    .B(net2916),
    .C(net1478),
    .Y(_13258_));
 AOI21x1_ASAP7_75t_R _42221_ (.A1(net2956),
    .A2(_09701_),
    .B(_13258_),
    .Y(_13259_));
 NAND3x1_ASAP7_75t_R _42222_ (.A(_13254_),
    .B(_13257_),
    .C(_13259_),
    .Y(_13260_));
 NOR2x1_ASAP7_75t_R _42223_ (.A(_13249_),
    .B(_13260_),
    .Y(_13261_));
 NAND2x2_ASAP7_75t_R _42224_ (.A(_13243_),
    .B(_13261_),
    .Y(_13262_));
 AOI211x1_ASAP7_75t_R _42225_ (.A1(_09627_),
    .A2(net1762),
    .B(_13229_),
    .C(_13262_),
    .Y(_13264_));
 TAPCELL_ASAP7_75t_R PHY_29 ();
 AO21x2_ASAP7_75t_R _42227_ (.A1(_09961_),
    .A2(_09992_),
    .B(_10217_),
    .Y(_13266_));
 OAI21x1_ASAP7_75t_R _42228_ (.A1(_10060_),
    .A2(_10059_),
    .B(_12468_),
    .Y(_13267_));
 NOR3x2_ASAP7_75t_R _42229_ (.B(_13267_),
    .C(_10032_),
    .Y(_13268_),
    .A(_13266_));
 AND2x2_ASAP7_75t_R _42230_ (.A(net2565),
    .B(net1017),
    .Y(_13269_));
 AO22x2_ASAP7_75t_R _42231_ (.A1(_10099_),
    .A2(_10126_),
    .B1(_10140_),
    .B2(_13269_),
    .Y(_13270_));
 AO21x2_ASAP7_75t_R _42232_ (.A1(net2382),
    .A2(_10126_),
    .B(_10112_),
    .Y(_13271_));
 INVx1_ASAP7_75t_R _42233_ (.A(_10266_),
    .Y(_13272_));
 OAI21x1_ASAP7_75t_R _42234_ (.A1(net1167),
    .A2(_13272_),
    .B(_10241_),
    .Y(_13273_));
 NOR3x2_ASAP7_75t_R _42235_ (.B(_13271_),
    .C(_13273_),
    .Y(_13275_),
    .A(_13270_));
 NAND2x2_ASAP7_75t_R _42236_ (.A(_13268_),
    .B(_13275_),
    .Y(_13276_));
 NOR2x1_ASAP7_75t_R _42237_ (.A(_13041_),
    .B(_11579_),
    .Y(_13277_));
 AND2x2_ASAP7_75t_R _42238_ (.A(_11251_),
    .B(_11559_),
    .Y(_13278_));
 NAND2x1_ASAP7_75t_R _42239_ (.A(_13277_),
    .B(_13278_),
    .Y(_13279_));
 NOR2x1_ASAP7_75t_R _42240_ (.A(_10040_),
    .B(_10015_),
    .Y(_13280_));
 NOR2x1_ASAP7_75t_R _42241_ (.A(_09965_),
    .B(_13280_),
    .Y(_13281_));
 OAI21x1_ASAP7_75t_R _42242_ (.A1(_10085_),
    .A2(_10246_),
    .B(_11222_),
    .Y(_13282_));
 INVx1_ASAP7_75t_R _42243_ (.A(_13282_),
    .Y(_13283_));
 NAND2x1_ASAP7_75t_R _42244_ (.A(_13281_),
    .B(_13283_),
    .Y(_13284_));
 NOR2x1_ASAP7_75t_R _42245_ (.A(_13279_),
    .B(_13284_),
    .Y(_13286_));
 OAI21x1_ASAP7_75t_R _42246_ (.A1(_10042_),
    .A2(_10246_),
    .B(_10165_),
    .Y(_13287_));
 OAI21x1_ASAP7_75t_R _42247_ (.A1(_09901_),
    .A2(_09988_),
    .B(_10211_),
    .Y(_13288_));
 NOR2x1_ASAP7_75t_R _42248_ (.A(_13287_),
    .B(_13288_),
    .Y(_13289_));
 OAI21x1_ASAP7_75t_R _42249_ (.A1(net1705),
    .A2(_10011_),
    .B(_10278_),
    .Y(_13290_));
 NOR2x1_ASAP7_75t_R _42250_ (.A(_10070_),
    .B(_10085_),
    .Y(_13291_));
 NOR2x1_ASAP7_75t_R _42251_ (.A(_13291_),
    .B(_11622_),
    .Y(_13292_));
 INVx1_ASAP7_75t_R _42252_ (.A(_13292_),
    .Y(_13293_));
 NOR2x1_ASAP7_75t_R _42253_ (.A(_13290_),
    .B(_13293_),
    .Y(_13294_));
 NAND2x1_ASAP7_75t_R _42254_ (.A(_13289_),
    .B(_13294_),
    .Y(_13295_));
 INVx1_ASAP7_75t_R _42255_ (.A(_13295_),
    .Y(_13297_));
 NAND2x1_ASAP7_75t_R _42256_ (.A(_13286_),
    .B(_13297_),
    .Y(_13298_));
 NOR2x1_ASAP7_75t_R _42257_ (.A(_13276_),
    .B(_13298_),
    .Y(_13299_));
 AO21x1_ASAP7_75t_R _42258_ (.A1(_10008_),
    .A2(net1757),
    .B(_10035_),
    .Y(_13300_));
 AND2x2_ASAP7_75t_R _42259_ (.A(_13300_),
    .B(_12320_),
    .Y(_13301_));
 OA21x2_ASAP7_75t_R _42260_ (.A1(_09913_),
    .A2(net2660),
    .B(_12451_),
    .Y(_13302_));
 AND3x1_ASAP7_75t_R _42261_ (.A(_13301_),
    .B(_11591_),
    .C(_13302_),
    .Y(_13303_));
 OAI21x1_ASAP7_75t_R _42262_ (.A1(_10107_),
    .A2(_10048_),
    .B(_12372_),
    .Y(_13304_));
 NAND2x1_ASAP7_75t_R _42263_ (.A(_10133_),
    .B(_11212_),
    .Y(_13305_));
 OAI21x1_ASAP7_75t_R _42264_ (.A1(net2444),
    .A2(net2662),
    .B(_13305_),
    .Y(_13306_));
 NOR2x1_ASAP7_75t_R _42265_ (.A(_13304_),
    .B(_13306_),
    .Y(_13308_));
 NAND2x1_ASAP7_75t_R _42266_ (.A(_11571_),
    .B(net2804),
    .Y(_13309_));
 OAI21x1_ASAP7_75t_R _42267_ (.A1(net2925),
    .A2(net2808),
    .B(_13309_),
    .Y(_13310_));
 NAND2x1_ASAP7_75t_R _42268_ (.A(_10080_),
    .B(_09943_),
    .Y(_13311_));
 OAI21x1_ASAP7_75t_R _42269_ (.A1(_10003_),
    .A2(net2662),
    .B(_13311_),
    .Y(_13312_));
 NOR2x2_ASAP7_75t_R _42270_ (.A(_13310_),
    .B(_13312_),
    .Y(_13313_));
 NAND2x1_ASAP7_75t_R _42271_ (.A(_13308_),
    .B(_13313_),
    .Y(_13314_));
 NAND2x1_ASAP7_75t_R _42272_ (.A(_12356_),
    .B(_10201_),
    .Y(_13315_));
 NOR2x1_ASAP7_75t_R _42273_ (.A(_13315_),
    .B(_13314_),
    .Y(_13316_));
 NAND2x2_ASAP7_75t_R _42274_ (.A(_13303_),
    .B(_13316_),
    .Y(_13317_));
 INVx1_ASAP7_75t_R _42275_ (.A(_13317_),
    .Y(_13319_));
 NAND2x2_ASAP7_75t_R _42276_ (.A(_13299_),
    .B(_13319_),
    .Y(_13320_));
 AO21x1_ASAP7_75t_R _42277_ (.A1(net2382),
    .A2(_09905_),
    .B(net3015),
    .Y(_13321_));
 OAI22x1_ASAP7_75t_R _42278_ (.A1(_13321_),
    .A2(_11593_),
    .B1(net1019),
    .B2(_11282_),
    .Y(_13322_));
 OA211x2_ASAP7_75t_R _42279_ (.A1(net2353),
    .A2(net1661),
    .B(_12380_),
    .C(_12348_),
    .Y(_13323_));
 NAND2x1_ASAP7_75t_R _42280_ (.A(_13322_),
    .B(_13323_),
    .Y(_13324_));
 NAND2x1_ASAP7_75t_R _42281_ (.A(_11261_),
    .B(_09947_),
    .Y(_13325_));
 NOR2x1_ASAP7_75t_R _42282_ (.A(_11580_),
    .B(_13325_),
    .Y(_13326_));
 AND3x1_ASAP7_75t_R _42283_ (.A(_13326_),
    .B(_10293_),
    .C(_11234_),
    .Y(_13327_));
 INVx1_ASAP7_75t_R _42284_ (.A(_13327_),
    .Y(_13328_));
 NOR2x1_ASAP7_75t_R _42285_ (.A(_13324_),
    .B(_13328_),
    .Y(_13330_));
 NOR2x1_ASAP7_75t_R _42286_ (.A(_10070_),
    .B(net2358),
    .Y(_13331_));
 AOI21x1_ASAP7_75t_R _42287_ (.A1(net3015),
    .A2(_13031_),
    .B(_13331_),
    .Y(_13332_));
 AOI21x1_ASAP7_75t_R _42288_ (.A1(net3015),
    .A2(_13075_),
    .B(_11637_),
    .Y(_13333_));
 NAND2x2_ASAP7_75t_R _42289_ (.A(_13332_),
    .B(_13333_),
    .Y(_13334_));
 AO21x1_ASAP7_75t_R _42290_ (.A1(_11656_),
    .A2(_09881_),
    .B(_11286_),
    .Y(_13335_));
 AO21x1_ASAP7_75t_R _42291_ (.A1(_10063_),
    .A2(net948),
    .B(_09901_),
    .Y(_13336_));
 NAND2x2_ASAP7_75t_R _42292_ (.A(_11628_),
    .B(_13336_),
    .Y(_13337_));
 NOR3x2_ASAP7_75t_R _42293_ (.B(_13335_),
    .C(_13337_),
    .Y(_13338_),
    .A(_13334_));
 OA21x2_ASAP7_75t_R _42294_ (.A1(_09883_),
    .A2(net2627),
    .B(_10030_),
    .Y(_13339_));
 NOR2x1_ASAP7_75t_R _42295_ (.A(net3309),
    .B(_10240_),
    .Y(_13341_));
 NOR2x1_ASAP7_75t_R _42296_ (.A(net2662),
    .B(net2357),
    .Y(_13342_));
 OR3x1_ASAP7_75t_R _42297_ (.A(_13339_),
    .B(_13341_),
    .C(_13342_),
    .Y(_13343_));
 NAND2x1_ASAP7_75t_R _42298_ (.A(_13074_),
    .B(_10107_),
    .Y(_13344_));
 AOI22x1_ASAP7_75t_R _42299_ (.A1(_13344_),
    .A2(_10099_),
    .B1(net2383),
    .B2(_10264_),
    .Y(_13345_));
 AO21x1_ASAP7_75t_R _42300_ (.A1(_10063_),
    .A2(_09928_),
    .B(net2253),
    .Y(_13346_));
 OA21x2_ASAP7_75t_R _42301_ (.A1(net2808),
    .A2(_10246_),
    .B(_13346_),
    .Y(_13347_));
 NAND2x1_ASAP7_75t_R _42302_ (.A(_13345_),
    .B(_13347_),
    .Y(_13348_));
 NOR2x1_ASAP7_75t_R _42303_ (.A(_13343_),
    .B(_13348_),
    .Y(_13349_));
 NAND2x2_ASAP7_75t_R _42304_ (.A(_13338_),
    .B(_13349_),
    .Y(_13350_));
 INVx2_ASAP7_75t_R _42305_ (.A(_13350_),
    .Y(_13352_));
 NAND2x2_ASAP7_75t_R _42306_ (.A(_13352_),
    .B(_13330_),
    .Y(_13353_));
 INVx1_ASAP7_75t_R _42307_ (.A(_10300_),
    .Y(_13354_));
 NOR3x2_ASAP7_75t_R _42308_ (.B(_13353_),
    .C(_13354_),
    .Y(_13355_),
    .A(_13320_));
 NAND2x2_ASAP7_75t_R _42309_ (.A(net1434),
    .B(_13355_),
    .Y(_13356_));
 NOR2x1_ASAP7_75t_R _42310_ (.A(_13262_),
    .B(_13229_),
    .Y(_13357_));
 NAND2x2_ASAP7_75t_R _42311_ (.A(_09628_),
    .B(_13357_),
    .Y(_13358_));
 INVx1_ASAP7_75t_R _42312_ (.A(_13273_),
    .Y(_13359_));
 NOR2x1_ASAP7_75t_R _42313_ (.A(_13271_),
    .B(_13270_),
    .Y(_13360_));
 NAND2x2_ASAP7_75t_R _42314_ (.A(_13359_),
    .B(_13360_),
    .Y(_13361_));
 INVx1_ASAP7_75t_R _42315_ (.A(_13268_),
    .Y(_13363_));
 NOR2x2_ASAP7_75t_R _42316_ (.A(_13361_),
    .B(_13363_),
    .Y(_13364_));
 INVx1_ASAP7_75t_R _42317_ (.A(_13286_),
    .Y(_13365_));
 NOR2x1_ASAP7_75t_R _42318_ (.A(_13295_),
    .B(_13365_),
    .Y(_13366_));
 NAND2x1_ASAP7_75t_R _42319_ (.A(_13364_),
    .B(_13366_),
    .Y(_13367_));
 NOR2x2_ASAP7_75t_R _42320_ (.A(_13317_),
    .B(_13367_),
    .Y(_13368_));
 INVx1_ASAP7_75t_R _42321_ (.A(_13324_),
    .Y(_13369_));
 NAND2x1_ASAP7_75t_R _42322_ (.A(_13327_),
    .B(_13369_),
    .Y(_13370_));
 NOR2x2_ASAP7_75t_R _42323_ (.A(_13350_),
    .B(_13370_),
    .Y(_13371_));
 NAND3x2_ASAP7_75t_R _42324_ (.B(_13371_),
    .C(_10300_),
    .Y(_13372_),
    .A(_13368_));
 NAND2x2_ASAP7_75t_R _42325_ (.A(_13358_),
    .B(_13372_),
    .Y(_13374_));
 NOR2x1_ASAP7_75t_R _42326_ (.A(_10453_),
    .B(_10363_),
    .Y(_13375_));
 NAND2x2_ASAP7_75t_R _42327_ (.A(net2727),
    .B(_13375_),
    .Y(_13376_));
 OA21x2_ASAP7_75t_R _42328_ (.A1(net3291),
    .A2(_10554_),
    .B(_10537_),
    .Y(_13377_));
 AOI211x1_ASAP7_75t_R _42329_ (.A1(_11341_),
    .A2(_10537_),
    .B(_13377_),
    .C(_12675_),
    .Y(_13378_));
 AO21x2_ASAP7_75t_R _42330_ (.A1(_11323_),
    .A2(net3335),
    .B(_10546_),
    .Y(_13379_));
 AO21x1_ASAP7_75t_R _42331_ (.A1(net1115),
    .A2(_10502_),
    .B(_10546_),
    .Y(_13380_));
 AO21x1_ASAP7_75t_R _42332_ (.A1(net3051),
    .A2(net1659),
    .B(_10546_),
    .Y(_13381_));
 AO21x1_ASAP7_75t_R _42333_ (.A1(_10505_),
    .A2(net1051),
    .B(_10546_),
    .Y(_13382_));
 AND4x1_ASAP7_75t_R _42334_ (.A(_13379_),
    .B(_13380_),
    .C(_13381_),
    .D(_13382_),
    .Y(_13383_));
 NAND2x1_ASAP7_75t_R _42335_ (.A(_13378_),
    .B(_13383_),
    .Y(_13385_));
 AO21x1_ASAP7_75t_R _42336_ (.A1(net1115),
    .A2(net3318),
    .B(net2228),
    .Y(_13386_));
 AO21x1_ASAP7_75t_R _42337_ (.A1(net3157),
    .A2(net1125),
    .B(net2228),
    .Y(_13387_));
 AO21x1_ASAP7_75t_R _42338_ (.A1(_10505_),
    .A2(net1517),
    .B(net2228),
    .Y(_13388_));
 AND3x1_ASAP7_75t_R _42339_ (.A(_13386_),
    .B(_13387_),
    .C(_13388_),
    .Y(_13389_));
 AO21x1_ASAP7_75t_R _42340_ (.A1(_10459_),
    .A2(_10410_),
    .B(_11355_),
    .Y(_13390_));
 OA211x2_ASAP7_75t_R _42341_ (.A1(_11323_),
    .A2(_11355_),
    .B(_11940_),
    .C(_13390_),
    .Y(_13391_));
 NAND2x1_ASAP7_75t_R _42342_ (.A(_13389_),
    .B(_13391_),
    .Y(_13392_));
 NOR2x1_ASAP7_75t_R _42343_ (.A(_13385_),
    .B(_13392_),
    .Y(_13393_));
 NOR2x1_ASAP7_75t_R _42344_ (.A(_10367_),
    .B(net966),
    .Y(_13394_));
 OA21x2_ASAP7_75t_R _42345_ (.A1(_13394_),
    .A2(_10597_),
    .B(_10601_),
    .Y(_13396_));
 NOR3x1_ASAP7_75t_R _42346_ (.A(_11530_),
    .B(_13396_),
    .C(_11919_),
    .Y(_13397_));
 OA211x2_ASAP7_75t_R _42347_ (.A1(_10367_),
    .A2(net3338),
    .B(_10589_),
    .C(net1885),
    .Y(_13398_));
 INVx1_ASAP7_75t_R _42348_ (.A(_13398_),
    .Y(_13399_));
 AO21x1_ASAP7_75t_R _42349_ (.A1(net3051),
    .A2(net1077),
    .B(net2227),
    .Y(_13400_));
 NAND3x1_ASAP7_75t_R _42350_ (.A(_13397_),
    .B(_13399_),
    .C(_13400_),
    .Y(_13401_));
 AO21x1_ASAP7_75t_R _42351_ (.A1(_11323_),
    .A2(net1125),
    .B(net1840),
    .Y(_13402_));
 AO21x1_ASAP7_75t_R _42352_ (.A1(net3051),
    .A2(net1659),
    .B(net1840),
    .Y(_13403_));
 AO21x1_ASAP7_75t_R _42353_ (.A1(net1115),
    .A2(_10502_),
    .B(net1840),
    .Y(_13404_));
 NAND2x1_ASAP7_75t_R _42354_ (.A(net3034),
    .B(_10579_),
    .Y(_13405_));
 AND4x1_ASAP7_75t_R _42355_ (.A(_13402_),
    .B(_13403_),
    .C(_13404_),
    .D(_13405_),
    .Y(_13407_));
 AO21x1_ASAP7_75t_R _42356_ (.A1(net1659),
    .A2(_11312_),
    .B(net2211),
    .Y(_13408_));
 AO21x1_ASAP7_75t_R _42357_ (.A1(net2463),
    .A2(net1306),
    .B(net2211),
    .Y(_13409_));
 OA211x2_ASAP7_75t_R _42358_ (.A1(net1144),
    .A2(net2211),
    .B(_13408_),
    .C(_13409_),
    .Y(_13410_));
 NAND2x1_ASAP7_75t_R _42359_ (.A(_13407_),
    .B(_13410_),
    .Y(_13411_));
 NOR2x1_ASAP7_75t_R _42360_ (.A(_13401_),
    .B(_13411_),
    .Y(_13412_));
 NAND2x1_ASAP7_75t_R _42361_ (.A(_13412_),
    .B(_13393_),
    .Y(_13413_));
 AO21x1_ASAP7_75t_R _42362_ (.A1(net2463),
    .A2(net1125),
    .B(net1881),
    .Y(_13414_));
 AO21x1_ASAP7_75t_R _42363_ (.A1(net2954),
    .A2(net1055),
    .B(net1881),
    .Y(_13415_));
 INVx1_ASAP7_75t_R _42364_ (.A(_12965_),
    .Y(_13416_));
 AND3x1_ASAP7_75t_R _42365_ (.A(_13414_),
    .B(_13415_),
    .C(_13416_),
    .Y(_13418_));
 NAND2x2_ASAP7_75t_R _42366_ (.A(_10367_),
    .B(_11488_),
    .Y(_13419_));
 AO21x1_ASAP7_75t_R _42367_ (.A1(_11364_),
    .A2(net3298),
    .B(net2329),
    .Y(_13420_));
 AND3x1_ASAP7_75t_R _42368_ (.A(_13419_),
    .B(_11957_),
    .C(_13420_),
    .Y(_13421_));
 NAND2x2_ASAP7_75t_R _42369_ (.A(_13418_),
    .B(_13421_),
    .Y(_13422_));
 AO21x1_ASAP7_75t_R _42370_ (.A1(net2957),
    .A2(_10410_),
    .B(_10358_),
    .Y(_13423_));
 AO21x1_ASAP7_75t_R _42371_ (.A1(net1115),
    .A2(net1306),
    .B(_10358_),
    .Y(_13424_));
 AND3x1_ASAP7_75t_R _42372_ (.A(_11971_),
    .B(_13424_),
    .C(_11969_),
    .Y(_13425_));
 NAND2x2_ASAP7_75t_R _42373_ (.A(_13423_),
    .B(_13425_),
    .Y(_13426_));
 NAND3x2_ASAP7_75t_R _42374_ (.B(_10345_),
    .C(_10351_),
    .Y(_13427_),
    .A(_11475_));
 NOR3x2_ASAP7_75t_R _42375_ (.B(_13426_),
    .C(_13427_),
    .Y(_13429_),
    .A(_13422_));
 AO21x1_ASAP7_75t_R _42376_ (.A1(_10502_),
    .A2(net3318),
    .B(net2020),
    .Y(_13430_));
 AO21x1_ASAP7_75t_R _42377_ (.A1(_10459_),
    .A2(net2954),
    .B(net2020),
    .Y(_13431_));
 AO21x1_ASAP7_75t_R _42378_ (.A1(_10421_),
    .A2(net1125),
    .B(net2020),
    .Y(_13432_));
 AND3x1_ASAP7_75t_R _42379_ (.A(_13430_),
    .B(_13431_),
    .C(_13432_),
    .Y(_13433_));
 AO21x1_ASAP7_75t_R _42380_ (.A1(_11323_),
    .A2(_10420_),
    .B(net2233),
    .Y(_13434_));
 OA211x2_ASAP7_75t_R _42381_ (.A1(net1306),
    .A2(net2233),
    .B(_13434_),
    .C(_12744_),
    .Y(_13435_));
 NAND2x1_ASAP7_75t_R _42382_ (.A(_13433_),
    .B(_13435_),
    .Y(_13436_));
 NAND2x1_ASAP7_75t_R _42383_ (.A(_10492_),
    .B(_11976_),
    .Y(_13437_));
 OA211x2_ASAP7_75t_R _42384_ (.A1(_10327_),
    .A2(net975),
    .B(_10483_),
    .C(net3319),
    .Y(_13438_));
 NOR2x1_ASAP7_75t_R _42385_ (.A(_13437_),
    .B(_13438_),
    .Y(_13440_));
 AO21x1_ASAP7_75t_R _42386_ (.A1(net1115),
    .A2(net1414),
    .B(net2249),
    .Y(_13441_));
 AO21x1_ASAP7_75t_R _42387_ (.A1(net3051),
    .A2(net1659),
    .B(net2249),
    .Y(_13442_));
 OA211x2_ASAP7_75t_R _42388_ (.A1(net1876),
    .A2(net2249),
    .B(_13441_),
    .C(_13442_),
    .Y(_13443_));
 NAND2x1_ASAP7_75t_R _42389_ (.A(_13440_),
    .B(_13443_),
    .Y(_13444_));
 NOR2x1_ASAP7_75t_R _42390_ (.A(_13436_),
    .B(_13444_),
    .Y(_13445_));
 NAND2x2_ASAP7_75t_R _42391_ (.A(_13429_),
    .B(_13445_),
    .Y(_13446_));
 NOR2x2_ASAP7_75t_R _42392_ (.A(_13413_),
    .B(_13446_),
    .Y(_13447_));
 NAND2x2_ASAP7_75t_R _42393_ (.A(_13376_),
    .B(_13447_),
    .Y(_13448_));
 INVx1_ASAP7_75t_R _42394_ (.A(_13448_),
    .Y(_13449_));
 AO21x1_ASAP7_75t_R _42395_ (.A1(_13356_),
    .A2(_13374_),
    .B(_13449_),
    .Y(_13451_));
 NAND2x2_ASAP7_75t_R _42396_ (.A(_13358_),
    .B(_13355_),
    .Y(_13452_));
 NAND2x2_ASAP7_75t_R _42397_ (.A(net1434),
    .B(_13372_),
    .Y(_13453_));
 AO21x1_ASAP7_75t_R _42398_ (.A1(_13452_),
    .A2(_13453_),
    .B(_13448_),
    .Y(_13454_));
 AOI211x1_ASAP7_75t_R _42399_ (.A1(_10626_),
    .A2(_10658_),
    .B(net3040),
    .C(net2025),
    .Y(_13455_));
 NOR2x1_ASAP7_75t_R _42400_ (.A(_10854_),
    .B(net3040),
    .Y(_13456_));
 AOI211x1_ASAP7_75t_R _42401_ (.A1(_12643_),
    .A2(_10774_),
    .B(_13455_),
    .C(_13456_),
    .Y(_13457_));
 AO21x1_ASAP7_75t_R _42402_ (.A1(_10767_),
    .A2(net1982),
    .B(_10755_),
    .Y(_13458_));
 AND2x2_ASAP7_75t_R _42403_ (.A(_13458_),
    .B(_12646_),
    .Y(_13459_));
 NAND3x2_ASAP7_75t_R _42404_ (.B(_10956_),
    .C(_13459_),
    .Y(_13460_),
    .A(_13457_));
 NAND2x1_ASAP7_75t_R _42405_ (.A(_12915_),
    .B(_11783_),
    .Y(_13462_));
 AO21x1_ASAP7_75t_R _42406_ (.A1(net1288),
    .A2(net3058),
    .B(_10725_),
    .Y(_13463_));
 OAI21x1_ASAP7_75t_R _42407_ (.A1(net1424),
    .A2(_10966_),
    .B(_13463_),
    .Y(_13464_));
 NOR2x1_ASAP7_75t_R _42408_ (.A(_13462_),
    .B(_13464_),
    .Y(_13465_));
 OA31x2_ASAP7_75t_R _42409_ (.A1(_10708_),
    .A2(_11851_),
    .A3(net3061),
    .B1(_12664_),
    .Y(_13466_));
 AO21x1_ASAP7_75t_R _42410_ (.A1(_11853_),
    .A2(_12664_),
    .B(_10971_),
    .Y(_13467_));
 NOR3x1_ASAP7_75t_R _42411_ (.A(_13466_),
    .B(_10974_),
    .C(_13467_),
    .Y(_13468_));
 NAND2x1_ASAP7_75t_R _42412_ (.A(_13465_),
    .B(_13468_),
    .Y(_13469_));
 NOR2x2_ASAP7_75t_R _42413_ (.A(_13460_),
    .B(_13469_),
    .Y(_13470_));
 AOI221x1_ASAP7_75t_R _42414_ (.A1(net1501),
    .A2(_10658_),
    .B1(_10740_),
    .B2(_10732_),
    .C(net3021),
    .Y(_13471_));
 OR3x2_ASAP7_75t_R _42415_ (.A(_11825_),
    .B(_12940_),
    .C(_13471_),
    .Y(_13473_));
 AO21x1_ASAP7_75t_R _42416_ (.A1(net1288),
    .A2(net3049),
    .B(net3045),
    .Y(_13474_));
 AO21x1_ASAP7_75t_R _42417_ (.A1(_10788_),
    .A2(_10700_),
    .B(net3045),
    .Y(_13475_));
 NAND2x1_ASAP7_75t_R _42418_ (.A(_13474_),
    .B(_13475_),
    .Y(_13476_));
 OR3x2_ASAP7_75t_R _42419_ (.A(_13476_),
    .B(_10688_),
    .C(_12923_),
    .Y(_13477_));
 AO21x1_ASAP7_75t_R _42420_ (.A1(net1492),
    .A2(_10740_),
    .B(_10696_),
    .Y(_13478_));
 OA21x2_ASAP7_75t_R _42421_ (.A1(_10696_),
    .A2(_10678_),
    .B(_13478_),
    .Y(_13479_));
 AOI21x1_ASAP7_75t_R _42422_ (.A1(_10701_),
    .A2(_10732_),
    .B(_10705_),
    .Y(_13480_));
 INVx1_ASAP7_75t_R _42423_ (.A(_10938_),
    .Y(_13481_));
 OA21x2_ASAP7_75t_R _42424_ (.A1(_13481_),
    .A2(_11798_),
    .B(_10713_),
    .Y(_13482_));
 NOR2x1_ASAP7_75t_R _42425_ (.A(_13480_),
    .B(_13482_),
    .Y(_13484_));
 NAND2x2_ASAP7_75t_R _42426_ (.A(_13479_),
    .B(_13484_),
    .Y(_13485_));
 NOR3x2_ASAP7_75t_R _42427_ (.B(_13477_),
    .C(_13485_),
    .Y(_13486_),
    .A(_13473_));
 NAND2x2_ASAP7_75t_R _42428_ (.A(_13470_),
    .B(_13486_),
    .Y(_13487_));
 AND3x1_ASAP7_75t_R _42429_ (.A(_10901_),
    .B(_10791_),
    .C(net1336),
    .Y(_13488_));
 AOI211x1_ASAP7_75t_R _42430_ (.A1(_10791_),
    .A2(_10733_),
    .B(_13488_),
    .C(_12594_),
    .Y(_13489_));
 NAND2x1_ASAP7_75t_R _42431_ (.A(_10791_),
    .B(_12643_),
    .Y(_13490_));
 AO21x1_ASAP7_75t_R _42432_ (.A1(_10783_),
    .A2(_11039_),
    .B(_10796_),
    .Y(_13491_));
 AND2x2_ASAP7_75t_R _42433_ (.A(_13491_),
    .B(_10804_),
    .Y(_13492_));
 NAND3x1_ASAP7_75t_R _42434_ (.A(_13489_),
    .B(_13490_),
    .C(_13492_),
    .Y(_13493_));
 AO21x1_ASAP7_75t_R _42435_ (.A1(_10783_),
    .A2(net3053),
    .B(_10810_),
    .Y(_13495_));
 NAND2x1_ASAP7_75t_R _42436_ (.A(_11008_),
    .B(_10809_),
    .Y(_13496_));
 NAND2x1_ASAP7_75t_R _42437_ (.A(net3061),
    .B(_10809_),
    .Y(_13497_));
 AND3x1_ASAP7_75t_R _42438_ (.A(_13495_),
    .B(_13496_),
    .C(_13497_),
    .Y(_13498_));
 AO221x1_ASAP7_75t_R _42439_ (.A1(_10740_),
    .A2(_10732_),
    .B1(_10684_),
    .B2(_10710_),
    .C(_10810_),
    .Y(_13499_));
 OA21x2_ASAP7_75t_R _42440_ (.A1(_10708_),
    .A2(_10996_),
    .B(_10992_),
    .Y(_13500_));
 AOI211x1_ASAP7_75t_R _42441_ (.A1(net1501),
    .A2(_10658_),
    .B(net3056),
    .C(_10732_),
    .Y(_13501_));
 AOI211x1_ASAP7_75t_R _42442_ (.A1(_10626_),
    .A2(_10658_),
    .B(net3056),
    .C(_10740_),
    .Y(_13502_));
 NOR3x1_ASAP7_75t_R _42443_ (.A(_13500_),
    .B(_13501_),
    .C(_13502_),
    .Y(_13503_));
 NAND3x1_ASAP7_75t_R _42444_ (.A(_13498_),
    .B(_13499_),
    .C(_13503_),
    .Y(_13504_));
 NOR2x1_ASAP7_75t_R _42445_ (.A(_13493_),
    .B(_13504_),
    .Y(_13506_));
 AO21x1_ASAP7_75t_R _42446_ (.A1(_10767_),
    .A2(net1862),
    .B(net3029),
    .Y(_13507_));
 AO21x1_ASAP7_75t_R _42447_ (.A1(_10745_),
    .A2(net1288),
    .B(_10826_),
    .Y(_13508_));
 AND4x1_ASAP7_75t_R _42448_ (.A(_13507_),
    .B(_12259_),
    .C(_13508_),
    .D(_12893_),
    .Y(_13509_));
 AO21x1_ASAP7_75t_R _42449_ (.A1(net1862),
    .A2(net1991),
    .B(net3054),
    .Y(_13510_));
 OA211x2_ASAP7_75t_R _42450_ (.A1(_10807_),
    .A2(net3054),
    .B(_13510_),
    .C(_10871_),
    .Y(_13511_));
 NAND2x1_ASAP7_75t_R _42451_ (.A(_13509_),
    .B(_13511_),
    .Y(_13512_));
 AO21x1_ASAP7_75t_R _42452_ (.A1(net1446),
    .A2(_10701_),
    .B(_10843_),
    .Y(_13513_));
 AO21x1_ASAP7_75t_R _42453_ (.A1(_11039_),
    .A2(net1982),
    .B(_10843_),
    .Y(_13514_));
 OA211x2_ASAP7_75t_R _42454_ (.A1(net3053),
    .A2(_10843_),
    .B(_13513_),
    .C(_13514_),
    .Y(_13515_));
 AO21x1_ASAP7_75t_R _42455_ (.A1(_10783_),
    .A2(net3053),
    .B(net3033),
    .Y(_13517_));
 AO21x1_ASAP7_75t_R _42456_ (.A1(net3049),
    .A2(net1492),
    .B(net3033),
    .Y(_13518_));
 OA211x2_ASAP7_75t_R _42457_ (.A1(net3033),
    .A2(_10671_),
    .B(_13517_),
    .C(_13518_),
    .Y(_13519_));
 NAND2x1_ASAP7_75t_R _42458_ (.A(_13515_),
    .B(_13519_),
    .Y(_13520_));
 NOR2x2_ASAP7_75t_R _42459_ (.A(_13512_),
    .B(_13520_),
    .Y(_13521_));
 NAND2x2_ASAP7_75t_R _42460_ (.A(_13506_),
    .B(_13521_),
    .Y(_13522_));
 NOR3x2_ASAP7_75t_R _42461_ (.B(_13522_),
    .C(_11885_),
    .Y(_13523_),
    .A(_13487_));
 XOR2x1_ASAP7_75t_R _42462_ (.A(_13523_),
    .Y(_13524_),
    .B(net2054));
 INVx1_ASAP7_75t_R _42463_ (.A(_13524_),
    .Y(_13525_));
 AOI21x1_ASAP7_75t_R _42464_ (.A1(_13451_),
    .A2(_13454_),
    .B(_13525_),
    .Y(_13526_));
 AO21x1_ASAP7_75t_R _42465_ (.A1(_13452_),
    .A2(_13453_),
    .B(_13449_),
    .Y(_13528_));
 AO21x1_ASAP7_75t_R _42466_ (.A1(_13356_),
    .A2(_13374_),
    .B(_13448_),
    .Y(_13529_));
 AOI21x1_ASAP7_75t_R _42467_ (.A1(_13528_),
    .A2(_13529_),
    .B(_13524_),
    .Y(_13530_));
 OAI21x1_ASAP7_75t_R _42468_ (.A1(_13526_),
    .A2(_13530_),
    .B(net392),
    .Y(_13531_));
 INVx1_ASAP7_75t_R _42469_ (.A(_13531_),
    .Y(_13532_));
 OAI21x1_ASAP7_75t_R _42470_ (.A1(_13191_),
    .A2(_13532_),
    .B(_00411_),
    .Y(_13533_));
 INVx1_ASAP7_75t_R _42471_ (.A(_13191_),
    .Y(_13534_));
 NAND3x1_ASAP7_75t_R _42472_ (.A(_13531_),
    .B(_17450_),
    .C(_13534_),
    .Y(_13535_));
 NAND2x1_ASAP7_75t_R _42473_ (.A(_13535_),
    .B(_13533_),
    .Y(_00103_));
 NAND2x2_ASAP7_75t_R _42474_ (.A(_00812_),
    .B(net389),
    .Y(_13536_));
 AO21x1_ASAP7_75t_R _42475_ (.A1(net3020),
    .A2(net3058),
    .B(_10696_),
    .Y(_13538_));
 NOR2x1_ASAP7_75t_R _42476_ (.A(_10696_),
    .B(_10693_),
    .Y(_13539_));
 INVx1_ASAP7_75t_R _42477_ (.A(_13539_),
    .Y(_13540_));
 AND3x1_ASAP7_75t_R _42478_ (.A(_13538_),
    .B(_13540_),
    .C(_11809_),
    .Y(_13541_));
 INVx1_ASAP7_75t_R _42479_ (.A(_10714_),
    .Y(_13542_));
 AO21x1_ASAP7_75t_R _42480_ (.A1(_10700_),
    .A2(_10656_),
    .B(_10705_),
    .Y(_13543_));
 AND3x1_ASAP7_75t_R _42481_ (.A(_13542_),
    .B(_12621_),
    .C(_13543_),
    .Y(_13544_));
 NAND2x2_ASAP7_75t_R _42482_ (.A(_13541_),
    .B(_13544_),
    .Y(_13545_));
 OA21x2_ASAP7_75t_R _42483_ (.A1(_10831_),
    .A2(_10733_),
    .B(_10642_),
    .Y(_13546_));
 OR4x2_ASAP7_75t_R _42484_ (.A(_10904_),
    .B(_13546_),
    .C(_10688_),
    .D(_12629_),
    .Y(_13547_));
 NOR2x1_ASAP7_75t_R _42485_ (.A(_10985_),
    .B(_12227_),
    .Y(_13549_));
 INVx1_ASAP7_75t_R _42486_ (.A(_13549_),
    .Y(_13550_));
 NOR3x2_ASAP7_75t_R _42487_ (.B(_13547_),
    .C(_13550_),
    .Y(_13551_),
    .A(_13545_));
 AO21x1_ASAP7_75t_R _42488_ (.A1(_10767_),
    .A2(net1862),
    .B(_10755_),
    .Y(_13552_));
 AO21x1_ASAP7_75t_R _42489_ (.A1(_10745_),
    .A2(net1288),
    .B(_10755_),
    .Y(_13553_));
 AO21x1_ASAP7_75t_R _42490_ (.A1(_10938_),
    .A2(_10694_),
    .B(net3041),
    .Y(_13554_));
 AND4x2_ASAP7_75t_R _42491_ (.A(_13552_),
    .B(_13553_),
    .C(_13554_),
    .D(_12649_),
    .Y(_13555_));
 OA21x2_ASAP7_75t_R _42492_ (.A1(_10782_),
    .A2(_11008_),
    .B(_12664_),
    .Y(_13556_));
 NOR2x1_ASAP7_75t_R _42493_ (.A(_10739_),
    .B(net1446),
    .Y(_13557_));
 NOR2x1_ASAP7_75t_R _42494_ (.A(net1982),
    .B(_10739_),
    .Y(_13558_));
 OR4x2_ASAP7_75t_R _42495_ (.A(_13556_),
    .B(_10741_),
    .C(_13557_),
    .D(_13558_),
    .Y(_13560_));
 NAND2x1_ASAP7_75t_R _42496_ (.A(_10737_),
    .B(_12213_),
    .Y(_13561_));
 OA21x2_ASAP7_75t_R _42497_ (.A1(_12643_),
    .A2(_10681_),
    .B(_10736_),
    .Y(_13562_));
 OA21x2_ASAP7_75t_R _42498_ (.A1(_10792_),
    .A2(_11043_),
    .B(_10736_),
    .Y(_13563_));
 NOR2x1_ASAP7_75t_R _42499_ (.A(net3020),
    .B(_10725_),
    .Y(_13564_));
 OR4x2_ASAP7_75t_R _42500_ (.A(_13561_),
    .B(_13562_),
    .C(_13563_),
    .D(_13564_),
    .Y(_13565_));
 NOR2x2_ASAP7_75t_R _42501_ (.A(_13560_),
    .B(_13565_),
    .Y(_13566_));
 NAND3x2_ASAP7_75t_R _42502_ (.B(_13555_),
    .C(_13566_),
    .Y(_13567_),
    .A(_13551_));
 AO21x1_ASAP7_75t_R _42503_ (.A1(net3053),
    .A2(net1982),
    .B(net3030),
    .Y(_13568_));
 AO21x1_ASAP7_75t_R _42504_ (.A1(net1446),
    .A2(_10807_),
    .B(net3030),
    .Y(_13569_));
 OA21x2_ASAP7_75t_R _42505_ (.A1(net3020),
    .A2(net3030),
    .B(_13569_),
    .Y(_13571_));
 NAND2x1_ASAP7_75t_R _42506_ (.A(_13568_),
    .B(_13571_),
    .Y(_13572_));
 INVx1_ASAP7_75t_R _42507_ (.A(_13572_),
    .Y(_13573_));
 AO21x1_ASAP7_75t_R _42508_ (.A1(net1446),
    .A2(_10788_),
    .B(_10864_),
    .Y(_13574_));
 NOR2x1_ASAP7_75t_R _42509_ (.A(net3047),
    .B(_10864_),
    .Y(_13575_));
 INVx1_ASAP7_75t_R _42510_ (.A(_13575_),
    .Y(_13576_));
 AND2x2_ASAP7_75t_R _42511_ (.A(_13574_),
    .B(_13576_),
    .Y(_13577_));
 AO21x1_ASAP7_75t_R _42512_ (.A1(_10783_),
    .A2(net1475),
    .B(net3054),
    .Y(_13578_));
 AO21x1_ASAP7_75t_R _42513_ (.A1(net1862),
    .A2(_10671_),
    .B(net3054),
    .Y(_13579_));
 AND3x1_ASAP7_75t_R _42514_ (.A(_13577_),
    .B(_13578_),
    .C(_13579_),
    .Y(_13580_));
 NAND2x1_ASAP7_75t_R _42515_ (.A(_13573_),
    .B(_13580_),
    .Y(_13582_));
 NAND2x1_ASAP7_75t_R _42516_ (.A(_10869_),
    .B(_11860_),
    .Y(_13583_));
 NAND2x1_ASAP7_75t_R _42517_ (.A(_13583_),
    .B(_12249_),
    .Y(_13584_));
 OA211x2_ASAP7_75t_R _42518_ (.A1(_10626_),
    .A2(_10658_),
    .B(_10847_),
    .C(net2119),
    .Y(_13585_));
 NAND2x1_ASAP7_75t_R _42519_ (.A(_12586_),
    .B(_13517_),
    .Y(_13586_));
 AOI21x1_ASAP7_75t_R _42520_ (.A1(net1288),
    .A2(_10788_),
    .B(_10843_),
    .Y(_13587_));
 OR4x2_ASAP7_75t_R _42521_ (.A(_13584_),
    .B(_13585_),
    .C(_13586_),
    .D(_13587_),
    .Y(_13588_));
 NOR2x2_ASAP7_75t_R _42522_ (.A(_13582_),
    .B(_13588_),
    .Y(_13589_));
 INVx1_ASAP7_75t_R _42523_ (.A(_12874_),
    .Y(_13590_));
 AOI211x1_ASAP7_75t_R _42524_ (.A1(_11833_),
    .A2(_10996_),
    .B(_13590_),
    .C(_11836_),
    .Y(_13591_));
 OA21x2_ASAP7_75t_R _42525_ (.A1(_10658_),
    .A2(_11007_),
    .B(_10787_),
    .Y(_13593_));
 AO21x1_ASAP7_75t_R _42526_ (.A1(net1446),
    .A2(_10788_),
    .B(_10785_),
    .Y(_13594_));
 AO21x1_ASAP7_75t_R _42527_ (.A1(net3058),
    .A2(_10656_),
    .B(_10785_),
    .Y(_13595_));
 AND2x2_ASAP7_75t_R _42528_ (.A(_13594_),
    .B(_13595_),
    .Y(_13596_));
 AND3x1_ASAP7_75t_R _42529_ (.A(_13591_),
    .B(_13593_),
    .C(_13596_),
    .Y(_13597_));
 NOR2x1_ASAP7_75t_R _42530_ (.A(_10814_),
    .B(_12610_),
    .Y(_13598_));
 AND2x2_ASAP7_75t_R _42531_ (.A(_10831_),
    .B(_10809_),
    .Y(_13599_));
 INVx1_ASAP7_75t_R _42532_ (.A(_13599_),
    .Y(_13600_));
 INVx1_ASAP7_75t_R _42533_ (.A(_11854_),
    .Y(_13601_));
 AND3x1_ASAP7_75t_R _42534_ (.A(_13598_),
    .B(_13600_),
    .C(_13601_),
    .Y(_13602_));
 AO21x1_ASAP7_75t_R _42535_ (.A1(_10767_),
    .A2(net1862),
    .B(net3056),
    .Y(_13604_));
 AO21x1_ASAP7_75t_R _42536_ (.A1(_10682_),
    .A2(net1475),
    .B(net3056),
    .Y(_13605_));
 AO21x1_ASAP7_75t_R _42537_ (.A1(net3020),
    .A2(net1288),
    .B(net3056),
    .Y(_13606_));
 NAND2x1_ASAP7_75t_R _42538_ (.A(net1345),
    .B(_10992_),
    .Y(_13607_));
 AND4x1_ASAP7_75t_R _42539_ (.A(_13604_),
    .B(_13605_),
    .C(_13606_),
    .D(_13607_),
    .Y(_13608_));
 AND2x2_ASAP7_75t_R _42540_ (.A(_13602_),
    .B(_13608_),
    .Y(_13609_));
 NAND2x1_ASAP7_75t_R _42541_ (.A(_13597_),
    .B(_13609_),
    .Y(_13610_));
 INVx1_ASAP7_75t_R _42542_ (.A(_13610_),
    .Y(_13611_));
 NAND2x2_ASAP7_75t_R _42543_ (.A(_13589_),
    .B(_13611_),
    .Y(_13612_));
 NOR3x2_ASAP7_75t_R _42544_ (.B(_13612_),
    .C(_11885_),
    .Y(_13613_),
    .A(_13567_));
 AO21x1_ASAP7_75t_R _42545_ (.A1(_09658_),
    .A2(_09631_),
    .B(_09730_),
    .Y(_13615_));
 AND2x2_ASAP7_75t_R _42546_ (.A(_12131_),
    .B(_13615_),
    .Y(_13616_));
 AO21x1_ASAP7_75t_R _42547_ (.A1(_09711_),
    .A2(_09798_),
    .B(_09730_),
    .Y(_13617_));
 AO21x1_ASAP7_75t_R _42548_ (.A1(_09611_),
    .A2(_09739_),
    .B(_09730_),
    .Y(_13618_));
 AND2x2_ASAP7_75t_R _42549_ (.A(_13617_),
    .B(_13618_),
    .Y(_13619_));
 OA21x2_ASAP7_75t_R _42550_ (.A1(_09580_),
    .A2(_09582_),
    .B(_09846_),
    .Y(_13620_));
 AOI21x1_ASAP7_75t_R _42551_ (.A1(_09738_),
    .A2(_13205_),
    .B(_09649_),
    .Y(_13621_));
 NOR2x1_ASAP7_75t_R _42552_ (.A(_13620_),
    .B(_13621_),
    .Y(_13622_));
 NAND3x1_ASAP7_75t_R _42553_ (.A(_13616_),
    .B(_13619_),
    .C(_13622_),
    .Y(_13623_));
 AO221x1_ASAP7_75t_R _42554_ (.A1(_09589_),
    .A2(_09573_),
    .B1(net1477),
    .B2(_09597_),
    .C(_09682_),
    .Y(_13624_));
 AO21x1_ASAP7_75t_R _42555_ (.A1(_09769_),
    .A2(net2104),
    .B(net2339),
    .Y(_13626_));
 AO21x1_ASAP7_75t_R _42556_ (.A1(net2940),
    .A2(net2327),
    .B(net2339),
    .Y(_13627_));
 AND2x2_ASAP7_75t_R _42557_ (.A(_13626_),
    .B(_13627_),
    .Y(_13628_));
 NAND3x1_ASAP7_75t_R _42558_ (.A(_13624_),
    .B(_13211_),
    .C(_13628_),
    .Y(_13629_));
 NOR2x1_ASAP7_75t_R _42559_ (.A(_13623_),
    .B(_13629_),
    .Y(_13630_));
 AO21x1_ASAP7_75t_R _42560_ (.A1(_09714_),
    .A2(net2104),
    .B(net2922),
    .Y(_13631_));
 AO21x1_ASAP7_75t_R _42561_ (.A1(net1561),
    .A2(net2937),
    .B(net2922),
    .Y(_13632_));
 NAND2x1_ASAP7_75t_R _42562_ (.A(_13631_),
    .B(_13632_),
    .Y(_13633_));
 AO21x1_ASAP7_75t_R _42563_ (.A1(_09658_),
    .A2(_09631_),
    .B(net2922),
    .Y(_13634_));
 OAI21x1_ASAP7_75t_R _42564_ (.A1(net2922),
    .A2(_09772_),
    .B(_13634_),
    .Y(_13635_));
 NOR2x1_ASAP7_75t_R _42565_ (.A(_13633_),
    .B(_13635_),
    .Y(_13637_));
 NAND2x1_ASAP7_75t_R _42566_ (.A(_12045_),
    .B(_13125_),
    .Y(_13638_));
 AOI211x1_ASAP7_75t_R _42567_ (.A1(_09589_),
    .A2(_09573_),
    .B(net2959),
    .C(net983),
    .Y(_13639_));
 INVx1_ASAP7_75t_R _42568_ (.A(_13639_),
    .Y(_13640_));
 NAND2x1_ASAP7_75t_R _42569_ (.A(_11748_),
    .B(_13640_),
    .Y(_13641_));
 NOR2x1_ASAP7_75t_R _42570_ (.A(_13638_),
    .B(_13641_),
    .Y(_13642_));
 NAND2x1_ASAP7_75t_R _42571_ (.A(_13637_),
    .B(_13642_),
    .Y(_13643_));
 OA21x2_ASAP7_75t_R _42572_ (.A1(_09761_),
    .A2(_11128_),
    .B(_11090_),
    .Y(_13644_));
 AOI211x1_ASAP7_75t_R _42573_ (.A1(_09589_),
    .A2(net1280),
    .B(net2000),
    .C(_09597_),
    .Y(_13645_));
 NOR3x1_ASAP7_75t_R _42574_ (.A(_13644_),
    .B(_13645_),
    .C(_12032_),
    .Y(_13646_));
 NAND2x1_ASAP7_75t_R _42575_ (.A(_11111_),
    .B(_09806_),
    .Y(_13648_));
 OAI21x1_ASAP7_75t_R _42576_ (.A1(_11675_),
    .A2(_11766_),
    .B(_09806_),
    .Y(_13649_));
 NAND2x2_ASAP7_75t_R _42577_ (.A(_13648_),
    .B(_13649_),
    .Y(_13650_));
 NOR2x2_ASAP7_75t_R _42578_ (.A(net1509),
    .B(_09817_),
    .Y(_13651_));
 AOI211x1_ASAP7_75t_R _42579_ (.A1(_00615_),
    .A2(net1278),
    .B(net1508),
    .C(_09674_),
    .Y(_13652_));
 NOR3x2_ASAP7_75t_R _42580_ (.B(_13651_),
    .C(_13652_),
    .Y(_13653_),
    .A(_13650_));
 NAND2x1_ASAP7_75t_R _42581_ (.A(_13646_),
    .B(_13653_),
    .Y(_13654_));
 NOR2x1_ASAP7_75t_R _42582_ (.A(_13643_),
    .B(_13654_),
    .Y(_13655_));
 NAND2x1_ASAP7_75t_R _42583_ (.A(_13630_),
    .B(_13655_),
    .Y(_13656_));
 NAND2x1_ASAP7_75t_R _42584_ (.A(_12090_),
    .B(_09747_),
    .Y(_13657_));
 NAND2x1_ASAP7_75t_R _42585_ (.A(_09716_),
    .B(_13234_),
    .Y(_13659_));
 NOR2x1_ASAP7_75t_R _42586_ (.A(_13657_),
    .B(_13659_),
    .Y(_13660_));
 NAND2x1_ASAP7_75t_R _42587_ (.A(_13232_),
    .B(_11051_),
    .Y(_13661_));
 AO21x1_ASAP7_75t_R _42588_ (.A1(_09658_),
    .A2(net2558),
    .B(_09692_),
    .Y(_13662_));
 OAI21x1_ASAP7_75t_R _42589_ (.A1(net2940),
    .A2(net2547),
    .B(_13662_),
    .Y(_13663_));
 NOR2x1_ASAP7_75t_R _42590_ (.A(_13661_),
    .B(_13663_),
    .Y(_13664_));
 NAND2x1_ASAP7_75t_R _42591_ (.A(_13660_),
    .B(_13664_),
    .Y(_13665_));
 OA21x2_ASAP7_75t_R _42592_ (.A1(_11736_),
    .A2(_09761_),
    .B(_09838_),
    .Y(_13666_));
 NOR2x2_ASAP7_75t_R _42593_ (.A(_13163_),
    .B(_13666_),
    .Y(_13667_));
 OA21x2_ASAP7_75t_R _42594_ (.A1(_11134_),
    .A2(_11167_),
    .B(net2927),
    .Y(_13668_));
 AOI211x1_ASAP7_75t_R _42595_ (.A1(_09589_),
    .A2(_09573_),
    .B(_09597_),
    .C(net2656),
    .Y(_13670_));
 NOR2x2_ASAP7_75t_R _42596_ (.A(_13668_),
    .B(_13670_),
    .Y(_13671_));
 AOI211x1_ASAP7_75t_R _42597_ (.A1(_09589_),
    .A2(net1278),
    .B(_09597_),
    .C(net2291),
    .Y(_13672_));
 NOR2x2_ASAP7_75t_R _42598_ (.A(_11722_),
    .B(_13672_),
    .Y(_13673_));
 NAND3x2_ASAP7_75t_R _42599_ (.B(_13671_),
    .C(_13673_),
    .Y(_13674_),
    .A(_13667_));
 NOR2x2_ASAP7_75t_R _42600_ (.A(_13665_),
    .B(_13674_),
    .Y(_13675_));
 AO21x1_ASAP7_75t_R _42601_ (.A1(net1289),
    .A2(_09644_),
    .B(_09672_),
    .Y(_13676_));
 AO21x1_ASAP7_75t_R _42602_ (.A1(net3243),
    .A2(net985),
    .B(_09672_),
    .Y(_13677_));
 AND2x2_ASAP7_75t_R _42603_ (.A(_13676_),
    .B(_13677_),
    .Y(_13678_));
 AO21x1_ASAP7_75t_R _42604_ (.A1(_09743_),
    .A2(_09769_),
    .B(net2605),
    .Y(_13679_));
 NAND2x1_ASAP7_75t_R _42605_ (.A(_11182_),
    .B(_09826_),
    .Y(_13681_));
 AND3x1_ASAP7_75t_R _42606_ (.A(_12553_),
    .B(_13679_),
    .C(_13681_),
    .Y(_13682_));
 NAND2x1_ASAP7_75t_R _42607_ (.A(_13678_),
    .B(_13682_),
    .Y(_13683_));
 AO21x1_ASAP7_75t_R _42608_ (.A1(_09611_),
    .A2(_09739_),
    .B(net2914),
    .Y(_13684_));
 AO21x1_ASAP7_75t_R _42609_ (.A1(net1518),
    .A2(net2828),
    .B(net2914),
    .Y(_13685_));
 NAND2x1_ASAP7_75t_R _42610_ (.A(_13684_),
    .B(_13685_),
    .Y(_13686_));
 AO21x1_ASAP7_75t_R _42611_ (.A1(_11161_),
    .A2(net1289),
    .B(net2914),
    .Y(_13687_));
 NAND2x1_ASAP7_75t_R _42612_ (.A(_09697_),
    .B(_13687_),
    .Y(_13688_));
 AO21x1_ASAP7_75t_R _42613_ (.A1(net2940),
    .A2(_09812_),
    .B(net2501),
    .Y(_13689_));
 AO21x1_ASAP7_75t_R _42614_ (.A1(net2503),
    .A2(net3243),
    .B(net2501),
    .Y(_13690_));
 NAND2x1_ASAP7_75t_R _42615_ (.A(_13689_),
    .B(_13690_),
    .Y(_13692_));
 OR3x1_ASAP7_75t_R _42616_ (.A(_13686_),
    .B(_13688_),
    .C(_13692_),
    .Y(_13693_));
 NOR2x1_ASAP7_75t_R _42617_ (.A(_13683_),
    .B(_13693_),
    .Y(_13694_));
 NAND2x1_ASAP7_75t_R _42618_ (.A(_13675_),
    .B(_13694_),
    .Y(_13695_));
 NOR2x2_ASAP7_75t_R _42619_ (.A(_13656_),
    .B(_13695_),
    .Y(_13696_));
 XOR2x2_ASAP7_75t_R _42620_ (.A(_10121_),
    .B(_13696_),
    .Y(_13697_));
 INVx2_ASAP7_75t_R _42621_ (.A(_13697_),
    .Y(_13698_));
 NOR2x2_ASAP7_75t_R _42622_ (.A(_13613_),
    .B(_13698_),
    .Y(_13699_));
 INVx1_ASAP7_75t_R _42623_ (.A(_13612_),
    .Y(_13700_));
 INVx1_ASAP7_75t_R _42624_ (.A(_13551_),
    .Y(_13701_));
 NAND2x1_ASAP7_75t_R _42625_ (.A(_13555_),
    .B(_13566_),
    .Y(_13703_));
 NOR2x2_ASAP7_75t_R _42626_ (.A(_13701_),
    .B(_13703_),
    .Y(_13704_));
 NAND3x2_ASAP7_75t_R _42627_ (.B(_13704_),
    .C(_10991_),
    .Y(_13705_),
    .A(_13700_));
 NOR2x2_ASAP7_75t_R _42628_ (.A(_13697_),
    .B(_13705_),
    .Y(_13706_));
 NAND2x1_ASAP7_75t_R _42629_ (.A(net961),
    .B(net1495),
    .Y(_13707_));
 AO21x1_ASAP7_75t_R _42630_ (.A1(_11323_),
    .A2(_13707_),
    .B(_10567_),
    .Y(_13708_));
 AO21x1_ASAP7_75t_R _42631_ (.A1(net1077),
    .A2(_10410_),
    .B(_10567_),
    .Y(_13709_));
 NAND2x1_ASAP7_75t_R _42632_ (.A(_11341_),
    .B(_10572_),
    .Y(_13710_));
 NAND3x1_ASAP7_75t_R _42633_ (.A(_13708_),
    .B(_13709_),
    .C(_13710_),
    .Y(_13711_));
 AOI21x1_ASAP7_75t_R _42634_ (.A1(net2561),
    .A2(net2695),
    .B(_10578_),
    .Y(_13712_));
 AOI21x1_ASAP7_75t_R _42635_ (.A1(net1051),
    .A2(_10505_),
    .B(_10578_),
    .Y(_13714_));
 NOR3x1_ASAP7_75t_R _42636_ (.A(_13712_),
    .B(_13714_),
    .C(_12996_),
    .Y(_13715_));
 INVx1_ASAP7_75t_R _42637_ (.A(_13715_),
    .Y(_13716_));
 NOR2x1_ASAP7_75t_R _42638_ (.A(_13711_),
    .B(_13716_),
    .Y(_13717_));
 OAI21x1_ASAP7_75t_R _42639_ (.A1(net3338),
    .A2(_11525_),
    .B(_11907_),
    .Y(_13718_));
 INVx1_ASAP7_75t_R _42640_ (.A(_13718_),
    .Y(_13719_));
 NAND2x1_ASAP7_75t_R _42641_ (.A(_10597_),
    .B(_10589_),
    .Y(_13720_));
 INVx1_ASAP7_75t_R _42642_ (.A(_13720_),
    .Y(_13721_));
 AOI211x1_ASAP7_75t_R _42643_ (.A1(_10367_),
    .A2(net3338),
    .B(_10586_),
    .C(net966),
    .Y(_13722_));
 NOR2x1_ASAP7_75t_R _42644_ (.A(_13721_),
    .B(_13722_),
    .Y(_13723_));
 NAND2x1_ASAP7_75t_R _42645_ (.A(_13719_),
    .B(_13723_),
    .Y(_13725_));
 AO21x1_ASAP7_75t_R _42646_ (.A1(_10382_),
    .A2(_10310_),
    .B(_10341_),
    .Y(_13726_));
 AOI21x1_ASAP7_75t_R _42647_ (.A1(_10604_),
    .A2(_13726_),
    .B(net2526),
    .Y(_13727_));
 INVx1_ASAP7_75t_R _42648_ (.A(_13727_),
    .Y(_13728_));
 AOI211x1_ASAP7_75t_R _42649_ (.A1(net975),
    .A2(_00576_),
    .B(net2526),
    .C(net3012),
    .Y(_13729_));
 OA21x2_ASAP7_75t_R _42650_ (.A1(_10385_),
    .A2(_13394_),
    .B(_10601_),
    .Y(_13730_));
 NOR2x1_ASAP7_75t_R _42651_ (.A(_13729_),
    .B(_13730_),
    .Y(_13731_));
 NAND2x1_ASAP7_75t_R _42652_ (.A(_13728_),
    .B(_13731_),
    .Y(_13732_));
 NOR2x1_ASAP7_75t_R _42653_ (.A(_13725_),
    .B(_13732_),
    .Y(_13733_));
 NAND2x1_ASAP7_75t_R _42654_ (.A(_13717_),
    .B(_13733_),
    .Y(_13734_));
 NOR2x1_ASAP7_75t_R _42655_ (.A(_11355_),
    .B(_11323_),
    .Y(_13736_));
 AOI221x1_ASAP7_75t_R _42656_ (.A1(_10367_),
    .A2(net3338),
    .B1(_10341_),
    .B2(net1514),
    .C(_11355_),
    .Y(_13737_));
 NOR2x1_ASAP7_75t_R _42657_ (.A(_13736_),
    .B(_13737_),
    .Y(_13738_));
 AO21x1_ASAP7_75t_R _42658_ (.A1(_10518_),
    .A2(net3157),
    .B(_10515_),
    .Y(_13739_));
 AO21x1_ASAP7_75t_R _42659_ (.A1(net2441),
    .A2(_11364_),
    .B(_10515_),
    .Y(_13740_));
 AND2x2_ASAP7_75t_R _42660_ (.A(_13739_),
    .B(_13740_),
    .Y(_13741_));
 NAND2x1_ASAP7_75t_R _42661_ (.A(_13738_),
    .B(_13741_),
    .Y(_13742_));
 INVx1_ASAP7_75t_R _42662_ (.A(_13742_),
    .Y(_13743_));
 NAND2x2_ASAP7_75t_R _42663_ (.A(_10576_),
    .B(_10547_),
    .Y(_13744_));
 NAND2x2_ASAP7_75t_R _42664_ (.A(_11341_),
    .B(_10547_),
    .Y(_13745_));
 NAND3x2_ASAP7_75t_R _42665_ (.B(_13744_),
    .C(_13745_),
    .Y(_13747_),
    .A(_13379_));
 AO21x1_ASAP7_75t_R _42666_ (.A1(net1143),
    .A2(net1051),
    .B(_10540_),
    .Y(_13748_));
 NAND2x1_ASAP7_75t_R _42667_ (.A(_13748_),
    .B(_11927_),
    .Y(_13749_));
 AO21x1_ASAP7_75t_R _42668_ (.A1(net2561),
    .A2(_10471_),
    .B(_10540_),
    .Y(_13750_));
 AO21x1_ASAP7_75t_R _42669_ (.A1(net3052),
    .A2(net1855),
    .B(_10540_),
    .Y(_13751_));
 NAND2x1_ASAP7_75t_R _42670_ (.A(_13750_),
    .B(_13751_),
    .Y(_13752_));
 NOR2x2_ASAP7_75t_R _42671_ (.A(_13749_),
    .B(_13752_),
    .Y(_13753_));
 INVx1_ASAP7_75t_R _42672_ (.A(_13753_),
    .Y(_13754_));
 NOR2x1_ASAP7_75t_R _42673_ (.A(_13747_),
    .B(_13754_),
    .Y(_13755_));
 NAND2x1_ASAP7_75t_R _42674_ (.A(_13743_),
    .B(_13755_),
    .Y(_13756_));
 NOR2x1_ASAP7_75t_R _42675_ (.A(_13734_),
    .B(_13756_),
    .Y(_13758_));
 OAI21x1_ASAP7_75t_R _42676_ (.A1(_10399_),
    .A2(_10551_),
    .B(_10406_),
    .Y(_13759_));
 NAND3x2_ASAP7_75t_R _42677_ (.B(_10422_),
    .C(_13759_),
    .Y(_13760_),
    .A(_13419_));
 AO21x1_ASAP7_75t_R _42678_ (.A1(_10382_),
    .A2(_10317_),
    .B(net965),
    .Y(_13761_));
 AOI21x1_ASAP7_75t_R _42679_ (.A1(_11383_),
    .A2(_13761_),
    .B(net2448),
    .Y(_13762_));
 INVx1_ASAP7_75t_R _42680_ (.A(_13762_),
    .Y(_13763_));
 NOR2x2_ASAP7_75t_R _42681_ (.A(_11364_),
    .B(net2450),
    .Y(_13764_));
 OA21x2_ASAP7_75t_R _42682_ (.A1(_11967_),
    .A2(_11349_),
    .B(_11481_),
    .Y(_13765_));
 NOR2x1_ASAP7_75t_R _42683_ (.A(_13764_),
    .B(_13765_),
    .Y(_13766_));
 NAND2x1_ASAP7_75t_R _42684_ (.A(_13763_),
    .B(_13766_),
    .Y(_13767_));
 NOR2x1_ASAP7_75t_R _42685_ (.A(_13760_),
    .B(_13767_),
    .Y(_13769_));
 NOR2x1_ASAP7_75t_R _42686_ (.A(_10336_),
    .B(_11954_),
    .Y(_13770_));
 AOI211x1_ASAP7_75t_R _42687_ (.A1(_10367_),
    .A2(_10316_),
    .B(_10336_),
    .C(_10341_),
    .Y(_13771_));
 NOR2x2_ASAP7_75t_R _42688_ (.A(_13770_),
    .B(_13771_),
    .Y(_13772_));
 NOR2x1_ASAP7_75t_R _42689_ (.A(_10358_),
    .B(_11954_),
    .Y(_13773_));
 AOI211x1_ASAP7_75t_R _42690_ (.A1(_10367_),
    .A2(_10316_),
    .B(_10358_),
    .C(net965),
    .Y(_13774_));
 NOR2x2_ASAP7_75t_R _42691_ (.A(_13773_),
    .B(_13774_),
    .Y(_13775_));
 AO31x2_ASAP7_75t_R _42692_ (.A1(_10505_),
    .A2(_10442_),
    .A3(net1511),
    .B(_10358_),
    .Y(_13776_));
 NAND3x2_ASAP7_75t_R _42693_ (.B(_13775_),
    .C(_13776_),
    .Y(_13777_),
    .A(_13772_));
 INVx1_ASAP7_75t_R _42694_ (.A(_13777_),
    .Y(_13778_));
 NAND2x2_ASAP7_75t_R _42695_ (.A(_13769_),
    .B(_13778_),
    .Y(_13780_));
 AO21x1_ASAP7_75t_R _42696_ (.A1(_10471_),
    .A2(net971),
    .B(_10454_),
    .Y(_13781_));
 NAND2x1_ASAP7_75t_R _42697_ (.A(net3019),
    .B(_10462_),
    .Y(_13782_));
 NAND3x1_ASAP7_75t_R _42698_ (.A(_11995_),
    .B(_13781_),
    .C(_13782_),
    .Y(_13783_));
 INVx1_ASAP7_75t_R _42699_ (.A(_12745_),
    .Y(_13784_));
 INVx1_ASAP7_75t_R _42700_ (.A(_11398_),
    .Y(_13785_));
 AO21x1_ASAP7_75t_R _42701_ (.A1(_10471_),
    .A2(_11306_),
    .B(_10468_),
    .Y(_13786_));
 NAND2x1_ASAP7_75t_R _42702_ (.A(_13785_),
    .B(_13786_),
    .Y(_13787_));
 INVx1_ASAP7_75t_R _42703_ (.A(_13787_),
    .Y(_13788_));
 NAND2x1_ASAP7_75t_R _42704_ (.A(_13784_),
    .B(_13788_),
    .Y(_13789_));
 NOR2x1_ASAP7_75t_R _42705_ (.A(_13783_),
    .B(_13789_),
    .Y(_13791_));
 AO21x1_ASAP7_75t_R _42706_ (.A1(_10485_),
    .A2(_10329_),
    .B(net2070),
    .Y(_13792_));
 NAND2x1_ASAP7_75t_R _42707_ (.A(_10484_),
    .B(_13792_),
    .Y(_13793_));
 AO21x1_ASAP7_75t_R _42708_ (.A1(_10449_),
    .A2(net2354),
    .B(net2070),
    .Y(_13794_));
 AO21x1_ASAP7_75t_R _42709_ (.A1(net2561),
    .A2(_10370_),
    .B(net2070),
    .Y(_13795_));
 NAND2x1_ASAP7_75t_R _42710_ (.A(_13794_),
    .B(_13795_),
    .Y(_13796_));
 NOR2x1_ASAP7_75t_R _42711_ (.A(_13793_),
    .B(_13796_),
    .Y(_13797_));
 AO21x1_ASAP7_75t_R _42712_ (.A1(net3052),
    .A2(_10471_),
    .B(net2249),
    .Y(_13798_));
 AO21x1_ASAP7_75t_R _42713_ (.A1(net3037),
    .A2(net1055),
    .B(net2249),
    .Y(_13799_));
 NAND2x1_ASAP7_75t_R _42714_ (.A(_11932_),
    .B(_11413_),
    .Y(_13800_));
 NAND3x1_ASAP7_75t_R _42715_ (.A(_13798_),
    .B(_13799_),
    .C(_13800_),
    .Y(_13802_));
 INVx1_ASAP7_75t_R _42716_ (.A(_13802_),
    .Y(_13803_));
 NAND2x1_ASAP7_75t_R _42717_ (.A(_13797_),
    .B(_13803_),
    .Y(_13804_));
 INVx1_ASAP7_75t_R _42718_ (.A(_13804_),
    .Y(_13805_));
 NAND2x1_ASAP7_75t_R _42719_ (.A(_13791_),
    .B(_13805_),
    .Y(_13806_));
 NOR2x2_ASAP7_75t_R _42720_ (.A(_13780_),
    .B(_13806_),
    .Y(_13807_));
 NAND2x2_ASAP7_75t_R _42721_ (.A(_13758_),
    .B(_13807_),
    .Y(_13808_));
 XOR2x1_ASAP7_75t_R _42722_ (.A(_13372_),
    .Y(_13809_),
    .B(_13808_));
 INVx1_ASAP7_75t_R _42723_ (.A(_13809_),
    .Y(_13810_));
 OAI21x1_ASAP7_75t_R _42724_ (.A1(_13699_),
    .A2(_13706_),
    .B(_13810_),
    .Y(_13811_));
 NOR2x1_ASAP7_75t_R _42725_ (.A(_13697_),
    .B(_13613_),
    .Y(_13813_));
 NOR2x1_ASAP7_75t_R _42726_ (.A(_13698_),
    .B(_13705_),
    .Y(_13814_));
 OAI21x1_ASAP7_75t_R _42727_ (.A1(_13813_),
    .A2(_13814_),
    .B(_13809_),
    .Y(_13815_));
 AO21x2_ASAP7_75t_R _42728_ (.A1(_13811_),
    .A2(_13815_),
    .B(net389),
    .Y(_13816_));
 INVx2_ASAP7_75t_R _42729_ (.A(_00520_),
    .Y(_13817_));
 AOI21x1_ASAP7_75t_R _42730_ (.A1(_13536_),
    .A2(_13816_),
    .B(_13817_),
    .Y(_13818_));
 NAND2x1_ASAP7_75t_R _42731_ (.A(_13816_),
    .B(_13536_),
    .Y(_13819_));
 NOR2x1_ASAP7_75t_R _42732_ (.A(_00520_),
    .B(_13819_),
    .Y(_13820_));
 NOR2x1_ASAP7_75t_R _42733_ (.A(_13818_),
    .B(_13820_),
    .Y(_00104_));
 AND2x2_ASAP7_75t_R _42734_ (.A(net389),
    .B(_00811_),
    .Y(_13821_));
 INVx1_ASAP7_75t_R _42735_ (.A(_13747_),
    .Y(_13823_));
 NAND2x1_ASAP7_75t_R _42736_ (.A(_13753_),
    .B(_13823_),
    .Y(_13824_));
 NOR2x1_ASAP7_75t_R _42737_ (.A(_13742_),
    .B(_13824_),
    .Y(_13825_));
 INVx1_ASAP7_75t_R _42738_ (.A(_13717_),
    .Y(_13826_));
 NOR3x1_ASAP7_75t_R _42739_ (.A(_13727_),
    .B(_13730_),
    .C(_13729_),
    .Y(_13827_));
 INVx1_ASAP7_75t_R _42740_ (.A(_13725_),
    .Y(_13828_));
 NAND2x1_ASAP7_75t_R _42741_ (.A(_13827_),
    .B(_13828_),
    .Y(_13829_));
 NOR2x1_ASAP7_75t_R _42742_ (.A(_13826_),
    .B(_13829_),
    .Y(_13830_));
 NAND2x1_ASAP7_75t_R _42743_ (.A(_13825_),
    .B(_13830_),
    .Y(_13831_));
 NOR2x1_ASAP7_75t_R _42744_ (.A(_12745_),
    .B(_13787_),
    .Y(_13832_));
 INVx1_ASAP7_75t_R _42745_ (.A(_13783_),
    .Y(_13834_));
 NAND2x1_ASAP7_75t_R _42746_ (.A(_13832_),
    .B(_13834_),
    .Y(_13835_));
 NOR2x1_ASAP7_75t_R _42747_ (.A(_13835_),
    .B(_13804_),
    .Y(_13836_));
 INVx1_ASAP7_75t_R _42748_ (.A(_13760_),
    .Y(_13837_));
 NOR3x1_ASAP7_75t_R _42749_ (.A(_13765_),
    .B(_13762_),
    .C(_13764_),
    .Y(_13838_));
 NAND2x1_ASAP7_75t_R _42750_ (.A(_13837_),
    .B(_13838_),
    .Y(_13839_));
 NOR2x2_ASAP7_75t_R _42751_ (.A(_13777_),
    .B(_13839_),
    .Y(_13840_));
 NAND2x2_ASAP7_75t_R _42752_ (.A(_13836_),
    .B(_13840_),
    .Y(_13841_));
 NOR2x2_ASAP7_75t_R _42753_ (.A(_13831_),
    .B(_13841_),
    .Y(_13842_));
 TAPCELL_ASAP7_75t_R PHY_28 ();
 XOR2x2_ASAP7_75t_R _42755_ (.A(_10884_),
    .B(_09867_),
    .Y(_13845_));
 NOR2x1_ASAP7_75t_R _42756_ (.A(net2594),
    .B(_13845_),
    .Y(_13846_));
 NAND2x1_ASAP7_75t_R _42757_ (.A(net2592),
    .B(_13845_),
    .Y(_13847_));
 INVx1_ASAP7_75t_R _42758_ (.A(_13847_),
    .Y(_13848_));
 OAI21x1_ASAP7_75t_R _42759_ (.A1(_13846_),
    .A2(_13848_),
    .B(_11300_),
    .Y(_13849_));
 NAND2x1_ASAP7_75t_R _42760_ (.A(_13808_),
    .B(_13845_),
    .Y(_13850_));
 XOR2x1_ASAP7_75t_R _42761_ (.A(net2932),
    .Y(_13851_),
    .B(_10306_));
 NAND2x1_ASAP7_75t_R _42762_ (.A(net2592),
    .B(_13851_),
    .Y(_13852_));
 AOI21x1_ASAP7_75t_R _42763_ (.A1(_13850_),
    .A2(_13852_),
    .B(_11300_),
    .Y(_13853_));
 INVx1_ASAP7_75t_R _42764_ (.A(_13853_),
    .Y(_13854_));
 TAPCELL_ASAP7_75t_R PHY_27 ();
 AOI21x1_ASAP7_75t_R _42766_ (.A1(_13849_),
    .A2(_13854_),
    .B(net389),
    .Y(_13857_));
 INVx1_ASAP7_75t_R _42767_ (.A(_00412_),
    .Y(_13858_));
 OAI21x1_ASAP7_75t_R _42768_ (.A1(_13821_),
    .A2(_13857_),
    .B(_13858_),
    .Y(_13859_));
 NAND2x1_ASAP7_75t_R _42769_ (.A(_13808_),
    .B(_13851_),
    .Y(_13860_));
 AOI21x1_ASAP7_75t_R _42770_ (.A1(_13860_),
    .A2(_13847_),
    .B(_11050_),
    .Y(_13861_));
 OAI21x1_ASAP7_75t_R _42771_ (.A1(_13861_),
    .A2(_13853_),
    .B(net392),
    .Y(_13862_));
 INVx1_ASAP7_75t_R _42772_ (.A(_13821_),
    .Y(_13863_));
 NAND3x1_ASAP7_75t_R _42773_ (.A(_13862_),
    .B(_00412_),
    .C(_13863_),
    .Y(_13864_));
 NAND2x1_ASAP7_75t_R _42774_ (.A(_13859_),
    .B(_13864_),
    .Y(_00065_));
 NOR2x2_ASAP7_75t_R _42775_ (.A(net393),
    .B(_00810_),
    .Y(_13865_));
 INVx1_ASAP7_75t_R _42776_ (.A(_13865_),
    .Y(_13866_));
 NOR2x1_ASAP7_75t_R _42777_ (.A(_11300_),
    .B(_11297_),
    .Y(_13867_));
 NOR2x1_ASAP7_75t_R _42778_ (.A(_11050_),
    .B(_11303_),
    .Y(_13868_));
 OAI21x1_ASAP7_75t_R _42779_ (.A1(_10364_),
    .A2(_10614_),
    .B(_13842_),
    .Y(_13869_));
 INVx1_ASAP7_75t_R _42780_ (.A(_13869_),
    .Y(_13870_));
 NOR3x1_ASAP7_75t_R _42781_ (.A(_10614_),
    .B(_13842_),
    .C(_10364_),
    .Y(_13871_));
 OAI21x1_ASAP7_75t_R _42782_ (.A1(_13870_),
    .A2(_13871_),
    .B(_11886_),
    .Y(_13872_));
 NAND3x2_ASAP7_75t_R _42783_ (.B(net3055),
    .C(_10611_),
    .Y(_13873_),
    .A(_10562_));
 INVx1_ASAP7_75t_R _42784_ (.A(_10480_),
    .Y(_13874_));
 NOR2x1_ASAP7_75t_R _42785_ (.A(_10509_),
    .B(_13874_),
    .Y(_13876_));
 NAND3x2_ASAP7_75t_R _42786_ (.B(_10402_),
    .C(_10393_),
    .Y(_13877_),
    .A(net3036));
 NAND3x2_ASAP7_75t_R _42787_ (.B(_10438_),
    .C(_10444_),
    .Y(_13878_),
    .A(_10428_));
 NOR2x2_ASAP7_75t_R _42788_ (.A(_13877_),
    .B(_13878_),
    .Y(_13879_));
 NAND2x2_ASAP7_75t_R _42789_ (.A(_13876_),
    .B(_13879_),
    .Y(_13880_));
 NOR2x2_ASAP7_75t_R _42790_ (.A(_13873_),
    .B(_13880_),
    .Y(_13881_));
 NOR2x1_ASAP7_75t_R _42791_ (.A(_13842_),
    .B(_13881_),
    .Y(_13882_));
 NOR3x1_ASAP7_75t_R _42792_ (.A(_10614_),
    .B(_13808_),
    .C(_10364_),
    .Y(_13883_));
 INVx1_ASAP7_75t_R _42793_ (.A(_11886_),
    .Y(_13884_));
 OAI21x1_ASAP7_75t_R _42794_ (.A1(_13882_),
    .A2(_13883_),
    .B(_13884_),
    .Y(_13885_));
 NAND2x2_ASAP7_75t_R _42795_ (.A(_13872_),
    .B(_13885_),
    .Y(_13887_));
 OAI21x1_ASAP7_75t_R _42796_ (.A1(_13867_),
    .A2(_13868_),
    .B(_13887_),
    .Y(_13888_));
 NAND3x2_ASAP7_75t_R _42797_ (.B(_13376_),
    .C(_13808_),
    .Y(_13889_),
    .A(_13881_));
 AOI21x1_ASAP7_75t_R _42798_ (.A1(net3050),
    .A2(_13889_),
    .B(_13884_),
    .Y(_13890_));
 INVx1_ASAP7_75t_R _42799_ (.A(_13882_),
    .Y(_13891_));
 NAND3x1_ASAP7_75t_R _42800_ (.A(_13881_),
    .B(_13376_),
    .C(_13842_),
    .Y(_13892_));
 AOI21x1_ASAP7_75t_R _42801_ (.A1(_13891_),
    .A2(_13892_),
    .B(_11886_),
    .Y(_13893_));
 NOR2x2_ASAP7_75t_R _42802_ (.A(_13890_),
    .B(_13893_),
    .Y(_13894_));
 OAI21x1_ASAP7_75t_R _42803_ (.A1(_11298_),
    .A2(_11304_),
    .B(_13894_),
    .Y(_13895_));
 AOI21x1_ASAP7_75t_R _42804_ (.A1(_13888_),
    .A2(_13895_),
    .B(net389),
    .Y(_13896_));
 INVx1_ASAP7_75t_R _42805_ (.A(_13896_),
    .Y(_13898_));
 AOI21x1_ASAP7_75t_R _42806_ (.A1(_13866_),
    .A2(_13898_),
    .B(_00519_),
    .Y(_13899_));
 INVx1_ASAP7_75t_R _42807_ (.A(_00519_),
    .Y(_13900_));
 NOR3x1_ASAP7_75t_R _42808_ (.A(_13896_),
    .B(_13900_),
    .C(_13865_),
    .Y(_13901_));
 NOR2x1_ASAP7_75t_R _42809_ (.A(_13901_),
    .B(_13899_),
    .Y(_00066_));
 AND2x2_ASAP7_75t_R _42810_ (.A(net389),
    .B(_00809_),
    .Y(_13902_));
 TAPCELL_ASAP7_75t_R PHY_26 ();
 NOR2x2_ASAP7_75t_R _42812_ (.A(net2850),
    .B(_11776_),
    .Y(_13904_));
 AND2x2_ASAP7_75t_R _42813_ (.A(_11776_),
    .B(net2850),
    .Y(_13905_));
 XOR2x2_ASAP7_75t_R _42814_ (.A(_11886_),
    .B(_11427_),
    .Y(_13906_));
 INVx2_ASAP7_75t_R _42815_ (.A(_13906_),
    .Y(_13908_));
 OAI21x1_ASAP7_75t_R _42816_ (.A1(_13904_),
    .A2(_13905_),
    .B(_13908_),
    .Y(_13909_));
 NOR2x2_ASAP7_75t_R _42817_ (.A(net2850),
    .B(_11779_),
    .Y(_13910_));
 AND2x2_ASAP7_75t_R _42818_ (.A(_11779_),
    .B(net2850),
    .Y(_13911_));
 OAI21x1_ASAP7_75t_R _42819_ (.A1(_13910_),
    .A2(_13911_),
    .B(net3334),
    .Y(_13912_));
 AOI21x1_ASAP7_75t_R _42820_ (.A1(_13909_),
    .A2(_13912_),
    .B(net389),
    .Y(_13913_));
 INVx2_ASAP7_75t_R _42821_ (.A(_00518_),
    .Y(_13914_));
 OAI21x1_ASAP7_75t_R _42822_ (.A1(_13902_),
    .A2(_13913_),
    .B(_13914_),
    .Y(_13915_));
 NOR2x1_ASAP7_75t_R _42823_ (.A(net393),
    .B(_00809_),
    .Y(_13916_));
 OAI21x1_ASAP7_75t_R _42824_ (.A1(_13904_),
    .A2(_13905_),
    .B(net3334),
    .Y(_13917_));
 OAI21x1_ASAP7_75t_R _42825_ (.A1(_13910_),
    .A2(_13911_),
    .B(_13908_),
    .Y(_13919_));
 AOI21x1_ASAP7_75t_R _42826_ (.A1(_13917_),
    .A2(_13919_),
    .B(net389),
    .Y(_13920_));
 OAI21x1_ASAP7_75t_R _42827_ (.A1(_13916_),
    .A2(_13920_),
    .B(_00518_),
    .Y(_13921_));
 NAND2x2_ASAP7_75t_R _42828_ (.A(_13915_),
    .B(_13921_),
    .Y(_00067_));
 NOR2x1_ASAP7_75t_R _42829_ (.A(net393),
    .B(_00808_),
    .Y(_13922_));
 XOR2x2_ASAP7_75t_R _42830_ (.A(_11557_),
    .B(_13808_),
    .Y(_13923_));
 XOR2x1_ASAP7_75t_R _42831_ (.A(_13923_),
    .Y(_13924_),
    .B(_12670_));
 XOR2x2_ASAP7_75t_R _42832_ (.A(_12112_),
    .B(_12384_),
    .Y(_13925_));
 XOR2x1_ASAP7_75t_R _42833_ (.A(_13925_),
    .Y(_13926_),
    .B(_12388_));
 NOR2x1_ASAP7_75t_R _42834_ (.A(_13926_),
    .B(_13924_),
    .Y(_13927_));
 NOR3x2_ASAP7_75t_R _42835_ (.B(_12667_),
    .C(_12656_),
    .Y(_13929_),
    .A(_12641_));
 INVx1_ASAP7_75t_R _42836_ (.A(_12618_),
    .Y(_13930_));
 NAND2x2_ASAP7_75t_R _42837_ (.A(_13929_),
    .B(_13930_),
    .Y(_13931_));
 XOR2x1_ASAP7_75t_R _42838_ (.A(_13923_),
    .Y(_13932_),
    .B(_13931_));
 XOR2x1_ASAP7_75t_R _42839_ (.A(_13925_),
    .Y(_13933_),
    .B(_12291_));
 NOR2x1_ASAP7_75t_R _42840_ (.A(_13933_),
    .B(_13932_),
    .Y(_13934_));
 OAI21x1_ASAP7_75t_R _42841_ (.A1(_13927_),
    .A2(_13934_),
    .B(net393),
    .Y(_13935_));
 INVx1_ASAP7_75t_R _42842_ (.A(_13935_),
    .Y(_13936_));
 OAI21x1_ASAP7_75t_R _42843_ (.A1(_13922_),
    .A2(_13936_),
    .B(_00517_),
    .Y(_13937_));
 INVx1_ASAP7_75t_R _42844_ (.A(_00517_),
    .Y(_13938_));
 INVx1_ASAP7_75t_R _42845_ (.A(_13922_),
    .Y(_13940_));
 NAND3x1_ASAP7_75t_R _42846_ (.A(_13935_),
    .B(_13938_),
    .C(_13940_),
    .Y(_13941_));
 NAND2x1_ASAP7_75t_R _42847_ (.A(_13941_),
    .B(_13937_),
    .Y(_00068_));
 NOR2x2_ASAP7_75t_R _42848_ (.A(net393),
    .B(_00807_),
    .Y(_13942_));
 XOR2x2_ASAP7_75t_R _42849_ (.A(_12126_),
    .B(_13808_),
    .Y(_13943_));
 XOR2x1_ASAP7_75t_R _42850_ (.A(_13943_),
    .Y(_13944_),
    .B(_12567_));
 NOR2x1_ASAP7_75t_R _42851_ (.A(_10877_),
    .B(_12670_),
    .Y(_13945_));
 NAND2x1_ASAP7_75t_R _42852_ (.A(_10877_),
    .B(_12670_),
    .Y(_13946_));
 INVx1_ASAP7_75t_R _42853_ (.A(_13946_),
    .Y(_13947_));
 OAI21x1_ASAP7_75t_R _42854_ (.A1(_13945_),
    .A2(_13947_),
    .B(_12944_),
    .Y(_13948_));
 NAND2x1_ASAP7_75t_R _42855_ (.A(_10878_),
    .B(_13931_),
    .Y(_13950_));
 INVx3_ASAP7_75t_R _42856_ (.A(_12944_),
    .Y(_13951_));
 NAND3x1_ASAP7_75t_R _42857_ (.A(_13950_),
    .B(_13946_),
    .C(_13951_),
    .Y(_13952_));
 NAND2x1_ASAP7_75t_R _42858_ (.A(_13948_),
    .B(_13952_),
    .Y(_13953_));
 NAND2x1_ASAP7_75t_R _42859_ (.A(_13944_),
    .B(_13953_),
    .Y(_13954_));
 NOR2x1_ASAP7_75t_R _42860_ (.A(_13953_),
    .B(_13944_),
    .Y(_13955_));
 INVx1_ASAP7_75t_R _42861_ (.A(_13955_),
    .Y(_13956_));
 AOI21x1_ASAP7_75t_R _42862_ (.A1(_13954_),
    .A2(_13956_),
    .B(net389),
    .Y(_13957_));
 OAI21x1_ASAP7_75t_R _42863_ (.A1(_13942_),
    .A2(_13957_),
    .B(_00516_),
    .Y(_13958_));
 XNOR2x1_ASAP7_75t_R _42864_ (.B(_13943_),
    .Y(_13959_),
    .A(_12567_));
 XOR2x1_ASAP7_75t_R _42865_ (.A(_12671_),
    .Y(_13961_),
    .B(_13951_));
 NOR2x1_ASAP7_75t_R _42866_ (.A(_13959_),
    .B(_13961_),
    .Y(_13962_));
 OAI21x1_ASAP7_75t_R _42867_ (.A1(_13955_),
    .A2(_13962_),
    .B(net392),
    .Y(_13963_));
 INVx1_ASAP7_75t_R _42868_ (.A(_13942_),
    .Y(_13964_));
 NAND3x1_ASAP7_75t_R _42869_ (.A(_13963_),
    .B(_17464_),
    .C(_13964_),
    .Y(_13965_));
 NAND2x1_ASAP7_75t_R _42870_ (.A(_13958_),
    .B(_13965_),
    .Y(_00069_));
 AND2x2_ASAP7_75t_R _42871_ (.A(net389),
    .B(_00806_),
    .Y(_13966_));
 INVx1_ASAP7_75t_R _42872_ (.A(_13134_),
    .Y(_13967_));
 NOR2x1_ASAP7_75t_R _42873_ (.A(_13114_),
    .B(_13103_),
    .Y(_13968_));
 NAND2x1_ASAP7_75t_R _42874_ (.A(_13967_),
    .B(_13968_),
    .Y(_13969_));
 INVx1_ASAP7_75t_R _42875_ (.A(_13162_),
    .Y(_13971_));
 NAND2x1_ASAP7_75t_R _42876_ (.A(_13171_),
    .B(_13168_),
    .Y(_13972_));
 NOR2x1_ASAP7_75t_R _42877_ (.A(_13971_),
    .B(_13972_),
    .Y(_13973_));
 INVx1_ASAP7_75t_R _42878_ (.A(_13153_),
    .Y(_13974_));
 NAND2x2_ASAP7_75t_R _42879_ (.A(_13973_),
    .B(_13974_),
    .Y(_13975_));
 NOR2x2_ASAP7_75t_R _42880_ (.A(_13969_),
    .B(_13975_),
    .Y(_13976_));
 NAND2x2_ASAP7_75t_R _42881_ (.A(_09628_),
    .B(_13976_),
    .Y(_13977_));
 NAND2x1_ASAP7_75t_R _42882_ (.A(_13096_),
    .B(_13977_),
    .Y(_13978_));
 INVx1_ASAP7_75t_R _42883_ (.A(_13096_),
    .Y(_13979_));
 NAND2x1_ASAP7_75t_R _42884_ (.A(_13175_),
    .B(_13979_),
    .Y(_13980_));
 INVx2_ASAP7_75t_R _42885_ (.A(_13523_),
    .Y(_13982_));
 AOI21x1_ASAP7_75t_R _42886_ (.A1(_13978_),
    .A2(_13980_),
    .B(_13982_),
    .Y(_13983_));
 NAND2x2_ASAP7_75t_R _42887_ (.A(_13096_),
    .B(_13175_),
    .Y(_13984_));
 NOR2x2_ASAP7_75t_R _42888_ (.A(_13096_),
    .B(_13175_),
    .Y(_13985_));
 INVx2_ASAP7_75t_R _42889_ (.A(_13985_),
    .Y(_13986_));
 AOI21x1_ASAP7_75t_R _42890_ (.A1(_13984_),
    .A2(_13986_),
    .B(_13523_),
    .Y(_13987_));
 XOR2x2_ASAP7_75t_R _42891_ (.A(_12944_),
    .B(_12761_),
    .Y(_13988_));
 OAI21x1_ASAP7_75t_R _42892_ (.A1(_13983_),
    .A2(_13987_),
    .B(_13988_),
    .Y(_13989_));
 AOI21x1_ASAP7_75t_R _42893_ (.A1(_13984_),
    .A2(_13986_),
    .B(_13982_),
    .Y(_13990_));
 NOR2x1_ASAP7_75t_R _42894_ (.A(_13523_),
    .B(_13177_),
    .Y(_13991_));
 INVx1_ASAP7_75t_R _42895_ (.A(_13988_),
    .Y(_13993_));
 OAI21x1_ASAP7_75t_R _42896_ (.A1(_13990_),
    .A2(_13991_),
    .B(_13993_),
    .Y(_13994_));
 AOI21x1_ASAP7_75t_R _42897_ (.A1(_13989_),
    .A2(_13994_),
    .B(net389),
    .Y(_13995_));
 INVx1_ASAP7_75t_R _42898_ (.A(_00515_),
    .Y(_13996_));
 OAI21x1_ASAP7_75t_R _42899_ (.A1(_13966_),
    .A2(_13995_),
    .B(_13996_),
    .Y(_13997_));
 NOR2x1_ASAP7_75t_R _42900_ (.A(net392),
    .B(_00806_),
    .Y(_13998_));
 OAI21x1_ASAP7_75t_R _42901_ (.A1(_13983_),
    .A2(_13987_),
    .B(_13993_),
    .Y(_13999_));
 OAI21x1_ASAP7_75t_R _42902_ (.A1(_13990_),
    .A2(_13991_),
    .B(_13988_),
    .Y(_14000_));
 AOI21x1_ASAP7_75t_R _42903_ (.A1(_13999_),
    .A2(_14000_),
    .B(net389),
    .Y(_14001_));
 OAI21x1_ASAP7_75t_R _42904_ (.A1(_13998_),
    .A2(_14001_),
    .B(_00515_),
    .Y(_14002_));
 NAND2x1_ASAP7_75t_R _42905_ (.A(_14002_),
    .B(_13997_),
    .Y(_00070_));
 OR2x2_ASAP7_75t_R _42906_ (.A(net393),
    .B(_00805_),
    .Y(_14004_));
 AOI21x1_ASAP7_75t_R _42907_ (.A1(_13374_),
    .A2(_13356_),
    .B(_13613_),
    .Y(_14005_));
 AOI21x1_ASAP7_75t_R _42908_ (.A1(_13452_),
    .A2(_13453_),
    .B(_13705_),
    .Y(_14006_));
 XOR2x2_ASAP7_75t_R _42909_ (.A(_13021_),
    .B(_13523_),
    .Y(_14007_));
 INVx2_ASAP7_75t_R _42910_ (.A(_14007_),
    .Y(_14008_));
 OAI21x1_ASAP7_75t_R _42911_ (.A1(_14005_),
    .A2(_14006_),
    .B(_14008_),
    .Y(_14009_));
 INVx1_ASAP7_75t_R _42912_ (.A(_14009_),
    .Y(_14010_));
 NOR2x1_ASAP7_75t_R _42913_ (.A(net1434),
    .B(_13372_),
    .Y(_14011_));
 NOR2x1_ASAP7_75t_R _42914_ (.A(_13358_),
    .B(_13355_),
    .Y(_14012_));
 OAI21x1_ASAP7_75t_R _42915_ (.A1(_14011_),
    .A2(_14012_),
    .B(_13613_),
    .Y(_14014_));
 NOR2x1_ASAP7_75t_R _42916_ (.A(_13358_),
    .B(_13372_),
    .Y(_14015_));
 NOR2x1_ASAP7_75t_R _42917_ (.A(net1435),
    .B(_13355_),
    .Y(_14016_));
 OAI21x1_ASAP7_75t_R _42918_ (.A1(_14015_),
    .A2(_14016_),
    .B(_13705_),
    .Y(_14017_));
 NAND3x2_ASAP7_75t_R _42919_ (.B(_14017_),
    .C(_14007_),
    .Y(_14018_),
    .A(_14014_));
 INVx1_ASAP7_75t_R _42920_ (.A(_14018_),
    .Y(_14019_));
 OAI21x1_ASAP7_75t_R _42921_ (.A1(_14010_),
    .A2(_14019_),
    .B(net393),
    .Y(_14020_));
 AOI21x1_ASAP7_75t_R _42922_ (.A1(_14004_),
    .A2(_14020_),
    .B(_00514_),
    .Y(_14021_));
 NAND2x1_ASAP7_75t_R _42923_ (.A(_00805_),
    .B(net389),
    .Y(_14022_));
 NAND3x1_ASAP7_75t_R _42924_ (.A(_14018_),
    .B(net393),
    .C(_14009_),
    .Y(_14023_));
 AOI21x1_ASAP7_75t_R _42925_ (.A1(_14022_),
    .A2(_14023_),
    .B(_17469_),
    .Y(_14025_));
 NOR2x1_ASAP7_75t_R _42926_ (.A(_14025_),
    .B(_14021_),
    .Y(_00071_));
 AND2x2_ASAP7_75t_R _42927_ (.A(net389),
    .B(_00804_),
    .Y(_14026_));
 XOR2x2_ASAP7_75t_R _42928_ (.A(_13448_),
    .B(net2514),
    .Y(_14027_));
 NOR2x2_ASAP7_75t_R _42929_ (.A(_13699_),
    .B(_13706_),
    .Y(_14028_));
 NAND2x1_ASAP7_75t_R _42930_ (.A(_14027_),
    .B(_14028_),
    .Y(_14029_));
 INVx2_ASAP7_75t_R _42931_ (.A(_14027_),
    .Y(_14030_));
 INVx2_ASAP7_75t_R _42932_ (.A(_14028_),
    .Y(_14031_));
 NAND2x1_ASAP7_75t_R _42933_ (.A(_14030_),
    .B(_14031_),
    .Y(_14032_));
 AOI21x1_ASAP7_75t_R _42934_ (.A1(_14029_),
    .A2(_14032_),
    .B(net389),
    .Y(_14033_));
 OAI21x1_ASAP7_75t_R _42935_ (.A1(_14026_),
    .A2(_14033_),
    .B(_17472_),
    .Y(_14035_));
 NOR2x1_ASAP7_75t_R _42936_ (.A(net392),
    .B(_00804_),
    .Y(_14036_));
 NAND2x1_ASAP7_75t_R _42937_ (.A(_14030_),
    .B(_14028_),
    .Y(_14037_));
 NAND2x1_ASAP7_75t_R _42938_ (.A(_14031_),
    .B(_14027_),
    .Y(_14038_));
 AOI21x1_ASAP7_75t_R _42939_ (.A1(_14037_),
    .A2(_14038_),
    .B(net389),
    .Y(_14039_));
 OAI21x1_ASAP7_75t_R _42940_ (.A1(_14036_),
    .A2(_14039_),
    .B(_00513_),
    .Y(_14040_));
 NAND2x1_ASAP7_75t_R _42941_ (.A(_14040_),
    .B(_14035_),
    .Y(_00072_));
 OR2x2_ASAP7_75t_R _42942_ (.A(net392),
    .B(_00803_),
    .Y(_14041_));
 INVx2_ASAP7_75t_R _42943_ (.A(_11048_),
    .Y(_14042_));
 XOR2x2_ASAP7_75t_R _42944_ (.A(_10884_),
    .B(net2310),
    .Y(_14043_));
 NAND2x2_ASAP7_75t_R _42945_ (.A(_14042_),
    .B(_14043_),
    .Y(_14045_));
 INVx2_ASAP7_75t_R _42946_ (.A(_14043_),
    .Y(_14046_));
 NAND2x2_ASAP7_75t_R _42947_ (.A(_11048_),
    .B(_14046_),
    .Y(_14047_));
 NAND2x2_ASAP7_75t_R _42948_ (.A(net3050),
    .B(_13889_),
    .Y(_14048_));
 INVx1_ASAP7_75t_R _42949_ (.A(_14048_),
    .Y(_14049_));
 AOI21x1_ASAP7_75t_R _42950_ (.A1(_14045_),
    .A2(_14047_),
    .B(_14049_),
    .Y(_14050_));
 NOR2x1_ASAP7_75t_R _42951_ (.A(_11048_),
    .B(_10884_),
    .Y(_14051_));
 AND2x2_ASAP7_75t_R _42952_ (.A(_10884_),
    .B(_11048_),
    .Y(_14052_));
 INVx4_ASAP7_75t_R _42953_ (.A(_13696_),
    .Y(_14053_));
 OAI21x1_ASAP7_75t_R _42954_ (.A1(_14051_),
    .A2(_14052_),
    .B(_14053_),
    .Y(_14054_));
 NOR2x1_ASAP7_75t_R _42955_ (.A(_14051_),
    .B(_14052_),
    .Y(_14056_));
 NAND2x1_ASAP7_75t_R _42956_ (.A(net2310),
    .B(_14056_),
    .Y(_14057_));
 AOI21x1_ASAP7_75t_R _42957_ (.A1(_14054_),
    .A2(_14057_),
    .B(_14048_),
    .Y(_14058_));
 OAI21x1_ASAP7_75t_R _42958_ (.A1(_14050_),
    .A2(_14058_),
    .B(net392),
    .Y(_14059_));
 AOI21x1_ASAP7_75t_R _42959_ (.A1(_14041_),
    .A2(_14059_),
    .B(_00413_),
    .Y(_14060_));
 NAND2x1_ASAP7_75t_R _42960_ (.A(_00803_),
    .B(net389),
    .Y(_14061_));
 AOI21x1_ASAP7_75t_R _42961_ (.A1(_14045_),
    .A2(_14047_),
    .B(_14048_),
    .Y(_14062_));
 AOI21x1_ASAP7_75t_R _42962_ (.A1(_14054_),
    .A2(_14057_),
    .B(_14049_),
    .Y(_14063_));
 OAI21x1_ASAP7_75t_R _42963_ (.A1(_14062_),
    .A2(_14063_),
    .B(net392),
    .Y(_14064_));
 AOI21x1_ASAP7_75t_R _42964_ (.A1(_14061_),
    .A2(_14064_),
    .B(_17475_),
    .Y(_14065_));
 NOR2x2_ASAP7_75t_R _42965_ (.A(_14065_),
    .B(_14060_),
    .Y(_00033_));
 OR2x2_ASAP7_75t_R _42966_ (.A(net392),
    .B(_00802_),
    .Y(_14067_));
 XNOR2x2_ASAP7_75t_R _42967_ (.A(_11426_),
    .B(_11296_),
    .Y(_14068_));
 OR2x2_ASAP7_75t_R _42968_ (.A(_09866_),
    .B(_13696_),
    .Y(_14069_));
 NAND3x2_ASAP7_75t_R _42969_ (.B(_09866_),
    .C(net1493),
    .Y(_14070_),
    .A(_13696_));
 NAND2x2_ASAP7_75t_R _42970_ (.A(_14069_),
    .B(_14070_),
    .Y(_14071_));
 XOR2x1_ASAP7_75t_R _42971_ (.A(_14068_),
    .Y(_14072_),
    .B(_14071_));
 NOR2x1_ASAP7_75t_R _42972_ (.A(_13887_),
    .B(_14072_),
    .Y(_14073_));
 XOR2x2_ASAP7_75t_R _42973_ (.A(_09867_),
    .B(_14053_),
    .Y(_14074_));
 NOR2x1_ASAP7_75t_R _42974_ (.A(_14068_),
    .B(_14074_),
    .Y(_14075_));
 XOR2x2_ASAP7_75t_R _42975_ (.A(_11296_),
    .B(_11426_),
    .Y(_14077_));
 NOR2x1_ASAP7_75t_R _42976_ (.A(_14077_),
    .B(_14071_),
    .Y(_14078_));
 OAI21x1_ASAP7_75t_R _42977_ (.A1(_14075_),
    .A2(_14078_),
    .B(_13887_),
    .Y(_14079_));
 INVx1_ASAP7_75t_R _42978_ (.A(_14079_),
    .Y(_14080_));
 OAI21x1_ASAP7_75t_R _42979_ (.A1(_14073_),
    .A2(_14080_),
    .B(net392),
    .Y(_14081_));
 AOI21x1_ASAP7_75t_R _42980_ (.A1(_14067_),
    .A2(_14081_),
    .B(_00414_),
    .Y(_14082_));
 NAND2x1_ASAP7_75t_R _42981_ (.A(_00802_),
    .B(net389),
    .Y(_14083_));
 XOR2x1_ASAP7_75t_R _42982_ (.A(_14071_),
    .Y(_14084_),
    .B(_14077_));
 NAND2x1_ASAP7_75t_R _42983_ (.A(_13894_),
    .B(_14084_),
    .Y(_14085_));
 NAND3x1_ASAP7_75t_R _42984_ (.A(_14085_),
    .B(net392),
    .C(_14079_),
    .Y(_14086_));
 AOI21x1_ASAP7_75t_R _42985_ (.A1(_14083_),
    .A2(_14086_),
    .B(_17478_),
    .Y(_14088_));
 NOR2x2_ASAP7_75t_R _42986_ (.A(_14082_),
    .B(_14088_),
    .Y(_00034_));
 AND2x2_ASAP7_75t_R _42987_ (.A(net389),
    .B(_00801_),
    .Y(_14089_));
 XNOR2x2_ASAP7_75t_R _42988_ (.A(_11666_),
    .B(_11193_),
    .Y(_14090_));
 NOR2x2_ASAP7_75t_R _42989_ (.A(net2850),
    .B(net3364),
    .Y(_14091_));
 AND2x2_ASAP7_75t_R _42990_ (.A(_14090_),
    .B(net2850),
    .Y(_14092_));
 XOR2x2_ASAP7_75t_R _42991_ (.A(net3336),
    .B(_11557_),
    .Y(_14093_));
 OAI21x1_ASAP7_75t_R _42992_ (.A1(_14091_),
    .A2(_14092_),
    .B(_14093_),
    .Y(_14094_));
 INVx2_ASAP7_75t_R _42993_ (.A(_14093_),
    .Y(_14095_));
 XOR2x1_ASAP7_75t_R _42994_ (.A(_14090_),
    .Y(_14096_),
    .B(net2850));
 NAND2x1_ASAP7_75t_R _42995_ (.A(_14095_),
    .B(_14096_),
    .Y(_14098_));
 AOI21x1_ASAP7_75t_R _42996_ (.A1(_14094_),
    .A2(_14098_),
    .B(net389),
    .Y(_14099_));
 INVx1_ASAP7_75t_R _42997_ (.A(_00512_),
    .Y(_14100_));
 OAI21x1_ASAP7_75t_R _42998_ (.A1(_14089_),
    .A2(_14099_),
    .B(_14100_),
    .Y(_14101_));
 NOR2x1_ASAP7_75t_R _42999_ (.A(net393),
    .B(_00801_),
    .Y(_14102_));
 OAI21x1_ASAP7_75t_R _43000_ (.A1(_14091_),
    .A2(_14092_),
    .B(_14095_),
    .Y(_14103_));
 NAND2x1_ASAP7_75t_R _43001_ (.A(_14096_),
    .B(net3363),
    .Y(_14104_));
 AOI21x1_ASAP7_75t_R _43002_ (.A1(_14103_),
    .A2(_14104_),
    .B(net389),
    .Y(_14105_));
 OAI21x1_ASAP7_75t_R _43003_ (.A1(_14102_),
    .A2(_14105_),
    .B(_00512_),
    .Y(_14106_));
 NAND2x1_ASAP7_75t_R _43004_ (.A(_14106_),
    .B(_14101_),
    .Y(_00035_));
 NOR2x1_ASAP7_75t_R _43005_ (.A(net393),
    .B(_00800_),
    .Y(_14108_));
 XOR2x2_ASAP7_75t_R _43006_ (.A(_11775_),
    .B(_14053_),
    .Y(_14109_));
 XOR2x2_ASAP7_75t_R _43007_ (.A(_12384_),
    .B(_12126_),
    .Y(_14110_));
 XOR2x1_ASAP7_75t_R _43008_ (.A(_14109_),
    .Y(_14111_),
    .B(_14110_));
 NOR2x1_ASAP7_75t_R _43009_ (.A(_14111_),
    .B(_13924_),
    .Y(_14112_));
 XOR2x2_ASAP7_75t_R _43010_ (.A(_11775_),
    .B(_13696_),
    .Y(_14113_));
 XOR2x1_ASAP7_75t_R _43011_ (.A(_14113_),
    .Y(_14114_),
    .B(_14110_));
 NOR2x1_ASAP7_75t_R _43012_ (.A(_14114_),
    .B(_13932_),
    .Y(_14115_));
 OAI21x1_ASAP7_75t_R _43013_ (.A1(_14112_),
    .A2(_14115_),
    .B(net393),
    .Y(_14116_));
 INVx1_ASAP7_75t_R _43014_ (.A(_14116_),
    .Y(_14117_));
 OAI21x1_ASAP7_75t_R _43015_ (.A1(_14108_),
    .A2(_14117_),
    .B(_00511_),
    .Y(_14119_));
 INVx1_ASAP7_75t_R _43016_ (.A(_00511_),
    .Y(_14120_));
 INVx1_ASAP7_75t_R _43017_ (.A(_14108_),
    .Y(_14121_));
 NAND3x1_ASAP7_75t_R _43018_ (.A(_14116_),
    .B(_14120_),
    .C(_14121_),
    .Y(_14122_));
 NAND2x1_ASAP7_75t_R _43019_ (.A(_14122_),
    .B(_14119_),
    .Y(_00036_));
 AND2x2_ASAP7_75t_R _43020_ (.A(net389),
    .B(_00799_),
    .Y(_14123_));
 XOR2x2_ASAP7_75t_R _43021_ (.A(_13943_),
    .B(_13951_),
    .Y(_14124_));
 XNOR2x1_ASAP7_75t_R _43022_ (.B(_12761_),
    .Y(_14125_),
    .A(_12486_));
 XOR2x2_ASAP7_75t_R _43023_ (.A(_12112_),
    .B(_14053_),
    .Y(_14126_));
 XOR2x2_ASAP7_75t_R _43024_ (.A(_14125_),
    .B(_14126_),
    .Y(_14127_));
 NAND2x1_ASAP7_75t_R _43025_ (.A(_14124_),
    .B(_14127_),
    .Y(_14129_));
 INVx2_ASAP7_75t_R _43026_ (.A(_14124_),
    .Y(_14130_));
 INVx2_ASAP7_75t_R _43027_ (.A(_14127_),
    .Y(_14131_));
 NAND2x1_ASAP7_75t_R _43028_ (.A(_14130_),
    .B(_14131_),
    .Y(_14132_));
 AOI21x1_ASAP7_75t_R _43029_ (.A1(_14129_),
    .A2(_14132_),
    .B(net389),
    .Y(_14133_));
 OAI21x1_ASAP7_75t_R _43030_ (.A1(_14123_),
    .A2(_14133_),
    .B(_17484_),
    .Y(_14134_));
 NOR2x1_ASAP7_75t_R _43031_ (.A(net393),
    .B(_00799_),
    .Y(_14135_));
 NAND2x1_ASAP7_75t_R _43032_ (.A(_14130_),
    .B(_14127_),
    .Y(_14136_));
 NAND2x1_ASAP7_75t_R _43033_ (.A(_14124_),
    .B(_14131_),
    .Y(_14137_));
 AOI21x1_ASAP7_75t_R _43034_ (.A1(_14136_),
    .A2(_14137_),
    .B(net389),
    .Y(_14138_));
 OAI21x1_ASAP7_75t_R _43035_ (.A1(_14135_),
    .A2(_14138_),
    .B(_00510_),
    .Y(_14140_));
 NAND2x1_ASAP7_75t_R _43036_ (.A(_14140_),
    .B(_14134_),
    .Y(_00037_));
 AND2x2_ASAP7_75t_R _43037_ (.A(net389),
    .B(_00798_),
    .Y(_14141_));
 AOI21x1_ASAP7_75t_R _43038_ (.A1(net2682),
    .A2(_13095_),
    .B(_12566_),
    .Y(_14142_));
 INVx1_ASAP7_75t_R _43039_ (.A(_14142_),
    .Y(_14143_));
 NAND3x1_ASAP7_75t_R _43040_ (.A(_13095_),
    .B(_12566_),
    .C(net2682),
    .Y(_14144_));
 AOI21x1_ASAP7_75t_R _43041_ (.A1(_14143_),
    .A2(_14144_),
    .B(_13982_),
    .Y(_14145_));
 INVx1_ASAP7_75t_R _43042_ (.A(_14145_),
    .Y(_14146_));
 AO21x1_ASAP7_75t_R _43043_ (.A1(_13095_),
    .A2(net2681),
    .B(_12781_),
    .Y(_14147_));
 NAND3x1_ASAP7_75t_R _43044_ (.A(_12781_),
    .B(_13095_),
    .C(net2681),
    .Y(_14148_));
 AOI21x1_ASAP7_75t_R _43045_ (.A1(_14147_),
    .A2(_14148_),
    .B(_13523_),
    .Y(_14150_));
 INVx1_ASAP7_75t_R _43046_ (.A(_14150_),
    .Y(_14151_));
 OAI21x1_ASAP7_75t_R _43047_ (.A1(_10364_),
    .A2(_13020_),
    .B(_12762_),
    .Y(_14152_));
 NAND2x1_ASAP7_75t_R _43048_ (.A(_13021_),
    .B(_12761_),
    .Y(_14153_));
 NAND2x1_ASAP7_75t_R _43049_ (.A(_14152_),
    .B(_14153_),
    .Y(_14154_));
 INVx1_ASAP7_75t_R _43050_ (.A(_14154_),
    .Y(_14155_));
 AOI21x1_ASAP7_75t_R _43051_ (.A1(_14146_),
    .A2(_14151_),
    .B(_14155_),
    .Y(_14156_));
 INVx1_ASAP7_75t_R _43052_ (.A(_14156_),
    .Y(_14157_));
 NAND3x1_ASAP7_75t_R _43053_ (.A(_14151_),
    .B(_14146_),
    .C(_14155_),
    .Y(_14158_));
 AOI21x1_ASAP7_75t_R _43054_ (.A1(_14157_),
    .A2(_14158_),
    .B(net389),
    .Y(_14159_));
 INVx1_ASAP7_75t_R _43055_ (.A(_00415_),
    .Y(_14161_));
 OAI21x1_ASAP7_75t_R _43056_ (.A1(_14141_),
    .A2(_14159_),
    .B(_14161_),
    .Y(_14162_));
 NOR3x1_ASAP7_75t_R _43057_ (.A(_14150_),
    .B(_14145_),
    .C(net3295),
    .Y(_14163_));
 OAI21x1_ASAP7_75t_R _43058_ (.A1(_14156_),
    .A2(_14163_),
    .B(net393),
    .Y(_14164_));
 INVx1_ASAP7_75t_R _43059_ (.A(_14141_),
    .Y(_14165_));
 NAND3x1_ASAP7_75t_R _43060_ (.A(_14164_),
    .B(_00415_),
    .C(_14165_),
    .Y(_14166_));
 NAND2x1_ASAP7_75t_R _43061_ (.A(_14162_),
    .B(_14166_),
    .Y(_00038_));
 AND2x2_ASAP7_75t_R _43062_ (.A(net389),
    .B(_00797_),
    .Y(_14167_));
 NAND2x2_ASAP7_75t_R _43063_ (.A(_13355_),
    .B(_13175_),
    .Y(_14168_));
 NAND2x1_ASAP7_75t_R _43064_ (.A(_13372_),
    .B(_13977_),
    .Y(_14169_));
 AOI21x1_ASAP7_75t_R _43065_ (.A1(_14168_),
    .A2(_14169_),
    .B(_13705_),
    .Y(_14171_));
 NAND2x1_ASAP7_75t_R _43066_ (.A(_13372_),
    .B(_13175_),
    .Y(_14172_));
 NAND2x2_ASAP7_75t_R _43067_ (.A(_13355_),
    .B(_13977_),
    .Y(_14173_));
 AOI21x1_ASAP7_75t_R _43068_ (.A1(_14172_),
    .A2(_14173_),
    .B(_13613_),
    .Y(_14174_));
 XNOR2x2_ASAP7_75t_R _43069_ (.A(_13021_),
    .B(_13448_),
    .Y(_14175_));
 INVx2_ASAP7_75t_R _43070_ (.A(_14175_),
    .Y(_14176_));
 OAI21x1_ASAP7_75t_R _43071_ (.A1(_14171_),
    .A2(_14174_),
    .B(_14176_),
    .Y(_14177_));
 AOI21x1_ASAP7_75t_R _43072_ (.A1(_14168_),
    .A2(_14169_),
    .B(_13613_),
    .Y(_14178_));
 AOI21x1_ASAP7_75t_R _43073_ (.A1(_14172_),
    .A2(_14173_),
    .B(_13705_),
    .Y(_14179_));
 OAI21x1_ASAP7_75t_R _43074_ (.A1(_14178_),
    .A2(_14179_),
    .B(_14175_),
    .Y(_14180_));
 AOI21x1_ASAP7_75t_R _43075_ (.A1(_14177_),
    .A2(_14180_),
    .B(net389),
    .Y(_14182_));
 OAI21x1_ASAP7_75t_R _43076_ (.A1(_14167_),
    .A2(_14182_),
    .B(_17490_),
    .Y(_14183_));
 NOR2x1_ASAP7_75t_R _43077_ (.A(net393),
    .B(_00797_),
    .Y(_14184_));
 OAI21x1_ASAP7_75t_R _43078_ (.A1(_14178_),
    .A2(_14179_),
    .B(_14176_),
    .Y(_14185_));
 OAI21x1_ASAP7_75t_R _43079_ (.A1(_14171_),
    .A2(_14174_),
    .B(_14175_),
    .Y(_14186_));
 AOI21x1_ASAP7_75t_R _43080_ (.A1(_14185_),
    .A2(_14186_),
    .B(net389),
    .Y(_14187_));
 OAI21x1_ASAP7_75t_R _43081_ (.A1(_14184_),
    .A2(_14187_),
    .B(_00416_),
    .Y(_14188_));
 NAND2x2_ASAP7_75t_R _43082_ (.A(_14183_),
    .B(_14188_),
    .Y(_00039_));
 AND2x2_ASAP7_75t_R _43083_ (.A(net389),
    .B(_00796_),
    .Y(_14189_));
 XOR2x1_ASAP7_75t_R _43084_ (.A(net1437),
    .Y(_14190_),
    .B(net2592));
 XOR2x1_ASAP7_75t_R _43085_ (.A(net2514),
    .Y(_14192_),
    .B(net1883));
 XOR2x1_ASAP7_75t_R _43086_ (.A(_14192_),
    .Y(_14193_),
    .B(_13449_));
 NAND2x1_ASAP7_75t_R _43087_ (.A(_14190_),
    .B(_14193_),
    .Y(_14194_));
 OR2x2_ASAP7_75t_R _43088_ (.A(_14193_),
    .B(_14190_),
    .Y(_14195_));
 AOI21x1_ASAP7_75t_R _43089_ (.A1(_14194_),
    .A2(_14195_),
    .B(net389),
    .Y(_14196_));
 OAI21x1_ASAP7_75t_R _43090_ (.A1(_14189_),
    .A2(_14196_),
    .B(_17493_),
    .Y(_14197_));
 NOR2x1_ASAP7_75t_R _43091_ (.A(net393),
    .B(_00796_),
    .Y(_14198_));
 XOR2x1_ASAP7_75t_R _43092_ (.A(net1437),
    .Y(_14199_),
    .B(_10883_));
 NAND2x1_ASAP7_75t_R _43093_ (.A(net2592),
    .B(_14199_),
    .Y(_14200_));
 XOR2x1_ASAP7_75t_R _43094_ (.A(net1436),
    .Y(_14201_),
    .B(net1883));
 NAND2x1_ASAP7_75t_R _43095_ (.A(_13808_),
    .B(_14201_),
    .Y(_14203_));
 AO21x1_ASAP7_75t_R _43096_ (.A1(_14200_),
    .A2(_14203_),
    .B(_14030_),
    .Y(_14204_));
 NAND3x1_ASAP7_75t_R _43097_ (.A(_14203_),
    .B(_14200_),
    .C(_14030_),
    .Y(_14205_));
 AOI21x1_ASAP7_75t_R _43098_ (.A1(_14204_),
    .A2(_14205_),
    .B(net389),
    .Y(_14206_));
 OAI21x1_ASAP7_75t_R _43099_ (.A1(_14198_),
    .A2(_14206_),
    .B(_00509_),
    .Y(_14207_));
 NAND2x1_ASAP7_75t_R _43100_ (.A(_14207_),
    .B(_14197_),
    .Y(_00040_));
 NOR2x1_ASAP7_75t_R _43101_ (.A(net393),
    .B(_00795_),
    .Y(_14208_));
 NOR2x1_ASAP7_75t_R _43102_ (.A(_14042_),
    .B(_13697_),
    .Y(_14209_));
 INVx1_ASAP7_75t_R _43103_ (.A(_14209_),
    .Y(_14210_));
 NAND2x1_ASAP7_75t_R _43104_ (.A(_14042_),
    .B(_13697_),
    .Y(_14211_));
 XNOR2x1_ASAP7_75t_R _43105_ (.B(_10615_),
    .Y(_14213_),
    .A(net2860));
 NAND3x1_ASAP7_75t_R _43106_ (.A(_14210_),
    .B(_14211_),
    .C(_14213_),
    .Y(_14214_));
 AO21x1_ASAP7_75t_R _43107_ (.A1(_14210_),
    .A2(_14211_),
    .B(_14213_),
    .Y(_14215_));
 AOI21x1_ASAP7_75t_R _43108_ (.A1(_14214_),
    .A2(_14215_),
    .B(net389),
    .Y(_14216_));
 NOR2x1_ASAP7_75t_R _43109_ (.A(_14208_),
    .B(_14216_),
    .Y(_14217_));
 XOR2x1_ASAP7_75t_R _43110_ (.A(_14217_),
    .Y(_00001_),
    .B(_00508_));
 XOR2x2_ASAP7_75t_R _43111_ (.A(_11886_),
    .B(_11193_),
    .Y(_14218_));
 XOR2x1_ASAP7_75t_R _43112_ (.A(_14218_),
    .Y(_14219_),
    .B(_14074_));
 NAND2x1_ASAP7_75t_R _43113_ (.A(_11430_),
    .B(_14219_),
    .Y(_14220_));
 XOR2x1_ASAP7_75t_R _43114_ (.A(_14218_),
    .Y(_14221_),
    .B(_14071_));
 AOI21x1_ASAP7_75t_R _43115_ (.A1(_11432_),
    .A2(_14221_),
    .B(net389),
    .Y(_14223_));
 AND2x2_ASAP7_75t_R _43116_ (.A(net389),
    .B(_00794_),
    .Y(_14224_));
 AOI21x1_ASAP7_75t_R _43117_ (.A1(_14220_),
    .A2(_14223_),
    .B(_14224_),
    .Y(_14225_));
 XNOR2x1_ASAP7_75t_R _43118_ (.B(_14225_),
    .Y(_00002_),
    .A(_00507_));
 AND2x2_ASAP7_75t_R _43119_ (.A(net389),
    .B(_00793_),
    .Y(_14226_));
 NOR2x2_ASAP7_75t_R _43120_ (.A(net2850),
    .B(_11297_),
    .Y(_14227_));
 AND2x2_ASAP7_75t_R _43121_ (.A(_11297_),
    .B(net2850),
    .Y(_14228_));
 XNOR2x2_ASAP7_75t_R _43122_ (.A(_11557_),
    .B(_11775_),
    .Y(_14229_));
 INVx1_ASAP7_75t_R _43123_ (.A(_14229_),
    .Y(_14230_));
 OAI21x1_ASAP7_75t_R _43124_ (.A1(_14227_),
    .A2(_14228_),
    .B(_14230_),
    .Y(_14231_));
 XOR2x1_ASAP7_75t_R _43125_ (.A(_11297_),
    .Y(_14233_),
    .B(net2850));
 NAND2x1_ASAP7_75t_R _43126_ (.A(_14229_),
    .B(_14233_),
    .Y(_14234_));
 AOI21x1_ASAP7_75t_R _43127_ (.A1(_14231_),
    .A2(_14234_),
    .B(net389),
    .Y(_14235_));
 INVx1_ASAP7_75t_R _43128_ (.A(_00506_),
    .Y(_14236_));
 OAI21x1_ASAP7_75t_R _43129_ (.A1(_14226_),
    .A2(_14235_),
    .B(_14236_),
    .Y(_14237_));
 NOR2x1_ASAP7_75t_R _43130_ (.A(net393),
    .B(_00793_),
    .Y(_14238_));
 OAI21x1_ASAP7_75t_R _43131_ (.A1(_14227_),
    .A2(_14228_),
    .B(_14229_),
    .Y(_14239_));
 NAND2x1_ASAP7_75t_R _43132_ (.A(_14233_),
    .B(_14230_),
    .Y(_14240_));
 AOI21x1_ASAP7_75t_R _43133_ (.A1(_14239_),
    .A2(_14240_),
    .B(net389),
    .Y(_14241_));
 OAI21x1_ASAP7_75t_R _43134_ (.A1(_14238_),
    .A2(_14241_),
    .B(_00506_),
    .Y(_14242_));
 NAND2x1_ASAP7_75t_R _43135_ (.A(_14242_),
    .B(_14237_),
    .Y(_00003_));
 NOR2x1_ASAP7_75t_R _43136_ (.A(_14109_),
    .B(_12390_),
    .Y(_14244_));
 NOR2x1_ASAP7_75t_R _43137_ (.A(_14113_),
    .B(_12293_),
    .Y(_14245_));
 NAND2x1_ASAP7_75t_R _43138_ (.A(_12126_),
    .B(_12112_),
    .Y(_14246_));
 NAND2x1_ASAP7_75t_R _43139_ (.A(_12001_),
    .B(_12196_),
    .Y(_14247_));
 AOI21x1_ASAP7_75t_R _43140_ (.A1(_14246_),
    .A2(_14247_),
    .B(_13931_),
    .Y(_14248_));
 AOI21x1_ASAP7_75t_R _43141_ (.A1(_12114_),
    .A2(_12197_),
    .B(_12670_),
    .Y(_14249_));
 NOR2x1_ASAP7_75t_R _43142_ (.A(_14248_),
    .B(_14249_),
    .Y(_14250_));
 OAI21x1_ASAP7_75t_R _43143_ (.A1(_14244_),
    .A2(_14245_),
    .B(_14250_),
    .Y(_14251_));
 NOR2x1_ASAP7_75t_R _43144_ (.A(_14113_),
    .B(_12390_),
    .Y(_14252_));
 NOR2x1_ASAP7_75t_R _43145_ (.A(_14109_),
    .B(_12293_),
    .Y(_14254_));
 NOR2x1_ASAP7_75t_R _43146_ (.A(_12126_),
    .B(_12112_),
    .Y(_14255_));
 NOR2x1_ASAP7_75t_R _43147_ (.A(_12001_),
    .B(_12196_),
    .Y(_14256_));
 OAI21x1_ASAP7_75t_R _43148_ (.A1(_14255_),
    .A2(_14256_),
    .B(_12670_),
    .Y(_14257_));
 NOR2x1_ASAP7_75t_R _43149_ (.A(_12001_),
    .B(_12112_),
    .Y(_14258_));
 NOR2x1_ASAP7_75t_R _43150_ (.A(_12126_),
    .B(_12196_),
    .Y(_14259_));
 OAI21x1_ASAP7_75t_R _43151_ (.A1(_14258_),
    .A2(_14259_),
    .B(_13931_),
    .Y(_14260_));
 NAND2x1_ASAP7_75t_R _43152_ (.A(_14257_),
    .B(_14260_),
    .Y(_14261_));
 OAI21x1_ASAP7_75t_R _43153_ (.A1(_14252_),
    .A2(_14254_),
    .B(_14261_),
    .Y(_14262_));
 AOI21x1_ASAP7_75t_R _43154_ (.A1(_14251_),
    .A2(_14262_),
    .B(net389),
    .Y(_14263_));
 CKINVDCx5p33_ASAP7_75t_R _43155_ (.A(_00505_),
    .Y(_14265_));
 NOR2x1_ASAP7_75t_R _43156_ (.A(net393),
    .B(_00792_),
    .Y(_14266_));
 NOR3x1_ASAP7_75t_R _43157_ (.A(_14263_),
    .B(_14265_),
    .C(_14266_),
    .Y(_14267_));
 OA21x2_ASAP7_75t_R _43158_ (.A1(_14263_),
    .A2(_14266_),
    .B(_14265_),
    .Y(_14268_));
 NOR2x1_ASAP7_75t_R _43159_ (.A(_14268_),
    .B(_14267_),
    .Y(_00004_));
 NOR2x1_ASAP7_75t_R _43160_ (.A(net392),
    .B(_00791_),
    .Y(_14269_));
 XOR2x1_ASAP7_75t_R _43161_ (.A(_14126_),
    .Y(_14270_),
    .B(_12855_));
 XOR2x2_ASAP7_75t_R _43162_ (.A(_12761_),
    .B(_12781_),
    .Y(_14271_));
 XOR2x1_ASAP7_75t_R _43163_ (.A(_14271_),
    .Y(_14272_),
    .B(_12944_));
 NAND2x1_ASAP7_75t_R _43164_ (.A(_14270_),
    .B(_14272_),
    .Y(_14273_));
 INVx1_ASAP7_75t_R _43165_ (.A(_14270_),
    .Y(_14275_));
 INVx1_ASAP7_75t_R _43166_ (.A(_14272_),
    .Y(_14276_));
 NAND2x1_ASAP7_75t_R _43167_ (.A(_14276_),
    .B(_14275_),
    .Y(_14277_));
 AOI21x1_ASAP7_75t_R _43168_ (.A1(_14273_),
    .A2(_14277_),
    .B(net389),
    .Y(_14278_));
 OAI21x1_ASAP7_75t_R _43169_ (.A1(_14269_),
    .A2(_14278_),
    .B(_00504_),
    .Y(_14279_));
 AND2x2_ASAP7_75t_R _43170_ (.A(net389),
    .B(_00791_),
    .Y(_14280_));
 XOR2x1_ASAP7_75t_R _43171_ (.A(_12855_),
    .Y(_14281_),
    .B(_13951_));
 XOR2x1_ASAP7_75t_R _43172_ (.A(_14271_),
    .Y(_14282_),
    .B(_14126_));
 NAND2x1_ASAP7_75t_R _43173_ (.A(_14281_),
    .B(_14282_),
    .Y(_14283_));
 INVx1_ASAP7_75t_R _43174_ (.A(_14281_),
    .Y(_14284_));
 INVx1_ASAP7_75t_R _43175_ (.A(_14282_),
    .Y(_14286_));
 NAND2x1_ASAP7_75t_R _43176_ (.A(_14286_),
    .B(_14284_),
    .Y(_14287_));
 AOI21x1_ASAP7_75t_R _43177_ (.A1(_14283_),
    .A2(_14287_),
    .B(net389),
    .Y(_14288_));
 INVx1_ASAP7_75t_R _43178_ (.A(_00504_),
    .Y(_14289_));
 OAI21x1_ASAP7_75t_R _43179_ (.A1(_14280_),
    .A2(_14288_),
    .B(_14289_),
    .Y(_14290_));
 NAND2x1_ASAP7_75t_R _43180_ (.A(_14290_),
    .B(_14279_),
    .Y(_00005_));
 XOR2x1_ASAP7_75t_R _43181_ (.A(_12567_),
    .Y(_14291_),
    .B(_13175_));
 NAND2x1_ASAP7_75t_R _43182_ (.A(_14008_),
    .B(_14291_),
    .Y(_14292_));
 OA21x2_ASAP7_75t_R _43183_ (.A1(_14291_),
    .A2(_14008_),
    .B(net392),
    .Y(_14293_));
 AND2x2_ASAP7_75t_R _43184_ (.A(net389),
    .B(_00790_),
    .Y(_14294_));
 AOI21x1_ASAP7_75t_R _43185_ (.A1(_14292_),
    .A2(_14293_),
    .B(_14294_),
    .Y(_14296_));
 INVx3_ASAP7_75t_R _43186_ (.A(_00503_),
    .Y(_14297_));
 XOR2x1_ASAP7_75t_R _43187_ (.A(_14296_),
    .Y(_00006_),
    .B(_14297_));
 NOR2x2_ASAP7_75t_R _43188_ (.A(net393),
    .B(_00789_),
    .Y(_14298_));
 AOI21x1_ASAP7_75t_R _43189_ (.A1(_13984_),
    .A2(_13986_),
    .B(_13705_),
    .Y(_14299_));
 AOI22x1_ASAP7_75t_R _43190_ (.A1(_13976_),
    .A2(_09628_),
    .B1(net2683),
    .B2(_13095_),
    .Y(_14300_));
 NOR2x1_ASAP7_75t_R _43191_ (.A(_13096_),
    .B(_13977_),
    .Y(_14301_));
 OAI21x1_ASAP7_75t_R _43192_ (.A1(_14300_),
    .A2(_14301_),
    .B(_13705_),
    .Y(_14302_));
 INVx1_ASAP7_75t_R _43193_ (.A(_14302_),
    .Y(_14303_));
 XOR2x2_ASAP7_75t_R _43194_ (.A(_13448_),
    .B(net1434),
    .Y(_14304_));
 OAI21x1_ASAP7_75t_R _43195_ (.A1(_14299_),
    .A2(_14303_),
    .B(_14304_),
    .Y(_14306_));
 OAI21x1_ASAP7_75t_R _43196_ (.A1(_14300_),
    .A2(_14301_),
    .B(_13613_),
    .Y(_14307_));
 INVx2_ASAP7_75t_R _43197_ (.A(_13984_),
    .Y(_14308_));
 OAI21x1_ASAP7_75t_R _43198_ (.A1(_13985_),
    .A2(_14308_),
    .B(_13705_),
    .Y(_14309_));
 AOI21x1_ASAP7_75t_R _43199_ (.A1(_14307_),
    .A2(_14309_),
    .B(_14304_),
    .Y(_14310_));
 INVx1_ASAP7_75t_R _43200_ (.A(_14310_),
    .Y(_14311_));
 AOI21x1_ASAP7_75t_R _43201_ (.A1(_14306_),
    .A2(_14311_),
    .B(net389),
    .Y(_14312_));
 OAI21x1_ASAP7_75t_R _43202_ (.A1(_14298_),
    .A2(_14312_),
    .B(_00502_),
    .Y(_14313_));
 OAI21x1_ASAP7_75t_R _43203_ (.A1(_13985_),
    .A2(_14308_),
    .B(_13613_),
    .Y(_14314_));
 INVx1_ASAP7_75t_R _43204_ (.A(_14304_),
    .Y(_14315_));
 AOI21x1_ASAP7_75t_R _43205_ (.A1(_14302_),
    .A2(_14314_),
    .B(_14315_),
    .Y(_14317_));
 OAI21x1_ASAP7_75t_R _43206_ (.A1(_14317_),
    .A2(_14310_),
    .B(net392),
    .Y(_14318_));
 INVx2_ASAP7_75t_R _43207_ (.A(_00502_),
    .Y(_14319_));
 INVx1_ASAP7_75t_R _43208_ (.A(_14298_),
    .Y(_14320_));
 NAND3x1_ASAP7_75t_R _43209_ (.A(_14318_),
    .B(_14319_),
    .C(_14320_),
    .Y(_14321_));
 NAND2x1_ASAP7_75t_R _43210_ (.A(_14321_),
    .B(_14313_),
    .Y(_00007_));
 NOR2x2_ASAP7_75t_R _43211_ (.A(net393),
    .B(_00788_),
    .Y(_14322_));
 AO21x1_ASAP7_75t_R _43212_ (.A1(_13356_),
    .A2(_13374_),
    .B(net2310),
    .Y(_14323_));
 AO21x1_ASAP7_75t_R _43213_ (.A1(_13452_),
    .A2(_13453_),
    .B(_14053_),
    .Y(_14324_));
 XOR2x1_ASAP7_75t_R _43214_ (.A(net2514),
    .Y(_14325_),
    .B(net2592));
 INVx1_ASAP7_75t_R _43215_ (.A(_14325_),
    .Y(_14327_));
 AOI21x1_ASAP7_75t_R _43216_ (.A1(_14323_),
    .A2(_14324_),
    .B(_14327_),
    .Y(_14328_));
 AO21x1_ASAP7_75t_R _43217_ (.A1(_13356_),
    .A2(_13374_),
    .B(_14053_),
    .Y(_14329_));
 AO21x1_ASAP7_75t_R _43218_ (.A1(_13452_),
    .A2(_13453_),
    .B(net2310),
    .Y(_14330_));
 AOI21x1_ASAP7_75t_R _43219_ (.A1(_14329_),
    .A2(_14330_),
    .B(_14325_),
    .Y(_14331_));
 OAI21x1_ASAP7_75t_R _43220_ (.A1(_14328_),
    .A2(_14331_),
    .B(net392),
    .Y(_14332_));
 INVx1_ASAP7_75t_R _43221_ (.A(_14332_),
    .Y(_14333_));
 OAI21x1_ASAP7_75t_R _43222_ (.A1(_14322_),
    .A2(_14333_),
    .B(_00501_),
    .Y(_14334_));
 INVx1_ASAP7_75t_R _43223_ (.A(_00501_),
    .Y(_14335_));
 INVx1_ASAP7_75t_R _43224_ (.A(_14322_),
    .Y(_14336_));
 NAND3x1_ASAP7_75t_R _43225_ (.A(_14332_),
    .B(_14335_),
    .C(_14336_),
    .Y(_14338_));
 NAND2x1_ASAP7_75t_R _43226_ (.A(_14338_),
    .B(_14334_),
    .Y(_00008_));
 XNOR2x1_ASAP7_75t_R _43227_ (.B(_10884_),
    .Y(_00153_),
    .A(_00508_));
 XNOR2x1_ASAP7_75t_R _43228_ (.B(_11296_),
    .Y(_00154_),
    .A(_00507_));
 XOR2x1_ASAP7_75t_R _43229_ (.A(_11666_),
    .Y(_00155_),
    .B(_14236_));
 XOR2x1_ASAP7_75t_R _43230_ (.A(_12384_),
    .Y(_00156_),
    .B(_14265_));
 XOR2x1_ASAP7_75t_R _43231_ (.A(_12486_),
    .Y(_00157_),
    .B(_00504_));
 XOR2x1_ASAP7_75t_R _43232_ (.A(_13096_),
    .Y(_00158_),
    .B(_14297_));
 XOR2x1_ASAP7_75t_R _43233_ (.A(_13372_),
    .Y(_00159_),
    .B(_14319_));
 XOR2x1_ASAP7_75t_R _43234_ (.A(_10121_),
    .Y(_00160_),
    .B(_00501_));
 XOR2x1_ASAP7_75t_R _43235_ (.A(net3368),
    .Y(_00249_),
    .B(_00398_));
 XOR2x1_ASAP7_75t_R _43236_ (.A(net3419),
    .Y(_00250_),
    .B(_09479_));
 XOR2x1_ASAP7_75t_R _43237_ (.A(_07049_),
    .Y(_00251_),
    .B(_17275_));
 XOR2x1_ASAP7_75t_R _43238_ (.A(_07697_),
    .Y(_00252_),
    .B(_17284_));
 XOR2x1_ASAP7_75t_R _43239_ (.A(_08169_),
    .Y(_00253_),
    .B(_00486_));
 XOR2x1_ASAP7_75t_R _43240_ (.A(_08504_),
    .Y(_00254_),
    .B(_00405_));
 XOR2x1_ASAP7_75t_R _43241_ (.A(_08849_),
    .Y(_00255_),
    .B(_00407_));
 XOR2x1_ASAP7_75t_R _43242_ (.A(_05427_),
    .Y(_00256_),
    .B(_17312_));
 XOR2x1_ASAP7_75t_R _43243_ (.A(_04612_),
    .Y(_00209_),
    .B(_00460_));
 XOR2x1_ASAP7_75t_R _43244_ (.A(_02091_),
    .Y(_00210_),
    .B(_00459_));
 XOR2x1_ASAP7_75t_R _43245_ (.A(net2523),
    .Y(_00211_),
    .B(_04947_));
 XOR2x1_ASAP7_75t_R _43246_ (.A(net2793),
    .Y(_00212_),
    .B(_04966_));
 XOR2x1_ASAP7_75t_R _43247_ (.A(_03539_),
    .Y(_00213_),
    .B(_00456_));
 XOR2x1_ASAP7_75t_R _43248_ (.A(_03881_),
    .Y(_00214_),
    .B(_05012_));
 XOR2x1_ASAP7_75t_R _43249_ (.A(_04126_),
    .Y(_00215_),
    .B(_00454_));
 XOR2x2_ASAP7_75t_R _43250_ (.A(net2392),
    .B(_05044_),
    .Y(_00216_));
 XOR2x1_ASAP7_75t_R _43251_ (.A(_21388_),
    .Y(_00177_),
    .B(net2129));
 XOR2x1_ASAP7_75t_R _43252_ (.A(_18852_),
    .Y(_00178_),
    .B(net1146));
 XOR2x2_ASAP7_75t_R _43253_ (.A(net3317),
    .B(_05848_),
    .Y(_00179_));
 XOR2x1_ASAP7_75t_R _43254_ (.A(_19961_),
    .Y(_00180_),
    .B(_06189_));
 XOR2x1_ASAP7_75t_R _43255_ (.A(_20352_),
    .Y(_00181_),
    .B(_05749_));
 XOR2x1_ASAP7_75t_R _43256_ (.A(_20544_),
    .Y(_00182_),
    .B(_00423_));
 XOR2x1_ASAP7_75t_R _43257_ (.A(_20899_),
    .Y(_00183_),
    .B(_00422_));
 XOR2x1_ASAP7_75t_R _43258_ (.A(_17905_),
    .Y(_00184_),
    .B(net3386));
 XOR2x1_ASAP7_75t_R _43259_ (.A(_09867_),
    .Y(_00145_),
    .B(_17475_));
 XOR2x1_ASAP7_75t_R _43260_ (.A(_11193_),
    .Y(_00146_),
    .B(_17478_));
 XOR2x1_ASAP7_75t_R _43261_ (.A(_11775_),
    .Y(_00147_),
    .B(_14100_));
 XOR2x1_ASAP7_75t_R _43262_ (.A(_12112_),
    .Y(_00148_),
    .B(_14120_));
 XOR2x1_ASAP7_75t_R _43263_ (.A(_12566_),
    .Y(_00149_),
    .B(_17484_));
 XOR2x1_ASAP7_75t_R _43264_ (.A(_13175_),
    .Y(_00150_),
    .B(_00415_));
 XOR2x2_ASAP7_75t_R _43265_ (.A(_13264_),
    .B(_00416_),
    .Y(_00151_));
 XOR2x1_ASAP7_75t_R _43266_ (.A(net2310),
    .Y(_00152_),
    .B(_00509_));
 XOR2x1_ASAP7_75t_R _43267_ (.A(_05693_),
    .Y(_00241_),
    .B(_09284_));
 XOR2x1_ASAP7_75t_R _43268_ (.A(net1929),
    .Y(_00242_),
    .B(_00491_));
 XOR2x1_ASAP7_75t_R _43269_ (.A(_07159_),
    .Y(_00243_),
    .B(_00393_));
 XOR2x1_ASAP7_75t_R _43270_ (.A(_07806_),
    .Y(_00244_),
    .B(_09358_));
 XOR2x1_ASAP7_75t_R _43271_ (.A(_08005_),
    .Y(_00245_),
    .B(_00395_));
 XOR2x1_ASAP7_75t_R _43272_ (.A(net1861),
    .Y(_00246_),
    .B(_00490_));
 XOR2x1_ASAP7_75t_R _43273_ (.A(net2472),
    .Y(_00247_),
    .B(_16132_));
 XOR2x1_ASAP7_75t_R _43274_ (.A(net1739),
    .Y(_00248_),
    .B(_09453_));
 XOR2x1_ASAP7_75t_R _43275_ (.A(_01094_),
    .Y(_00201_),
    .B(_15661_));
 XOR2x1_ASAP7_75t_R _43276_ (.A(_02357_),
    .Y(_00202_),
    .B(_15784_));
 XOR2x1_ASAP7_75t_R _43277_ (.A(_02786_),
    .Y(_00203_),
    .B(_00466_));
 XOR2x1_ASAP7_75t_R _43278_ (.A(net2700),
    .Y(_00204_),
    .B(_04824_));
 XOR2x1_ASAP7_75t_R _43279_ (.A(net2803),
    .Y(_00205_),
    .B(_00464_));
 XOR2x1_ASAP7_75t_R _43280_ (.A(net2596),
    .Y(_00206_),
    .B(_00463_));
 XOR2x2_ASAP7_75t_R _43281_ (.A(_04201_),
    .B(_00462_),
    .Y(_00207_));
 XOR2x1_ASAP7_75t_R _43282_ (.A(net1886),
    .Y(_00208_),
    .B(_04902_));
 XOR2x1_ASAP7_75t_R _43283_ (.A(_18192_),
    .Y(_00169_),
    .B(_16287_));
 XOR2x1_ASAP7_75t_R _43284_ (.A(net1309),
    .Y(_00170_),
    .B(_16262_));
 XOR2x1_ASAP7_75t_R _43285_ (.A(_19574_),
    .Y(_00171_),
    .B(net3486));
 XOR2x1_ASAP7_75t_R _43286_ (.A(_19962_),
    .Y(_00172_),
    .B(_16276_));
 XOR2x1_ASAP7_75t_R _43287_ (.A(_20448_),
    .Y(_00173_),
    .B(net3502));
 XOR2x1_ASAP7_75t_R _43288_ (.A(_20624_),
    .Y(_00174_),
    .B(_16270_));
 XOR2x1_ASAP7_75t_R _43289_ (.A(_20967_),
    .Y(_00175_),
    .B(_00430_));
 XOR2x1_ASAP7_75t_R _43290_ (.A(_21292_),
    .Y(_00176_),
    .B(_16291_));
 XOR2x1_ASAP7_75t_R _43291_ (.A(_10615_),
    .Y(_00137_),
    .B(_00412_));
 XOR2x1_ASAP7_75t_R _43292_ (.A(net3337),
    .Y(_00138_),
    .B(_00519_));
 XOR2x1_ASAP7_75t_R _43293_ (.A(_11557_),
    .Y(_00139_),
    .B(_13914_));
 XOR2x1_ASAP7_75t_R _43294_ (.A(net2581),
    .Y(_00140_),
    .B(_13938_));
 XOR2x1_ASAP7_75t_R _43295_ (.A(_12761_),
    .Y(_00141_),
    .B(_17464_));
 XOR2x1_ASAP7_75t_R _43296_ (.A(_13021_),
    .Y(_00142_),
    .B(_00515_));
 XOR2x1_ASAP7_75t_R _43297_ (.A(_13448_),
    .Y(_00143_),
    .B(_17469_));
 XOR2x1_ASAP7_75t_R _43298_ (.A(net2593),
    .Y(_00144_),
    .B(_00513_));
 XOR2x1_ASAP7_75t_R _43299_ (.A(_06026_),
    .Y(_00225_),
    .B(_14603_));
 XOR2x1_ASAP7_75t_R _43300_ (.A(_06552_),
    .Y(_00226_),
    .B(_00495_));
 XOR2x1_ASAP7_75t_R _43301_ (.A(_07271_),
    .Y(_00227_),
    .B(_00389_));
 XNOR2x1_ASAP7_75t_R _43302_ (.B(net3418),
    .Y(_00228_),
    .A(_00390_));
 XOR2x1_ASAP7_75t_R _43303_ (.A(_08086_),
    .Y(_00229_),
    .B(_00391_));
 XOR2x1_ASAP7_75t_R _43304_ (.A(_08338_),
    .Y(_00230_),
    .B(_00494_));
 XOR2x1_ASAP7_75t_R _43305_ (.A(net1948),
    .Y(_00231_),
    .B(_17214_));
 XOR2x2_ASAP7_75t_R _43306_ (.A(net1964),
    .B(_17220_),
    .Y(_00232_));
 XOR2x2_ASAP7_75t_R _43307_ (.A(_01754_),
    .B(_14601_),
    .Y(_00193_));
 XOR2x1_ASAP7_75t_R _43308_ (.A(net2573),
    .Y(_00194_),
    .B(_00475_));
 XOR2x1_ASAP7_75t_R _43309_ (.A(net3268),
    .Y(_00195_),
    .B(_04670_));
 XOR2x1_ASAP7_75t_R _43310_ (.A(net3176),
    .Y(_00196_),
    .B(_04697_));
 XOR2x2_ASAP7_75t_R _43311_ (.A(_03466_),
    .B(_00472_),
    .Y(_00197_));
 XOR2x1_ASAP7_75t_R _43312_ (.A(_03960_),
    .Y(_00198_),
    .B(_00471_));
 XOR2x1_ASAP7_75t_R _43313_ (.A(_04282_),
    .Y(_00199_),
    .B(_00470_));
 XNOR2x1_ASAP7_75t_R _43314_ (.B(net3260),
    .Y(_00200_),
    .A(_00469_));
 XOR2x1_ASAP7_75t_R _43315_ (.A(_18507_),
    .Y(_00161_),
    .B(_15432_));
 XOR2x1_ASAP7_75t_R _43316_ (.A(_19252_),
    .Y(_00162_),
    .B(_15425_));
 XOR2x1_ASAP7_75t_R _43317_ (.A(_19560_),
    .Y(_00163_),
    .B(_15427_));
 XOR2x1_ASAP7_75t_R _43318_ (.A(_20049_),
    .Y(_00164_),
    .B(_15433_));
 XOR2x1_ASAP7_75t_R _43319_ (.A(net2537),
    .Y(_00165_),
    .B(_15400_));
 XOR2x1_ASAP7_75t_R _43320_ (.A(_20734_),
    .Y(_00166_),
    .B(_00439_));
 XOR2x1_ASAP7_75t_R _43321_ (.A(_21046_),
    .Y(_00167_),
    .B(_15402_));
 XOR2x1_ASAP7_75t_R _43322_ (.A(_21382_),
    .Y(_00168_),
    .B(_15411_));
 XOR2x2_ASAP7_75t_R _43323_ (.A(_11048_),
    .B(_10897_),
    .Y(_00129_));
 XOR2x1_ASAP7_75t_R _43324_ (.A(_11886_),
    .Y(_00130_),
    .B(_00410_));
 XOR2x1_ASAP7_75t_R _43325_ (.A(net2850),
    .Y(_00131_),
    .B(_00524_));
 XOR2x1_ASAP7_75t_R _43326_ (.A(_12670_),
    .Y(_00132_),
    .B(_00523_));
 XOR2x1_ASAP7_75t_R _43327_ (.A(_12944_),
    .Y(_00133_),
    .B(_00522_));
 XOR2x1_ASAP7_75t_R _43328_ (.A(_13523_),
    .Y(_00134_),
    .B(_00521_));
 XOR2x1_ASAP7_75t_R _43329_ (.A(_13613_),
    .Y(_00135_),
    .B(_00411_));
 XOR2x1_ASAP7_75t_R _43330_ (.A(net2516),
    .Y(_00136_),
    .B(_13817_));
 XOR2x1_ASAP7_75t_R _43331_ (.A(_09271_),
    .Y(_00217_),
    .B(_08779_));
 XOR2x1_ASAP7_75t_R _43332_ (.A(_07381_),
    .Y(_00218_),
    .B(_06930_));
 XOR2x1_ASAP7_75t_R _43333_ (.A(_07499_),
    .Y(_00219_),
    .B(_17139_));
 XOR2x1_ASAP7_75t_R _43334_ (.A(_07917_),
    .Y(_00220_),
    .B(_17145_));
 XOR2x1_ASAP7_75t_R _43335_ (.A(_08266_),
    .Y(_00221_),
    .B(_00387_));
 XOR2x1_ASAP7_75t_R _43336_ (.A(_08601_),
    .Y(_00222_),
    .B(_00498_));
 XOR2x1_ASAP7_75t_R _43337_ (.A(_09022_),
    .Y(_00223_),
    .B(_14360_));
 XOR2x1_ASAP7_75t_R _43338_ (.A(_06729_),
    .Y(_00224_),
    .B(_17171_));
 XOR2x2_ASAP7_75t_R _43339_ (.A(_04753_),
    .B(_08757_),
    .Y(_00185_));
 XOR2x1_ASAP7_75t_R _43340_ (.A(_02588_),
    .Y(_00186_),
    .B(_00483_));
 XOR2x1_ASAP7_75t_R _43341_ (.A(net2675),
    .Y(_00187_),
    .B(_02902_));
 XOR2x1_ASAP7_75t_R _43342_ (.A(_03710_),
    .Y(_00188_),
    .B(_00481_));
 XOR2x1_ASAP7_75t_R _43343_ (.A(_04041_),
    .Y(_00189_),
    .B(_00480_));
 XOR2x1_ASAP7_75t_R _43344_ (.A(net3141),
    .Y(_00190_),
    .B(_04052_));
 XOR2x2_ASAP7_75t_R _43345_ (.A(net3340),
    .B(_14358_),
    .Y(_00191_));
 XNOR2x1_ASAP7_75t_R _43346_ (.B(net2710),
    .Y(_00192_),
    .A(_00477_));
 XOR2x1_ASAP7_75t_R _43347_ (.A(_21582_),
    .Y(_00233_),
    .B(net3514));
 XOR2x2_ASAP7_75t_R _43348_ (.A(_19675_),
    .B(_14620_),
    .Y(_00234_));
 XOR2x1_ASAP7_75t_R _43349_ (.A(_19763_),
    .Y(_00235_),
    .B(net3526));
 XOR2x1_ASAP7_75t_R _43350_ (.A(_20267_),
    .Y(_00236_),
    .B(net3531));
 XOR2x1_ASAP7_75t_R _43351_ (.A(_20818_),
    .Y(_00237_),
    .B(_14682_));
 XOR2x1_ASAP7_75t_R _43352_ (.A(_21123_),
    .Y(_00238_),
    .B(_14643_));
 XOR2x1_ASAP7_75t_R _43353_ (.A(_21212_),
    .Y(_00239_),
    .B(_14758_));
 XOR2x2_ASAP7_75t_R _43354_ (.A(net2885),
    .B(_00445_),
    .Y(_00240_));
 BUFx4_ASAP7_75t_R clkbuf_leaf_0_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_0_clk));
 INVx1_ASAP7_75t_R _43356_ (.A(_00526_),
    .Y(\u0.r0.rcnt[2] ));
 INVx1_ASAP7_75t_R _43357_ (.A(_22101_),
    .Y(\u0.r0.rcnt[1] ));
 INVx2_ASAP7_75t_R _43358_ (.A(\u0.r0.rcnt_next[0] ),
    .Y(\u0.r0.rcnt[0] ));
 INVx1_ASAP7_75t_R _43359_ (.A(_00527_),
    .Y(net259));
 INVx1_ASAP7_75t_R _43360_ (.A(_00657_),
    .Y(net290));
 INVx1_ASAP7_75t_R _43361_ (.A(_00658_),
    .Y(net289));
 INVx1_ASAP7_75t_R _43362_ (.A(_00659_),
    .Y(net288));
 INVx1_ASAP7_75t_R _43363_ (.A(_00660_),
    .Y(net287));
 INVx1_ASAP7_75t_R _43364_ (.A(_00661_),
    .Y(net286));
 INVx1_ASAP7_75t_R _43365_ (.A(_00662_),
    .Y(net285));
 INVx1_ASAP7_75t_R _43366_ (.A(_00663_),
    .Y(net284));
 INVx1_ASAP7_75t_R _43367_ (.A(_00664_),
    .Y(net283));
 INVx1_ASAP7_75t_R _43368_ (.A(_00665_),
    .Y(net382));
 INVx1_ASAP7_75t_R _43369_ (.A(_00666_),
    .Y(net381));
 INVx1_ASAP7_75t_R _43370_ (.A(_00667_),
    .Y(net380));
 INVx1_ASAP7_75t_R _43371_ (.A(_00668_),
    .Y(net379));
 INVx1_ASAP7_75t_R _43372_ (.A(_00669_),
    .Y(net378));
 INVx1_ASAP7_75t_R _43373_ (.A(_00670_),
    .Y(net377));
 INVx1_ASAP7_75t_R _43374_ (.A(_00671_),
    .Y(net375));
 INVx1_ASAP7_75t_R _43375_ (.A(_00672_),
    .Y(net374));
 INVx1_ASAP7_75t_R _43376_ (.A(_00673_),
    .Y(net347));
 INVx1_ASAP7_75t_R _43377_ (.A(_00674_),
    .Y(net346));
 INVx1_ASAP7_75t_R _43378_ (.A(_00675_),
    .Y(net345));
 INVx1_ASAP7_75t_R _43379_ (.A(_00676_),
    .Y(net344));
 INVx1_ASAP7_75t_R _43380_ (.A(_00677_),
    .Y(net342));
 INVx1_ASAP7_75t_R _43381_ (.A(_00678_),
    .Y(net341));
 INVx1_ASAP7_75t_R _43382_ (.A(_00679_),
    .Y(net340));
 INVx1_ASAP7_75t_R _43383_ (.A(_00680_),
    .Y(net339));
 INVx1_ASAP7_75t_R _43384_ (.A(_00681_),
    .Y(net312));
 INVx1_ASAP7_75t_R _43385_ (.A(_00682_),
    .Y(net311));
 INVx1_ASAP7_75t_R _43386_ (.A(_00683_),
    .Y(net309));
 INVx1_ASAP7_75t_R _43387_ (.A(_00684_),
    .Y(net308));
 INVx1_ASAP7_75t_R _43388_ (.A(_00685_),
    .Y(net307));
 INVx1_ASAP7_75t_R _43389_ (.A(_00686_),
    .Y(net306));
 INVx1_ASAP7_75t_R _43390_ (.A(_00687_),
    .Y(net305));
 INVx1_ASAP7_75t_R _43391_ (.A(_00688_),
    .Y(net304));
 INVx1_ASAP7_75t_R _43392_ (.A(_00689_),
    .Y(net281));
 INVx1_ASAP7_75t_R _43393_ (.A(_00690_),
    .Y(net280));
 INVx1_ASAP7_75t_R _43394_ (.A(_00691_),
    .Y(net279));
 INVx1_ASAP7_75t_R _43395_ (.A(_00692_),
    .Y(net278));
 INVx1_ASAP7_75t_R _43396_ (.A(_00693_),
    .Y(net277));
 INVx1_ASAP7_75t_R _43397_ (.A(_00694_),
    .Y(net276));
 INVx1_ASAP7_75t_R _43398_ (.A(_00695_),
    .Y(net275));
 INVx1_ASAP7_75t_R _43399_ (.A(_00696_),
    .Y(net274));
 INVx1_ASAP7_75t_R _43400_ (.A(_00697_),
    .Y(net373));
 INVx1_ASAP7_75t_R _43401_ (.A(_00698_),
    .Y(net372));
 INVx1_ASAP7_75t_R _43402_ (.A(_00699_),
    .Y(net371));
 INVx1_ASAP7_75t_R _43403_ (.A(_00700_),
    .Y(net370));
 INVx1_ASAP7_75t_R _43404_ (.A(_00701_),
    .Y(net369));
 INVx1_ASAP7_75t_R _43405_ (.A(_00702_),
    .Y(net368));
 INVx1_ASAP7_75t_R _43406_ (.A(_00703_),
    .Y(net367));
 INVx1_ASAP7_75t_R _43407_ (.A(_00704_),
    .Y(net366));
 INVx1_ASAP7_75t_R _43408_ (.A(_00705_),
    .Y(net338));
 INVx1_ASAP7_75t_R _43409_ (.A(_00706_),
    .Y(net337));
 INVx1_ASAP7_75t_R _43410_ (.A(_00707_),
    .Y(net336));
 INVx1_ASAP7_75t_R _43411_ (.A(_00708_),
    .Y(net335));
 INVx1_ASAP7_75t_R _43412_ (.A(_00709_),
    .Y(net334));
 INVx1_ASAP7_75t_R _43413_ (.A(_00710_),
    .Y(net333));
 INVx1_ASAP7_75t_R _43414_ (.A(_00711_),
    .Y(net331));
 INVx1_ASAP7_75t_R _43415_ (.A(_00712_),
    .Y(net330));
 INVx1_ASAP7_75t_R _43416_ (.A(_00713_),
    .Y(net303));
 INVx1_ASAP7_75t_R _43417_ (.A(_00714_),
    .Y(net302));
 INVx1_ASAP7_75t_R _43418_ (.A(_00715_),
    .Y(net301));
 INVx1_ASAP7_75t_R _43419_ (.A(_00716_),
    .Y(net300));
 INVx1_ASAP7_75t_R _43420_ (.A(_00717_),
    .Y(net298));
 INVx1_ASAP7_75t_R _43421_ (.A(_00718_),
    .Y(net297));
 INVx1_ASAP7_75t_R _43422_ (.A(_00719_),
    .Y(net296));
 INVx1_ASAP7_75t_R _43423_ (.A(_00720_),
    .Y(net295));
 INVx1_ASAP7_75t_R _43424_ (.A(_00721_),
    .Y(net273));
 INVx1_ASAP7_75t_R _43425_ (.A(_00722_),
    .Y(net272));
 INVx1_ASAP7_75t_R _43426_ (.A(_00723_),
    .Y(net270));
 INVx1_ASAP7_75t_R _43427_ (.A(_00724_),
    .Y(net269));
 INVx1_ASAP7_75t_R _43428_ (.A(_00725_),
    .Y(net268));
 INVx1_ASAP7_75t_R _43429_ (.A(_00726_),
    .Y(net267));
 INVx1_ASAP7_75t_R _43430_ (.A(_00727_),
    .Y(net266));
 INVx1_ASAP7_75t_R _43431_ (.A(_00728_),
    .Y(net265));
 INVx1_ASAP7_75t_R _43432_ (.A(_00729_),
    .Y(net364));
 INVx1_ASAP7_75t_R _43433_ (.A(_00730_),
    .Y(net363));
 INVx1_ASAP7_75t_R _43434_ (.A(_00731_),
    .Y(net362));
 INVx1_ASAP7_75t_R _43435_ (.A(_00732_),
    .Y(net361));
 INVx1_ASAP7_75t_R _43436_ (.A(_00733_),
    .Y(net360));
 INVx1_ASAP7_75t_R _43437_ (.A(_00734_),
    .Y(net359));
 INVx1_ASAP7_75t_R _43438_ (.A(_00735_),
    .Y(net358));
 INVx1_ASAP7_75t_R _43439_ (.A(_00736_),
    .Y(net357));
 INVx1_ASAP7_75t_R _43440_ (.A(_00737_),
    .Y(net329));
 INVx1_ASAP7_75t_R _43441_ (.A(_00738_),
    .Y(net328));
 INVx1_ASAP7_75t_R _43442_ (.A(_00739_),
    .Y(net327));
 INVx1_ASAP7_75t_R _43443_ (.A(_00740_),
    .Y(net326));
 INVx1_ASAP7_75t_R _43444_ (.A(_00741_),
    .Y(net325));
 INVx1_ASAP7_75t_R _43445_ (.A(_00742_),
    .Y(net324));
 INVx1_ASAP7_75t_R _43446_ (.A(_00743_),
    .Y(net323));
 INVx1_ASAP7_75t_R _43447_ (.A(_00744_),
    .Y(net322));
 INVx1_ASAP7_75t_R _43448_ (.A(_00745_),
    .Y(net294));
 INVx1_ASAP7_75t_R _43449_ (.A(_00746_),
    .Y(net293));
 INVx1_ASAP7_75t_R _43450_ (.A(_00747_),
    .Y(net292));
 INVx1_ASAP7_75t_R _43451_ (.A(_00748_),
    .Y(net291));
 INVx1_ASAP7_75t_R _43452_ (.A(_00749_),
    .Y(net282));
 INVx1_ASAP7_75t_R _43453_ (.A(_00750_),
    .Y(net271));
 INVx1_ASAP7_75t_R _43454_ (.A(_00751_),
    .Y(net387));
 INVx1_ASAP7_75t_R _43455_ (.A(_00752_),
    .Y(net376));
 INVx1_ASAP7_75t_R _43456_ (.A(_00753_),
    .Y(net264));
 INVx1_ASAP7_75t_R _43457_ (.A(_00754_),
    .Y(net263));
 INVx1_ASAP7_75t_R _43458_ (.A(_00755_),
    .Y(net262));
 INVx1_ASAP7_75t_R _43459_ (.A(_00756_),
    .Y(net261));
 INVx1_ASAP7_75t_R _43460_ (.A(_00757_),
    .Y(net386));
 INVx1_ASAP7_75t_R _43461_ (.A(_00758_),
    .Y(net385));
 INVx1_ASAP7_75t_R _43462_ (.A(_00759_),
    .Y(net384));
 INVx1_ASAP7_75t_R _43463_ (.A(_00760_),
    .Y(net383));
 INVx1_ASAP7_75t_R _43464_ (.A(_00761_),
    .Y(net356));
 INVx1_ASAP7_75t_R _43465_ (.A(_00762_),
    .Y(net355));
 INVx1_ASAP7_75t_R _43466_ (.A(_00763_),
    .Y(net353));
 INVx1_ASAP7_75t_R _43467_ (.A(_00764_),
    .Y(net352));
 INVx1_ASAP7_75t_R _43468_ (.A(_00765_),
    .Y(net351));
 INVx1_ASAP7_75t_R _43469_ (.A(_00766_),
    .Y(net350));
 INVx1_ASAP7_75t_R _43470_ (.A(_00767_),
    .Y(net349));
 INVx1_ASAP7_75t_R _43471_ (.A(_00768_),
    .Y(net348));
 INVx1_ASAP7_75t_R _43472_ (.A(_00769_),
    .Y(net320));
 INVx1_ASAP7_75t_R _43473_ (.A(_00770_),
    .Y(net319));
 INVx1_ASAP7_75t_R _43474_ (.A(_00771_),
    .Y(net318));
 INVx2_ASAP7_75t_R _43475_ (.A(_00772_),
    .Y(net317));
 INVx1_ASAP7_75t_R _43476_ (.A(_00773_),
    .Y(net316));
 INVx1_ASAP7_75t_R _43477_ (.A(_00774_),
    .Y(net315));
 INVx1_ASAP7_75t_R _43478_ (.A(_00775_),
    .Y(net314));
 INVx1_ASAP7_75t_R _43479_ (.A(_00776_),
    .Y(net313));
 INVx1_ASAP7_75t_R _43480_ (.A(_00777_),
    .Y(net365));
 INVx1_ASAP7_75t_R _43481_ (.A(_00778_),
    .Y(net354));
 INVx1_ASAP7_75t_R _43482_ (.A(_00779_),
    .Y(net343));
 INVx1_ASAP7_75t_R _43483_ (.A(_00780_),
    .Y(net332));
 INVx1_ASAP7_75t_R _43484_ (.A(_00781_),
    .Y(net321));
 INVx1_ASAP7_75t_R _43485_ (.A(_00782_),
    .Y(net310));
 INVx1_ASAP7_75t_R _43486_ (.A(_00783_),
    .Y(net299));
 INVx1_ASAP7_75t_R _43487_ (.A(_00784_),
    .Y(net260));
 TAPCELL_ASAP7_75t_R PHY_25 ();
 NOR2x1_ASAP7_75t_R _43489_ (.A(net404),
    .B(_00915_),
    .Y(_14366_));
 AO21x1_ASAP7_75t_R _43490_ (.A1(net404),
    .A2(net3964),
    .B(_14366_),
    .Y(_00930_));
 NOR2x1_ASAP7_75t_R _43491_ (.A(net404),
    .B(_00914_),
    .Y(_14367_));
 AO21x1_ASAP7_75t_R _43492_ (.A1(net404),
    .A2(net3867),
    .B(_14367_),
    .Y(_00931_));
 NOR2x1_ASAP7_75t_R _43493_ (.A(net404),
    .B(_00913_),
    .Y(_14368_));
 AO21x1_ASAP7_75t_R _43494_ (.A1(net404),
    .A2(net3758),
    .B(_14368_),
    .Y(_00932_));
 NOR2x1_ASAP7_75t_R _43495_ (.A(net404),
    .B(_00912_),
    .Y(_14369_));
 AO21x1_ASAP7_75t_R _43496_ (.A1(net404),
    .A2(net3993),
    .B(_14369_),
    .Y(_00933_));
 NOR2x1_ASAP7_75t_R _43497_ (.A(net404),
    .B(_00911_),
    .Y(_14370_));
 AO21x1_ASAP7_75t_R _43498_ (.A1(net404),
    .A2(net3642),
    .B(_14370_),
    .Y(_00934_));
 NOR2x1_ASAP7_75t_R _43499_ (.A(net403),
    .B(_00910_),
    .Y(_14371_));
 AO21x1_ASAP7_75t_R _43500_ (.A1(net403),
    .A2(net4027),
    .B(_14371_),
    .Y(_00935_));
 NOR2x1_ASAP7_75t_R _43501_ (.A(net404),
    .B(_00909_),
    .Y(_14372_));
 AO21x1_ASAP7_75t_R _43502_ (.A1(net404),
    .A2(net3571),
    .B(_14372_),
    .Y(_00936_));
 TAPCELL_ASAP7_75t_R PHY_24 ();
 NOR2x1_ASAP7_75t_R _43504_ (.A(net404),
    .B(_00908_),
    .Y(_14374_));
 AO21x1_ASAP7_75t_R _43505_ (.A1(net404),
    .A2(net3621),
    .B(_14374_),
    .Y(_00937_));
 NOR2x1_ASAP7_75t_R _43506_ (.A(net129),
    .B(_00907_),
    .Y(_14376_));
 AO21x1_ASAP7_75t_R _43507_ (.A1(net3839),
    .A2(net3565),
    .B(_14376_),
    .Y(_00938_));
 NOR2x1_ASAP7_75t_R _43508_ (.A(net404),
    .B(_00906_),
    .Y(_14377_));
 AO21x1_ASAP7_75t_R _43509_ (.A1(net404),
    .A2(net3574),
    .B(_14377_),
    .Y(_00939_));
 TAPCELL_ASAP7_75t_R PHY_23 ();
 TAPCELL_ASAP7_75t_R PHY_22 ();
 NOR2x1_ASAP7_75t_R _43512_ (.A(net404),
    .B(_00905_),
    .Y(_14380_));
 AO21x1_ASAP7_75t_R _43513_ (.A1(net404),
    .A2(net3586),
    .B(_14380_),
    .Y(_00940_));
 NOR2x1_ASAP7_75t_R _43514_ (.A(net129),
    .B(_00904_),
    .Y(_14381_));
 AO21x1_ASAP7_75t_R _43515_ (.A1(net129),
    .A2(net3764),
    .B(_14381_),
    .Y(_00941_));
 NOR2x1_ASAP7_75t_R _43516_ (.A(net129),
    .B(_00903_),
    .Y(_14383_));
 AO21x1_ASAP7_75t_R _43517_ (.A1(net129),
    .A2(net3701),
    .B(_14383_),
    .Y(_00942_));
 NOR2x1_ASAP7_75t_R _43518_ (.A(net129),
    .B(_00902_),
    .Y(_14384_));
 AO21x1_ASAP7_75t_R _43519_ (.A1(net129),
    .A2(net3755),
    .B(_14384_),
    .Y(_00943_));
 NOR2x1_ASAP7_75t_R _43520_ (.A(net129),
    .B(_00901_),
    .Y(_14385_));
 AO21x1_ASAP7_75t_R _43521_ (.A1(net129),
    .A2(net3737),
    .B(_14385_),
    .Y(_00944_));
 NOR2x1_ASAP7_75t_R _43522_ (.A(net405),
    .B(_00900_),
    .Y(_14386_));
 AO21x1_ASAP7_75t_R _43523_ (.A1(net405),
    .A2(net3725),
    .B(_14386_),
    .Y(_00945_));
 NOR2x1_ASAP7_75t_R _43524_ (.A(net404),
    .B(_00899_),
    .Y(_14387_));
 AO21x1_ASAP7_75t_R _43525_ (.A1(net405),
    .A2(net3713),
    .B(_14387_),
    .Y(_00946_));
 TAPCELL_ASAP7_75t_R PHY_21 ();
 NOR2x1_ASAP7_75t_R _43527_ (.A(net404),
    .B(_00898_),
    .Y(_14390_));
 AO21x1_ASAP7_75t_R _43528_ (.A1(net404),
    .A2(net3665),
    .B(_14390_),
    .Y(_00947_));
 NOR2x1_ASAP7_75t_R _43529_ (.A(net405),
    .B(_00897_),
    .Y(_14391_));
 AO21x1_ASAP7_75t_R _43530_ (.A1(net405),
    .A2(net3731),
    .B(_14391_),
    .Y(_00948_));
 NOR2x1_ASAP7_75t_R _43531_ (.A(net405),
    .B(_00896_),
    .Y(_14392_));
 AO21x1_ASAP7_75t_R _43532_ (.A1(net405),
    .A2(net3752),
    .B(_14392_),
    .Y(_00949_));
 TAPCELL_ASAP7_75t_R PHY_20 ();
 NOR2x1_ASAP7_75t_R _43534_ (.A(net404),
    .B(_00895_),
    .Y(_14394_));
 AO21x1_ASAP7_75t_R _43535_ (.A1(net404),
    .A2(net3722),
    .B(_14394_),
    .Y(_00950_));
 NOR2x1_ASAP7_75t_R _43536_ (.A(net404),
    .B(_00894_),
    .Y(_14396_));
 AO21x1_ASAP7_75t_R _43537_ (.A1(net404),
    .A2(net3710),
    .B(_14396_),
    .Y(_00951_));
 NOR2x1_ASAP7_75t_R _43538_ (.A(net404),
    .B(_00893_),
    .Y(_14397_));
 AO21x1_ASAP7_75t_R _43539_ (.A1(net404),
    .A2(net3577),
    .B(_14397_),
    .Y(_00952_));
 NOR2x1_ASAP7_75t_R _43540_ (.A(net404),
    .B(_00892_),
    .Y(_14398_));
 AO21x1_ASAP7_75t_R _43541_ (.A1(net404),
    .A2(net3686),
    .B(_14398_),
    .Y(_00953_));
 NOR2x1_ASAP7_75t_R _43542_ (.A(net404),
    .B(_00891_),
    .Y(_14399_));
 AO21x1_ASAP7_75t_R _43543_ (.A1(net404),
    .A2(net3870),
    .B(_14399_),
    .Y(_00954_));
 NOR2x1_ASAP7_75t_R _43544_ (.A(net404),
    .B(_00890_),
    .Y(_14400_));
 AO21x1_ASAP7_75t_R _43545_ (.A1(net404),
    .A2(net3952),
    .B(_14400_),
    .Y(_00955_));
 NOR2x1_ASAP7_75t_R _43546_ (.A(net404),
    .B(_00889_),
    .Y(_14402_));
 AO21x1_ASAP7_75t_R _43547_ (.A1(net404),
    .A2(net3767),
    .B(_14402_),
    .Y(_00956_));
 TAPCELL_ASAP7_75t_R PHY_19 ();
 NOR2x1_ASAP7_75t_R _43549_ (.A(net404),
    .B(_00888_),
    .Y(_14404_));
 AO21x1_ASAP7_75t_R _43550_ (.A1(net404),
    .A2(net3928),
    .B(_14404_),
    .Y(_00957_));
 NOR2x1_ASAP7_75t_R _43551_ (.A(net404),
    .B(_00887_),
    .Y(_14405_));
 AO21x1_ASAP7_75t_R _43552_ (.A1(net404),
    .A2(net3800),
    .B(_14405_),
    .Y(_00958_));
 NOR2x1_ASAP7_75t_R _43553_ (.A(net404),
    .B(_00886_),
    .Y(_14406_));
 AO21x1_ASAP7_75t_R _43554_ (.A1(net404),
    .A2(net3934),
    .B(_14406_),
    .Y(_00959_));
 TAPCELL_ASAP7_75t_R PHY_18 ();
 NOR2x1_ASAP7_75t_R _43556_ (.A(net404),
    .B(_00885_),
    .Y(_14409_));
 AO21x1_ASAP7_75t_R _43557_ (.A1(net404),
    .A2(net3779),
    .B(_14409_),
    .Y(_00960_));
 NOR2x1_ASAP7_75t_R _43558_ (.A(net404),
    .B(_00884_),
    .Y(_14410_));
 AO21x1_ASAP7_75t_R _43559_ (.A1(net404),
    .A2(net3773),
    .B(_14410_),
    .Y(_00961_));
 NOR2x1_ASAP7_75t_R _43560_ (.A(net401),
    .B(_00883_),
    .Y(_14411_));
 AO21x1_ASAP7_75t_R _43561_ (.A1(net401),
    .A2(net3749),
    .B(_14411_),
    .Y(_00962_));
 NOR2x1_ASAP7_75t_R _43562_ (.A(net401),
    .B(_00882_),
    .Y(_14412_));
 AO21x1_ASAP7_75t_R _43563_ (.A1(net401),
    .A2(net3716),
    .B(_14412_),
    .Y(_00963_));
 NOR2x1_ASAP7_75t_R _43564_ (.A(net401),
    .B(_00881_),
    .Y(_14413_));
 AO21x1_ASAP7_75t_R _43565_ (.A1(net401),
    .A2(net3734),
    .B(_14413_),
    .Y(_00964_));
 NOR2x1_ASAP7_75t_R _43566_ (.A(net401),
    .B(_00880_),
    .Y(_14415_));
 AO21x1_ASAP7_75t_R _43567_ (.A1(net401),
    .A2(net3639),
    .B(_14415_),
    .Y(_00965_));
 NOR2x1_ASAP7_75t_R _43568_ (.A(net404),
    .B(_00879_),
    .Y(_14416_));
 AO21x1_ASAP7_75t_R _43569_ (.A1(net404),
    .A2(net3976),
    .B(_14416_),
    .Y(_00966_));
 TAPCELL_ASAP7_75t_R PHY_17 ();
 NOR2x1_ASAP7_75t_R _43571_ (.A(net404),
    .B(_00878_),
    .Y(_14418_));
 AO21x1_ASAP7_75t_R _43572_ (.A1(net404),
    .A2(net4029),
    .B(_14418_),
    .Y(_00967_));
 NOR2x1_ASAP7_75t_R _43573_ (.A(net401),
    .B(_00877_),
    .Y(_14419_));
 AO21x1_ASAP7_75t_R _43574_ (.A1(net401),
    .A2(net3740),
    .B(_14419_),
    .Y(_00968_));
 NOR2x1_ASAP7_75t_R _43575_ (.A(net401),
    .B(_00876_),
    .Y(_14421_));
 AO21x1_ASAP7_75t_R _43576_ (.A1(net401),
    .A2(net3719),
    .B(_14421_),
    .Y(_00969_));
 TAPCELL_ASAP7_75t_R PHY_16 ();
 NOR2x1_ASAP7_75t_R _43578_ (.A(net401),
    .B(_00875_),
    .Y(_14423_));
 AO21x1_ASAP7_75t_R _43579_ (.A1(net401),
    .A2(net3692),
    .B(_14423_),
    .Y(_00970_));
 NOR2x1_ASAP7_75t_R _43580_ (.A(net401),
    .B(_00874_),
    .Y(_14424_));
 AO21x1_ASAP7_75t_R _43581_ (.A1(net401),
    .A2(net3680),
    .B(_14424_),
    .Y(_00971_));
 NOR2x1_ASAP7_75t_R _43582_ (.A(net401),
    .B(_00873_),
    .Y(_14425_));
 AO21x1_ASAP7_75t_R _43583_ (.A1(net401),
    .A2(net3698),
    .B(_14425_),
    .Y(_00972_));
 NOR2x1_ASAP7_75t_R _43584_ (.A(net401),
    .B(_00872_),
    .Y(_14426_));
 AO21x1_ASAP7_75t_R _43585_ (.A1(net401),
    .A2(net3645),
    .B(_14426_),
    .Y(_00973_));
 NOR2x1_ASAP7_75t_R _43586_ (.A(net401),
    .B(_00871_),
    .Y(_14428_));
 AO21x1_ASAP7_75t_R _43587_ (.A1(net401),
    .A2(net3636),
    .B(_14428_),
    .Y(_00974_));
 NOR2x1_ASAP7_75t_R _43588_ (.A(net401),
    .B(_00870_),
    .Y(_14429_));
 AO21x1_ASAP7_75t_R _43589_ (.A1(net401),
    .A2(net3624),
    .B(_14429_),
    .Y(_00975_));
 NOR2x1_ASAP7_75t_R _43590_ (.A(net403),
    .B(_00869_),
    .Y(_14430_));
 AO21x1_ASAP7_75t_R _43591_ (.A1(net403),
    .A2(net3902),
    .B(_14430_),
    .Y(_00976_));
 TAPCELL_ASAP7_75t_R PHY_15 ();
 NOR2x1_ASAP7_75t_R _43593_ (.A(net404),
    .B(_00868_),
    .Y(_14432_));
 AO21x1_ASAP7_75t_R _43594_ (.A1(net404),
    .A2(net4002),
    .B(_14432_),
    .Y(_00977_));
 NOR2x1_ASAP7_75t_R _43595_ (.A(net401),
    .B(_00867_),
    .Y(_14434_));
 AO21x1_ASAP7_75t_R _43596_ (.A1(net401),
    .A2(net3683),
    .B(_14434_),
    .Y(_00978_));
 NOR2x1_ASAP7_75t_R _43597_ (.A(net401),
    .B(_00866_),
    .Y(_14435_));
 AO21x1_ASAP7_75t_R _43598_ (.A1(net401),
    .A2(net3668),
    .B(_14435_),
    .Y(_00979_));
 TAPCELL_ASAP7_75t_R PHY_14 ();
 NOR2x1_ASAP7_75t_R _43600_ (.A(net401),
    .B(_00865_),
    .Y(_14437_));
 AO21x1_ASAP7_75t_R _43601_ (.A1(net401),
    .A2(net3609),
    .B(_14437_),
    .Y(_00980_));
 NOR2x1_ASAP7_75t_R _43602_ (.A(net402),
    .B(_00864_),
    .Y(_14438_));
 AO21x1_ASAP7_75t_R _43603_ (.A1(net402),
    .A2(net3695),
    .B(_14438_),
    .Y(_00981_));
 NOR2x1_ASAP7_75t_R _43604_ (.A(net401),
    .B(_00863_),
    .Y(_14439_));
 AO21x1_ASAP7_75t_R _43605_ (.A1(net401),
    .A2(net3943),
    .B(_14439_),
    .Y(_00982_));
 NOR2x1_ASAP7_75t_R _43606_ (.A(net402),
    .B(_00862_),
    .Y(_14441_));
 AO21x1_ASAP7_75t_R _43607_ (.A1(net402),
    .A2(net3594),
    .B(_14441_),
    .Y(_00983_));
 NOR2x1_ASAP7_75t_R _43608_ (.A(net401),
    .B(_00861_),
    .Y(_14442_));
 AO21x1_ASAP7_75t_R _43609_ (.A1(net401),
    .A2(net3633),
    .B(_14442_),
    .Y(_00984_));
 NOR2x1_ASAP7_75t_R _43610_ (.A(net402),
    .B(_00860_),
    .Y(_14443_));
 AO21x1_ASAP7_75t_R _43611_ (.A1(net402),
    .A2(net3580),
    .B(_14443_),
    .Y(_00985_));
 NOR2x1_ASAP7_75t_R _43612_ (.A(net401),
    .B(_00859_),
    .Y(_14444_));
 AO21x1_ASAP7_75t_R _43613_ (.A1(net401),
    .A2(net3746),
    .B(_14444_),
    .Y(_00986_));
 TAPCELL_ASAP7_75t_R PHY_13 ();
 NOR2x1_ASAP7_75t_R _43615_ (.A(net401),
    .B(_00858_),
    .Y(_14447_));
 AO21x1_ASAP7_75t_R _43616_ (.A1(net401),
    .A2(net3707),
    .B(_14447_),
    .Y(_00987_));
 NOR2x1_ASAP7_75t_R _43617_ (.A(net401),
    .B(_00857_),
    .Y(_14448_));
 AO21x1_ASAP7_75t_R _43618_ (.A1(net401),
    .A2(net3648),
    .B(_14448_),
    .Y(_00988_));
 NOR2x1_ASAP7_75t_R _43619_ (.A(net401),
    .B(_00856_),
    .Y(_14449_));
 AO21x1_ASAP7_75t_R _43620_ (.A1(net401),
    .A2(net3704),
    .B(_14449_),
    .Y(_00989_));
 TAPCELL_ASAP7_75t_R PHY_12 ();
 NOR2x1_ASAP7_75t_R _43622_ (.A(net401),
    .B(_00855_),
    .Y(_14451_));
 AO21x1_ASAP7_75t_R _43623_ (.A1(net401),
    .A2(net3618),
    .B(_14451_),
    .Y(_00990_));
 NOR2x1_ASAP7_75t_R _43624_ (.A(net401),
    .B(_00854_),
    .Y(_14452_));
 AO21x1_ASAP7_75t_R _43625_ (.A1(net401),
    .A2(net3955),
    .B(_14452_),
    .Y(_00991_));
 NOR2x1_ASAP7_75t_R _43626_ (.A(net401),
    .B(_00853_),
    .Y(_14454_));
 AO21x1_ASAP7_75t_R _43627_ (.A1(net401),
    .A2(net3689),
    .B(_14454_),
    .Y(_00992_));
 NOR2x1_ASAP7_75t_R _43628_ (.A(net401),
    .B(_00852_),
    .Y(_14455_));
 AO21x1_ASAP7_75t_R _43629_ (.A1(net401),
    .A2(net3656),
    .B(_14455_),
    .Y(_00993_));
 NOR2x1_ASAP7_75t_R _43630_ (.A(net402),
    .B(_00851_),
    .Y(_14456_));
 AO21x1_ASAP7_75t_R _43631_ (.A1(net402),
    .A2(net3583),
    .B(_14456_),
    .Y(_00994_));
 NOR2x1_ASAP7_75t_R _43632_ (.A(net402),
    .B(_00850_),
    .Y(_14457_));
 AO21x1_ASAP7_75t_R _43633_ (.A1(net402),
    .A2(net3615),
    .B(_14457_),
    .Y(_00995_));
 NOR2x1_ASAP7_75t_R _43634_ (.A(net402),
    .B(_00849_),
    .Y(_14458_));
 AO21x1_ASAP7_75t_R _43635_ (.A1(net402),
    .A2(net3671),
    .B(_14458_),
    .Y(_00996_));
 TAPCELL_ASAP7_75t_R PHY_11 ();
 NOR2x1_ASAP7_75t_R _43637_ (.A(net402),
    .B(_00848_),
    .Y(_14461_));
 AO21x1_ASAP7_75t_R _43638_ (.A1(net402),
    .A2(net3849),
    .B(_14461_),
    .Y(_00997_));
 NOR2x1_ASAP7_75t_R _43639_ (.A(net402),
    .B(_00847_),
    .Y(_14462_));
 AO21x1_ASAP7_75t_R _43640_ (.A1(net402),
    .A2(net3836),
    .B(_14462_),
    .Y(_00998_));
 NOR2x1_ASAP7_75t_R _43641_ (.A(net402),
    .B(_00846_),
    .Y(_14463_));
 AO21x1_ASAP7_75t_R _43642_ (.A1(net402),
    .A2(net3788),
    .B(_14463_),
    .Y(_00999_));
 TAPCELL_ASAP7_75t_R PHY_10 ();
 NOR2x1_ASAP7_75t_R _43644_ (.A(net402),
    .B(_00845_),
    .Y(_14465_));
 AO21x1_ASAP7_75t_R _43645_ (.A1(net402),
    .A2(net3806),
    .B(_14465_),
    .Y(_01000_));
 NOR2x1_ASAP7_75t_R _43646_ (.A(net402),
    .B(_00844_),
    .Y(_14467_));
 AO21x1_ASAP7_75t_R _43647_ (.A1(net402),
    .A2(net3899),
    .B(_14467_),
    .Y(_01001_));
 NOR2x1_ASAP7_75t_R _43648_ (.A(net402),
    .B(_00843_),
    .Y(_14468_));
 AO21x1_ASAP7_75t_R _43649_ (.A1(net402),
    .A2(net3662),
    .B(_14468_),
    .Y(_01002_));
 NOR2x1_ASAP7_75t_R _43650_ (.A(net402),
    .B(_00842_),
    .Y(_14469_));
 AO21x1_ASAP7_75t_R _43651_ (.A1(net402),
    .A2(net3845),
    .B(_14469_),
    .Y(_01003_));
 NOR2x1_ASAP7_75t_R _43652_ (.A(net402),
    .B(_00841_),
    .Y(_14470_));
 AO21x1_ASAP7_75t_R _43653_ (.A1(net402),
    .A2(net3913),
    .B(_14470_),
    .Y(_01004_));
 NOR2x1_ASAP7_75t_R _43654_ (.A(net129),
    .B(_00840_),
    .Y(_14471_));
 AO21x1_ASAP7_75t_R _43655_ (.A1(net129),
    .A2(net3743),
    .B(_14471_),
    .Y(_01005_));
 NOR2x1_ASAP7_75t_R _43656_ (.A(net129),
    .B(_00839_),
    .Y(_14473_));
 AO21x1_ASAP7_75t_R _43657_ (.A1(net405),
    .A2(net3728),
    .B(_14473_),
    .Y(_01006_));
 TAPCELL_ASAP7_75t_R PHY_9 ();
 NOR2x1_ASAP7_75t_R _43659_ (.A(net402),
    .B(_00838_),
    .Y(_14475_));
 AO21x1_ASAP7_75t_R _43660_ (.A1(net402),
    .A2(net3606),
    .B(_14475_),
    .Y(_01007_));
 NOR2x1_ASAP7_75t_R _43661_ (.A(net402),
    .B(_00837_),
    .Y(_14476_));
 AO21x1_ASAP7_75t_R _43662_ (.A1(net402),
    .A2(net3812),
    .B(_14476_),
    .Y(_01008_));
 NOR2x1_ASAP7_75t_R _43663_ (.A(net402),
    .B(_00836_),
    .Y(_14477_));
 AO21x1_ASAP7_75t_R _43664_ (.A1(net402),
    .A2(net3776),
    .B(_14477_),
    .Y(_01009_));
 TAPCELL_ASAP7_75t_R PHY_8 ();
 NOR2x1_ASAP7_75t_R _43666_ (.A(net402),
    .B(_00835_),
    .Y(_14480_));
 AO21x1_ASAP7_75t_R _43667_ (.A1(net402),
    .A2(net3630),
    .B(_14480_),
    .Y(_01010_));
 NOR2x1_ASAP7_75t_R _43668_ (.A(net402),
    .B(_00834_),
    .Y(_14481_));
 AO21x1_ASAP7_75t_R _43669_ (.A1(net402),
    .A2(net3653),
    .B(_14481_),
    .Y(_01011_));
 NOR2x1_ASAP7_75t_R _43670_ (.A(net402),
    .B(_00833_),
    .Y(_14482_));
 AO21x1_ASAP7_75t_R _43671_ (.A1(net402),
    .A2(net3827),
    .B(_14482_),
    .Y(_01012_));
 NOR2x1_ASAP7_75t_R _43672_ (.A(net402),
    .B(_00832_),
    .Y(_14483_));
 AO21x1_ASAP7_75t_R _43673_ (.A1(net402),
    .A2(net3612),
    .B(_14483_),
    .Y(_01013_));
 NOR2x1_ASAP7_75t_R _43674_ (.A(net402),
    .B(_00831_),
    .Y(_14484_));
 AO21x1_ASAP7_75t_R _43675_ (.A1(net402),
    .A2(net3597),
    .B(_14484_),
    .Y(_01014_));
 NOR2x1_ASAP7_75t_R _43676_ (.A(net402),
    .B(_00830_),
    .Y(_14486_));
 AO21x1_ASAP7_75t_R _43677_ (.A1(net402),
    .A2(net3797),
    .B(_14486_),
    .Y(_01015_));
 NOR2x1_ASAP7_75t_R _43678_ (.A(net402),
    .B(_00829_),
    .Y(_14487_));
 AO21x1_ASAP7_75t_R _43679_ (.A1(net402),
    .A2(net3878),
    .B(_14487_),
    .Y(_01016_));
 TAPCELL_ASAP7_75t_R PHY_7 ();
 NOR2x1_ASAP7_75t_R _43681_ (.A(net402),
    .B(_00828_),
    .Y(_14489_));
 AO21x1_ASAP7_75t_R _43682_ (.A1(net402),
    .A2(net3842),
    .B(_14489_),
    .Y(_01017_));
 NOR2x1_ASAP7_75t_R _43683_ (.A(net402),
    .B(_00827_),
    .Y(_14490_));
 AO21x1_ASAP7_75t_R _43684_ (.A1(net402),
    .A2(net3627),
    .B(_14490_),
    .Y(_01018_));
 NOR2x1_ASAP7_75t_R _43685_ (.A(net402),
    .B(_00826_),
    .Y(_14492_));
 AO21x1_ASAP7_75t_R _43686_ (.A1(net402),
    .A2(net3589),
    .B(_14492_),
    .Y(_01019_));
 TAPCELL_ASAP7_75t_R PHY_6 ();
 NOR2x1_ASAP7_75t_R _43688_ (.A(net402),
    .B(_00825_),
    .Y(_14494_));
 AO21x1_ASAP7_75t_R _43689_ (.A1(net402),
    .A2(net3674),
    .B(_14494_),
    .Y(_01020_));
 NOR2x1_ASAP7_75t_R _43690_ (.A(net402),
    .B(_00824_),
    .Y(_14495_));
 AO21x1_ASAP7_75t_R _43691_ (.A1(net402),
    .A2(net3905),
    .B(_14495_),
    .Y(_01021_));
 NOR2x1_ASAP7_75t_R _43692_ (.A(net402),
    .B(_00823_),
    .Y(_14496_));
 AO21x1_ASAP7_75t_R _43693_ (.A1(net402),
    .A2(net3677),
    .B(_14496_),
    .Y(_01022_));
 NOR2x1_ASAP7_75t_R _43694_ (.A(net402),
    .B(_00822_),
    .Y(_14497_));
 AO21x1_ASAP7_75t_R _43695_ (.A1(net402),
    .A2(net3600),
    .B(_14497_),
    .Y(_01023_));
 NOR2x1_ASAP7_75t_R _43696_ (.A(net402),
    .B(_00821_),
    .Y(_14499_));
 AO21x1_ASAP7_75t_R _43697_ (.A1(net402),
    .A2(net3858),
    .B(_14499_),
    .Y(_01024_));
 NOR2x1_ASAP7_75t_R _43698_ (.A(net402),
    .B(_00820_),
    .Y(_14500_));
 AO21x1_ASAP7_75t_R _43699_ (.A1(net402),
    .A2(net3603),
    .B(_14500_),
    .Y(_01025_));
 NOR2x1_ASAP7_75t_R _43700_ (.A(net403),
    .B(_00819_),
    .Y(_14501_));
 AO21x1_ASAP7_75t_R _43701_ (.A1(net403),
    .A2(net3818),
    .B(_14501_),
    .Y(_01026_));
 TAPCELL_ASAP7_75t_R PHY_5 ();
 NOR2x1_ASAP7_75t_R _43703_ (.A(net403),
    .B(_00818_),
    .Y(_14503_));
 AO21x1_ASAP7_75t_R _43704_ (.A1(net403),
    .A2(net3791),
    .B(_14503_),
    .Y(_01027_));
 NOR2x1_ASAP7_75t_R _43705_ (.A(net403),
    .B(_00817_),
    .Y(_14505_));
 AO21x1_ASAP7_75t_R _43706_ (.A1(net403),
    .A2(net3949),
    .B(_14505_),
    .Y(_01028_));
 NOR2x1_ASAP7_75t_R _43707_ (.A(net403),
    .B(_00816_),
    .Y(_14506_));
 AO21x1_ASAP7_75t_R _43708_ (.A1(net403),
    .A2(net3919),
    .B(_14506_),
    .Y(_01029_));
 TAPCELL_ASAP7_75t_R PHY_4 ();
 NOR2x1_ASAP7_75t_R _43710_ (.A(net403),
    .B(_00815_),
    .Y(_14508_));
 AO21x1_ASAP7_75t_R _43711_ (.A1(net403),
    .A2(net3958),
    .B(_14508_),
    .Y(_01030_));
 NOR2x1_ASAP7_75t_R _43712_ (.A(net403),
    .B(_00814_),
    .Y(_14509_));
 AO21x1_ASAP7_75t_R _43713_ (.A1(net403),
    .A2(net3961),
    .B(_14509_),
    .Y(_01031_));
 NOR2x1_ASAP7_75t_R _43714_ (.A(net403),
    .B(_00813_),
    .Y(_14510_));
 AO21x1_ASAP7_75t_R _43715_ (.A1(net403),
    .A2(net3925),
    .B(_14510_),
    .Y(_01032_));
 NOR2x1_ASAP7_75t_R _43716_ (.A(net405),
    .B(_00812_),
    .Y(_14512_));
 AO21x1_ASAP7_75t_R _43717_ (.A1(net405),
    .A2(net3988),
    .B(_14512_),
    .Y(_01033_));
 NOR2x1_ASAP7_75t_R _43718_ (.A(net403),
    .B(_00811_),
    .Y(_14513_));
 AO21x1_ASAP7_75t_R _43719_ (.A1(net403),
    .A2(net3896),
    .B(_14513_),
    .Y(_01034_));
 NOR2x1_ASAP7_75t_R _43720_ (.A(net403),
    .B(_00810_),
    .Y(_14514_));
 AO21x1_ASAP7_75t_R _43721_ (.A1(net403),
    .A2(net3833),
    .B(_14514_),
    .Y(_01035_));
 NOR2x1_ASAP7_75t_R _43722_ (.A(net403),
    .B(_00809_),
    .Y(_14515_));
 AO21x1_ASAP7_75t_R _43723_ (.A1(net403),
    .A2(net3922),
    .B(_14515_),
    .Y(_01036_));
 TAPCELL_ASAP7_75t_R PHY_3 ();
 NOR2x1_ASAP7_75t_R _43725_ (.A(net402),
    .B(_00808_),
    .Y(_14518_));
 AO21x1_ASAP7_75t_R _43726_ (.A1(net402),
    .A2(net3568),
    .B(_14518_),
    .Y(_01037_));
 NOR2x1_ASAP7_75t_R _43727_ (.A(net403),
    .B(_00807_),
    .Y(_14519_));
 AO21x1_ASAP7_75t_R _43728_ (.A1(net403),
    .A2(net3937),
    .B(_14519_),
    .Y(_01038_));
 NOR2x1_ASAP7_75t_R _43729_ (.A(net403),
    .B(_00806_),
    .Y(_14520_));
 AO21x1_ASAP7_75t_R _43730_ (.A1(net403),
    .A2(net3884),
    .B(_14520_),
    .Y(_01039_));
 TAPCELL_ASAP7_75t_R PHY_2 ();
 NOR2x1_ASAP7_75t_R _43732_ (.A(net405),
    .B(_00805_),
    .Y(_14522_));
 AO21x1_ASAP7_75t_R _43733_ (.A1(net405),
    .A2(net3985),
    .B(_14522_),
    .Y(_01040_));
 NOR2x1_ASAP7_75t_R _43734_ (.A(net403),
    .B(_00804_),
    .Y(_14523_));
 AO21x1_ASAP7_75t_R _43735_ (.A1(net403),
    .A2(net3809),
    .B(_14523_),
    .Y(_01041_));
 NOR2x1_ASAP7_75t_R _43736_ (.A(net403),
    .B(_00803_),
    .Y(_14525_));
 AO21x1_ASAP7_75t_R _43737_ (.A1(net403),
    .A2(net3782),
    .B(_14525_),
    .Y(_01042_));
 NOR2x1_ASAP7_75t_R _43738_ (.A(net403),
    .B(_00802_),
    .Y(_14526_));
 AO21x1_ASAP7_75t_R _43739_ (.A1(net403),
    .A2(net3803),
    .B(_14526_),
    .Y(_01043_));
 NOR2x1_ASAP7_75t_R _43740_ (.A(net403),
    .B(_00801_),
    .Y(_14527_));
 AO21x1_ASAP7_75t_R _43741_ (.A1(net403),
    .A2(net3931),
    .B(_14527_),
    .Y(_01044_));
 NOR2x1_ASAP7_75t_R _43742_ (.A(net403),
    .B(_00800_),
    .Y(_14528_));
 AO21x1_ASAP7_75t_R _43743_ (.A1(net403),
    .A2(net3946),
    .B(_14528_),
    .Y(_01045_));
 NOR2x1_ASAP7_75t_R _43744_ (.A(net405),
    .B(_00799_),
    .Y(_14529_));
 AO21x1_ASAP7_75t_R _43745_ (.A1(net405),
    .A2(net3996),
    .B(_14529_),
    .Y(_01046_));
 TAPCELL_ASAP7_75t_R PHY_1 ();
 NOR2x1_ASAP7_75t_R _43747_ (.A(net403),
    .B(_00798_),
    .Y(_14532_));
 AO21x1_ASAP7_75t_R _43748_ (.A1(net403),
    .A2(net3973),
    .B(_14532_),
    .Y(_01047_));
 NOR2x1_ASAP7_75t_R _43749_ (.A(net404),
    .B(_00797_),
    .Y(_14533_));
 AO21x1_ASAP7_75t_R _43750_ (.A1(net404),
    .A2(net4094),
    .B(_14533_),
    .Y(_01048_));
 NOR2x1_ASAP7_75t_R _43751_ (.A(net405),
    .B(_00796_),
    .Y(_14534_));
 AO21x1_ASAP7_75t_R _43752_ (.A1(net405),
    .A2(net3979),
    .B(_14534_),
    .Y(_01049_));
 NOR2x1_ASAP7_75t_R _43753_ (.A(net403),
    .B(_00795_),
    .Y(_14535_));
 AO21x1_ASAP7_75t_R _43754_ (.A1(net403),
    .A2(net3887),
    .B(_14535_),
    .Y(_01050_));
 NOR2x1_ASAP7_75t_R _43755_ (.A(net403),
    .B(_00794_),
    .Y(_14537_));
 AO21x1_ASAP7_75t_R _43756_ (.A1(net403),
    .A2(net3852),
    .B(_14537_),
    .Y(_01051_));
 NOR2x1_ASAP7_75t_R _43757_ (.A(net403),
    .B(_00793_),
    .Y(_14538_));
 AO21x1_ASAP7_75t_R _43758_ (.A1(net403),
    .A2(net3761),
    .B(_14538_),
    .Y(_01052_));
 NOR2x1_ASAP7_75t_R _43759_ (.A(net403),
    .B(_00792_),
    .Y(_14539_));
 AO21x1_ASAP7_75t_R _43760_ (.A1(net403),
    .A2(net3821),
    .B(_14539_),
    .Y(_01053_));
 NOR2x1_ASAP7_75t_R _43761_ (.A(net403),
    .B(_00791_),
    .Y(_14540_));
 AO21x1_ASAP7_75t_R _43762_ (.A1(net403),
    .A2(net3785),
    .B(_14540_),
    .Y(_01054_));
 NOR2x1_ASAP7_75t_R _43763_ (.A(net403),
    .B(_00790_),
    .Y(_14541_));
 AO21x1_ASAP7_75t_R _43764_ (.A1(net403),
    .A2(net3910),
    .B(_14541_),
    .Y(_01055_));
 NOR2x1_ASAP7_75t_R _43765_ (.A(net403),
    .B(_00789_),
    .Y(_14543_));
 AO21x1_ASAP7_75t_R _43766_ (.A1(net403),
    .A2(net3830),
    .B(_14543_),
    .Y(_01056_));
 NOR2x1_ASAP7_75t_R _43767_ (.A(net403),
    .B(_00788_),
    .Y(_14544_));
 AO21x1_ASAP7_75t_R _43768_ (.A1(net403),
    .A2(net3824),
    .B(_14544_),
    .Y(_01057_));
 TAPCELL_ASAP7_75t_R PHY_0 ();
 AO21x1_ASAP7_75t_R _43770_ (.A1(_22105_),
    .A2(_00919_),
    .B(net401),
    .Y(_00922_));
 INVx1_ASAP7_75t_R _43771_ (.A(_00417_),
    .Y(_14546_));
 XOR2x2_ASAP7_75t_R _43772_ (.A(_00525_),
    .B(_00918_),
    .Y(_14547_));
 AND3x1_ASAP7_75t_R _43773_ (.A(_14547_),
    .B(_22105_),
    .C(_00919_),
    .Y(_14548_));
 AO21x1_ASAP7_75t_R _43774_ (.A1(_14546_),
    .A2(_00919_),
    .B(_14548_),
    .Y(_14549_));
 AND2x2_ASAP7_75t_R _43775_ (.A(_14549_),
    .B(net399),
    .Y(_00923_));
 INVx1_ASAP7_75t_R _43776_ (.A(_00419_),
    .Y(_14551_));
 INVx1_ASAP7_75t_R _43777_ (.A(_00919_),
    .Y(_14552_));
 NOR2x1_ASAP7_75t_R _43778_ (.A(_14552_),
    .B(_14547_),
    .Y(_14553_));
 AND3x1_ASAP7_75t_R _43779_ (.A(_14547_),
    .B(_14546_),
    .C(_00919_),
    .Y(_14554_));
 AO21x1_ASAP7_75t_R _43780_ (.A1(_14551_),
    .A2(_14553_),
    .B(_14554_),
    .Y(_14555_));
 AND2x2_ASAP7_75t_R _43781_ (.A(_14555_),
    .B(net399),
    .Y(_00924_));
 INVx1_ASAP7_75t_R _43782_ (.A(_00418_),
    .Y(_14556_));
 AO21x1_ASAP7_75t_R _43783_ (.A1(_14556_),
    .A2(_14553_),
    .B(_14548_),
    .Y(_14557_));
 AND2x2_ASAP7_75t_R _43784_ (.A(_14557_),
    .B(net398),
    .Y(_00925_));
 NOR2x2_ASAP7_75t_R _43785_ (.A(_00919_),
    .B(_14547_),
    .Y(_14559_));
 AO21x1_ASAP7_75t_R _43786_ (.A1(_22105_),
    .A2(_14559_),
    .B(_14548_),
    .Y(_14560_));
 OA21x2_ASAP7_75t_R _43787_ (.A1(_14560_),
    .A2(_14554_),
    .B(net398),
    .Y(_00926_));
 AO21x1_ASAP7_75t_R _43788_ (.A1(_14546_),
    .A2(_14559_),
    .B(_14554_),
    .Y(_14561_));
 AND2x2_ASAP7_75t_R _43789_ (.A(_14561_),
    .B(net399),
    .Y(_00927_));
 AND3x1_ASAP7_75t_R _43790_ (.A(_14559_),
    .B(net399),
    .C(_14551_),
    .Y(_00928_));
 AND3x1_ASAP7_75t_R _43791_ (.A(_14559_),
    .B(net399),
    .C(_14556_),
    .Y(_00929_));
 AND2x2_ASAP7_75t_R _43792_ (.A(_22107_),
    .B(_17523_),
    .Y(_14562_));
 INVx1_ASAP7_75t_R _43793_ (.A(_14562_),
    .Y(_14563_));
 AND4x1_ASAP7_75t_R _43794_ (.A(_14563_),
    .B(net398),
    .C(net3815),
    .D(_00420_),
    .Y(_01061_));
 NOR2x1_ASAP7_75t_R _43795_ (.A(net401),
    .B(\u0.r0.rcnt[0] ),
    .Y(_01062_));
 NOR2x1_ASAP7_75t_R _43796_ (.A(net401),
    .B(_00916_),
    .Y(_01063_));
 NOR2x1_ASAP7_75t_R _43797_ (.A(net401),
    .B(_00919_),
    .Y(_01064_));
 AND2x2_ASAP7_75t_R _43798_ (.A(_14547_),
    .B(net398),
    .Y(_01065_));
 NAND2x1_ASAP7_75t_R _43799_ (.A(net398),
    .B(_14562_),
    .Y(_14565_));
 OA211x2_ASAP7_75t_R _43800_ (.A1(net3839),
    .A2(_00787_),
    .B(_14565_),
    .C(net3815),
    .Y(_01058_));
 INVx1_ASAP7_75t_R _43801_ (.A(_17523_),
    .Y(_14566_));
 OAI21x1_ASAP7_75t_R _43802_ (.A1(_00786_),
    .A2(_00787_),
    .B(net398),
    .Y(_14567_));
 AO21x1_ASAP7_75t_R _43803_ (.A1(_14566_),
    .A2(_22107_),
    .B(_14567_),
    .Y(_14568_));
 AND2x2_ASAP7_75t_R _43804_ (.A(_14568_),
    .B(net3815),
    .Y(_01059_));
 XOR2x1_ASAP7_75t_R _43805_ (.A(_00785_),
    .Y(_14570_),
    .B(_00920_));
 OA211x2_ASAP7_75t_R _43806_ (.A1(net3839),
    .A2(_14570_),
    .B(_14565_),
    .C(net3815),
    .Y(_01060_));
 HAxp5_ASAP7_75t_R _43807_ (.A(\u0.r0.rcnt_next[0] ),
    .B(_22101_),
    .CON(_00417_),
    .SN(_00916_));
 HAxp5_ASAP7_75t_R _43808_ (.A(\u0.r0.rcnt_next[0] ),
    .B(\u0.r0.rcnt[1] ),
    .CON(_00418_),
    .SN(_22102_));
 HAxp5_ASAP7_75t_R _43809_ (.A(\u0.r0.rcnt[0] ),
    .B(_22101_),
    .CON(_00419_),
    .SN(_22103_));
 HAxp5_ASAP7_75t_R _43810_ (.A(\u0.r0.rcnt[0] ),
    .B(\u0.r0.rcnt[1] ),
    .CON(_00917_),
    .SN(_22104_));
 HAxp5_ASAP7_75t_R _43811_ (.A(\u0.r0.rcnt[2] ),
    .B(_22105_),
    .CON(_00918_),
    .SN(_00919_));
 HAxp5_ASAP7_75t_R _43812_ (.A(_22106_),
    .B(_22107_),
    .CON(_00920_),
    .SN(_00420_));
 DFFLQNx2_ASAP7_75t_R _43813_ (.QN(_00397_),
    .CLK(net935),
    .D(_00922_));
 DFFLQNx2_ASAP7_75t_R _43814_ (.QN(_00399_),
    .CLK(net934),
    .D(_00923_));
 DFFLQNx2_ASAP7_75t_R _43815_ (.QN(_00401_),
    .CLK(net933),
    .D(_00924_));
 DFFLQNx2_ASAP7_75t_R _43816_ (.QN(_00402_),
    .CLK(net932),
    .D(_00925_));
 DFFLQNx2_ASAP7_75t_R _43817_ (.QN(_00403_),
    .CLK(net931),
    .D(_00926_));
 DFFLQNx2_ASAP7_75t_R _43818_ (.QN(_00404_),
    .CLK(net930),
    .D(_00927_));
 DFFLQNx2_ASAP7_75t_R _43819_ (.QN(_00406_),
    .CLK(net929),
    .D(_00928_));
 DFFLQNx2_ASAP7_75t_R _43820_ (.QN(_00408_),
    .CLK(net928),
    .D(_00929_));
 DFFLQNx2_ASAP7_75t_R _43821_ (.QN(_00915_),
    .CLK(net927),
    .D(net3965));
 DFFLQNx2_ASAP7_75t_R _43822_ (.QN(_00914_),
    .CLK(net926),
    .D(net3868));
 DFFLQNx2_ASAP7_75t_R _43823_ (.QN(_00913_),
    .CLK(net925),
    .D(net3759));
 DFFLQNx2_ASAP7_75t_R _43824_ (.QN(_00912_),
    .CLK(net924),
    .D(net3994));
 DFFLQNx2_ASAP7_75t_R _43825_ (.QN(_00911_),
    .CLK(net923),
    .D(net3643));
 DFFLQNx2_ASAP7_75t_R _43826_ (.QN(_00910_),
    .CLK(net922),
    .D(_00935_));
 DFFLQNx2_ASAP7_75t_R _43827_ (.QN(_00909_),
    .CLK(net921),
    .D(net3572));
 DFFLQNx2_ASAP7_75t_R _43828_ (.QN(_00908_),
    .CLK(net920),
    .D(net3622));
 DFFLQNx2_ASAP7_75t_R _43829_ (.QN(_00907_),
    .CLK(net919),
    .D(net3566));
 DFFLQNx2_ASAP7_75t_R _43830_ (.QN(_00906_),
    .CLK(net918),
    .D(net3575));
 DFFLQNx2_ASAP7_75t_R _43831_ (.QN(_00905_),
    .CLK(net917),
    .D(net3587));
 DFFLQNx2_ASAP7_75t_R _43832_ (.QN(_00904_),
    .CLK(net916),
    .D(net3765));
 DFFLQNx2_ASAP7_75t_R _43833_ (.QN(_00903_),
    .CLK(net915),
    .D(net3702));
 DFFLQNx2_ASAP7_75t_R _43834_ (.QN(_00902_),
    .CLK(net914),
    .D(net3756));
 DFFLQNx2_ASAP7_75t_R _43835_ (.QN(_00901_),
    .CLK(net913),
    .D(net3738));
 DFFLQNx2_ASAP7_75t_R _43836_ (.QN(_00900_),
    .CLK(net912),
    .D(net3726));
 DFFLQNx2_ASAP7_75t_R _43837_ (.QN(_00899_),
    .CLK(net911),
    .D(net3714));
 DFFLQNx2_ASAP7_75t_R _43838_ (.QN(_00898_),
    .CLK(net910),
    .D(net3666));
 DFFLQNx2_ASAP7_75t_R _43839_ (.QN(_00897_),
    .CLK(net909),
    .D(net3732));
 DFFLQNx2_ASAP7_75t_R _43840_ (.QN(_00896_),
    .CLK(net908),
    .D(net3753));
 DFFLQNx2_ASAP7_75t_R _43841_ (.QN(_00895_),
    .CLK(net907),
    .D(net3723));
 DFFLQNx2_ASAP7_75t_R _43842_ (.QN(_00894_),
    .CLK(net906),
    .D(net3711));
 DFFLQNx2_ASAP7_75t_R _43843_ (.QN(_00893_),
    .CLK(net905),
    .D(net3578));
 DFFLQNx2_ASAP7_75t_R _43844_ (.QN(_00892_),
    .CLK(net904),
    .D(net3687));
 DFFLQNx2_ASAP7_75t_R _43845_ (.QN(_00891_),
    .CLK(net903),
    .D(net3871));
 DFFLQNx2_ASAP7_75t_R _43846_ (.QN(_00890_),
    .CLK(net902),
    .D(net3953));
 DFFLQNx2_ASAP7_75t_R _43847_ (.QN(_00889_),
    .CLK(net901),
    .D(net3768));
 DFFLQNx2_ASAP7_75t_R _43848_ (.QN(_00888_),
    .CLK(net900),
    .D(net3929));
 DFFLQNx2_ASAP7_75t_R _43849_ (.QN(_00887_),
    .CLK(net899),
    .D(net3801));
 DFFLQNx2_ASAP7_75t_R _43850_ (.QN(_00886_),
    .CLK(net898),
    .D(net3935));
 DFFLQNx2_ASAP7_75t_R _43851_ (.QN(_00885_),
    .CLK(net897),
    .D(net3780));
 DFFLQNx2_ASAP7_75t_R _43852_ (.QN(_00884_),
    .CLK(net896),
    .D(net3774));
 DFFLQNx2_ASAP7_75t_R _43853_ (.QN(_00883_),
    .CLK(net895),
    .D(net3750));
 DFFLQNx2_ASAP7_75t_R _43854_ (.QN(_00882_),
    .CLK(net894),
    .D(net3717));
 DFFLQNx2_ASAP7_75t_R _43855_ (.QN(_00881_),
    .CLK(net893),
    .D(net3735));
 DFFLQNx2_ASAP7_75t_R _43856_ (.QN(_00880_),
    .CLK(net892),
    .D(net3640));
 DFFLQNx2_ASAP7_75t_R _43857_ (.QN(_00879_),
    .CLK(net891),
    .D(net3977));
 DFFLQNx2_ASAP7_75t_R _43858_ (.QN(_00878_),
    .CLK(net890),
    .D(_00967_));
 DFFLQNx2_ASAP7_75t_R _43859_ (.QN(_00877_),
    .CLK(net889),
    .D(net3741));
 DFFLQNx2_ASAP7_75t_R _43860_ (.QN(_00876_),
    .CLK(net888),
    .D(net3720));
 DFFLQNx2_ASAP7_75t_R _43861_ (.QN(_00875_),
    .CLK(net887),
    .D(net3693));
 DFFLQNx2_ASAP7_75t_R _43862_ (.QN(_00874_),
    .CLK(net886),
    .D(net3681));
 DFFLQNx2_ASAP7_75t_R _43863_ (.QN(_00873_),
    .CLK(net885),
    .D(net3699));
 DFFLQNx2_ASAP7_75t_R _43864_ (.QN(_00872_),
    .CLK(net884),
    .D(net3646));
 DFFLQNx2_ASAP7_75t_R _43865_ (.QN(_00871_),
    .CLK(net883),
    .D(net3637));
 DFFLQNx2_ASAP7_75t_R _43866_ (.QN(_00870_),
    .CLK(net882),
    .D(net3625));
 DFFLQNx2_ASAP7_75t_R _43867_ (.QN(_00869_),
    .CLK(net881),
    .D(net3903));
 DFFLQNx2_ASAP7_75t_R _43868_ (.QN(_00868_),
    .CLK(net880),
    .D(net4003));
 DFFLQNx2_ASAP7_75t_R _43869_ (.QN(_00867_),
    .CLK(net879),
    .D(net3684));
 DFFLQNx2_ASAP7_75t_R _43870_ (.QN(_00866_),
    .CLK(net878),
    .D(net3669));
 DFFLQNx2_ASAP7_75t_R _43871_ (.QN(_00865_),
    .CLK(net877),
    .D(net3610));
 DFFLQNx2_ASAP7_75t_R _43872_ (.QN(_00864_),
    .CLK(net876),
    .D(net3696));
 DFFLQNx2_ASAP7_75t_R _43873_ (.QN(_00863_),
    .CLK(net875),
    .D(net3944));
 DFFLQNx2_ASAP7_75t_R _43874_ (.QN(_00862_),
    .CLK(net874),
    .D(net3595));
 DFFLQNx2_ASAP7_75t_R _43875_ (.QN(_00861_),
    .CLK(net873),
    .D(net3634));
 DFFLQNx2_ASAP7_75t_R _43876_ (.QN(_00860_),
    .CLK(net872),
    .D(net3581));
 DFFLQNx2_ASAP7_75t_R _43877_ (.QN(_00859_),
    .CLK(net871),
    .D(net3747));
 DFFLQNx2_ASAP7_75t_R _43878_ (.QN(_00858_),
    .CLK(net870),
    .D(net3708));
 DFFLQNx2_ASAP7_75t_R _43879_ (.QN(_00857_),
    .CLK(net869),
    .D(net3649));
 DFFLQNx2_ASAP7_75t_R _43880_ (.QN(_00856_),
    .CLK(net868),
    .D(net3705));
 DFFLQNx2_ASAP7_75t_R _43881_ (.QN(_00855_),
    .CLK(net867),
    .D(net3619));
 DFFLQNx2_ASAP7_75t_R _43882_ (.QN(_00854_),
    .CLK(net866),
    .D(net3956));
 DFFLQNx2_ASAP7_75t_R _43883_ (.QN(_00853_),
    .CLK(net865),
    .D(net3690));
 DFFLQNx2_ASAP7_75t_R _43884_ (.QN(_00852_),
    .CLK(net864),
    .D(net3657));
 DFFLQNx2_ASAP7_75t_R _43885_ (.QN(_00851_),
    .CLK(net863),
    .D(net3584));
 DFFLQNx2_ASAP7_75t_R _43886_ (.QN(_00850_),
    .CLK(net862),
    .D(net3616));
 DFFLQNx2_ASAP7_75t_R _43887_ (.QN(_00849_),
    .CLK(net861),
    .D(net3672));
 DFFLQNx2_ASAP7_75t_R _43888_ (.QN(_00848_),
    .CLK(net860),
    .D(net3850));
 DFFLQNx2_ASAP7_75t_R _43889_ (.QN(_00847_),
    .CLK(net859),
    .D(net3837));
 DFFLQNx2_ASAP7_75t_R _43890_ (.QN(_00846_),
    .CLK(net858),
    .D(net3789));
 DFFLQNx2_ASAP7_75t_R _43891_ (.QN(_00845_),
    .CLK(net857),
    .D(net3807));
 DFFLQNx2_ASAP7_75t_R _43892_ (.QN(_00844_),
    .CLK(net856),
    .D(net3900));
 DFFLQNx2_ASAP7_75t_R _43893_ (.QN(_00843_),
    .CLK(net855),
    .D(net3663));
 DFFLQNx2_ASAP7_75t_R _43894_ (.QN(_00842_),
    .CLK(net854),
    .D(net3846));
 DFFLQNx2_ASAP7_75t_R _43895_ (.QN(_00841_),
    .CLK(net853),
    .D(net3914));
 DFFLQNx2_ASAP7_75t_R _43896_ (.QN(_00840_),
    .CLK(net852),
    .D(net3744));
 DFFLQNx2_ASAP7_75t_R _43897_ (.QN(_00839_),
    .CLK(net851),
    .D(net3729));
 DFFLQNx2_ASAP7_75t_R _43898_ (.QN(_00838_),
    .CLK(net850),
    .D(net3607));
 DFFLQNx2_ASAP7_75t_R _43899_ (.QN(_00837_),
    .CLK(net849),
    .D(net3813));
 DFFLQNx2_ASAP7_75t_R _43900_ (.QN(_00836_),
    .CLK(net848),
    .D(net3777));
 DFFLQNx2_ASAP7_75t_R _43901_ (.QN(_00835_),
    .CLK(net847),
    .D(net3631));
 DFFLQNx2_ASAP7_75t_R _43902_ (.QN(_00834_),
    .CLK(net846),
    .D(net3654));
 DFFLQNx2_ASAP7_75t_R _43903_ (.QN(_00833_),
    .CLK(net845),
    .D(net3828));
 DFFLQNx2_ASAP7_75t_R _43904_ (.QN(_00832_),
    .CLK(net844),
    .D(net3613));
 DFFLQNx2_ASAP7_75t_R _43905_ (.QN(_00831_),
    .CLK(net843),
    .D(net3598));
 DFFLQNx2_ASAP7_75t_R _43906_ (.QN(_00830_),
    .CLK(net842),
    .D(net3798));
 DFFLQNx2_ASAP7_75t_R _43907_ (.QN(_00829_),
    .CLK(net841),
    .D(net3879));
 DFFLQNx2_ASAP7_75t_R _43908_ (.QN(_00828_),
    .CLK(net840),
    .D(net3843));
 DFFLQNx2_ASAP7_75t_R _43909_ (.QN(_00827_),
    .CLK(net839),
    .D(net3628));
 DFFLQNx2_ASAP7_75t_R _43910_ (.QN(_00826_),
    .CLK(net838),
    .D(net3590));
 DFFLQNx2_ASAP7_75t_R _43911_ (.QN(_00825_),
    .CLK(net837),
    .D(net3675));
 DFFLQNx2_ASAP7_75t_R _43912_ (.QN(_00824_),
    .CLK(net836),
    .D(net3906));
 DFFLQNx2_ASAP7_75t_R _43913_ (.QN(_00823_),
    .CLK(net835),
    .D(net3678));
 DFFLQNx2_ASAP7_75t_R _43914_ (.QN(_00822_),
    .CLK(net834),
    .D(net3601));
 DFFLQNx2_ASAP7_75t_R _43915_ (.QN(_00821_),
    .CLK(net833),
    .D(net3859));
 DFFLQNx2_ASAP7_75t_R _43916_ (.QN(_00820_),
    .CLK(net832),
    .D(net3604));
 DFFLQNx2_ASAP7_75t_R _43917_ (.QN(_00819_),
    .CLK(net831),
    .D(net3819));
 DFFLQNx2_ASAP7_75t_R _43918_ (.QN(_00818_),
    .CLK(net830),
    .D(net3792));
 DFFLQNx2_ASAP7_75t_R _43919_ (.QN(_00817_),
    .CLK(net829),
    .D(net3950));
 DFFLQNx2_ASAP7_75t_R _43920_ (.QN(_00816_),
    .CLK(net828),
    .D(net3920));
 DFFLQNx2_ASAP7_75t_R _43921_ (.QN(_00815_),
    .CLK(net827),
    .D(net3959));
 DFFLQNx2_ASAP7_75t_R _43922_ (.QN(_00814_),
    .CLK(net826),
    .D(net3962));
 DFFLQNx2_ASAP7_75t_R _43923_ (.QN(_00813_),
    .CLK(net825),
    .D(net3926));
 DFFLQNx2_ASAP7_75t_R _43924_ (.QN(_00812_),
    .CLK(net824),
    .D(net3989));
 DFFLQNx2_ASAP7_75t_R _43925_ (.QN(_00811_),
    .CLK(net823),
    .D(net3897));
 DFFLQNx2_ASAP7_75t_R _43926_ (.QN(_00810_),
    .CLK(net822),
    .D(net3834));
 DFFLQNx2_ASAP7_75t_R _43927_ (.QN(_00809_),
    .CLK(net821),
    .D(net3923));
 DFFLQNx2_ASAP7_75t_R _43928_ (.QN(_00808_),
    .CLK(net820),
    .D(net3569));
 DFFLQNx2_ASAP7_75t_R _43929_ (.QN(_00807_),
    .CLK(net819),
    .D(net3938));
 DFFLQNx2_ASAP7_75t_R _43930_ (.QN(_00806_),
    .CLK(net818),
    .D(net3885));
 DFFLQNx2_ASAP7_75t_R _43931_ (.QN(_00805_),
    .CLK(net817),
    .D(net3986));
 DFFLQNx2_ASAP7_75t_R _43932_ (.QN(_00804_),
    .CLK(net816),
    .D(net3810));
 DFFLQNx2_ASAP7_75t_R _43933_ (.QN(_00803_),
    .CLK(net815),
    .D(net3783));
 DFFLQNx2_ASAP7_75t_R _43934_ (.QN(_00802_),
    .CLK(net814),
    .D(net3804));
 DFFLQNx2_ASAP7_75t_R _43935_ (.QN(_00801_),
    .CLK(net813),
    .D(net3932));
 DFFLQNx2_ASAP7_75t_R _43936_ (.QN(_00800_),
    .CLK(net812),
    .D(net3947));
 DFFLQNx2_ASAP7_75t_R _43937_ (.QN(_00799_),
    .CLK(net811),
    .D(net3997));
 DFFLQNx2_ASAP7_75t_R _43938_ (.QN(_00798_),
    .CLK(net810),
    .D(net3974));
 DFFLQNx2_ASAP7_75t_R _43939_ (.QN(_00797_),
    .CLK(net809),
    .D(_01048_));
 DFFLQNx2_ASAP7_75t_R _43940_ (.QN(_00796_),
    .CLK(net808),
    .D(net3980));
 DFFLQNx2_ASAP7_75t_R _43941_ (.QN(_00795_),
    .CLK(net807),
    .D(net3888));
 DFFLQNx2_ASAP7_75t_R _43942_ (.QN(_00794_),
    .CLK(net806),
    .D(net3853));
 DFFLQNx2_ASAP7_75t_R _43943_ (.QN(_00793_),
    .CLK(net805),
    .D(net3762));
 DFFLQNx2_ASAP7_75t_R _43944_ (.QN(_00792_),
    .CLK(net804),
    .D(net3822));
 DFFLQNx2_ASAP7_75t_R _43945_ (.QN(_00791_),
    .CLK(net803),
    .D(net3786));
 DFFLQNx2_ASAP7_75t_R _43946_ (.QN(_00790_),
    .CLK(net802),
    .D(net3911));
 DFFLQNx2_ASAP7_75t_R _43947_ (.QN(_00789_),
    .CLK(net801),
    .D(net3831));
 DFFLQNx2_ASAP7_75t_R _43948_ (.QN(_00788_),
    .CLK(net800),
    .D(net3825));
 DFFLQNx2_ASAP7_75t_R _43949_ (.QN(_00787_),
    .CLK(net799),
    .D(net3840));
 DFFLQNx2_ASAP7_75t_R _43950_ (.QN(_00786_),
    .CLK(net798),
    .D(net3816));
 DFFLQNx2_ASAP7_75t_R _43951_ (.QN(_00785_),
    .CLK(net797),
    .D(_01060_));
 DFFLQNx2_ASAP7_75t_R _43952_ (.QN(_00784_),
    .CLK(net796),
    .D(_00233_));
 DFFLQNx3_ASAP7_75t_R _43953_ (.CLK(net795),
    .D(_00234_),
    .QN(_00783_));
 DFFLQNx2_ASAP7_75t_R _43954_ (.QN(_00782_),
    .CLK(net794),
    .D(_00235_));
 DFFLQNx2_ASAP7_75t_R _43955_ (.QN(_00781_),
    .CLK(net793),
    .D(_00236_));
 DFFLQNx3_ASAP7_75t_R _43956_ (.CLK(net792),
    .D(_00237_),
    .QN(_00780_));
 DFFLQNx2_ASAP7_75t_R _43957_ (.QN(_00779_),
    .CLK(net791),
    .D(_00238_));
 DFFLQNx3_ASAP7_75t_R _43958_ (.CLK(net790),
    .D(_00239_),
    .QN(_00778_));
 DFFLQNx3_ASAP7_75t_R _43959_ (.CLK(net789),
    .D(_00240_),
    .QN(_00777_));
 DFFLQNx3_ASAP7_75t_R _43960_ (.CLK(net788),
    .D(_00185_),
    .QN(_00776_));
 DFFLQNx3_ASAP7_75t_R _43961_ (.CLK(net787),
    .D(_00186_),
    .QN(_00775_));
 DFFLQNx3_ASAP7_75t_R _43962_ (.CLK(net786),
    .D(_00187_),
    .QN(_00774_));
 DFFLQNx2_ASAP7_75t_R _43963_ (.QN(_00773_),
    .CLK(net785),
    .D(_00188_));
 DFFLQNx2_ASAP7_75t_R _43964_ (.QN(_00772_),
    .CLK(net784),
    .D(_00189_));
 DFFLQNx2_ASAP7_75t_R _43965_ (.QN(_00771_),
    .CLK(net783),
    .D(_00190_));
 DFFLQNx3_ASAP7_75t_R _43966_ (.CLK(net782),
    .D(_00191_),
    .QN(_00770_));
 DFFLQNx2_ASAP7_75t_R _43967_ (.QN(_00769_),
    .CLK(net781),
    .D(_00192_));
 DFFLQNx3_ASAP7_75t_R _43968_ (.CLK(net780),
    .D(_00217_),
    .QN(_00768_));
 DFFLQNx3_ASAP7_75t_R _43969_ (.CLK(net779),
    .D(_00218_),
    .QN(_00767_));
 DFFLQNx3_ASAP7_75t_R _43970_ (.CLK(net778),
    .D(_00219_),
    .QN(_00766_));
 DFFLQNx3_ASAP7_75t_R _43971_ (.CLK(net777),
    .D(_00220_),
    .QN(_00765_));
 DFFLQNx2_ASAP7_75t_R _43972_ (.QN(_00764_),
    .CLK(net776),
    .D(_00221_));
 DFFLQNx3_ASAP7_75t_R _43973_ (.CLK(net775),
    .D(_00222_),
    .QN(_00763_));
 DFFLQNx3_ASAP7_75t_R _43974_ (.CLK(net774),
    .D(_00223_),
    .QN(_00762_));
 DFFLQNx3_ASAP7_75t_R _43975_ (.CLK(net773),
    .D(_00224_),
    .QN(_00761_));
 DFFLQNx2_ASAP7_75t_R _43976_ (.QN(_00760_),
    .CLK(net772),
    .D(_00129_));
 DFFLQNx2_ASAP7_75t_R _43977_ (.QN(_00759_),
    .CLK(net771),
    .D(_00130_));
 DFFLQNx1_ASAP7_75t_R _43978_ (.CLK(net770),
    .D(_00131_),
    .QN(_00758_));
 DFFLQNx3_ASAP7_75t_R _43979_ (.CLK(net769),
    .D(_00132_),
    .QN(_00757_));
 DFFLQNx3_ASAP7_75t_R _43980_ (.CLK(net768),
    .D(_00133_),
    .QN(_00756_));
 DFFLQNx3_ASAP7_75t_R _43981_ (.CLK(net767),
    .D(_00134_),
    .QN(_00755_));
 DFFLQNx3_ASAP7_75t_R _43982_ (.CLK(net766),
    .D(_00135_),
    .QN(_00754_));
 DFFLQNx3_ASAP7_75t_R _43983_ (.CLK(net765),
    .D(_00136_),
    .QN(_00753_));
 DFFLQNx2_ASAP7_75t_R _43984_ (.QN(_00752_),
    .CLK(net764),
    .D(_00161_));
 DFFLQNx3_ASAP7_75t_R _43985_ (.CLK(net763),
    .D(_00162_),
    .QN(_00751_));
 DFFLQNx3_ASAP7_75t_R _43986_ (.CLK(net762),
    .D(_00163_),
    .QN(_00750_));
 DFFLQNx2_ASAP7_75t_R _43987_ (.QN(_00749_),
    .CLK(net761),
    .D(_00164_));
 DFFLQNx1_ASAP7_75t_R _43988_ (.CLK(net760),
    .D(_00165_),
    .QN(_00748_));
 DFFLQNx2_ASAP7_75t_R _43989_ (.QN(_00747_),
    .CLK(net759),
    .D(_00166_));
 DFFLQNx2_ASAP7_75t_R _43990_ (.QN(_00746_),
    .CLK(net758),
    .D(_00167_));
 DFFLQNx3_ASAP7_75t_R _43991_ (.CLK(net757),
    .D(_00168_),
    .QN(_00745_));
 DFFLQNx1_ASAP7_75t_R _43992_ (.CLK(net756),
    .D(_00193_),
    .QN(_00744_));
 DFFLQNx2_ASAP7_75t_R _43993_ (.QN(_00743_),
    .CLK(net755),
    .D(_00194_));
 DFFLQNx3_ASAP7_75t_R _43994_ (.CLK(net754),
    .D(_00195_),
    .QN(_00742_));
 DFFLQNx2_ASAP7_75t_R _43995_ (.QN(_00741_),
    .CLK(net753),
    .D(_00196_));
 DFFLQNx3_ASAP7_75t_R _43996_ (.CLK(net752),
    .D(_00197_),
    .QN(_00740_));
 DFFLQNx2_ASAP7_75t_R _43997_ (.QN(_00739_),
    .CLK(net751),
    .D(_00198_));
 DFFLQNx2_ASAP7_75t_R _43998_ (.QN(_00738_),
    .CLK(net750),
    .D(_00199_));
 DFFLQNx2_ASAP7_75t_R _43999_ (.QN(_00737_),
    .CLK(net749),
    .D(_00200_));
 DFFLQNx3_ASAP7_75t_R _44000_ (.CLK(net748),
    .D(_00225_),
    .QN(_00736_));
 DFFLQNx3_ASAP7_75t_R _44001_ (.CLK(net747),
    .D(_00226_),
    .QN(_00735_));
 DFFLQNx3_ASAP7_75t_R _44002_ (.CLK(net746),
    .D(_00227_),
    .QN(_00734_));
 DFFLQNx3_ASAP7_75t_R _44003_ (.CLK(net745),
    .D(_00228_),
    .QN(_00733_));
 DFFLQNx3_ASAP7_75t_R _44004_ (.CLK(net744),
    .D(_00229_),
    .QN(_00732_));
 DFFLQNx2_ASAP7_75t_R _44005_ (.QN(_00731_),
    .CLK(net743),
    .D(_00230_));
 DFFLQNx3_ASAP7_75t_R _44006_ (.CLK(net742),
    .D(_00231_),
    .QN(_00730_));
 DFFLQNx3_ASAP7_75t_R _44007_ (.CLK(net741),
    .D(_00232_),
    .QN(_00729_));
 DFFLQNx3_ASAP7_75t_R _44008_ (.CLK(net740),
    .D(_00137_),
    .QN(_00728_));
 DFFLQNx3_ASAP7_75t_R _44009_ (.CLK(net739),
    .D(_00138_),
    .QN(_00727_));
 DFFLQNx3_ASAP7_75t_R _44010_ (.CLK(net738),
    .D(_00139_),
    .QN(_00726_));
 DFFLQNx2_ASAP7_75t_R _44011_ (.QN(_00725_),
    .CLK(net737),
    .D(_00140_));
 DFFLQNx3_ASAP7_75t_R _44012_ (.CLK(net736),
    .D(_00141_),
    .QN(_00724_));
 DFFLQNx1_ASAP7_75t_R _44013_ (.CLK(net735),
    .D(_00142_),
    .QN(_00723_));
 DFFLQNx3_ASAP7_75t_R _44014_ (.CLK(net734),
    .D(_00143_),
    .QN(_00722_));
 DFFLQNx3_ASAP7_75t_R _44015_ (.CLK(net733),
    .D(_00144_),
    .QN(_00721_));
 DFFLQNx3_ASAP7_75t_R _44016_ (.CLK(net732),
    .D(_00169_),
    .QN(_00720_));
 DFFLQNx3_ASAP7_75t_R _44017_ (.CLK(net731),
    .D(_00170_),
    .QN(_00719_));
 DFFLQNx3_ASAP7_75t_R _44018_ (.CLK(net730),
    .D(_00171_),
    .QN(_00718_));
 DFFLQNx2_ASAP7_75t_R _44019_ (.QN(_00717_),
    .CLK(net729),
    .D(_00172_));
 DFFLQNx3_ASAP7_75t_R _44020_ (.CLK(net728),
    .D(_00173_),
    .QN(_00716_));
 DFFLQNx3_ASAP7_75t_R _44021_ (.CLK(net727),
    .D(_00174_),
    .QN(_00715_));
 DFFLQNx3_ASAP7_75t_R _44022_ (.CLK(net726),
    .D(_00175_),
    .QN(_00714_));
 DFFLQNx3_ASAP7_75t_R _44023_ (.CLK(net725),
    .D(_00176_),
    .QN(_00713_));
 DFFLQNx3_ASAP7_75t_R _44024_ (.CLK(net724),
    .D(_00201_),
    .QN(_00712_));
 DFFLQNx2_ASAP7_75t_R _44025_ (.QN(_00711_),
    .CLK(net723),
    .D(_00202_));
 DFFLQNx1_ASAP7_75t_R _44026_ (.CLK(net722),
    .D(_00203_),
    .QN(_00710_));
 DFFLQNx2_ASAP7_75t_R _44027_ (.QN(_00709_),
    .CLK(net721),
    .D(_00204_));
 DFFLQNx2_ASAP7_75t_R _44028_ (.QN(_00708_),
    .CLK(net720),
    .D(_00205_));
 DFFLQNx3_ASAP7_75t_R _44029_ (.CLK(net719),
    .D(_00206_),
    .QN(_00707_));
 DFFLQNx3_ASAP7_75t_R _44030_ (.CLK(net718),
    .D(_00207_),
    .QN(_00706_));
 DFFLQNx2_ASAP7_75t_R _44031_ (.QN(_00705_),
    .CLK(net717),
    .D(_00208_));
 DFFLQNx3_ASAP7_75t_R _44032_ (.CLK(net716),
    .D(_00241_),
    .QN(_00704_));
 DFFLQNx3_ASAP7_75t_R _44033_ (.CLK(net715),
    .D(_00242_),
    .QN(_00703_));
 DFFLQNx3_ASAP7_75t_R _44034_ (.CLK(net714),
    .D(_00243_),
    .QN(_00702_));
 DFFLQNx3_ASAP7_75t_R _44035_ (.CLK(net713),
    .D(_00244_),
    .QN(_00701_));
 DFFLQNx3_ASAP7_75t_R _44036_ (.CLK(net712),
    .D(_00245_),
    .QN(_00700_));
 DFFLQNx2_ASAP7_75t_R _44037_ (.QN(_00699_),
    .CLK(net711),
    .D(_00246_));
 DFFLQNx3_ASAP7_75t_R _44038_ (.CLK(net710),
    .D(_00247_),
    .QN(_00698_));
 DFFLQNx3_ASAP7_75t_R _44039_ (.CLK(net709),
    .D(_00248_),
    .QN(_00697_));
 DFFLQNx3_ASAP7_75t_R _44040_ (.CLK(net708),
    .D(_00145_),
    .QN(_00696_));
 DFFLQNx3_ASAP7_75t_R _44041_ (.CLK(net707),
    .D(_00146_),
    .QN(_00695_));
 DFFLQNx3_ASAP7_75t_R _44042_ (.CLK(net706),
    .D(_00147_),
    .QN(_00694_));
 DFFLQNx2_ASAP7_75t_R _44043_ (.QN(_00693_),
    .CLK(net705),
    .D(_00148_));
 DFFLQNx3_ASAP7_75t_R _44044_ (.CLK(net704),
    .D(_00149_),
    .QN(_00692_));
 DFFLQNx3_ASAP7_75t_R _44045_ (.CLK(net703),
    .D(_00150_),
    .QN(_00691_));
 DFFLQNx3_ASAP7_75t_R _44046_ (.CLK(net702),
    .D(_00151_),
    .QN(_00690_));
 DFFLQNx3_ASAP7_75t_R _44047_ (.CLK(net701),
    .D(_00152_),
    .QN(_00689_));
 DFFLQNx3_ASAP7_75t_R _44048_ (.CLK(net700),
    .D(_00177_),
    .QN(_00688_));
 DFFLQNx3_ASAP7_75t_R _44049_ (.CLK(net699),
    .D(_00178_),
    .QN(_00687_));
 DFFLQNx3_ASAP7_75t_R _44050_ (.CLK(net698),
    .D(_00179_),
    .QN(_00686_));
 DFFLQNx3_ASAP7_75t_R _44051_ (.CLK(net697),
    .D(_00180_),
    .QN(_00685_));
 DFFLQNx1_ASAP7_75t_R _44052_ (.CLK(net696),
    .D(_00181_),
    .QN(_00684_));
 DFFLQNx3_ASAP7_75t_R _44053_ (.CLK(net695),
    .D(_00182_),
    .QN(_00683_));
 DFFLQNx3_ASAP7_75t_R _44054_ (.CLK(net694),
    .D(_00183_),
    .QN(_00682_));
 DFFLQNx3_ASAP7_75t_R _44055_ (.CLK(net693),
    .D(_00184_),
    .QN(_00681_));
 DFFLQNx3_ASAP7_75t_R _44056_ (.CLK(net692),
    .D(_00209_),
    .QN(_00680_));
 DFFLQNx3_ASAP7_75t_R _44057_ (.CLK(net691),
    .D(_00210_),
    .QN(_00679_));
 DFFLQNx2_ASAP7_75t_R _44058_ (.QN(_00678_),
    .CLK(net690),
    .D(_00211_));
 DFFLQNx3_ASAP7_75t_R _44059_ (.CLK(net689),
    .D(_00212_),
    .QN(_00677_));
 DFFLQNx3_ASAP7_75t_R _44060_ (.CLK(net688),
    .D(_00213_),
    .QN(_00676_));
 DFFLQNx2_ASAP7_75t_R _44061_ (.QN(_00675_),
    .CLK(net687),
    .D(_00214_));
 DFFLQNx3_ASAP7_75t_R _44062_ (.CLK(net686),
    .D(_00215_),
    .QN(_00674_));
 DFFLQNx3_ASAP7_75t_R _44063_ (.CLK(net685),
    .D(_00216_),
    .QN(_00673_));
 DFFLQNx3_ASAP7_75t_R _44064_ (.CLK(net684),
    .D(_00249_),
    .QN(_00672_));
 DFFLQNx1_ASAP7_75t_R _44065_ (.CLK(net683),
    .D(_00250_),
    .QN(_00671_));
 DFFLQNx3_ASAP7_75t_R _44066_ (.CLK(net682),
    .D(_00251_),
    .QN(_00670_));
 DFFLQNx3_ASAP7_75t_R _44067_ (.CLK(net681),
    .D(_00252_),
    .QN(_00669_));
 DFFLQNx3_ASAP7_75t_R _44068_ (.CLK(net680),
    .D(_00253_),
    .QN(_00668_));
 DFFLQNx3_ASAP7_75t_R _44069_ (.CLK(net679),
    .D(_00254_),
    .QN(_00667_));
 DFFLQNx1_ASAP7_75t_R _44070_ (.CLK(net678),
    .D(_00255_),
    .QN(_00666_));
 DFFLQNx3_ASAP7_75t_R _44071_ (.CLK(net677),
    .D(_00256_),
    .QN(_00665_));
 DFFLQNx3_ASAP7_75t_R _44072_ (.CLK(net676),
    .D(_00153_),
    .QN(_00664_));
 DFFLQNx3_ASAP7_75t_R _44073_ (.CLK(net675),
    .D(_00154_),
    .QN(_00663_));
 DFFLQNx3_ASAP7_75t_R _44074_ (.CLK(net674),
    .D(_00155_),
    .QN(_00662_));
 DFFLQNx3_ASAP7_75t_R _44075_ (.CLK(net673),
    .D(_00156_),
    .QN(_00661_));
 DFFLQNx3_ASAP7_75t_R _44076_ (.CLK(net672),
    .D(_00157_),
    .QN(_00660_));
 DFFLQNx1_ASAP7_75t_R _44077_ (.CLK(net671),
    .D(_00158_),
    .QN(_00659_));
 DFFLQNx3_ASAP7_75t_R _44078_ (.CLK(net670),
    .D(_00159_),
    .QN(_00658_));
 DFFLQNx2_ASAP7_75t_R _44079_ (.QN(_00657_),
    .CLK(net669),
    .D(_00160_));
 DFFLQNx3_ASAP7_75t_R _44080_ (.CLK(net668),
    .D(_00001_),
    .QN(_00656_));
 DFFLQNx3_ASAP7_75t_R _44081_ (.CLK(net667),
    .D(_00002_),
    .QN(_00655_));
 DFFLQNx2_ASAP7_75t_R _44082_ (.QN(_00654_),
    .CLK(net666),
    .D(_00003_));
 DFFLQNx2_ASAP7_75t_R _44083_ (.QN(_00653_),
    .CLK(net665),
    .D(_00004_));
 DFFLQNx2_ASAP7_75t_R _44084_ (.QN(_00652_),
    .CLK(net664),
    .D(_00005_));
 DFFLQNx2_ASAP7_75t_R _44085_ (.QN(_00651_),
    .CLK(net663),
    .D(_00006_));
 DFFLQNx2_ASAP7_75t_R _44086_ (.QN(_00650_),
    .CLK(net662),
    .D(_00007_));
 DFFLQNx2_ASAP7_75t_R _44087_ (.QN(_00649_),
    .CLK(net661),
    .D(_00008_));
 DFFLQNx3_ASAP7_75t_R _44088_ (.CLK(net660),
    .D(_00033_),
    .QN(_00648_));
 DFFLQNx3_ASAP7_75t_R _44089_ (.CLK(net659),
    .D(_00034_),
    .QN(_00647_));
 DFFLQNx2_ASAP7_75t_R _44090_ (.QN(_00646_),
    .CLK(net658),
    .D(_00035_));
 DFFLQNx2_ASAP7_75t_R _44091_ (.QN(_00645_),
    .CLK(net657),
    .D(_00036_));
 DFFLQNx2_ASAP7_75t_R _44092_ (.QN(_00644_),
    .CLK(net656),
    .D(_00037_));
 DFFLQNx2_ASAP7_75t_R _44093_ (.QN(_00643_),
    .CLK(net655),
    .D(_00038_));
 DFFLQNx2_ASAP7_75t_R _44094_ (.QN(_00642_),
    .CLK(net654),
    .D(_00039_));
 DFFLQNx2_ASAP7_75t_R _44095_ (.QN(_00641_),
    .CLK(net653),
    .D(_00040_));
 DFFLQNx3_ASAP7_75t_R _44096_ (.CLK(net652),
    .D(_00065_),
    .QN(_00640_));
 DFFLQNx3_ASAP7_75t_R _44097_ (.CLK(net651),
    .D(_00066_),
    .QN(_00639_));
 DFFLQNx2_ASAP7_75t_R _44098_ (.QN(_00638_),
    .CLK(net650),
    .D(_00067_));
 DFFLQNx2_ASAP7_75t_R _44099_ (.QN(_00637_),
    .CLK(net649),
    .D(_00068_));
 DFFLQNx2_ASAP7_75t_R _44100_ (.QN(_00636_),
    .CLK(net648),
    .D(_00069_));
 DFFLQNx2_ASAP7_75t_R _44101_ (.QN(_00635_),
    .CLK(net647),
    .D(_00070_));
 DFFLQNx2_ASAP7_75t_R _44102_ (.QN(_00634_),
    .CLK(net646),
    .D(_00071_));
 DFFLQNx2_ASAP7_75t_R _44103_ (.QN(_00633_),
    .CLK(net645),
    .D(_00072_));
 DFFLQNx3_ASAP7_75t_R _44104_ (.CLK(net644),
    .D(_00097_),
    .QN(_00632_));
 DFFLQNx3_ASAP7_75t_R _44105_ (.CLK(net643),
    .D(_00098_),
    .QN(_00631_));
 DFFLQNx2_ASAP7_75t_R _44106_ (.QN(_00630_),
    .CLK(net642),
    .D(_00099_));
 DFFLQNx3_ASAP7_75t_R _44107_ (.CLK(net641),
    .D(_00100_),
    .QN(_00629_));
 DFFLQNx2_ASAP7_75t_R _44108_ (.QN(_00628_),
    .CLK(net640),
    .D(_00101_));
 DFFLQNx2_ASAP7_75t_R _44109_ (.QN(_00627_),
    .CLK(net639),
    .D(_00102_));
 DFFLQNx2_ASAP7_75t_R _44110_ (.QN(_00626_),
    .CLK(net638),
    .D(_00103_));
 DFFLQNx2_ASAP7_75t_R _44111_ (.QN(_00625_),
    .CLK(net637),
    .D(_00104_));
 DFFLQNx3_ASAP7_75t_R _44112_ (.CLK(net636),
    .D(_00009_),
    .QN(_00624_));
 DFFLQNx3_ASAP7_75t_R _44113_ (.CLK(net635),
    .D(_00010_),
    .QN(_00623_));
 DFFLQNx2_ASAP7_75t_R _44114_ (.QN(_00622_),
    .CLK(net634),
    .D(_00011_));
 DFFLQNx2_ASAP7_75t_R _44115_ (.QN(_00621_),
    .CLK(net633),
    .D(_00012_));
 DFFLQNx2_ASAP7_75t_R _44116_ (.QN(_00620_),
    .CLK(net632),
    .D(_00013_));
 DFFLQNx2_ASAP7_75t_R _44117_ (.QN(_00619_),
    .CLK(net631),
    .D(_00014_));
 DFFLQNx2_ASAP7_75t_R _44118_ (.QN(_00618_),
    .CLK(net630),
    .D(_00015_));
 DFFLQNx2_ASAP7_75t_R _44119_ (.QN(_00617_),
    .CLK(net629),
    .D(_00016_));
 DFFLQNx3_ASAP7_75t_R _44120_ (.CLK(net628),
    .D(_00041_),
    .QN(_00616_));
 DFFLQNx3_ASAP7_75t_R _44121_ (.CLK(net627),
    .D(_00042_),
    .QN(_00615_));
 DFFLQNx2_ASAP7_75t_R _44122_ (.QN(_00614_),
    .CLK(net626),
    .D(_00043_));
 DFFLQNx2_ASAP7_75t_R _44123_ (.QN(_00613_),
    .CLK(net625),
    .D(_00044_));
 DFFLQNx2_ASAP7_75t_R _44124_ (.QN(_00612_),
    .CLK(net624),
    .D(_00045_));
 DFFLQNx2_ASAP7_75t_R _44125_ (.QN(_00611_),
    .CLK(net623),
    .D(_00046_));
 DFFLQNx2_ASAP7_75t_R _44126_ (.QN(_00610_),
    .CLK(net622),
    .D(_00047_));
 DFFLQNx2_ASAP7_75t_R _44127_ (.QN(_00609_),
    .CLK(net621),
    .D(_00048_));
 DFFLQNx3_ASAP7_75t_R _44128_ (.CLK(net620),
    .D(_00073_),
    .QN(_00608_));
 DFFLQNx3_ASAP7_75t_R _44129_ (.CLK(net619),
    .D(_00074_),
    .QN(_00607_));
 DFFLQNx2_ASAP7_75t_R _44130_ (.QN(_00606_),
    .CLK(net618),
    .D(_00075_));
 DFFLQNx2_ASAP7_75t_R _44131_ (.QN(_00605_),
    .CLK(net617),
    .D(_00076_));
 DFFLQNx2_ASAP7_75t_R _44132_ (.QN(_00604_),
    .CLK(net616),
    .D(_00077_));
 DFFLQNx2_ASAP7_75t_R _44133_ (.QN(_00603_),
    .CLK(net615),
    .D(_00078_));
 DFFLQNx2_ASAP7_75t_R _44134_ (.QN(_00602_),
    .CLK(net614),
    .D(_00079_));
 DFFLQNx2_ASAP7_75t_R _44135_ (.QN(_00601_),
    .CLK(net613),
    .D(_00080_));
 DFFLQNx3_ASAP7_75t_R _44136_ (.CLK(net612),
    .D(_00105_),
    .QN(_00600_));
 DFFLQNx3_ASAP7_75t_R _44137_ (.CLK(net611),
    .D(_00106_),
    .QN(_00599_));
 DFFLQNx2_ASAP7_75t_R _44138_ (.QN(_00598_),
    .CLK(net610),
    .D(_00107_));
 DFFLQNx2_ASAP7_75t_R _44139_ (.QN(_00597_),
    .CLK(net609),
    .D(_00108_));
 DFFLQNx2_ASAP7_75t_R _44140_ (.QN(_00596_),
    .CLK(net608),
    .D(_00109_));
 DFFLQNx2_ASAP7_75t_R _44141_ (.QN(_00595_),
    .CLK(net607),
    .D(_00110_));
 DFFLQNx2_ASAP7_75t_R _44142_ (.QN(_00594_),
    .CLK(net606),
    .D(_00111_));
 DFFLQNx2_ASAP7_75t_R _44143_ (.QN(_00593_),
    .CLK(net605),
    .D(_00112_));
 DFFLQNx3_ASAP7_75t_R _44144_ (.CLK(net604),
    .D(_00017_),
    .QN(_00592_));
 DFFLQNx3_ASAP7_75t_R _44145_ (.CLK(net603),
    .D(_00018_),
    .QN(_00591_));
 DFFLQNx2_ASAP7_75t_R _44146_ (.QN(_00590_),
    .CLK(net602),
    .D(_00019_));
 DFFLQNx2_ASAP7_75t_R _44147_ (.QN(_00589_),
    .CLK(net601),
    .D(_00020_));
 DFFLQNx2_ASAP7_75t_R _44148_ (.QN(_00588_),
    .CLK(net600),
    .D(_00021_));
 DFFLQNx2_ASAP7_75t_R _44149_ (.QN(_00587_),
    .CLK(net599),
    .D(_00022_));
 DFFLQNx2_ASAP7_75t_R _44150_ (.QN(_00586_),
    .CLK(net598),
    .D(_00023_));
 DFFLQNx2_ASAP7_75t_R _44151_ (.QN(_00585_),
    .CLK(net597),
    .D(_00024_));
 DFFLQNx3_ASAP7_75t_R _44152_ (.CLK(net596),
    .D(_00049_),
    .QN(_00584_));
 DFFLQNx3_ASAP7_75t_R _44153_ (.CLK(net595),
    .D(_00050_),
    .QN(_00583_));
 DFFLQNx2_ASAP7_75t_R _44154_ (.QN(_00582_),
    .CLK(net594),
    .D(_00051_));
 DFFLQNx2_ASAP7_75t_R _44155_ (.QN(_00581_),
    .CLK(net593),
    .D(_00052_));
 DFFLQNx2_ASAP7_75t_R _44156_ (.QN(_00580_),
    .CLK(net592),
    .D(_00053_));
 DFFLQNx2_ASAP7_75t_R _44157_ (.QN(_00579_),
    .CLK(net591),
    .D(_00054_));
 DFFLQNx2_ASAP7_75t_R _44158_ (.QN(_00578_),
    .CLK(net590),
    .D(_00055_));
 DFFLQNx2_ASAP7_75t_R _44159_ (.QN(_00577_),
    .CLK(net589),
    .D(_00056_));
 DFFLQNx3_ASAP7_75t_R _44160_ (.CLK(net588),
    .D(_00081_),
    .QN(_00576_));
 DFFLQNx3_ASAP7_75t_R _44161_ (.CLK(net587),
    .D(_00082_),
    .QN(_00575_));
 DFFLQNx2_ASAP7_75t_R _44162_ (.QN(_00574_),
    .CLK(net586),
    .D(_00083_));
 DFFLQNx2_ASAP7_75t_R _44163_ (.QN(_00573_),
    .CLK(net585),
    .D(_00084_));
 DFFLQNx2_ASAP7_75t_R _44164_ (.QN(_00572_),
    .CLK(net584),
    .D(_00085_));
 DFFLQNx2_ASAP7_75t_R _44165_ (.QN(_00571_),
    .CLK(net583),
    .D(_00086_));
 DFFLQNx2_ASAP7_75t_R _44166_ (.QN(_00570_),
    .CLK(net582),
    .D(_00087_));
 DFFLQNx2_ASAP7_75t_R _44167_ (.QN(_00569_),
    .CLK(net581),
    .D(_00088_));
 DFFLQNx3_ASAP7_75t_R _44168_ (.CLK(net580),
    .D(_00113_),
    .QN(_00568_));
 DFFLQNx3_ASAP7_75t_R _44169_ (.CLK(net579),
    .D(_00114_),
    .QN(_00567_));
 DFFLQNx2_ASAP7_75t_R _44170_ (.QN(_00566_),
    .CLK(net578),
    .D(_00115_));
 DFFLQNx2_ASAP7_75t_R _44171_ (.QN(_00565_),
    .CLK(net577),
    .D(_00116_));
 DFFLQNx2_ASAP7_75t_R _44172_ (.QN(_00564_),
    .CLK(net576),
    .D(_00117_));
 DFFLQNx2_ASAP7_75t_R _44173_ (.QN(_00563_),
    .CLK(net575),
    .D(_00118_));
 DFFLQNx2_ASAP7_75t_R _44174_ (.QN(_00562_),
    .CLK(net574),
    .D(_00119_));
 DFFLQNx2_ASAP7_75t_R _44175_ (.QN(_00561_),
    .CLK(net573),
    .D(_00120_));
 DFFLQNx3_ASAP7_75t_R _44176_ (.CLK(net572),
    .D(_00025_),
    .QN(_00560_));
 DFFLQNx3_ASAP7_75t_R _44177_ (.CLK(net571),
    .D(_00026_),
    .QN(_00559_));
 DFFLQNx2_ASAP7_75t_R _44178_ (.QN(_00558_),
    .CLK(net570),
    .D(_00027_));
 DFFLQNx2_ASAP7_75t_R _44179_ (.QN(_00557_),
    .CLK(net569),
    .D(_00028_));
 DFFLQNx2_ASAP7_75t_R _44180_ (.QN(_00556_),
    .CLK(net568),
    .D(_00029_));
 DFFLQNx2_ASAP7_75t_R _44181_ (.QN(_00555_),
    .CLK(net567),
    .D(_00030_));
 DFFLQNx2_ASAP7_75t_R _44182_ (.QN(_00554_),
    .CLK(net566),
    .D(_00031_));
 DFFLQNx2_ASAP7_75t_R _44183_ (.QN(_00553_),
    .CLK(net565),
    .D(_00032_));
 DFFLQNx3_ASAP7_75t_R _44184_ (.CLK(net564),
    .D(_00057_),
    .QN(_00552_));
 DFFLQNx3_ASAP7_75t_R _44185_ (.CLK(net563),
    .D(_00058_),
    .QN(_00551_));
 DFFLQNx2_ASAP7_75t_R _44186_ (.QN(_00550_),
    .CLK(net562),
    .D(_00059_));
 DFFLQNx2_ASAP7_75t_R _44187_ (.QN(_00549_),
    .CLK(net561),
    .D(_00060_));
 DFFLQNx2_ASAP7_75t_R _44188_ (.QN(_00548_),
    .CLK(net560),
    .D(_00061_));
 DFFLQNx2_ASAP7_75t_R _44189_ (.QN(_00547_),
    .CLK(net559),
    .D(_00062_));
 DFFLQNx2_ASAP7_75t_R _44190_ (.QN(_00546_),
    .CLK(net558),
    .D(_00063_));
 DFFLQNx2_ASAP7_75t_R _44191_ (.QN(_00545_),
    .CLK(net557),
    .D(_00064_));
 DFFLQNx3_ASAP7_75t_R _44192_ (.CLK(net556),
    .D(_00089_),
    .QN(_00544_));
 DFFLQNx3_ASAP7_75t_R _44193_ (.CLK(net555),
    .D(_00090_),
    .QN(_00543_));
 DFFLQNx2_ASAP7_75t_R _44194_ (.QN(_00542_),
    .CLK(net554),
    .D(_00091_));
 DFFLQNx2_ASAP7_75t_R _44195_ (.QN(_00541_),
    .CLK(net553),
    .D(_00092_));
 DFFLQNx2_ASAP7_75t_R _44196_ (.QN(_00540_),
    .CLK(net552),
    .D(_00093_));
 DFFLQNx2_ASAP7_75t_R _44197_ (.QN(_00539_),
    .CLK(net551),
    .D(_00094_));
 DFFLQNx2_ASAP7_75t_R _44198_ (.QN(_00538_),
    .CLK(net550),
    .D(_00095_));
 DFFLQNx2_ASAP7_75t_R _44199_ (.QN(_00537_),
    .CLK(net549),
    .D(_00096_));
 DFFLQNx3_ASAP7_75t_R _44200_ (.CLK(net548),
    .D(_00121_),
    .QN(_00536_));
 DFFLQNx3_ASAP7_75t_R _44201_ (.CLK(net547),
    .D(_00122_),
    .QN(_00535_));
 DFFLQNx2_ASAP7_75t_R _44202_ (.QN(_00534_),
    .CLK(net546),
    .D(_00123_));
 DFFLQNx2_ASAP7_75t_R _44203_ (.QN(_00533_),
    .CLK(net545),
    .D(_00124_));
 DFFLQNx2_ASAP7_75t_R _44204_ (.QN(_00532_),
    .CLK(net544),
    .D(_00125_));
 DFFLQNx2_ASAP7_75t_R _44205_ (.QN(_00531_),
    .CLK(net543),
    .D(_00126_));
 DFFLQNx2_ASAP7_75t_R _44206_ (.QN(_00530_),
    .CLK(net542),
    .D(_00127_));
 DFFLQNx2_ASAP7_75t_R _44207_ (.QN(_00529_),
    .CLK(net541),
    .D(_00128_));
 DFFLQNx2_ASAP7_75t_R _44208_ (.QN(_00528_),
    .CLK(net540),
    .D(net405));
 DFFLQNx3_ASAP7_75t_R _44209_ (.CLK(net539),
    .D(_00000_),
    .QN(_00527_));
 DFFLQNx2_ASAP7_75t_R _44210_ (.QN(_22106_),
    .CLK(net538),
    .D(_01061_));
 DFFLQNx2_ASAP7_75t_R _44211_ (.QN(\u0.r0.rcnt_next[0] ),
    .CLK(net537),
    .D(_01062_));
 DFFLQNx2_ASAP7_75t_R _44212_ (.QN(_22101_),
    .CLK(net536),
    .D(_01063_));
 DFFLQNx3_ASAP7_75t_R _44213_ (.CLK(net535),
    .D(_01064_),
    .QN(_00526_));
 DFFLQNx1_ASAP7_75t_R _44214_ (.CLK(net534),
    .D(_01065_),
    .QN(_00525_));
 DFFLQNx2_ASAP7_75t_R _44215_ (.QN(_00409_),
    .CLK(net533),
    .D(_00257_));
 DFFLQNx2_ASAP7_75t_R _44216_ (.QN(_00410_),
    .CLK(net532),
    .D(_00268_));
 DFFLQNx2_ASAP7_75t_R _44217_ (.QN(_00524_),
    .CLK(net531),
    .D(_00279_));
 DFFLQNx2_ASAP7_75t_R _44218_ (.QN(_00523_),
    .CLK(net530),
    .D(_00282_));
 DFFLQNx2_ASAP7_75t_R _44219_ (.QN(_00522_),
    .CLK(net529),
    .D(_00283_));
 DFFLQNx2_ASAP7_75t_R _44220_ (.QN(_00521_),
    .CLK(net528),
    .D(_00284_));
 DFFLQNx2_ASAP7_75t_R _44221_ (.QN(_00411_),
    .CLK(net527),
    .D(_00285_));
 DFFLQNx2_ASAP7_75t_R _44222_ (.QN(_00520_),
    .CLK(net526),
    .D(_00286_));
 DFFLQNx2_ASAP7_75t_R _44223_ (.QN(_00412_),
    .CLK(net525),
    .D(_00287_));
 DFFLQNx2_ASAP7_75t_R _44224_ (.QN(_00519_),
    .CLK(net524),
    .D(_00288_));
 DFFLQNx2_ASAP7_75t_R _44225_ (.QN(_00518_),
    .CLK(net523),
    .D(_00258_));
 DFFLQNx2_ASAP7_75t_R _44226_ (.QN(_00517_),
    .CLK(net522),
    .D(_00259_));
 DFFLQNx2_ASAP7_75t_R _44227_ (.QN(_00516_),
    .CLK(net521),
    .D(_00260_));
 DFFLQNx2_ASAP7_75t_R _44228_ (.QN(_00515_),
    .CLK(net520),
    .D(_00261_));
 DFFLQNx2_ASAP7_75t_R _44229_ (.QN(_00514_),
    .CLK(net519),
    .D(_00262_));
 DFFLQNx2_ASAP7_75t_R _44230_ (.QN(_00513_),
    .CLK(net518),
    .D(_00263_));
 DFFLQNx2_ASAP7_75t_R _44231_ (.QN(_00413_),
    .CLK(net517),
    .D(_00264_));
 DFFLQNx2_ASAP7_75t_R _44232_ (.QN(_00414_),
    .CLK(net516),
    .D(_00265_));
 DFFLQNx2_ASAP7_75t_R _44233_ (.QN(_00512_),
    .CLK(net515),
    .D(_00266_));
 DFFLQNx2_ASAP7_75t_R _44234_ (.QN(_00511_),
    .CLK(net514),
    .D(_00267_));
 DFFLQNx2_ASAP7_75t_R _44235_ (.QN(_00510_),
    .CLK(net513),
    .D(_00269_));
 DFFLQNx2_ASAP7_75t_R _44236_ (.QN(_00415_),
    .CLK(net512),
    .D(_00270_));
 DFFLQNx2_ASAP7_75t_R _44237_ (.QN(_00416_),
    .CLK(net511),
    .D(_00271_));
 DFFLQNx2_ASAP7_75t_R _44238_ (.QN(_00509_),
    .CLK(net510),
    .D(_00272_));
 DFFLQNx2_ASAP7_75t_R _44239_ (.QN(_00508_),
    .CLK(net509),
    .D(_00273_));
 DFFLQNx2_ASAP7_75t_R _44240_ (.QN(_00507_),
    .CLK(net508),
    .D(_00274_));
 DFFLQNx2_ASAP7_75t_R _44241_ (.QN(_00506_),
    .CLK(net507),
    .D(_00275_));
 DFFLQNx2_ASAP7_75t_R _44242_ (.QN(_00505_),
    .CLK(net506),
    .D(_00276_));
 DFFLQNx2_ASAP7_75t_R _44243_ (.QN(_00504_),
    .CLK(net505),
    .D(_00277_));
 DFFLQNx2_ASAP7_75t_R _44244_ (.QN(_00503_),
    .CLK(net504),
    .D(_00278_));
 DFFLQNx2_ASAP7_75t_R _44245_ (.QN(_00502_),
    .CLK(net503),
    .D(_00280_));
 DFFLQNx2_ASAP7_75t_R _44246_ (.QN(_00501_),
    .CLK(net502),
    .D(_00281_));
 DFFLQNx2_ASAP7_75t_R _44247_ (.QN(_00500_),
    .CLK(net501),
    .D(_00289_));
 DFFLQNx2_ASAP7_75t_R _44248_ (.QN(_00499_),
    .CLK(net500),
    .D(_00300_));
 DFFLQNx2_ASAP7_75t_R _44249_ (.QN(_00385_),
    .CLK(net499),
    .D(_00311_));
 DFFLQNx2_ASAP7_75t_R _44250_ (.QN(_00386_),
    .CLK(net498),
    .D(_00314_));
 DFFLQNx2_ASAP7_75t_R _44251_ (.QN(_00387_),
    .CLK(net497),
    .D(_00315_));
 DFFLQNx2_ASAP7_75t_R _44252_ (.QN(_00498_),
    .CLK(net496),
    .D(_00316_));
 DFFLQNx2_ASAP7_75t_R _44253_ (.QN(_00497_),
    .CLK(net495),
    .D(_00317_));
 DFFLQNx2_ASAP7_75t_R _44254_ (.QN(_00388_),
    .CLK(net494),
    .D(_00318_));
 DFFLQNx2_ASAP7_75t_R _44255_ (.QN(_00496_),
    .CLK(net493),
    .D(_00319_));
 DFFLQNx2_ASAP7_75t_R _44256_ (.QN(_00495_),
    .CLK(net492),
    .D(_00320_));
 DFFLQNx2_ASAP7_75t_R _44257_ (.QN(_00389_),
    .CLK(net491),
    .D(_00290_));
 DFFLQNx2_ASAP7_75t_R _44258_ (.QN(_00390_),
    .CLK(net490),
    .D(_00291_));
 DFFLQNx2_ASAP7_75t_R _44259_ (.QN(_00391_),
    .CLK(net489),
    .D(_00292_));
 DFFLQNx2_ASAP7_75t_R _44260_ (.QN(_00494_),
    .CLK(net488),
    .D(_00293_));
 DFFLQNx2_ASAP7_75t_R _44261_ (.QN(_00493_),
    .CLK(net487),
    .D(_00294_));
 DFFLQNx2_ASAP7_75t_R _44262_ (.QN(_00392_),
    .CLK(net486),
    .D(_00295_));
 DFFLQNx2_ASAP7_75t_R _44263_ (.QN(_00492_),
    .CLK(net485),
    .D(_00296_));
 DFFLQNx2_ASAP7_75t_R _44264_ (.QN(_00491_),
    .CLK(net484),
    .D(_00297_));
 DFFLQNx2_ASAP7_75t_R _44265_ (.QN(_00393_),
    .CLK(net483),
    .D(_00298_));
 DFFLQNx2_ASAP7_75t_R _44266_ (.QN(_00394_),
    .CLK(net482),
    .D(_00299_));
 DFFLQNx2_ASAP7_75t_R _44267_ (.QN(_00395_),
    .CLK(net481),
    .D(_00301_));
 DFFLQNx2_ASAP7_75t_R _44268_ (.QN(_00490_),
    .CLK(net480),
    .D(_00302_));
 DFFLQNx2_ASAP7_75t_R _44269_ (.QN(_00489_),
    .CLK(net479),
    .D(_00303_));
 DFFLQNx2_ASAP7_75t_R _44270_ (.QN(_00396_),
    .CLK(net478),
    .D(_00304_));
 DFFLQNx2_ASAP7_75t_R _44271_ (.QN(_00398_),
    .CLK(net477),
    .D(_00305_));
 DFFLQNx2_ASAP7_75t_R _44272_ (.QN(_00400_),
    .CLK(net476),
    .D(_00306_));
 DFFLQNx2_ASAP7_75t_R _44273_ (.QN(_00488_),
    .CLK(net475),
    .D(_00307_));
 DFFLQNx2_ASAP7_75t_R _44274_ (.QN(_00487_),
    .CLK(net474),
    .D(_00308_));
 DFFLQNx2_ASAP7_75t_R _44275_ (.QN(_00486_),
    .CLK(net473),
    .D(_00309_));
 DFFLQNx2_ASAP7_75t_R _44276_ (.QN(_00405_),
    .CLK(net472),
    .D(_00310_));
 DFFLQNx2_ASAP7_75t_R _44277_ (.QN(_00407_),
    .CLK(net471),
    .D(_00312_));
 DFFLQNx2_ASAP7_75t_R _44278_ (.QN(_00485_),
    .CLK(net470),
    .D(_00313_));
 DFFLQNx2_ASAP7_75t_R _44279_ (.QN(_00484_),
    .CLK(net469),
    .D(_00321_));
 DFFLQNx2_ASAP7_75t_R _44280_ (.QN(_00483_),
    .CLK(net468),
    .D(_00332_));
 DFFLQNx2_ASAP7_75t_R _44281_ (.QN(_00482_),
    .CLK(net467),
    .D(_00343_));
 DFFLQNx2_ASAP7_75t_R _44282_ (.QN(_00481_),
    .CLK(net466),
    .D(_00346_));
 DFFLQNx2_ASAP7_75t_R _44283_ (.QN(_00480_),
    .CLK(net465),
    .D(_00347_));
 DFFLQNx2_ASAP7_75t_R _44284_ (.QN(_00479_),
    .CLK(net464),
    .D(_00348_));
 DFFLQNx2_ASAP7_75t_R _44285_ (.QN(_00478_),
    .CLK(net463),
    .D(_00349_));
 DFFLQNx2_ASAP7_75t_R _44286_ (.QN(_00477_),
    .CLK(net462),
    .D(_00350_));
 DFFLQNx2_ASAP7_75t_R _44287_ (.QN(_00476_),
    .CLK(net461),
    .D(_00351_));
 DFFLQNx2_ASAP7_75t_R _44288_ (.QN(_00475_),
    .CLK(net460),
    .D(_00352_));
 DFFLQNx2_ASAP7_75t_R _44289_ (.QN(_00474_),
    .CLK(net459),
    .D(_00322_));
 DFFLQNx2_ASAP7_75t_R _44290_ (.QN(_00473_),
    .CLK(net458),
    .D(_00323_));
 DFFLQNx2_ASAP7_75t_R _44291_ (.QN(_00472_),
    .CLK(net457),
    .D(_00324_));
 DFFLQNx2_ASAP7_75t_R _44292_ (.QN(_00471_),
    .CLK(net456),
    .D(_00325_));
 DFFLQNx2_ASAP7_75t_R _44293_ (.QN(_00470_),
    .CLK(net455),
    .D(_00326_));
 DFFLQNx2_ASAP7_75t_R _44294_ (.QN(_00469_),
    .CLK(net454),
    .D(_00327_));
 DFFLQNx2_ASAP7_75t_R _44295_ (.QN(_00468_),
    .CLK(net453),
    .D(_00328_));
 DFFLQNx2_ASAP7_75t_R _44296_ (.QN(_00467_),
    .CLK(net452),
    .D(_00329_));
 DFFLQNx2_ASAP7_75t_R _44297_ (.QN(_00466_),
    .CLK(net451),
    .D(_00330_));
 DFFLQNx2_ASAP7_75t_R _44298_ (.QN(_00465_),
    .CLK(net450),
    .D(net3941));
 DFFLQNx2_ASAP7_75t_R _44299_ (.QN(_00464_),
    .CLK(net449),
    .D(_00333_));
 DFFLQNx2_ASAP7_75t_R _44300_ (.QN(_00463_),
    .CLK(net448),
    .D(_00334_));
 DFFLQNx2_ASAP7_75t_R _44301_ (.QN(_00462_),
    .CLK(net447),
    .D(_00335_));
 DFFLQNx2_ASAP7_75t_R _44302_ (.QN(_00461_),
    .CLK(net446),
    .D(_00336_));
 DFFLQNx2_ASAP7_75t_R _44303_ (.QN(_00460_),
    .CLK(net445),
    .D(_00337_));
 DFFLQNx2_ASAP7_75t_R _44304_ (.QN(_00459_),
    .CLK(net444),
    .D(_00338_));
 DFFLQNx2_ASAP7_75t_R _44305_ (.QN(_00458_),
    .CLK(net443),
    .D(_00339_));
 DFFLQNx2_ASAP7_75t_R _44306_ (.QN(_00457_),
    .CLK(net442),
    .D(_00340_));
 DFFLQNx2_ASAP7_75t_R _44307_ (.QN(_00456_),
    .CLK(net441),
    .D(_00341_));
 DFFLQNx2_ASAP7_75t_R _44308_ (.QN(_00455_),
    .CLK(net440),
    .D(_00342_));
 DFFLQNx2_ASAP7_75t_R _44309_ (.QN(_00454_),
    .CLK(net439),
    .D(_00344_));
 DFFLQNx2_ASAP7_75t_R _44310_ (.QN(_00453_),
    .CLK(net438),
    .D(_00345_));
 DFFLQNx3_ASAP7_75t_R _44311_ (.CLK(net437),
    .D(_00353_),
    .QN(_00452_));
 DFFLQNx3_ASAP7_75t_R _44312_ (.CLK(net436),
    .D(_00364_),
    .QN(_00451_));
 DFFLQNx3_ASAP7_75t_R _44313_ (.CLK(net435),
    .D(_00375_),
    .QN(_00450_));
 DFFLQNx2_ASAP7_75t_R _44314_ (.QN(_00449_),
    .CLK(net434),
    .D(_00378_));
 DFFLQNx2_ASAP7_75t_R _44315_ (.QN(_00448_),
    .CLK(net433),
    .D(_00379_));
 DFFLQNx2_ASAP7_75t_R _44316_ (.QN(_00447_),
    .CLK(net432),
    .D(_00380_));
 DFFLQNx2_ASAP7_75t_R _44317_ (.QN(_00446_),
    .CLK(net431),
    .D(_00381_));
 DFFLQNx2_ASAP7_75t_R _44318_ (.QN(_00445_),
    .CLK(net430),
    .D(_00382_));
 DFFLQNx3_ASAP7_75t_R _44319_ (.CLK(net429),
    .D(_00383_),
    .QN(_00444_));
 DFFLQNx3_ASAP7_75t_R _44320_ (.CLK(net428),
    .D(_00384_),
    .QN(_00443_));
 DFFLQNx2_ASAP7_75t_R _44321_ (.QN(_00442_),
    .CLK(net427),
    .D(_00354_));
 DFFLQNx2_ASAP7_75t_R _44322_ (.QN(_00441_),
    .CLK(net426),
    .D(_00355_));
 DFFLQNx2_ASAP7_75t_R _44323_ (.QN(_00440_),
    .CLK(net425),
    .D(_00356_));
 DFFLQNx2_ASAP7_75t_R _44324_ (.QN(_00439_),
    .CLK(net424),
    .D(_00357_));
 DFFLQNx2_ASAP7_75t_R _44325_ (.QN(_00438_),
    .CLK(net423),
    .D(_00358_));
 DFFLQNx2_ASAP7_75t_R _44326_ (.QN(_00437_),
    .CLK(net422),
    .D(_00359_));
 DFFLQNx3_ASAP7_75t_R _44327_ (.CLK(net421),
    .D(_00360_),
    .QN(_00436_));
 DFFLQNx3_ASAP7_75t_R _44328_ (.CLK(net420),
    .D(_00361_),
    .QN(_00435_));
 DFFLQNx3_ASAP7_75t_R _44329_ (.CLK(net419),
    .D(_00362_),
    .QN(_00434_));
 DFFLQNx3_ASAP7_75t_R _44330_ (.CLK(net418),
    .D(_00363_),
    .QN(_00433_));
 DFFLQNx2_ASAP7_75t_R _44331_ (.QN(_00432_),
    .CLK(net417),
    .D(_00365_));
 DFFLQNx2_ASAP7_75t_R _44332_ (.QN(_00431_),
    .CLK(net416),
    .D(_00366_));
 DFFLQNx3_ASAP7_75t_R _44333_ (.CLK(net415),
    .D(_00367_),
    .QN(_00430_));
 DFFLQNx3_ASAP7_75t_R _44334_ (.CLK(net414),
    .D(_00368_),
    .QN(_00429_));
 DFFLQNx3_ASAP7_75t_R _44335_ (.CLK(net413),
    .D(_00369_),
    .QN(_00428_));
 DFFLQNx3_ASAP7_75t_R _44336_ (.CLK(net412),
    .D(_00370_),
    .QN(_00427_));
 DFFLQNx2_ASAP7_75t_R _44337_ (.QN(_00426_),
    .CLK(net411),
    .D(net3865));
 DFFLQNx2_ASAP7_75t_R _44338_ (.QN(_00425_),
    .CLK(net410),
    .D(_00372_));
 DFFLQNx2_ASAP7_75t_R _44339_ (.QN(_00424_),
    .CLK(net409),
    .D(_00373_));
 DFFLQNx2_ASAP7_75t_R _44340_ (.QN(_00423_),
    .CLK(net408),
    .D(_00374_));
 DFFLQNx2_ASAP7_75t_R _44341_ (.QN(_00422_),
    .CLK(net407),
    .D(_00376_));
 DFFLQNx3_ASAP7_75t_R _44342_ (.CLK(net406),
    .D(_00377_),
    .QN(_00421_));
 INVx1_ASAP7_75t_R _98_129 (.A(clknet_leaf_7_clk),
    .Y(net534));
 INVx1_ASAP7_75t_R _98_130 (.A(clknet_leaf_7_clk),
    .Y(net535));
 INVx1_ASAP7_75t_R _98_131 (.A(clknet_leaf_7_clk),
    .Y(net536));
 INVx1_ASAP7_75t_R _98_132 (.A(clknet_leaf_7_clk),
    .Y(net537));
 INVx1_ASAP7_75t_R _98_133 (.A(clknet_leaf_4_clk),
    .Y(net538));
 INVx1_ASAP7_75t_R _98_134 (.A(clknet_leaf_4_clk),
    .Y(net539));
 INVx1_ASAP7_75t_R _98_135 (.A(clknet_leaf_2_clk),
    .Y(net540));
 INVx1_ASAP7_75t_R _98_136 (.A(clknet_leaf_17_clk),
    .Y(net541));
 INVx1_ASAP7_75t_R _98_137 (.A(clknet_leaf_17_clk),
    .Y(net542));
 INVx1_ASAP7_75t_R _98_138 (.A(clknet_leaf_0_clk),
    .Y(net543));
 INVx1_ASAP7_75t_R _98_139 (.A(clknet_leaf_17_clk),
    .Y(net544));
 INVx1_ASAP7_75t_R _98_140 (.A(clknet_leaf_1_clk),
    .Y(net545));
 INVx1_ASAP7_75t_R _98_141 (.A(clknet_leaf_17_clk),
    .Y(net546));
 INVx1_ASAP7_75t_R _98_142 (.A(clknet_leaf_17_clk),
    .Y(net547));
 INVx1_ASAP7_75t_R _98_143 (.A(clknet_leaf_17_clk),
    .Y(net548));
 INVx1_ASAP7_75t_R _98_144 (.A(clknet_leaf_4_clk),
    .Y(net549));
 INVx1_ASAP7_75t_R _98_145 (.A(clknet_leaf_4_clk),
    .Y(net550));
 INVx1_ASAP7_75t_R _98_146 (.A(clknet_leaf_3_clk),
    .Y(net551));
 INVx1_ASAP7_75t_R _98_147 (.A(clknet_leaf_3_clk),
    .Y(net552));
 INVx1_ASAP7_75t_R _148 (.A(clknet_leaf_4_clk),
    .Y(net553));
 INVx1_ASAP7_75t_R _148_149 (.A(clknet_leaf_2_clk),
    .Y(net554));
 INVx1_ASAP7_75t_R _148_150 (.A(clknet_leaf_2_clk),
    .Y(net555));
 INVx1_ASAP7_75t_R _148_151 (.A(clknet_leaf_4_clk),
    .Y(net556));
 INVx1_ASAP7_75t_R _148_152 (.A(clknet_leaf_2_clk),
    .Y(net557));
 INVx1_ASAP7_75t_R _148_153 (.A(clknet_leaf_2_clk),
    .Y(net558));
 INVx1_ASAP7_75t_R _148_154 (.A(clknet_leaf_2_clk),
    .Y(net559));
 INVx1_ASAP7_75t_R _148_155 (.A(clknet_leaf_3_clk),
    .Y(net560));
 INVx1_ASAP7_75t_R _148_156 (.A(clknet_leaf_3_clk),
    .Y(net561));
 INVx1_ASAP7_75t_R _148_157 (.A(clknet_leaf_7_clk),
    .Y(net562));
 INVx1_ASAP7_75t_R _148_158 (.A(clknet_leaf_7_clk),
    .Y(net563));
 INVx1_ASAP7_75t_R _148_159 (.A(clknet_leaf_2_clk),
    .Y(net564));
 INVx1_ASAP7_75t_R _148_160 (.A(clknet_leaf_1_clk),
    .Y(net565));
 INVx1_ASAP7_75t_R _148_161 (.A(clknet_leaf_0_clk),
    .Y(net566));
 INVx1_ASAP7_75t_R _148_162 (.A(clknet_leaf_1_clk),
    .Y(net567));
 INVx1_ASAP7_75t_R _148_163 (.A(clknet_leaf_1_clk),
    .Y(net568));
 INVx1_ASAP7_75t_R _148_164 (.A(clknet_leaf_0_clk),
    .Y(net569));
 INVx1_ASAP7_75t_R _148_165 (.A(clknet_leaf_0_clk),
    .Y(net570));
 INVx1_ASAP7_75t_R _148_166 (.A(clknet_leaf_0_clk),
    .Y(net571));
 INVx1_ASAP7_75t_R _148_167 (.A(clknet_leaf_0_clk),
    .Y(net572));
 INVx1_ASAP7_75t_R _148_168 (.A(clknet_leaf_11_clk),
    .Y(net573));
 INVx1_ASAP7_75t_R _148_169 (.A(clknet_leaf_12_clk),
    .Y(net574));
 INVx1_ASAP7_75t_R _148_170 (.A(clknet_leaf_11_clk),
    .Y(net575));
 INVx1_ASAP7_75t_R _148_171 (.A(clknet_leaf_12_clk),
    .Y(net576));
 INVx1_ASAP7_75t_R _148_172 (.A(clknet_leaf_7_clk),
    .Y(net577));
 INVx1_ASAP7_75t_R _148_173 (.A(clknet_leaf_15_clk),
    .Y(net578));
 INVx1_ASAP7_75t_R _148_174 (.A(clknet_leaf_15_clk),
    .Y(net579));
 INVx1_ASAP7_75t_R _148_175 (.A(clknet_leaf_15_clk),
    .Y(net580));
 INVx1_ASAP7_75t_R _148_176 (.A(clknet_leaf_12_clk),
    .Y(net581));
 INVx1_ASAP7_75t_R _148_177 (.A(clknet_leaf_15_clk),
    .Y(net582));
 INVx1_ASAP7_75t_R _148_178 (.A(clknet_leaf_12_clk),
    .Y(net583));
 INVx1_ASAP7_75t_R _148_179 (.A(clknet_leaf_11_clk),
    .Y(net584));
 INVx1_ASAP7_75t_R _148_180 (.A(clknet_leaf_10_clk),
    .Y(net585));
 INVx1_ASAP7_75t_R _148_181 (.A(clknet_leaf_12_clk),
    .Y(net586));
 INVx1_ASAP7_75t_R _148_182 (.A(clknet_leaf_12_clk),
    .Y(net587));
 INVx1_ASAP7_75t_R _148_183 (.A(clknet_leaf_13_clk),
    .Y(net588));
 INVx1_ASAP7_75t_R _148_184 (.A(clknet_leaf_9_clk),
    .Y(net589));
 INVx1_ASAP7_75t_R _148_185 (.A(clknet_leaf_8_clk),
    .Y(net590));
 INVx1_ASAP7_75t_R _148_186 (.A(clknet_leaf_9_clk),
    .Y(net591));
 INVx1_ASAP7_75t_R _148_187 (.A(clknet_leaf_8_clk),
    .Y(net592));
 INVx1_ASAP7_75t_R _148_188 (.A(clknet_leaf_9_clk),
    .Y(net593));
 INVx1_ASAP7_75t_R _148_189 (.A(clknet_leaf_9_clk),
    .Y(net594));
 INVx1_ASAP7_75t_R _148_190 (.A(clknet_leaf_9_clk),
    .Y(net595));
 INVx1_ASAP7_75t_R _148_191 (.A(clknet_leaf_9_clk),
    .Y(net596));
 INVx1_ASAP7_75t_R _148_192 (.A(clknet_leaf_12_clk),
    .Y(net597));
 INVx1_ASAP7_75t_R _148_193 (.A(clknet_leaf_11_clk),
    .Y(net598));
 INVx1_ASAP7_75t_R _148_194 (.A(clknet_leaf_11_clk),
    .Y(net599));
 INVx1_ASAP7_75t_R _148_195 (.A(clknet_leaf_10_clk),
    .Y(net600));
 INVx1_ASAP7_75t_R _148_196 (.A(clknet_leaf_10_clk),
    .Y(net601));
 INVx1_ASAP7_75t_R _148_197 (.A(clknet_leaf_10_clk),
    .Y(net602));
 INVx1_ASAP7_75t_R _198 (.A(clknet_leaf_10_clk),
    .Y(net603));
 INVx1_ASAP7_75t_R _198_199 (.A(clknet_leaf_12_clk),
    .Y(net604));
 INVx1_ASAP7_75t_R _198_200 (.A(clknet_leaf_7_clk),
    .Y(net605));
 INVx1_ASAP7_75t_R _198_201 (.A(clknet_leaf_11_clk),
    .Y(net606));
 INVx1_ASAP7_75t_R _198_202 (.A(clknet_leaf_6_clk),
    .Y(net607));
 INVx1_ASAP7_75t_R _198_203 (.A(clknet_leaf_6_clk),
    .Y(net608));
 INVx1_ASAP7_75t_R _198_204 (.A(clknet_leaf_6_clk),
    .Y(net609));
 INVx1_ASAP7_75t_R _198_205 (.A(clknet_leaf_9_clk),
    .Y(net610));
 INVx1_ASAP7_75t_R _198_206 (.A(clknet_leaf_9_clk),
    .Y(net611));
 INVx1_ASAP7_75t_R _198_207 (.A(clknet_leaf_9_clk),
    .Y(net612));
 INVx1_ASAP7_75t_R _198_208 (.A(clknet_leaf_6_clk),
    .Y(net613));
 INVx1_ASAP7_75t_R _198_209 (.A(clknet_leaf_7_clk),
    .Y(net614));
 INVx1_ASAP7_75t_R _198_210 (.A(clknet_leaf_6_clk),
    .Y(net615));
 INVx1_ASAP7_75t_R _198_211 (.A(clknet_leaf_4_clk),
    .Y(net616));
 INVx1_ASAP7_75t_R _198_212 (.A(clknet_leaf_4_clk),
    .Y(net617));
 INVx1_ASAP7_75t_R _198_213 (.A(clknet_leaf_4_clk),
    .Y(net618));
 INVx1_ASAP7_75t_R _198_214 (.A(clknet_leaf_4_clk),
    .Y(net619));
 INVx1_ASAP7_75t_R _198_215 (.A(clknet_leaf_4_clk),
    .Y(net620));
 INVx1_ASAP7_75t_R _198_216 (.A(clknet_leaf_7_clk),
    .Y(net621));
 INVx1_ASAP7_75t_R _198_217 (.A(clknet_leaf_6_clk),
    .Y(net622));
 INVx1_ASAP7_75t_R _198_218 (.A(clknet_leaf_1_clk),
    .Y(net623));
 INVx1_ASAP7_75t_R _198_219 (.A(clknet_leaf_6_clk),
    .Y(net624));
 INVx1_ASAP7_75t_R _198_220 (.A(clknet_leaf_2_clk),
    .Y(net625));
 INVx1_ASAP7_75t_R _198_221 (.A(clknet_leaf_1_clk),
    .Y(net626));
 INVx1_ASAP7_75t_R _198_222 (.A(clknet_leaf_15_clk),
    .Y(net627));
 INVx1_ASAP7_75t_R _198_223 (.A(clknet_leaf_15_clk),
    .Y(net628));
 INVx1_ASAP7_75t_R _198_224 (.A(clknet_leaf_8_clk),
    .Y(net629));
 INVx1_ASAP7_75t_R _198_225 (.A(clknet_leaf_8_clk),
    .Y(net630));
 INVx1_ASAP7_75t_R _198_226 (.A(clknet_leaf_8_clk),
    .Y(net631));
 INVx1_ASAP7_75t_R _198_227 (.A(clknet_leaf_8_clk),
    .Y(net632));
 INVx1_ASAP7_75t_R _198_228 (.A(clknet_leaf_9_clk),
    .Y(net633));
 INVx1_ASAP7_75t_R _198_229 (.A(clknet_leaf_9_clk),
    .Y(net634));
 INVx1_ASAP7_75t_R _198_230 (.A(clknet_leaf_9_clk),
    .Y(net635));
 INVx1_ASAP7_75t_R _198_231 (.A(clknet_leaf_8_clk),
    .Y(net636));
 INVx1_ASAP7_75t_R _198_232 (.A(clknet_leaf_15_clk),
    .Y(net637));
 INVx1_ASAP7_75t_R _198_233 (.A(clknet_leaf_16_clk),
    .Y(net638));
 INVx1_ASAP7_75t_R _198_234 (.A(clknet_leaf_15_clk),
    .Y(net639));
 INVx1_ASAP7_75t_R _198_235 (.A(clknet_leaf_15_clk),
    .Y(net640));
 INVx1_ASAP7_75t_R _198_236 (.A(clknet_leaf_16_clk),
    .Y(net641));
 INVx1_ASAP7_75t_R _198_237 (.A(clknet_leaf_7_clk),
    .Y(net642));
 INVx1_ASAP7_75t_R _198_238 (.A(clknet_leaf_7_clk),
    .Y(net643));
 INVx1_ASAP7_75t_R _198_239 (.A(clknet_leaf_7_clk),
    .Y(net644));
 INVx1_ASAP7_75t_R _198_240 (.A(clknet_leaf_14_clk),
    .Y(net645));
 INVx1_ASAP7_75t_R _198_241 (.A(clknet_leaf_15_clk),
    .Y(net646));
 INVx1_ASAP7_75t_R _198_242 (.A(clknet_leaf_16_clk),
    .Y(net647));
 INVx1_ASAP7_75t_R _198_243 (.A(clknet_leaf_16_clk),
    .Y(net648));
 INVx1_ASAP7_75t_R _198_244 (.A(clknet_leaf_15_clk),
    .Y(net649));
 INVx1_ASAP7_75t_R _198_245 (.A(clknet_leaf_14_clk),
    .Y(net650));
 INVx1_ASAP7_75t_R _198_246 (.A(clknet_leaf_14_clk),
    .Y(net651));
 INVx1_ASAP7_75t_R _198_247 (.A(clknet_leaf_14_clk),
    .Y(net652));
 INVx1_ASAP7_75t_R _248 (.A(clknet_leaf_15_clk),
    .Y(net653));
 INVx1_ASAP7_75t_R _248_249 (.A(clknet_leaf_17_clk),
    .Y(net654));
 INVx1_ASAP7_75t_R _248_250 (.A(clknet_leaf_16_clk),
    .Y(net655));
 INVx1_ASAP7_75t_R _248_251 (.A(clknet_leaf_15_clk),
    .Y(net656));
 INVx1_ASAP7_75t_R _248_252 (.A(clknet_leaf_16_clk),
    .Y(net657));
 INVx1_ASAP7_75t_R _248_253 (.A(clknet_leaf_17_clk),
    .Y(net658));
 INVx1_ASAP7_75t_R _248_254 (.A(clknet_leaf_17_clk),
    .Y(net659));
 INVx1_ASAP7_75t_R _248_255 (.A(clknet_leaf_17_clk),
    .Y(net660));
 INVx1_ASAP7_75t_R _248_256 (.A(clknet_leaf_13_clk),
    .Y(net661));
 INVx1_ASAP7_75t_R _248_257 (.A(clknet_leaf_14_clk),
    .Y(net662));
 INVx1_ASAP7_75t_R _248_258 (.A(clknet_leaf_13_clk),
    .Y(net663));
 INVx1_ASAP7_75t_R _248_259 (.A(clknet_leaf_14_clk),
    .Y(net664));
 INVx1_ASAP7_75t_R _248_260 (.A(clknet_leaf_14_clk),
    .Y(net665));
 INVx1_ASAP7_75t_R _248_261 (.A(clknet_leaf_13_clk),
    .Y(net666));
 INVx1_ASAP7_75t_R _248_262 (.A(clknet_leaf_13_clk),
    .Y(net667));
 INVx1_ASAP7_75t_R _248_263 (.A(clknet_leaf_14_clk),
    .Y(net668));
 INVx1_ASAP7_75t_R _248_264 (.A(clknet_leaf_13_clk),
    .Y(net669));
 INVx1_ASAP7_75t_R _248_265 (.A(clknet_leaf_13_clk),
    .Y(net670));
 INVx1_ASAP7_75t_R _248_266 (.A(clknet_leaf_14_clk),
    .Y(net671));
 INVx1_ASAP7_75t_R _248_267 (.A(clknet_leaf_13_clk),
    .Y(net672));
 INVx1_ASAP7_75t_R _248_268 (.A(clknet_leaf_14_clk),
    .Y(net673));
 INVx1_ASAP7_75t_R _248_269 (.A(clknet_leaf_13_clk),
    .Y(net674));
 INVx1_ASAP7_75t_R _248_270 (.A(clknet_leaf_13_clk),
    .Y(net675));
 INVx1_ASAP7_75t_R _248_271 (.A(clknet_leaf_14_clk),
    .Y(net676));
 INVx1_ASAP7_75t_R _248_272 (.A(clknet_leaf_9_clk),
    .Y(net677));
 INVx1_ASAP7_75t_R _248_273 (.A(clknet_leaf_9_clk),
    .Y(net678));
 INVx1_ASAP7_75t_R _248_274 (.A(clknet_leaf_5_clk),
    .Y(net679));
 INVx1_ASAP7_75t_R _248_275 (.A(clknet_leaf_8_clk),
    .Y(net680));
 INVx1_ASAP7_75t_R _248_276 (.A(clknet_leaf_5_clk),
    .Y(net681));
 INVx1_ASAP7_75t_R _248_277 (.A(clknet_leaf_9_clk),
    .Y(net682));
 INVx1_ASAP7_75t_R _248_278 (.A(clknet_leaf_9_clk),
    .Y(net683));
 INVx1_ASAP7_75t_R _248_279 (.A(clknet_leaf_8_clk),
    .Y(net684));
 INVx1_ASAP7_75t_R _248_280 (.A(clknet_leaf_10_clk),
    .Y(net685));
 INVx1_ASAP7_75t_R _248_281 (.A(clknet_leaf_12_clk),
    .Y(net686));
 INVx1_ASAP7_75t_R _248_282 (.A(clknet_leaf_11_clk),
    .Y(net687));
 INVx1_ASAP7_75t_R _248_283 (.A(clknet_leaf_10_clk),
    .Y(net688));
 INVx1_ASAP7_75t_R _248_284 (.A(clknet_leaf_10_clk),
    .Y(net689));
 INVx1_ASAP7_75t_R _248_285 (.A(clknet_leaf_10_clk),
    .Y(net690));
 INVx1_ASAP7_75t_R _248_286 (.A(clknet_leaf_10_clk),
    .Y(net691));
 INVx1_ASAP7_75t_R _248_287 (.A(clknet_leaf_12_clk),
    .Y(net692));
 INVx1_ASAP7_75t_R _248_288 (.A(clknet_leaf_0_clk),
    .Y(net693));
 INVx1_ASAP7_75t_R _248_289 (.A(clknet_leaf_0_clk),
    .Y(net694));
 INVx1_ASAP7_75t_R _248_290 (.A(clknet_leaf_0_clk),
    .Y(net695));
 INVx1_ASAP7_75t_R _248_291 (.A(clknet_leaf_0_clk),
    .Y(net696));
 INVx1_ASAP7_75t_R _248_292 (.A(clknet_leaf_0_clk),
    .Y(net697));
 INVx1_ASAP7_75t_R _248_293 (.A(clknet_leaf_17_clk),
    .Y(net698));
 INVx1_ASAP7_75t_R _248_294 (.A(clknet_leaf_0_clk),
    .Y(net699));
 INVx1_ASAP7_75t_R _248_295 (.A(clknet_leaf_0_clk),
    .Y(net700));
 INVx1_ASAP7_75t_R _248_296 (.A(clknet_leaf_14_clk),
    .Y(net701));
 INVx1_ASAP7_75t_R _248_297 (.A(clknet_leaf_16_clk),
    .Y(net702));
 INVx1_ASAP7_75t_R _298 (.A(clknet_leaf_16_clk),
    .Y(net703));
 INVx1_ASAP7_75t_R _298_299 (.A(clknet_leaf_16_clk),
    .Y(net704));
 INVx1_ASAP7_75t_R _298_300 (.A(clknet_leaf_16_clk),
    .Y(net705));
 INVx1_ASAP7_75t_R _298_301 (.A(clknet_leaf_16_clk),
    .Y(net706));
 INVx1_ASAP7_75t_R _298_302 (.A(clknet_leaf_13_clk),
    .Y(net707));
 INVx1_ASAP7_75t_R _298_303 (.A(clknet_leaf_13_clk),
    .Y(net708));
 INVx1_ASAP7_75t_R _298_304 (.A(clknet_leaf_5_clk),
    .Y(net709));
 INVx1_ASAP7_75t_R _298_305 (.A(clknet_leaf_5_clk),
    .Y(net710));
 INVx1_ASAP7_75t_R _298_306 (.A(clknet_leaf_4_clk),
    .Y(net711));
 INVx1_ASAP7_75t_R _298_307 (.A(clknet_leaf_5_clk),
    .Y(net712));
 INVx1_ASAP7_75t_R _298_308 (.A(clknet_leaf_5_clk),
    .Y(net713));
 INVx1_ASAP7_75t_R _298_309 (.A(clknet_leaf_5_clk),
    .Y(net714));
 INVx1_ASAP7_75t_R _298_310 (.A(clknet_leaf_9_clk),
    .Y(net715));
 INVx1_ASAP7_75t_R _298_311 (.A(clknet_leaf_8_clk),
    .Y(net716));
 INVx1_ASAP7_75t_R _298_312 (.A(clknet_leaf_9_clk),
    .Y(net717));
 INVx1_ASAP7_75t_R _298_313 (.A(clknet_leaf_10_clk),
    .Y(net718));
 INVx1_ASAP7_75t_R _298_314 (.A(clknet_leaf_9_clk),
    .Y(net719));
 INVx1_ASAP7_75t_R _298_315 (.A(clknet_leaf_8_clk),
    .Y(net720));
 INVx1_ASAP7_75t_R _298_316 (.A(clknet_leaf_9_clk),
    .Y(net721));
 INVx1_ASAP7_75t_R _298_317 (.A(clknet_leaf_10_clk),
    .Y(net722));
 INVx1_ASAP7_75t_R _298_318 (.A(clknet_leaf_11_clk),
    .Y(net723));
 INVx1_ASAP7_75t_R _298_319 (.A(clknet_leaf_10_clk),
    .Y(net724));
 INVx1_ASAP7_75t_R _298_320 (.A(clknet_leaf_2_clk),
    .Y(net725));
 INVx1_ASAP7_75t_R _298_321 (.A(clknet_leaf_2_clk),
    .Y(net726));
 INVx1_ASAP7_75t_R _298_322 (.A(clknet_leaf_3_clk),
    .Y(net727));
 INVx1_ASAP7_75t_R _298_323 (.A(clknet_leaf_3_clk),
    .Y(net728));
 INVx1_ASAP7_75t_R _298_324 (.A(clknet_leaf_3_clk),
    .Y(net729));
 INVx1_ASAP7_75t_R _298_325 (.A(clknet_leaf_2_clk),
    .Y(net730));
 INVx1_ASAP7_75t_R _298_326 (.A(clknet_leaf_2_clk),
    .Y(net731));
 INVx1_ASAP7_75t_R _298_327 (.A(clknet_leaf_3_clk),
    .Y(net732));
 INVx1_ASAP7_75t_R _298_328 (.A(clknet_leaf_14_clk),
    .Y(net733));
 INVx1_ASAP7_75t_R _298_329 (.A(clknet_leaf_16_clk),
    .Y(net734));
 INVx1_ASAP7_75t_R _298_330 (.A(clknet_leaf_16_clk),
    .Y(net735));
 INVx1_ASAP7_75t_R _298_331 (.A(clknet_leaf_16_clk),
    .Y(net736));
 INVx1_ASAP7_75t_R _298_332 (.A(clknet_leaf_15_clk),
    .Y(net737));
 INVx1_ASAP7_75t_R _298_333 (.A(clknet_leaf_16_clk),
    .Y(net738));
 INVx1_ASAP7_75t_R _298_334 (.A(clknet_leaf_13_clk),
    .Y(net739));
 INVx1_ASAP7_75t_R _298_335 (.A(clknet_leaf_13_clk),
    .Y(net740));
 INVx1_ASAP7_75t_R _298_336 (.A(clknet_leaf_9_clk),
    .Y(net741));
 INVx1_ASAP7_75t_R _298_337 (.A(clknet_leaf_5_clk),
    .Y(net742));
 INVx1_ASAP7_75t_R _298_338 (.A(clknet_leaf_5_clk),
    .Y(net743));
 INVx1_ASAP7_75t_R _298_339 (.A(clknet_leaf_4_clk),
    .Y(net744));
 INVx1_ASAP7_75t_R _298_340 (.A(clknet_leaf_3_clk),
    .Y(net745));
 INVx1_ASAP7_75t_R _298_341 (.A(clknet_leaf_4_clk),
    .Y(net746));
 INVx1_ASAP7_75t_R _298_342 (.A(clknet_leaf_5_clk),
    .Y(net747));
 INVx1_ASAP7_75t_R _298_343 (.A(clknet_leaf_8_clk),
    .Y(net748));
 INVx1_ASAP7_75t_R _298_344 (.A(clknet_leaf_11_clk),
    .Y(net749));
 INVx1_ASAP7_75t_R _298_345 (.A(clknet_leaf_11_clk),
    .Y(net750));
 INVx1_ASAP7_75t_R _298_346 (.A(clknet_leaf_10_clk),
    .Y(net751));
 INVx1_ASAP7_75t_R _298_347 (.A(clknet_leaf_10_clk),
    .Y(net752));
 INVx1_ASAP7_75t_R _348 (.A(clknet_leaf_10_clk),
    .Y(net753));
 INVx1_ASAP7_75t_R _348_349 (.A(clknet_leaf_12_clk),
    .Y(net754));
 INVx1_ASAP7_75t_R _348_350 (.A(clknet_leaf_11_clk),
    .Y(net755));
 INVx1_ASAP7_75t_R _348_351 (.A(clknet_leaf_10_clk),
    .Y(net756));
 INVx1_ASAP7_75t_R _348_352 (.A(clknet_leaf_3_clk),
    .Y(net757));
 INVx1_ASAP7_75t_R _348_353 (.A(clknet_leaf_3_clk),
    .Y(net758));
 INVx1_ASAP7_75t_R _348_354 (.A(clknet_leaf_3_clk),
    .Y(net759));
 INVx1_ASAP7_75t_R _348_355 (.A(clknet_leaf_3_clk),
    .Y(net760));
 INVx1_ASAP7_75t_R _348_356 (.A(clknet_leaf_3_clk),
    .Y(net761));
 INVx1_ASAP7_75t_R _348_357 (.A(clknet_leaf_2_clk),
    .Y(net762));
 INVx1_ASAP7_75t_R _348_358 (.A(clknet_leaf_2_clk),
    .Y(net763));
 INVx1_ASAP7_75t_R _348_359 (.A(clknet_leaf_3_clk),
    .Y(net764));
 INVx1_ASAP7_75t_R _348_360 (.A(clknet_leaf_16_clk),
    .Y(net765));
 INVx1_ASAP7_75t_R _348_361 (.A(clknet_leaf_16_clk),
    .Y(net766));
 INVx1_ASAP7_75t_R _348_362 (.A(clknet_leaf_17_clk),
    .Y(net767));
 INVx1_ASAP7_75t_R _348_363 (.A(clknet_leaf_16_clk),
    .Y(net768));
 INVx1_ASAP7_75t_R _348_364 (.A(clknet_leaf_16_clk),
    .Y(net769));
 INVx1_ASAP7_75t_R _348_365 (.A(clknet_leaf_13_clk),
    .Y(net770));
 INVx1_ASAP7_75t_R _348_366 (.A(clknet_leaf_13_clk),
    .Y(net771));
 INVx1_ASAP7_75t_R _348_367 (.A(clknet_leaf_13_clk),
    .Y(net772));
 INVx1_ASAP7_75t_R _348_368 (.A(clknet_leaf_5_clk),
    .Y(net773));
 INVx1_ASAP7_75t_R _348_369 (.A(clknet_leaf_5_clk),
    .Y(net774));
 INVx1_ASAP7_75t_R _348_370 (.A(clknet_leaf_5_clk),
    .Y(net775));
 INVx1_ASAP7_75t_R _348_371 (.A(clknet_leaf_6_clk),
    .Y(net776));
 INVx1_ASAP7_75t_R _348_372 (.A(clknet_leaf_5_clk),
    .Y(net777));
 INVx1_ASAP7_75t_R _348_373 (.A(clknet_leaf_9_clk),
    .Y(net778));
 INVx1_ASAP7_75t_R _348_374 (.A(clknet_leaf_9_clk),
    .Y(net779));
 INVx1_ASAP7_75t_R _348_375 (.A(clknet_leaf_8_clk),
    .Y(net780));
 INVx1_ASAP7_75t_R _348_376 (.A(clknet_leaf_12_clk),
    .Y(net781));
 INVx1_ASAP7_75t_R _348_377 (.A(clknet_leaf_12_clk),
    .Y(net782));
 INVx1_ASAP7_75t_R _348_378 (.A(clknet_leaf_12_clk),
    .Y(net783));
 INVx1_ASAP7_75t_R _348_379 (.A(clknet_leaf_12_clk),
    .Y(net784));
 INVx1_ASAP7_75t_R _348_380 (.A(clknet_leaf_10_clk),
    .Y(net785));
 INVx1_ASAP7_75t_R _348_381 (.A(clknet_leaf_12_clk),
    .Y(net786));
 INVx1_ASAP7_75t_R _348_382 (.A(clknet_leaf_12_clk),
    .Y(net787));
 INVx1_ASAP7_75t_R _348_383 (.A(clknet_leaf_12_clk),
    .Y(net788));
 INVx1_ASAP7_75t_R _348_384 (.A(clknet_leaf_0_clk),
    .Y(net789));
 INVx1_ASAP7_75t_R _348_385 (.A(clknet_leaf_2_clk),
    .Y(net790));
 INVx1_ASAP7_75t_R _348_386 (.A(clknet_leaf_0_clk),
    .Y(net791));
 INVx1_ASAP7_75t_R _348_387 (.A(clknet_leaf_0_clk),
    .Y(net792));
 INVx1_ASAP7_75t_R _348_388 (.A(clknet_leaf_0_clk),
    .Y(net793));
 INVx1_ASAP7_75t_R _348_389 (.A(clknet_leaf_15_clk),
    .Y(net794));
 INVx1_ASAP7_75t_R _348_390 (.A(clknet_leaf_17_clk),
    .Y(net795));
 INVx1_ASAP7_75t_R _348_391 (.A(clknet_leaf_1_clk),
    .Y(net796));
 INVx1_ASAP7_75t_R _348_392 (.A(clknet_leaf_4_clk),
    .Y(net797));
 INVx1_ASAP7_75t_R _348_393 (.A(clknet_leaf_4_clk),
    .Y(net798));
 INVx1_ASAP7_75t_R _348_394 (.A(clknet_leaf_4_clk),
    .Y(net799));
 INVx1_ASAP7_75t_R _348_395 (.A(clknet_leaf_13_clk),
    .Y(net800));
 INVx1_ASAP7_75t_R _348_396 (.A(clknet_leaf_13_clk),
    .Y(net801));
 INVx1_ASAP7_75t_R _348_397 (.A(clknet_leaf_14_clk),
    .Y(net802));
 INVx1_ASAP7_75t_R _398 (.A(clknet_leaf_14_clk),
    .Y(net803));
 INVx1_ASAP7_75t_R _398_399 (.A(clknet_leaf_14_clk),
    .Y(net804));
 INVx1_ASAP7_75t_R _398_400 (.A(clknet_leaf_13_clk),
    .Y(net805));
 INVx1_ASAP7_75t_R _398_401 (.A(clknet_leaf_13_clk),
    .Y(net806));
 INVx1_ASAP7_75t_R _398_402 (.A(clknet_leaf_13_clk),
    .Y(net807));
 INVx1_ASAP7_75t_R _398_403 (.A(clknet_leaf_1_clk),
    .Y(net808));
 INVx1_ASAP7_75t_R _398_404 (.A(clknet_leaf_17_clk),
    .Y(net809));
 INVx1_ASAP7_75t_R _398_405 (.A(clknet_leaf_17_clk),
    .Y(net810));
 INVx1_ASAP7_75t_R _398_406 (.A(clknet_leaf_0_clk),
    .Y(net811));
 INVx1_ASAP7_75t_R _398_407 (.A(clknet_leaf_16_clk),
    .Y(net812));
 INVx1_ASAP7_75t_R _398_408 (.A(clknet_leaf_16_clk),
    .Y(net813));
 INVx1_ASAP7_75t_R _398_409 (.A(clknet_leaf_14_clk),
    .Y(net814));
 INVx1_ASAP7_75t_R _398_410 (.A(clknet_leaf_14_clk),
    .Y(net815));
 INVx1_ASAP7_75t_R _398_411 (.A(clknet_leaf_14_clk),
    .Y(net816));
 INVx1_ASAP7_75t_R _398_412 (.A(clknet_leaf_1_clk),
    .Y(net817));
 INVx1_ASAP7_75t_R _398_413 (.A(clknet_leaf_16_clk),
    .Y(net818));
 INVx1_ASAP7_75t_R _398_414 (.A(clknet_leaf_16_clk),
    .Y(net819));
 INVx1_ASAP7_75t_R _398_415 (.A(clknet_leaf_4_clk),
    .Y(net820));
 INVx1_ASAP7_75t_R _398_416 (.A(clknet_leaf_16_clk),
    .Y(net821));
 INVx1_ASAP7_75t_R _398_417 (.A(clknet_leaf_13_clk),
    .Y(net822));
 INVx1_ASAP7_75t_R _398_418 (.A(clknet_leaf_13_clk),
    .Y(net823));
 INVx1_ASAP7_75t_R _398_419 (.A(clknet_leaf_1_clk),
    .Y(net824));
 INVx1_ASAP7_75t_R _398_420 (.A(clknet_leaf_16_clk),
    .Y(net825));
 INVx1_ASAP7_75t_R _398_421 (.A(clknet_leaf_17_clk),
    .Y(net826));
 INVx1_ASAP7_75t_R _398_422 (.A(clknet_leaf_17_clk),
    .Y(net827));
 INVx1_ASAP7_75t_R _398_423 (.A(clknet_leaf_16_clk),
    .Y(net828));
 INVx1_ASAP7_75t_R _398_424 (.A(clknet_leaf_16_clk),
    .Y(net829));
 INVx1_ASAP7_75t_R _398_425 (.A(clknet_leaf_13_clk),
    .Y(net830));
 INVx1_ASAP7_75t_R _398_426 (.A(clknet_leaf_13_clk),
    .Y(net831));
 INVx1_ASAP7_75t_R _398_427 (.A(clknet_leaf_9_clk),
    .Y(net832));
 INVx1_ASAP7_75t_R _398_428 (.A(clknet_leaf_5_clk),
    .Y(net833));
 INVx1_ASAP7_75t_R _398_429 (.A(clknet_leaf_4_clk),
    .Y(net834));
 INVx1_ASAP7_75t_R _398_430 (.A(clknet_leaf_8_clk),
    .Y(net835));
 INVx1_ASAP7_75t_R _398_431 (.A(clknet_leaf_5_clk),
    .Y(net836));
 INVx1_ASAP7_75t_R _398_432 (.A(clknet_leaf_8_clk),
    .Y(net837));
 INVx1_ASAP7_75t_R _398_433 (.A(clknet_leaf_9_clk),
    .Y(net838));
 INVx1_ASAP7_75t_R _398_434 (.A(clknet_leaf_8_clk),
    .Y(net839));
 INVx1_ASAP7_75t_R _398_435 (.A(clknet_leaf_5_clk),
    .Y(net840));
 INVx1_ASAP7_75t_R _398_436 (.A(clknet_leaf_5_clk),
    .Y(net841));
 INVx1_ASAP7_75t_R _398_437 (.A(clknet_leaf_5_clk),
    .Y(net842));
 INVx1_ASAP7_75t_R _398_438 (.A(clknet_leaf_4_clk),
    .Y(net843));
 INVx1_ASAP7_75t_R _398_439 (.A(clknet_leaf_4_clk),
    .Y(net844));
 INVx1_ASAP7_75t_R _398_440 (.A(clknet_leaf_5_clk),
    .Y(net845));
 INVx1_ASAP7_75t_R _398_441 (.A(clknet_leaf_8_clk),
    .Y(net846));
 INVx1_ASAP7_75t_R _398_442 (.A(clknet_leaf_8_clk),
    .Y(net847));
 INVx1_ASAP7_75t_R _398_443 (.A(clknet_leaf_6_clk),
    .Y(net848));
 INVx1_ASAP7_75t_R _398_444 (.A(clknet_leaf_5_clk),
    .Y(net849));
 INVx1_ASAP7_75t_R _398_445 (.A(clknet_leaf_4_clk),
    .Y(net850));
 INVx1_ASAP7_75t_R _398_446 (.A(clknet_leaf_3_clk),
    .Y(net851));
 INVx1_ASAP7_75t_R _398_447 (.A(clknet_leaf_3_clk),
    .Y(net852));
 INVx1_ASAP7_75t_R _448 (.A(clknet_leaf_5_clk),
    .Y(net853));
 INVx1_ASAP7_75t_R _448_449 (.A(clknet_leaf_5_clk),
    .Y(net854));
 INVx1_ASAP7_75t_R _448_450 (.A(clknet_leaf_8_clk),
    .Y(net855));
 INVx1_ASAP7_75t_R _448_451 (.A(clknet_leaf_5_clk),
    .Y(net856));
 INVx1_ASAP7_75t_R _448_452 (.A(clknet_leaf_6_clk),
    .Y(net857));
 INVx1_ASAP7_75t_R _448_453 (.A(clknet_leaf_5_clk),
    .Y(net858));
 INVx1_ASAP7_75t_R _448_454 (.A(clknet_leaf_5_clk),
    .Y(net859));
 INVx1_ASAP7_75t_R _448_455 (.A(clknet_leaf_5_clk),
    .Y(net860));
 INVx1_ASAP7_75t_R _448_456 (.A(clknet_leaf_8_clk),
    .Y(net861));
 INVx1_ASAP7_75t_R _448_457 (.A(clknet_leaf_9_clk),
    .Y(net862));
 INVx1_ASAP7_75t_R _448_458 (.A(clknet_leaf_9_clk),
    .Y(net863));
 INVx1_ASAP7_75t_R _448_459 (.A(clknet_leaf_10_clk),
    .Y(net864));
 INVx1_ASAP7_75t_R _448_460 (.A(clknet_leaf_12_clk),
    .Y(net865));
 INVx1_ASAP7_75t_R _448_461 (.A(clknet_leaf_11_clk),
    .Y(net866));
 INVx1_ASAP7_75t_R _448_462 (.A(clknet_leaf_10_clk),
    .Y(net867));
 INVx1_ASAP7_75t_R _448_463 (.A(clknet_leaf_10_clk),
    .Y(net868));
 INVx1_ASAP7_75t_R _448_464 (.A(clknet_leaf_10_clk),
    .Y(net869));
 INVx1_ASAP7_75t_R _448_465 (.A(clknet_leaf_12_clk),
    .Y(net870));
 INVx1_ASAP7_75t_R _448_466 (.A(clknet_leaf_12_clk),
    .Y(net871));
 INVx1_ASAP7_75t_R _448_467 (.A(clknet_leaf_9_clk),
    .Y(net872));
 INVx1_ASAP7_75t_R _448_468 (.A(clknet_leaf_10_clk),
    .Y(net873));
 INVx1_ASAP7_75t_R _448_469 (.A(clknet_leaf_9_clk),
    .Y(net874));
 INVx1_ASAP7_75t_R _448_470 (.A(clknet_leaf_8_clk),
    .Y(net875));
 INVx1_ASAP7_75t_R _448_471 (.A(clknet_leaf_9_clk),
    .Y(net876));
 INVx1_ASAP7_75t_R _448_472 (.A(clknet_leaf_10_clk),
    .Y(net877));
 INVx1_ASAP7_75t_R _448_473 (.A(clknet_leaf_10_clk),
    .Y(net878));
 INVx1_ASAP7_75t_R _448_474 (.A(clknet_leaf_10_clk),
    .Y(net879));
 INVx1_ASAP7_75t_R _448_475 (.A(clknet_leaf_14_clk),
    .Y(net880));
 INVx1_ASAP7_75t_R _448_476 (.A(clknet_leaf_13_clk),
    .Y(net881));
 INVx1_ASAP7_75t_R _448_477 (.A(clknet_leaf_10_clk),
    .Y(net882));
 INVx1_ASAP7_75t_R _448_478 (.A(clknet_leaf_10_clk),
    .Y(net883));
 INVx1_ASAP7_75t_R _448_479 (.A(clknet_leaf_10_clk),
    .Y(net884));
 INVx1_ASAP7_75t_R _448_480 (.A(clknet_leaf_12_clk),
    .Y(net885));
 INVx1_ASAP7_75t_R _448_481 (.A(clknet_leaf_12_clk),
    .Y(net886));
 INVx1_ASAP7_75t_R _448_482 (.A(clknet_leaf_12_clk),
    .Y(net887));
 INVx1_ASAP7_75t_R _448_483 (.A(clknet_leaf_12_clk),
    .Y(net888));
 INVx1_ASAP7_75t_R _448_484 (.A(clknet_leaf_12_clk),
    .Y(net889));
 INVx1_ASAP7_75t_R _448_485 (.A(clknet_leaf_15_clk),
    .Y(net890));
 INVx1_ASAP7_75t_R _448_486 (.A(clknet_leaf_14_clk),
    .Y(net891));
 INVx1_ASAP7_75t_R _448_487 (.A(clknet_leaf_10_clk),
    .Y(net892));
 INVx1_ASAP7_75t_R _448_488 (.A(clknet_leaf_12_clk),
    .Y(net893));
 INVx1_ASAP7_75t_R _448_489 (.A(clknet_leaf_12_clk),
    .Y(net894));
 INVx1_ASAP7_75t_R _448_490 (.A(clknet_leaf_12_clk),
    .Y(net895));
 INVx1_ASAP7_75t_R _448_491 (.A(clknet_leaf_0_clk),
    .Y(net896));
 INVx1_ASAP7_75t_R _448_492 (.A(clknet_leaf_0_clk),
    .Y(net897));
 INVx1_ASAP7_75t_R _448_493 (.A(clknet_leaf_17_clk),
    .Y(net898));
 INVx1_ASAP7_75t_R _448_494 (.A(clknet_leaf_0_clk),
    .Y(net899));
 INVx1_ASAP7_75t_R _448_495 (.A(clknet_leaf_0_clk),
    .Y(net900));
 INVx1_ASAP7_75t_R _448_496 (.A(clknet_leaf_0_clk),
    .Y(net901));
 INVx1_ASAP7_75t_R _448_497 (.A(clknet_leaf_17_clk),
    .Y(net902));
 INVx1_ASAP7_75t_R _498 (.A(clknet_leaf_0_clk),
    .Y(net903));
 INVx1_ASAP7_75t_R _498_499 (.A(clknet_leaf_3_clk),
    .Y(net904));
 INVx1_ASAP7_75t_R _498_500 (.A(clknet_leaf_2_clk),
    .Y(net905));
 INVx1_ASAP7_75t_R _498_501 (.A(clknet_leaf_3_clk),
    .Y(net906));
 INVx1_ASAP7_75t_R _498_502 (.A(clknet_leaf_3_clk),
    .Y(net907));
 INVx1_ASAP7_75t_R _498_503 (.A(clknet_leaf_3_clk),
    .Y(net908));
 INVx1_ASAP7_75t_R _498_504 (.A(clknet_leaf_3_clk),
    .Y(net909));
 INVx1_ASAP7_75t_R _498_505 (.A(clknet_leaf_3_clk),
    .Y(net910));
 INVx1_ASAP7_75t_R _498_506 (.A(clknet_leaf_3_clk),
    .Y(net911));
 INVx1_ASAP7_75t_R _498_507 (.A(clknet_leaf_3_clk),
    .Y(net912));
 INVx1_ASAP7_75t_R _498_508 (.A(clknet_leaf_3_clk),
    .Y(net913));
 INVx1_ASAP7_75t_R _498_509 (.A(clknet_leaf_3_clk),
    .Y(net914));
 INVx1_ASAP7_75t_R _498_510 (.A(clknet_leaf_3_clk),
    .Y(net915));
 INVx1_ASAP7_75t_R _498_511 (.A(clknet_leaf_3_clk),
    .Y(net916));
 INVx1_ASAP7_75t_R _498_512 (.A(clknet_leaf_2_clk),
    .Y(net917));
 INVx1_ASAP7_75t_R _498_513 (.A(clknet_leaf_2_clk),
    .Y(net918));
 INVx1_ASAP7_75t_R _498_514 (.A(clknet_leaf_4_clk),
    .Y(net919));
 INVx1_ASAP7_75t_R _498_515 (.A(clknet_leaf_2_clk),
    .Y(net920));
 INVx1_ASAP7_75t_R _498_516 (.A(clknet_leaf_2_clk),
    .Y(net921));
 INVx1_ASAP7_75t_R _498_517 (.A(clknet_leaf_17_clk),
    .Y(net922));
 INVx1_ASAP7_75t_R _498_518 (.A(clknet_leaf_2_clk),
    .Y(net923));
 INVx1_ASAP7_75t_R _498_519 (.A(clknet_leaf_15_clk),
    .Y(net924));
 INVx1_ASAP7_75t_R _498_520 (.A(clknet_leaf_0_clk),
    .Y(net925));
 INVx1_ASAP7_75t_R _498_521 (.A(clknet_leaf_0_clk),
    .Y(net926));
 INVx1_ASAP7_75t_R _498_522 (.A(clknet_leaf_0_clk),
    .Y(net927));
 INVx1_ASAP7_75t_R _498_523 (.A(clknet_leaf_8_clk),
    .Y(net928));
 INVx1_ASAP7_75t_R _498_524 (.A(clknet_leaf_7_clk),
    .Y(net929));
 INVx1_ASAP7_75t_R _498_525 (.A(clknet_leaf_1_clk),
    .Y(net930));
 INVx1_ASAP7_75t_R _498_526 (.A(clknet_leaf_8_clk),
    .Y(net931));
 INVx1_ASAP7_75t_R _498_527 (.A(clknet_leaf_6_clk),
    .Y(net932));
 INVx1_ASAP7_75t_R _498_528 (.A(clknet_leaf_11_clk),
    .Y(net933));
 INVx1_ASAP7_75t_R _498_529 (.A(clknet_leaf_7_clk),
    .Y(net934));
 INVx1_ASAP7_75t_R _498_530 (.A(clknet_leaf_7_clk),
    .Y(net935));
 BUFx4_ASAP7_75t_R clkbuf_leaf_1_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_1_clk));
 BUFx4_ASAP7_75t_R clkbuf_leaf_2_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_2_clk));
 BUFx4_ASAP7_75t_R clkbuf_leaf_3_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_3_clk));
 BUFx4_ASAP7_75t_R clkbuf_leaf_4_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_4_clk));
 BUFx4_ASAP7_75t_R clkbuf_leaf_5_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_5_clk));
 BUFx4_ASAP7_75t_R clkbuf_leaf_6_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_6_clk));
 BUFx4_ASAP7_75t_R clkbuf_leaf_7_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_7_clk));
 BUFx4_ASAP7_75t_R clkbuf_leaf_8_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_8_clk));
 BUFx4_ASAP7_75t_R clkbuf_leaf_9_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_9_clk));
 BUFx4_ASAP7_75t_R clkbuf_leaf_10_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_10_clk));
 BUFx4_ASAP7_75t_R clkbuf_leaf_11_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_11_clk));
 BUFx4_ASAP7_75t_R clkbuf_leaf_12_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_12_clk));
 BUFx4_ASAP7_75t_R clkbuf_leaf_13_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_13_clk));
 BUFx4_ASAP7_75t_R clkbuf_leaf_14_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_14_clk));
 BUFx4_ASAP7_75t_R clkbuf_leaf_15_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_15_clk));
 BUFx4_ASAP7_75t_R clkbuf_leaf_16_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_16_clk));
 BUFx4_ASAP7_75t_R clkbuf_leaf_17_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_17_clk));
 BUFx4_ASAP7_75t_R clkbuf_0_clk (.A(clk),
    .Y(clknet_0_clk));
 BUFx4_ASAP7_75t_R clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Y(clknet_1_0__leaf_clk));
 BUFx4_ASAP7_75t_R clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Y(clknet_1_1__leaf_clk));
 BUFx6f_ASAP7_75t_R split531 (.A(_17685_),
    .Y(net936));
 BUFx10_ASAP7_75t_R split532 (.A(_18296_),
    .Y(net937));
 BUFx12f_ASAP7_75t_R split533 (.A(_01318_),
    .Y(net938));
 BUFx6f_ASAP7_75t_R split534 (.A(net1348),
    .Y(net939));
 BUFx6f_ASAP7_75t_R split535 (.A(_01148_),
    .Y(net940));
 BUFx10_ASAP7_75t_R split536 (.A(_17563_),
    .Y(net941));
 BUFx3_ASAP7_75t_R rebuffer537 (.A(_09890_),
    .Y(net942));
 BUFx2_ASAP7_75t_R rebuffer538 (.A(net942),
    .Y(net943));
 BUFx2_ASAP7_75t_R rebuffer539 (.A(net942),
    .Y(net944));
 BUFx6f_ASAP7_75t_R rebuffer540 (.A(_09890_),
    .Y(net945));
 BUFx2_ASAP7_75t_R rebuffer541 (.A(net945),
    .Y(net946));
 BUFx6f_ASAP7_75t_R rebuffer542 (.A(net945),
    .Y(net947));
 BUFx6f_ASAP7_75t_R rebuffer543 (.A(net947),
    .Y(net948));
 BUFx6f_ASAP7_75t_R rebuffer544 (.A(net945),
    .Y(net949));
 BUFx6f_ASAP7_75t_R rebuffer545 (.A(_01765_),
    .Y(net950));
 BUFx2_ASAP7_75t_R rebuffer546 (.A(net950),
    .Y(net951));
 BUFx2_ASAP7_75t_R rebuffer547 (.A(net950),
    .Y(net952));
 BUFx2_ASAP7_75t_R rebuffer548 (.A(net950),
    .Y(net953));
 BUFx2_ASAP7_75t_R rebuffer549 (.A(_01765_),
    .Y(net954));
 BUFx2_ASAP7_75t_R rebuffer550 (.A(_01765_),
    .Y(net955));
 BUFx3_ASAP7_75t_R rebuffer551 (.A(_10310_),
    .Y(net956));
 BUFx2_ASAP7_75t_R rebuffer552 (.A(_10310_),
    .Y(net957));
 BUFx2_ASAP7_75t_R rebuffer553 (.A(net957),
    .Y(net958));
 BUFx2_ASAP7_75t_R rebuffer554 (.A(net958),
    .Y(net959));
 BUFx3_ASAP7_75t_R rebuffer555 (.A(_10310_),
    .Y(net960));
 BUFx2_ASAP7_75t_R rebuffer556 (.A(net960),
    .Y(net961));
 BUFx6f_ASAP7_75t_R rebuffer557 (.A(net2739),
    .Y(net962));
 BUFx3_ASAP7_75t_R rebuffer558 (.A(_05737_),
    .Y(net963));
 BUFx10_ASAP7_75t_R split559 (.A(_05131_),
    .Y(net964));
 BUFx2_ASAP7_75t_R rebuffer560 (.A(_10348_),
    .Y(net965));
 BUFx2_ASAP7_75t_R rebuffer561 (.A(_10348_),
    .Y(net966));
 BUFx2_ASAP7_75t_R rebuffer562 (.A(net966),
    .Y(net967));
 BUFx12f_ASAP7_75t_R rebuffer563 (.A(_10348_),
    .Y(net968));
 BUFx2_ASAP7_75t_R rebuffer564 (.A(net968),
    .Y(net969));
 BUFx2_ASAP7_75t_R rebuffer565 (.A(net968),
    .Y(net970));
 BUFx2_ASAP7_75t_R rebuffer566 (.A(net968),
    .Y(net971));
 BUFx6f_ASAP7_75t_R rebuffer567 (.A(net968),
    .Y(net972));
 BUFx2_ASAP7_75t_R rebuffer568 (.A(_10348_),
    .Y(net973));
 BUFx6f_ASAP7_75t_R split569 (.A(_17958_),
    .Y(net974));
 BUFx10_ASAP7_75t_R split570 (.A(net1372),
    .Y(net975));
 BUFx6f_ASAP7_75t_R rebuffer571 (.A(_09881_),
    .Y(net976));
 BUFx6f_ASAP7_75t_R rebuffer572 (.A(net976),
    .Y(net977));
 BUFx2_ASAP7_75t_R rebuffer573 (.A(net976),
    .Y(net978));
 BUFx2_ASAP7_75t_R rebuffer574 (.A(net976),
    .Y(net979));
 BUFx6f_ASAP7_75t_R split575 (.A(_05805_),
    .Y(net980));
 BUFx6f_ASAP7_75t_R rebuffer576 (.A(_09607_),
    .Y(net981));
 BUFx2_ASAP7_75t_R rebuffer577 (.A(net981),
    .Y(net982));
 BUFx2_ASAP7_75t_R rebuffer578 (.A(net982),
    .Y(net983));
 BUFx2_ASAP7_75t_R rebuffer579 (.A(net981),
    .Y(net984));
 BUFx2_ASAP7_75t_R rebuffer580 (.A(net984),
    .Y(net985));
 BUFx2_ASAP7_75t_R rebuffer581 (.A(net985),
    .Y(net986));
 BUFx2_ASAP7_75t_R rebuffer582 (.A(net984),
    .Y(net987));
 BUFx2_ASAP7_75t_R rebuffer583 (.A(net2798),
    .Y(net988));
 BUFx6f_ASAP7_75t_R split584 (.A(_00584_),
    .Y(net989));
 BUFx10_ASAP7_75t_R split585 (.A(_05135_),
    .Y(net990));
 BUFx6f_ASAP7_75t_R split586 (.A(_21938_),
    .Y(net991));
 BUFx6f_ASAP7_75t_R split587 (.A(_05105_),
    .Y(net992));
 BUFx2_ASAP7_75t_R rebuffer588 (.A(_21879_),
    .Y(net993));
 BUFx2_ASAP7_75t_R rebuffer589 (.A(net993),
    .Y(net994));
 BUFx2_ASAP7_75t_R rebuffer590 (.A(_21879_),
    .Y(net995));
 BUFx2_ASAP7_75t_R rebuffer591 (.A(net995),
    .Y(net996));
 BUFx6f_ASAP7_75t_R rebuffer592 (.A(_17685_),
    .Y(net997));
 BUFx6f_ASAP7_75t_R rebuffer593 (.A(_17685_),
    .Y(net998));
 BUFx6f_ASAP7_75t_R rebuffer594 (.A(net998),
    .Y(net999));
 BUFx6f_ASAP7_75t_R split595 (.A(_00583_),
    .Y(net1000));
 BUFx2_ASAP7_75t_R rebuffer596 (.A(_17536_),
    .Y(net1001));
 BUFx2_ASAP7_75t_R rebuffer597 (.A(net1001),
    .Y(net1002));
 BUFx12f_ASAP7_75t_R rebuffer598 (.A(_17536_),
    .Y(net1003));
 BUFx2_ASAP7_75t_R rebuffer599 (.A(net1003),
    .Y(net1004));
 BUFx2_ASAP7_75t_R rebuffer600 (.A(net1003),
    .Y(net1005));
 BUFx6f_ASAP7_75t_R rebuffer601 (.A(net1003),
    .Y(net1006));
 BUFx2_ASAP7_75t_R rebuffer602 (.A(net1003),
    .Y(net1007));
 BUFx2_ASAP7_75t_R rebuffer603 (.A(net1007),
    .Y(net1008));
 BUFx2_ASAP7_75t_R rebuffer604 (.A(_18514_),
    .Y(net1009));
 BUFx2_ASAP7_75t_R rebuffer605 (.A(net1069),
    .Y(net1010));
 BUFx2_ASAP7_75t_R rebuffer606 (.A(_18514_),
    .Y(net1011));
 BUFx2_ASAP7_75t_R rebuffer607 (.A(_05936_),
    .Y(net1012));
 BUFx2_ASAP7_75t_R rebuffer608 (.A(_00655_),
    .Y(net1013));
 BUFx2_ASAP7_75t_R rebuffer609 (.A(_00655_),
    .Y(net1014));
 BUFx6f_ASAP7_75t_R rebuffer610 (.A(_00655_),
    .Y(net1015));
 BUFx2_ASAP7_75t_R rebuffer611 (.A(net1015),
    .Y(net1016));
 BUFx12f_ASAP7_75t_R rebuffer612 (.A(_00655_),
    .Y(net1017));
 BUFx2_ASAP7_75t_R rebuffer613 (.A(net1017),
    .Y(net1018));
 BUFx4f_ASAP7_75t_R rebuffer614 (.A(_00655_),
    .Y(net1019));
 BUFx2_ASAP7_75t_R rebuffer615 (.A(net1019),
    .Y(net1020));
 BUFx2_ASAP7_75t_R rebuffer616 (.A(net1019),
    .Y(net1021));
 BUFx2_ASAP7_75t_R rebuffer617 (.A(net1021),
    .Y(net1022));
 BUFx2_ASAP7_75t_R rebuffer618 (.A(net1021),
    .Y(net1023));
 BUFx2_ASAP7_75t_R rebuffer619 (.A(net1023),
    .Y(net1024));
 BUFx2_ASAP7_75t_R rebuffer620 (.A(_01513_),
    .Y(net1025));
 BUFx2_ASAP7_75t_R rebuffer621 (.A(net1025),
    .Y(net1026));
 BUFx2_ASAP7_75t_R rebuffer622 (.A(net2470),
    .Y(net1027));
 BUFx6f_ASAP7_75t_R rebuffer623 (.A(net2470),
    .Y(net1028));
 BUFx2_ASAP7_75t_R rebuffer624 (.A(net1028),
    .Y(net1029));
 BUFx6f_ASAP7_75t_R split625 (.A(_17582_),
    .Y(net1030));
 BUFx3_ASAP7_75t_R rebuffer626 (.A(_05455_),
    .Y(net1031));
 BUFx2_ASAP7_75t_R rebuffer627 (.A(net1031),
    .Y(net1032));
 BUFx2_ASAP7_75t_R rebuffer628 (.A(net1032),
    .Y(net1033));
 BUFx12f_ASAP7_75t_R rebuffer629 (.A(_05455_),
    .Y(net1034));
 BUFx2_ASAP7_75t_R rebuffer630 (.A(net1034),
    .Y(net1035));
 BUFx4f_ASAP7_75t_R rebuffer631 (.A(net1035),
    .Y(net1036));
 BUFx6f_ASAP7_75t_R split632 (.A(_06429_),
    .Y(net1037));
 BUFx6f_ASAP7_75t_R split633 (.A(_02259_),
    .Y(net1038));
 BUFx2_ASAP7_75t_R rebuffer634 (.A(_21907_),
    .Y(net1039));
 BUFx12f_ASAP7_75t_R rebuffer635 (.A(_21907_),
    .Y(net1040));
 BUFx2_ASAP7_75t_R rebuffer636 (.A(net1040),
    .Y(net1041));
 BUFx2_ASAP7_75t_R rebuffer637 (.A(net1041),
    .Y(net1042));
 BUFx2_ASAP7_75t_R rebuffer638 (.A(net1040),
    .Y(net1043));
 BUFx2_ASAP7_75t_R rebuffer639 (.A(net1040),
    .Y(net1044));
 BUFx2_ASAP7_75t_R rebuffer640 (.A(net1044),
    .Y(net1045));
 BUFx2_ASAP7_75t_R rebuffer641 (.A(net1040),
    .Y(net1046));
 BUFx4f_ASAP7_75t_R split642 (.A(_06145_),
    .Y(net1047));
 BUFx10_ASAP7_75t_R split643 (.A(_21922_),
    .Y(net1048));
 BUFx10_ASAP7_75t_R split644 (.A(net1168),
    .Y(net1049));
 BUFx2_ASAP7_75t_R rebuffer645 (.A(_17999_),
    .Y(net1050));
 BUFx6f_ASAP7_75t_R rebuffer646 (.A(_10442_),
    .Y(net1051));
 BUFx2_ASAP7_75t_R rebuffer647 (.A(net1051),
    .Y(net1052));
 BUFx2_ASAP7_75t_R rebuffer648 (.A(net1051),
    .Y(net1053));
 BUFx2_ASAP7_75t_R rebuffer649 (.A(net1051),
    .Y(net1054));
 BUFx4f_ASAP7_75t_R rebuffer650 (.A(_10442_),
    .Y(net1055));
 BUFx2_ASAP7_75t_R rebuffer651 (.A(net1055),
    .Y(net1056));
 BUFx2_ASAP7_75t_R rebuffer652 (.A(_00647_),
    .Y(net1057));
 BUFx12f_ASAP7_75t_R rebuffer653 (.A(_00647_),
    .Y(net1058));
 BUFx2_ASAP7_75t_R rebuffer654 (.A(net3204),
    .Y(net1059));
 BUFx2_ASAP7_75t_R rebuffer655 (.A(net1058),
    .Y(net1060));
 BUFx2_ASAP7_75t_R rebuffer656 (.A(net1060),
    .Y(net1061));
 BUFx2_ASAP7_75t_R rebuffer657 (.A(net1061),
    .Y(net1062));
 BUFx2_ASAP7_75t_R rebuffer658 (.A(net3204),
    .Y(net1063));
 BUFx12f_ASAP7_75t_R rebuffer659 (.A(_00647_),
    .Y(net1064));
 BUFx2_ASAP7_75t_R rebuffer660 (.A(_09933_),
    .Y(net1065));
 BUFx2_ASAP7_75t_R rebuffer661 (.A(net1065),
    .Y(net1066));
 BUFx3_ASAP7_75t_R rebuffer662 (.A(net1065),
    .Y(net1067));
 BUFx4f_ASAP7_75t_R split663 (.A(_17999_),
    .Y(net1068));
 BUFx3_ASAP7_75t_R split664 (.A(_18514_),
    .Y(net1069));
 BUFx12f_ASAP7_75t_R rebuffer665 (.A(_17960_),
    .Y(net1070));
 BUFx2_ASAP7_75t_R rebuffer666 (.A(net1070),
    .Y(net1071));
 BUFx4f_ASAP7_75t_R rebuffer667 (.A(net1070),
    .Y(net1072));
 BUFx2_ASAP7_75t_R rebuffer668 (.A(net1072),
    .Y(net1073));
 BUFx2_ASAP7_75t_R rebuffer669 (.A(net1072),
    .Y(net1074));
 BUFx2_ASAP7_75t_R rebuffer670 (.A(net1070),
    .Y(net1075));
 BUFx6f_ASAP7_75t_R split671 (.A(_01194_),
    .Y(net1076));
 BUFx6f_ASAP7_75t_R rebuffer672 (.A(_10394_),
    .Y(net1077));
 BUFx2_ASAP7_75t_R rebuffer673 (.A(net1077),
    .Y(net1078));
 BUFx6f_ASAP7_75t_R rebuffer674 (.A(_10394_),
    .Y(net1079));
 BUFx2_ASAP7_75t_R rebuffer675 (.A(net1079),
    .Y(net1080));
 BUFx6f_ASAP7_75t_R split676 (.A(_17645_),
    .Y(net1081));
 BUFx10_ASAP7_75t_R split677 (.A(_17596_),
    .Y(net1082));
 BUFx6f_ASAP7_75t_R split678 (.A(_06574_),
    .Y(net1083));
 BUFx6f_ASAP7_75t_R rebuffer679 (.A(_05532_),
    .Y(net1084));
 BUFx2_ASAP7_75t_R rebuffer680 (.A(net1084),
    .Y(net1085));
 BUFx2_ASAP7_75t_R rebuffer681 (.A(net2610),
    .Y(net1086));
 BUFx6f_ASAP7_75t_R split682 (.A(net1681),
    .Y(net1087));
 BUFx3_ASAP7_75t_R rebuffer683 (.A(_17534_),
    .Y(net1088));
 BUFx2_ASAP7_75t_R rebuffer684 (.A(net1088),
    .Y(net1089));
 BUFx6f_ASAP7_75t_R split685 (.A(_10396_),
    .Y(net1090));
 BUFx10_ASAP7_75t_R split686 (.A(_05070_),
    .Y(net1091));
 BUFx6f_ASAP7_75t_R rebuffer687 (.A(_06037_),
    .Y(net1092));
 BUFx6f_ASAP7_75t_R rebuffer688 (.A(net1092),
    .Y(net1093));
 BUFx2_ASAP7_75t_R rebuffer689 (.A(net1093),
    .Y(net1094));
 BUFx2_ASAP7_75t_R rebuffer690 (.A(net1094),
    .Y(net1095));
 BUFx6f_ASAP7_75t_R rebuffer691 (.A(_06037_),
    .Y(net1096));
 BUFx10_ASAP7_75t_R split692 (.A(_17815_),
    .Y(net1097));
 BUFx6f_ASAP7_75t_R split693 (.A(_17593_),
    .Y(net1098));
 BUFx12f_ASAP7_75t_R rebuffer694 (.A(_09596_),
    .Y(net1099));
 BUFx2_ASAP7_75t_R rebuffer695 (.A(net1099),
    .Y(net1100));
 BUFx2_ASAP7_75t_R rebuffer696 (.A(net1100),
    .Y(net1101));
 BUFx6f_ASAP7_75t_R split697 (.A(_09798_),
    .Y(net1102));
 BUFx6f_ASAP7_75t_R split698 (.A(_17570_),
    .Y(net1103));
 BUFx6f_ASAP7_75t_R split699 (.A(_01496_),
    .Y(net1104));
 BUFx6f_ASAP7_75t_R rebuffer700 (.A(_00615_),
    .Y(net1105));
 BUFx2_ASAP7_75t_R rebuffer701 (.A(net1105),
    .Y(net1106));
 BUFx12f_ASAP7_75t_R rebuffer702 (.A(net1105),
    .Y(net1107));
 BUFx2_ASAP7_75t_R rebuffer703 (.A(net1107),
    .Y(net1108));
 BUFx2_ASAP7_75t_R rebuffer704 (.A(net1107),
    .Y(net1109));
 BUFx2_ASAP7_75t_R rebuffer705 (.A(net1109),
    .Y(net1110));
 BUFx12f_ASAP7_75t_R rebuffer706 (.A(_00615_),
    .Y(net1111));
 BUFx2_ASAP7_75t_R rebuffer707 (.A(net1111),
    .Y(net1112));
 BUFx2_ASAP7_75t_R rebuffer708 (.A(net1111),
    .Y(net1113));
 BUFx6f_ASAP7_75t_R split709 (.A(_10333_),
    .Y(net1114));
 BUFx10_ASAP7_75t_R split710 (.A(_10365_),
    .Y(net1115));
 BUFx6f_ASAP7_75t_R split711 (.A(net1357),
    .Y(net1116));
 BUFx6f_ASAP7_75t_R split712 (.A(net1642),
    .Y(net1117));
 BUFx6f_ASAP7_75t_R split713 (.A(_05825_),
    .Y(net1118));
 BUFx6f_ASAP7_75t_R split714 (.A(_01384_),
    .Y(net1119));
 BUFx6f_ASAP7_75t_R split715 (.A(_00639_),
    .Y(net1120));
 BUFx6f_ASAP7_75t_R split716 (.A(_18014_),
    .Y(net1121));
 BUFx6f_ASAP7_75t_R split717 (.A(_01128_),
    .Y(net1122));
 BUFx10_ASAP7_75t_R split718 (.A(net1533),
    .Y(net1123));
 BUFx6f_ASAP7_75t_R split719 (.A(_05490_),
    .Y(net1124));
 BUFx6f_ASAP7_75t_R split720 (.A(_10451_),
    .Y(net1125));
 BUFx2_ASAP7_75t_R rebuffer721 (.A(_01775_),
    .Y(net1126));
 BUFx12f_ASAP7_75t_R rebuffer722 (.A(_01775_),
    .Y(net1127));
 BUFx2_ASAP7_75t_R rebuffer723 (.A(net1127),
    .Y(net1128));
 BUFx2_ASAP7_75t_R rebuffer724 (.A(net1128),
    .Y(net1129));
 BUFx2_ASAP7_75t_R rebuffer725 (.A(net1127),
    .Y(net1130));
 BUFx2_ASAP7_75t_R rebuffer726 (.A(net1130),
    .Y(net1131));
 BUFx2_ASAP7_75t_R rebuffer727 (.A(net1127),
    .Y(net1132));
 BUFx2_ASAP7_75t_R rebuffer728 (.A(_01775_),
    .Y(net1133));
 BUFx6f_ASAP7_75t_R rebuffer729 (.A(_01111_),
    .Y(net1134));
 BUFx2_ASAP7_75t_R rebuffer730 (.A(net1134),
    .Y(net1135));
 BUFx2_ASAP7_75t_R rebuffer731 (.A(net1135),
    .Y(net1136));
 BUFx2_ASAP7_75t_R rebuffer732 (.A(_01111_),
    .Y(net1137));
 BUFx6f_ASAP7_75t_R split733 (.A(_01892_),
    .Y(net1138));
 BUFx6f_ASAP7_75t_R split734 (.A(net1405),
    .Y(net1139));
 BUFx6f_ASAP7_75t_R split735 (.A(_05165_),
    .Y(net1140));
 BUFx2_ASAP7_75t_R rebuffer736 (.A(_01318_),
    .Y(net1141));
 BUFx6f_ASAP7_75t_R rebuffer737 (.A(_01318_),
    .Y(net1142));
 BUFx4f_ASAP7_75t_R rebuffer738 (.A(_10408_),
    .Y(net1143));
 BUFx3_ASAP7_75t_R rebuffer739 (.A(net1143),
    .Y(net1144));
 BUFx6f_ASAP7_75t_R rebuffer740 (.A(_17999_),
    .Y(net1145));
 BUFx12_ASAP7_75t_R split741 (.A(net1621),
    .Y(net1146));
 BUFx12f_ASAP7_75t_R rebuffer742 (.A(_00624_),
    .Y(net1147));
 BUFx2_ASAP7_75t_R rebuffer743 (.A(net1147),
    .Y(net1148));
 BUFx2_ASAP7_75t_R rebuffer744 (.A(net1148),
    .Y(net1149));
 BUFx2_ASAP7_75t_R rebuffer745 (.A(net1148),
    .Y(net1150));
 BUFx6f_ASAP7_75t_R rebuffer746 (.A(net1147),
    .Y(net1151));
 BUFx2_ASAP7_75t_R rebuffer747 (.A(net1151),
    .Y(net1152));
 BUFx2_ASAP7_75t_R rebuffer748 (.A(net1152),
    .Y(net1153));
 BUFx2_ASAP7_75t_R rebuffer749 (.A(net1153),
    .Y(net1154));
 BUFx2_ASAP7_75t_R rebuffer750 (.A(net1151),
    .Y(net1155));
 BUFx2_ASAP7_75t_R rebuffer751 (.A(_00624_),
    .Y(net1156));
 BUFx6f_ASAP7_75t_R split752 (.A(_01825_),
    .Y(net1157));
 BUFx12_ASAP7_75t_R split753 (.A(_01246_),
    .Y(net1158));
 BUFx12f_ASAP7_75t_R rebuffer754 (.A(_00656_),
    .Y(net1159));
 BUFx3_ASAP7_75t_R rebuffer755 (.A(net1159),
    .Y(net1160));
 BUFx12f_ASAP7_75t_R rebuffer756 (.A(net1159),
    .Y(net1161));
 BUFx2_ASAP7_75t_R rebuffer757 (.A(net1161),
    .Y(net1162));
 BUFx2_ASAP7_75t_R rebuffer758 (.A(net1162),
    .Y(net1163));
 BUFx3_ASAP7_75t_R rebuffer759 (.A(net1161),
    .Y(net1164));
 BUFx2_ASAP7_75t_R rebuffer760 (.A(net1164),
    .Y(net1165));
 BUFx2_ASAP7_75t_R rebuffer761 (.A(net1164),
    .Y(net1166));
 BUFx2_ASAP7_75t_R rebuffer762 (.A(net1166),
    .Y(net1167));
 BUFx2_ASAP7_75t_R rebuffer763 (.A(_00552_),
    .Y(net1168));
 BUFx12f_ASAP7_75t_R rebuffer764 (.A(_00552_),
    .Y(net1169));
 BUFx12f_ASAP7_75t_R rebuffer765 (.A(net1169),
    .Y(net1170));
 BUFx2_ASAP7_75t_R rebuffer766 (.A(net1170),
    .Y(net1171));
 BUFx2_ASAP7_75t_R rebuffer767 (.A(net1171),
    .Y(net1172));
 BUFx2_ASAP7_75t_R rebuffer768 (.A(net1170),
    .Y(net1173));
 BUFx12f_ASAP7_75t_R rebuffer769 (.A(_05778_),
    .Y(net1174));
 BUFx2_ASAP7_75t_R rebuffer770 (.A(net1174),
    .Y(net1175));
 BUFx6f_ASAP7_75t_R rebuffer771 (.A(net1175),
    .Y(net1176));
 BUFx2_ASAP7_75t_R rebuffer772 (.A(net1176),
    .Y(net1177));
 BUFx2_ASAP7_75t_R rebuffer773 (.A(net1176),
    .Y(net1178));
 BUFx2_ASAP7_75t_R rebuffer774 (.A(_05778_),
    .Y(net1179));
 BUFx2_ASAP7_75t_R rebuffer775 (.A(net1179),
    .Y(net1180));
 BUFx2_ASAP7_75t_R rebuffer776 (.A(_05778_),
    .Y(net1181));
 BUFx2_ASAP7_75t_R rebuffer777 (.A(net1181),
    .Y(net1182));
 BUFx2_ASAP7_75t_R rebuffer778 (.A(net1181),
    .Y(net1183));
 BUFx12f_ASAP7_75t_R rebuffer779 (.A(_00560_),
    .Y(net1184));
 BUFx2_ASAP7_75t_R rebuffer780 (.A(net2770),
    .Y(net1185));
 BUFx3_ASAP7_75t_R rebuffer781 (.A(net1185),
    .Y(net1186));
 BUFx2_ASAP7_75t_R rebuffer782 (.A(net2770),
    .Y(net1187));
 BUFx12f_ASAP7_75t_R rebuffer783 (.A(net1184),
    .Y(net1188));
 BUFx2_ASAP7_75t_R rebuffer784 (.A(net1188),
    .Y(net1189));
 BUFx2_ASAP7_75t_R rebuffer785 (.A(net1184),
    .Y(net1190));
 BUFx2_ASAP7_75t_R rebuffer786 (.A(net1184),
    .Y(net1191));
 BUFx2_ASAP7_75t_R rebuffer787 (.A(net2770),
    .Y(net1192));
 BUFx2_ASAP7_75t_R rebuffer788 (.A(net2770),
    .Y(net1193));
 BUFx4f_ASAP7_75t_R rebuffer789 (.A(net1193),
    .Y(net1194));
 BUFx6f_ASAP7_75t_R rebuffer790 (.A(_01127_),
    .Y(net1195));
 BUFx6f_ASAP7_75t_R rebuffer791 (.A(_01127_),
    .Y(net1196));
 BUFx3_ASAP7_75t_R rebuffer792 (.A(net1196),
    .Y(net1197));
 BUFx6f_ASAP7_75t_R rebuffer793 (.A(_18295_),
    .Y(net1198));
 BUFx2_ASAP7_75t_R rebuffer794 (.A(net1198),
    .Y(net1199));
 BUFx2_ASAP7_75t_R rebuffer795 (.A(_00584_),
    .Y(net1200));
 BUFx12f_ASAP7_75t_R rebuffer796 (.A(_00584_),
    .Y(net1201));
 BUFx2_ASAP7_75t_R rebuffer797 (.A(net1201),
    .Y(net1202));
 BUFx6f_ASAP7_75t_R rebuffer798 (.A(net1201),
    .Y(net1203));
 BUFx2_ASAP7_75t_R rebuffer799 (.A(net1203),
    .Y(net1204));
 BUFx3_ASAP7_75t_R rebuffer800 (.A(_05460_),
    .Y(net1205));
 BUFx2_ASAP7_75t_R rebuffer801 (.A(net1205),
    .Y(net1206));
 BUFx6f_ASAP7_75t_R rebuffer802 (.A(net1205),
    .Y(net1207));
 BUFx6f_ASAP7_75t_R rebuffer803 (.A(_05460_),
    .Y(net1208));
 BUFx2_ASAP7_75t_R rebuffer804 (.A(net1208),
    .Y(net1209));
 BUFx2_ASAP7_75t_R rebuffer805 (.A(net1209),
    .Y(net1210));
 BUFx2_ASAP7_75t_R rebuffer806 (.A(net1209),
    .Y(net1211));
 BUFx2_ASAP7_75t_R rebuffer807 (.A(net1208),
    .Y(net1212));
 BUFx2_ASAP7_75t_R rebuffer808 (.A(net1212),
    .Y(net1213));
 BUFx2_ASAP7_75t_R rebuffer809 (.A(_06278_),
    .Y(net1214));
 BUFx3_ASAP7_75t_R rebuffer810 (.A(_06278_),
    .Y(net1215));
 BUFx2_ASAP7_75t_R rebuffer811 (.A(net1215),
    .Y(net1216));
 BUFx6f_ASAP7_75t_R split812 (.A(_06085_),
    .Y(net1217));
 BUFx6f_ASAP7_75t_R rebuffer813 (.A(_09586_),
    .Y(net1218));
 BUFx2_ASAP7_75t_R rebuffer814 (.A(net1218),
    .Y(net1219));
 BUFx2_ASAP7_75t_R rebuffer815 (.A(net1219),
    .Y(net1220));
 BUFx12f_ASAP7_75t_R rebuffer816 (.A(_00543_),
    .Y(net1221));
 BUFx12f_ASAP7_75t_R rebuffer817 (.A(net1221),
    .Y(net1222));
 BUFx6f_ASAP7_75t_R rebuffer818 (.A(net1222),
    .Y(net1223));
 BUFx2_ASAP7_75t_R rebuffer819 (.A(net1223),
    .Y(net1224));
 BUFx12f_ASAP7_75t_R rebuffer820 (.A(net1221),
    .Y(net1225));
 BUFx2_ASAP7_75t_R rebuffer821 (.A(net1225),
    .Y(net1226));
 BUFx2_ASAP7_75t_R rebuffer822 (.A(net1225),
    .Y(net1227));
 BUFx2_ASAP7_75t_R rebuffer823 (.A(net1225),
    .Y(net1228));
 BUFx2_ASAP7_75t_R rebuffer824 (.A(net1228),
    .Y(net1229));
 BUFx2_ASAP7_75t_R rebuffer825 (.A(net1815),
    .Y(net1230));
 BUFx2_ASAP7_75t_R rebuffer826 (.A(net1815),
    .Y(net1231));
 BUFx3_ASAP7_75t_R rebuffer827 (.A(_17946_),
    .Y(net1232));
 BUFx2_ASAP7_75t_R rebuffer828 (.A(_17946_),
    .Y(net1233));
 BUFx2_ASAP7_75t_R rebuffer829 (.A(_17946_),
    .Y(net1234));
 BUFx12f_ASAP7_75t_R rebuffer830 (.A(_17946_),
    .Y(net1235));
 BUFx2_ASAP7_75t_R rebuffer831 (.A(_17946_),
    .Y(net1236));
 BUFx6f_ASAP7_75t_R split832 (.A(_05073_),
    .Y(net1237));
 BUFx3_ASAP7_75t_R rebuffer833 (.A(_01524_),
    .Y(net1238));
 BUFx2_ASAP7_75t_R rebuffer834 (.A(net1238),
    .Y(net1239));
 BUFx2_ASAP7_75t_R rebuffer835 (.A(_01524_),
    .Y(net1240));
 BUFx4f_ASAP7_75t_R rebuffer836 (.A(_01524_),
    .Y(net1241));
 BUFx2_ASAP7_75t_R rebuffer837 (.A(net1241),
    .Y(net1242));
 BUFx2_ASAP7_75t_R rebuffer838 (.A(net1242),
    .Y(net1243));
 BUFx3_ASAP7_75t_R rebuffer839 (.A(_01825_),
    .Y(net1244));
 BUFx4f_ASAP7_75t_R rebuffer840 (.A(_01825_),
    .Y(net1245));
 BUFx6f_ASAP7_75t_R split841 (.A(_09738_),
    .Y(net1246));
 BUFx12f_ASAP7_75t_R rebuffer842 (.A(_09878_),
    .Y(net1247));
 BUFx2_ASAP7_75t_R rebuffer843 (.A(net1247),
    .Y(net1248));
 BUFx4f_ASAP7_75t_R rebuffer844 (.A(net1247),
    .Y(net1249));
 BUFx3_ASAP7_75t_R rebuffer845 (.A(_09878_),
    .Y(net1250));
 BUFx2_ASAP7_75t_R rebuffer846 (.A(net1250),
    .Y(net1251));
 BUFx2_ASAP7_75t_R rebuffer847 (.A(net1250),
    .Y(net1252));
 BUFx6f_ASAP7_75t_R split848 (.A(_01797_),
    .Y(net1253));
 BUFx6f_ASAP7_75t_R split849 (.A(_18239_),
    .Y(net1254));
 BUFx3_ASAP7_75t_R rebuffer850 (.A(_21937_),
    .Y(net1255));
 BUFx6f_ASAP7_75t_R rebuffer851 (.A(net1255),
    .Y(net1256));
 BUFx2_ASAP7_75t_R rebuffer852 (.A(net1256),
    .Y(net1257));
 BUFx2_ASAP7_75t_R rebuffer853 (.A(net1256),
    .Y(net1258));
 BUFx2_ASAP7_75t_R rebuffer854 (.A(_21937_),
    .Y(net1259));
 BUFx2_ASAP7_75t_R rebuffer855 (.A(_06153_),
    .Y(net1260));
 BUFx2_ASAP7_75t_R rebuffer856 (.A(_06153_),
    .Y(net1261));
 BUFx2_ASAP7_75t_R rebuffer857 (.A(net1261),
    .Y(net1262));
 BUFx10_ASAP7_75t_R split858 (.A(_00640_),
    .Y(net1263));
 BUFx2_ASAP7_75t_R rebuffer859 (.A(_10318_),
    .Y(net1264));
 BUFx2_ASAP7_75t_R rebuffer860 (.A(net1264),
    .Y(net1265));
 BUFx6f_ASAP7_75t_R split861 (.A(_01188_),
    .Y(net1266));
 BUFx6f_ASAP7_75t_R split862 (.A(_05503_),
    .Y(net1267));
 BUFx2_ASAP7_75t_R rebuffer863 (.A(_10339_),
    .Y(net1268));
 BUFx2_ASAP7_75t_R rebuffer864 (.A(net1268),
    .Y(net1269));
 BUFx2_ASAP7_75t_R rebuffer865 (.A(net1269),
    .Y(net1270));
 BUFx2_ASAP7_75t_R rebuffer866 (.A(net1270),
    .Y(net1271));
 BUFx2_ASAP7_75t_R rebuffer867 (.A(net1270),
    .Y(net1272));
 BUFx2_ASAP7_75t_R rebuffer868 (.A(net3032),
    .Y(net1273));
 BUFx3_ASAP7_75t_R rebuffer869 (.A(_01115_),
    .Y(net1274));
 BUFx2_ASAP7_75t_R rebuffer870 (.A(_01115_),
    .Y(net1275));
 BUFx6f_ASAP7_75t_R split871 (.A(_00631_),
    .Y(net1276));
 BUFx6f_ASAP7_75t_R split872 (.A(net1682),
    .Y(net1277));
 BUFx6f_ASAP7_75t_R rebuffer873 (.A(_00616_),
    .Y(net1278));
 BUFx2_ASAP7_75t_R rebuffer874 (.A(net1278),
    .Y(net1279));
 BUFx2_ASAP7_75t_R rebuffer875 (.A(net1279),
    .Y(net1280));
 BUFx2_ASAP7_75t_R rebuffer876 (.A(net1280),
    .Y(net1281));
 BUFx6f_ASAP7_75t_R rebuffer877 (.A(_00616_),
    .Y(net1282));
 BUFx2_ASAP7_75t_R rebuffer878 (.A(net1282),
    .Y(net1283));
 BUFx2_ASAP7_75t_R rebuffer879 (.A(net1282),
    .Y(net1284));
 BUFx2_ASAP7_75t_R rebuffer880 (.A(net1284),
    .Y(net1285));
 BUFx2_ASAP7_75t_R rebuffer881 (.A(net1285),
    .Y(net1286));
 BUFx2_ASAP7_75t_R rebuffer882 (.A(net1282),
    .Y(net1287));
 BUFx6f_ASAP7_75t_R split883 (.A(_10628_),
    .Y(net1288));
 BUFx3_ASAP7_75t_R rebuffer884 (.A(_09636_),
    .Y(net1289));
 BUFx2_ASAP7_75t_R rebuffer885 (.A(net1289),
    .Y(net1290));
 BUFx2_ASAP7_75t_R rebuffer886 (.A(net1289),
    .Y(net1291));
 BUFx2_ASAP7_75t_R rebuffer887 (.A(net1291),
    .Y(net1292));
 BUFx3_ASAP7_75t_R rebuffer888 (.A(_01194_),
    .Y(net1293));
 BUFx2_ASAP7_75t_R rebuffer889 (.A(_01194_),
    .Y(net1294));
 BUFx2_ASAP7_75t_R rebuffer890 (.A(net2507),
    .Y(net1295));
 BUFx2_ASAP7_75t_R rebuffer891 (.A(net2507),
    .Y(net1296));
 BUFx2_ASAP7_75t_R rebuffer892 (.A(net2507),
    .Y(net1297));
 BUFx2_ASAP7_75t_R rebuffer893 (.A(_01768_),
    .Y(net1298));
 BUFx5_ASAP7_75t_R rebuffer894 (.A(_01768_),
    .Y(net1299));
 BUFx2_ASAP7_75t_R rebuffer895 (.A(net1299),
    .Y(net1300));
 BUFx2_ASAP7_75t_R rebuffer896 (.A(net1299),
    .Y(net1301));
 BUFx2_ASAP7_75t_R rebuffer897 (.A(net1299),
    .Y(net1302));
 BUFx2_ASAP7_75t_R rebuffer898 (.A(_05089_),
    .Y(net1303));
 BUFx2_ASAP7_75t_R rebuffer899 (.A(net1303),
    .Y(net1304));
 BUFx2_ASAP7_75t_R rebuffer900 (.A(_05089_),
    .Y(net1305));
 BUFx6f_ASAP7_75t_R split901 (.A(_10471_),
    .Y(net1306));
 BUFx6f_ASAP7_75t_R split902 (.A(_18532_),
    .Y(net1307));
 BUFx6f_ASAP7_75t_R rebuffer903 (.A(_18968_),
    .Y(net1308));
 BUFx2_ASAP7_75t_R rebuffer904 (.A(net1308),
    .Y(net1309));
 BUFx12f_ASAP7_75t_R rebuffer905 (.A(_00583_),
    .Y(net1310));
 BUFx12f_ASAP7_75t_R rebuffer906 (.A(net1310),
    .Y(net1311));
 BUFx2_ASAP7_75t_R rebuffer907 (.A(net1311),
    .Y(net1312));
 BUFx2_ASAP7_75t_R rebuffer908 (.A(net1311),
    .Y(net1313));
 BUFx2_ASAP7_75t_R rebuffer909 (.A(net1310),
    .Y(net1314));
 BUFx3_ASAP7_75t_R rebuffer910 (.A(net1314),
    .Y(net1315));
 BUFx2_ASAP7_75t_R rebuffer911 (.A(net3332),
    .Y(net1316));
 BUFx2_ASAP7_75t_R rebuffer912 (.A(net1316),
    .Y(net1317));
 BUFx6f_ASAP7_75t_R split913 (.A(net1581),
    .Y(net1318));
 BUFx12f_ASAP7_75t_R rebuffer914 (.A(_00623_),
    .Y(net1319));
 BUFx2_ASAP7_75t_R rebuffer915 (.A(net3438),
    .Y(net1320));
 BUFx2_ASAP7_75t_R rebuffer916 (.A(net3438),
    .Y(net1321));
 BUFx2_ASAP7_75t_R rebuffer917 (.A(net3438),
    .Y(net1322));
 BUFx2_ASAP7_75t_R rebuffer918 (.A(net1319),
    .Y(net1323));
 BUFx2_ASAP7_75t_R rebuffer919 (.A(net1323),
    .Y(net1324));
 BUFx2_ASAP7_75t_R rebuffer920 (.A(net1323),
    .Y(net1325));
 BUFx6f_ASAP7_75t_R rebuffer921 (.A(_00623_),
    .Y(net1326));
 BUFx12f_ASAP7_75t_R rebuffer922 (.A(_01124_),
    .Y(net1327));
 BUFx2_ASAP7_75t_R rebuffer923 (.A(net1327),
    .Y(net1328));
 BUFx2_ASAP7_75t_R rebuffer924 (.A(net1327),
    .Y(net1329));
 BUFx2_ASAP7_75t_R rebuffer925 (.A(net1329),
    .Y(net1330));
 BUFx2_ASAP7_75t_R rebuffer926 (.A(net1330),
    .Y(net1331));
 BUFx2_ASAP7_75t_R rebuffer927 (.A(net1329),
    .Y(net1332));
 BUFx2_ASAP7_75t_R rebuffer928 (.A(net1332),
    .Y(net1333));
 BUFx2_ASAP7_75t_R rebuffer929 (.A(_01124_),
    .Y(net1334));
 BUFx6f_ASAP7_75t_R split930 (.A(_18411_),
    .Y(net1335));
 BUFx6f_ASAP7_75t_R rebuffer931 (.A(_10618_),
    .Y(net1336));
 BUFx2_ASAP7_75t_R rebuffer932 (.A(net1336),
    .Y(net1337));
 BUFx12f_ASAP7_75t_R rebuffer933 (.A(_10618_),
    .Y(net1338));
 BUFx2_ASAP7_75t_R rebuffer934 (.A(net1338),
    .Y(net1339));
 BUFx3_ASAP7_75t_R rebuffer935 (.A(net1339),
    .Y(net1340));
 BUFx6f_ASAP7_75t_R split936 (.A(_00591_),
    .Y(net1341));
 BUFx4f_ASAP7_75t_R rebuffer937 (.A(net2147),
    .Y(net1342));
 BUFx2_ASAP7_75t_R rebuffer938 (.A(_10650_),
    .Y(net1343));
 BUFx3_ASAP7_75t_R rebuffer939 (.A(net1343),
    .Y(net1344));
 BUFx2_ASAP7_75t_R rebuffer940 (.A(net1344),
    .Y(net1345));
 BUFx2_ASAP7_75t_R rebuffer941 (.A(net1344),
    .Y(net1346));
 BUFx2_ASAP7_75t_R rebuffer942 (.A(net1343),
    .Y(net1347));
 BUFx4f_ASAP7_75t_R rebuffer943 (.A(_17956_),
    .Y(net1348));
 BUFx2_ASAP7_75t_R rebuffer944 (.A(net1348),
    .Y(net1349));
 BUFx2_ASAP7_75t_R rebuffer945 (.A(net1348),
    .Y(net1350));
 BUFx2_ASAP7_75t_R rebuffer946 (.A(_09904_),
    .Y(net1351));
 BUFx2_ASAP7_75t_R rebuffer947 (.A(net1351),
    .Y(net1352));
 BUFx12f_ASAP7_75t_R rebuffer948 (.A(_09904_),
    .Y(net1353));
 BUFx4f_ASAP7_75t_R rebuffer949 (.A(_09904_),
    .Y(net1354));
 BUFx4f_ASAP7_75t_R rebuffer950 (.A(net1354),
    .Y(net1355));
 BUFx2_ASAP7_75t_R rebuffer951 (.A(net1355),
    .Y(net1356));
 BUFx2_ASAP7_75t_R rebuffer952 (.A(_00599_),
    .Y(net1357));
 BUFx6f_ASAP7_75t_R rebuffer953 (.A(_00599_),
    .Y(net1358));
 BUFx3_ASAP7_75t_R rebuffer954 (.A(net1358),
    .Y(net1359));
 BUFx2_ASAP7_75t_R rebuffer955 (.A(net1359),
    .Y(net1360));
 BUFx2_ASAP7_75t_R rebuffer956 (.A(net1359),
    .Y(net1361));
 BUFx2_ASAP7_75t_R rebuffer957 (.A(net1361),
    .Y(net1362));
 BUFx3_ASAP7_75t_R rebuffer958 (.A(_00599_),
    .Y(net1363));
 BUFx2_ASAP7_75t_R rebuffer959 (.A(net1363),
    .Y(net1364));
 BUFx12f_ASAP7_75t_R rebuffer960 (.A(_17924_),
    .Y(net1365));
 BUFx2_ASAP7_75t_R rebuffer961 (.A(net1365),
    .Y(net1366));
 BUFx2_ASAP7_75t_R rebuffer962 (.A(net1365),
    .Y(net1367));
 BUFx2_ASAP7_75t_R rebuffer963 (.A(net1365),
    .Y(net1368));
 BUFx3_ASAP7_75t_R rebuffer964 (.A(net1368),
    .Y(net1369));
 BUFx2_ASAP7_75t_R rebuffer965 (.A(net1365),
    .Y(net1370));
 BUFx2_ASAP7_75t_R rebuffer966 (.A(_17924_),
    .Y(net1371));
 BUFx2_ASAP7_75t_R rebuffer967 (.A(_00575_),
    .Y(net1372));
 BUFx2_ASAP7_75t_R rebuffer968 (.A(_00575_),
    .Y(net1373));
 BUFx12f_ASAP7_75t_R rebuffer969 (.A(_00575_),
    .Y(net1374));
 BUFx2_ASAP7_75t_R rebuffer970 (.A(net3084),
    .Y(net1375));
 BUFx2_ASAP7_75t_R rebuffer971 (.A(net3084),
    .Y(net1376));
 BUFx2_ASAP7_75t_R rebuffer972 (.A(net3084),
    .Y(net1377));
 BUFx2_ASAP7_75t_R rebuffer973 (.A(net1377),
    .Y(net1378));
 BUFx2_ASAP7_75t_R rebuffer974 (.A(net3084),
    .Y(net1379));
 BUFx6f_ASAP7_75t_R rebuffer975 (.A(_17563_),
    .Y(net1380));
 BUFx6f_ASAP7_75t_R rebuffer976 (.A(_17563_),
    .Y(net1381));
 BUFx2_ASAP7_75t_R rebuffer977 (.A(net1381),
    .Y(net1382));
 BUFx2_ASAP7_75t_R rebuffer978 (.A(net1381),
    .Y(net1383));
 BUFx6f_ASAP7_75t_R rebuffer979 (.A(_09684_),
    .Y(net1384));
 BUFx6f_ASAP7_75t_R rebuffer980 (.A(_09684_),
    .Y(net1385));
 BUFx2_ASAP7_75t_R rebuffer981 (.A(net1385),
    .Y(net1386));
 BUFx6f_ASAP7_75t_R split982 (.A(_09711_),
    .Y(net1387));
 BUFx6f_ASAP7_75t_R split983 (.A(_18594_),
    .Y(net1388));
 BUFx3_ASAP7_75t_R rebuffer984 (.A(_00608_),
    .Y(net1389));
 BUFx2_ASAP7_75t_R rebuffer985 (.A(net1389),
    .Y(net1390));
 BUFx2_ASAP7_75t_R rebuffer986 (.A(net1389),
    .Y(net1391));
 BUFx2_ASAP7_75t_R rebuffer987 (.A(net1391),
    .Y(net1392));
 BUFx12f_ASAP7_75t_R rebuffer988 (.A(_00608_),
    .Y(net1393));
 BUFx2_ASAP7_75t_R rebuffer989 (.A(net1393),
    .Y(net1394));
 BUFx12f_ASAP7_75t_R rebuffer990 (.A(net1393),
    .Y(net1395));
 BUFx2_ASAP7_75t_R rebuffer991 (.A(net2990),
    .Y(net1396));
 BUFx4f_ASAP7_75t_R rebuffer992 (.A(net1393),
    .Y(net1397));
 BUFx2_ASAP7_75t_R rebuffer993 (.A(net2990),
    .Y(net1398));
 BUFx2_ASAP7_75t_R rebuffer994 (.A(_01555_),
    .Y(net1399));
 BUFx2_ASAP7_75t_R rebuffer995 (.A(net1399),
    .Y(net1400));
 BUFx3_ASAP7_75t_R rebuffer996 (.A(_05105_),
    .Y(net1401));
 BUFx3_ASAP7_75t_R rebuffer997 (.A(net1401),
    .Y(net1402));
 BUFx6f_ASAP7_75t_R rebuffer998 (.A(_05105_),
    .Y(net1403));
 BUFx10_ASAP7_75t_R split999 (.A(_18575_),
    .Y(net1404));
 BUFx2_ASAP7_75t_R rebuffer1000 (.A(_00551_),
    .Y(net1405));
 BUFx4f_ASAP7_75t_R rebuffer1001 (.A(_00551_),
    .Y(net1406));
 BUFx12f_ASAP7_75t_R rebuffer1002 (.A(_00551_),
    .Y(net1407));
 BUFx2_ASAP7_75t_R rebuffer1003 (.A(net1407),
    .Y(net1408));
 BUFx2_ASAP7_75t_R rebuffer1004 (.A(net1407),
    .Y(net1409));
 BUFx2_ASAP7_75t_R rebuffer1005 (.A(net1407),
    .Y(net1410));
 BUFx6f_ASAP7_75t_R rebuffer1006 (.A(net1407),
    .Y(net1411));
 BUFx2_ASAP7_75t_R rebuffer1007 (.A(net1407),
    .Y(net1412));
 BUFx4f_ASAP7_75t_R split1008 (.A(_01815_),
    .Y(net1413));
 BUFx6f_ASAP7_75t_R split1009 (.A(_10370_),
    .Y(net1414));
 BUFx3_ASAP7_75t_R rebuffer1010 (.A(_00536_),
    .Y(net1415));
 BUFx12f_ASAP7_75t_R rebuffer1011 (.A(_00536_),
    .Y(net1416));
 BUFx2_ASAP7_75t_R rebuffer1012 (.A(net1416),
    .Y(net1417));
 BUFx2_ASAP7_75t_R rebuffer1013 (.A(net1417),
    .Y(net1418));
 BUFx2_ASAP7_75t_R rebuffer1014 (.A(net1418),
    .Y(net1419));
 BUFx3_ASAP7_75t_R rebuffer1015 (.A(net1418),
    .Y(net1420));
 BUFx2_ASAP7_75t_R rebuffer1016 (.A(_00536_),
    .Y(net1421));
 BUFx2_ASAP7_75t_R rebuffer1017 (.A(net1421),
    .Y(net1422));
 BUFx2_ASAP7_75t_R rebuffer1018 (.A(net1422),
    .Y(net1423));
 BUFx2_ASAP7_75t_R rebuffer1019 (.A(net1423),
    .Y(net1424));
 BUFx2_ASAP7_75t_R rebuffer1020 (.A(net1421),
    .Y(net1425));
 BUFx6f_ASAP7_75t_R rebuffer1021 (.A(_01108_),
    .Y(net1426));
 BUFx6f_ASAP7_75t_R rebuffer1022 (.A(net1426),
    .Y(net1427));
 BUFx2_ASAP7_75t_R rebuffer1023 (.A(net1427),
    .Y(net1428));
 BUFx2_ASAP7_75t_R rebuffer1024 (.A(net1427),
    .Y(net1429));
 BUFx3_ASAP7_75t_R rebuffer1025 (.A(net1426),
    .Y(net1430));
 BUFx2_ASAP7_75t_R rebuffer1026 (.A(_01108_),
    .Y(net1431));
 BUFx2_ASAP7_75t_R rebuffer1027 (.A(net1431),
    .Y(net1432));
 BUFx2_ASAP7_75t_R rebuffer1028 (.A(net1431),
    .Y(net1433));
 BUFx6f_ASAP7_75t_R rebuffer1029 (.A(_13264_),
    .Y(net1434));
 BUFx2_ASAP7_75t_R rebuffer1030 (.A(net1434),
    .Y(net1435));
 BUFx2_ASAP7_75t_R rebuffer1031 (.A(net1434),
    .Y(net1436));
 BUFx3_ASAP7_75t_R rebuffer1032 (.A(net1434),
    .Y(net1437));
 BUFx2_ASAP7_75t_R rebuffer1033 (.A(net2569),
    .Y(net1438));
 BUFx2_ASAP7_75t_R rebuffer1034 (.A(net2569),
    .Y(net1439));
 BUFx2_ASAP7_75t_R rebuffer1035 (.A(net1439),
    .Y(net1440));
 BUFx2_ASAP7_75t_R rebuffer1036 (.A(net1440),
    .Y(net1441));
 BUFx2_ASAP7_75t_R rebuffer1037 (.A(net1880),
    .Y(net1442));
 BUFx2_ASAP7_75t_R rebuffer1038 (.A(net1880),
    .Y(net1443));
 BUFx2_ASAP7_75t_R rebuffer1039 (.A(net1880),
    .Y(net1444));
 BUFx2_ASAP7_75t_R rebuffer1040 (.A(net1444),
    .Y(net1445));
 BUFx6f_ASAP7_75t_R split1041 (.A(_10757_),
    .Y(net1446));
 BUFx12f_ASAP7_75t_R rebuffer1042 (.A(_00600_),
    .Y(net1447));
 BUFx3_ASAP7_75t_R rebuffer1043 (.A(net1447),
    .Y(net1448));
 BUFx2_ASAP7_75t_R rebuffer1044 (.A(net1448),
    .Y(net1449));
 BUFx2_ASAP7_75t_R rebuffer1045 (.A(net1449),
    .Y(net1450));
 BUFx2_ASAP7_75t_R rebuffer1046 (.A(net1448),
    .Y(net1451));
 BUFx2_ASAP7_75t_R rebuffer1047 (.A(net1451),
    .Y(net1452));
 BUFx2_ASAP7_75t_R rebuffer1048 (.A(net1451),
    .Y(net1453));
 BUFx12f_ASAP7_75t_R rebuffer1049 (.A(net1447),
    .Y(net1454));
 BUFx2_ASAP7_75t_R rebuffer1050 (.A(net1454),
    .Y(net1455));
 BUFx2_ASAP7_75t_R rebuffer1051 (.A(net1454),
    .Y(net1456));
 BUFx6f_ASAP7_75t_R split1052 (.A(_01612_),
    .Y(net1457));
 BUFx2_ASAP7_75t_R split1053 (.A(_01825_),
    .Y(net1458));
 BUFx2_ASAP7_75t_R rebuffer1054 (.A(_01773_),
    .Y(net1459));
 BUFx2_ASAP7_75t_R rebuffer1055 (.A(net1459),
    .Y(net1460));
 BUFx2_ASAP7_75t_R rebuffer1056 (.A(net1459),
    .Y(net1461));
 BUFx2_ASAP7_75t_R rebuffer1057 (.A(net2299),
    .Y(net1462));
 BUFx2_ASAP7_75t_R rebuffer1058 (.A(net2299),
    .Y(net1463));
 BUFx2_ASAP7_75t_R rebuffer1059 (.A(net1463),
    .Y(net1464));
 BUFx2_ASAP7_75t_R rebuffer1060 (.A(net2299),
    .Y(net1465));
 BUFx2_ASAP7_75t_R rebuffer1061 (.A(net1465),
    .Y(net1466));
 BUFx3_ASAP7_75t_R rebuffer1062 (.A(_00567_),
    .Y(net1467));
 BUFx2_ASAP7_75t_R rebuffer1063 (.A(net1467),
    .Y(net1468));
 BUFx3_ASAP7_75t_R rebuffer1064 (.A(_00567_),
    .Y(net1469));
 BUFx2_ASAP7_75t_R rebuffer1065 (.A(net1469),
    .Y(net1470));
 BUFx6f_ASAP7_75t_R rebuffer1066 (.A(_00567_),
    .Y(net1471));
 BUFx2_ASAP7_75t_R rebuffer1067 (.A(_00567_),
    .Y(net1472));
 BUFx2_ASAP7_75t_R rebuffer1068 (.A(net1472),
    .Y(net1473));
 BUFx2_ASAP7_75t_R rebuffer1069 (.A(_00567_),
    .Y(net1474));
 BUFx6f_ASAP7_75t_R split1070 (.A(_10771_),
    .Y(net1475));
 BUFx16f_ASAP7_75t_R rebuffer1071 (.A(_09579_),
    .Y(net1476));
 BUFx2_ASAP7_75t_R rebuffer1072 (.A(net1476),
    .Y(net1477));
 BUFx2_ASAP7_75t_R rebuffer1073 (.A(net1477),
    .Y(net1478));
 BUFx2_ASAP7_75t_R rebuffer1074 (.A(net1477),
    .Y(net1479));
 BUFx2_ASAP7_75t_R rebuffer1075 (.A(_09579_),
    .Y(net1480));
 BUFx2_ASAP7_75t_R rebuffer1076 (.A(_09579_),
    .Y(net1481));
 BUFx4f_ASAP7_75t_R rebuffer1077 (.A(_18296_),
    .Y(net1482));
 BUFx6f_ASAP7_75t_R rebuffer1078 (.A(_18296_),
    .Y(net1483));
 BUFx2_ASAP7_75t_R rebuffer1079 (.A(net1483),
    .Y(net1484));
 BUFx12f_ASAP7_75t_R rebuffer1080 (.A(_05056_),
    .Y(net1485));
 BUFx2_ASAP7_75t_R rebuffer1081 (.A(net1485),
    .Y(net1486));
 BUFx2_ASAP7_75t_R rebuffer1082 (.A(net1485),
    .Y(net1487));
 BUFx2_ASAP7_75t_R rebuffer1083 (.A(_05056_),
    .Y(net1488));
 BUFx2_ASAP7_75t_R rebuffer1084 (.A(net1488),
    .Y(net1489));
 BUFx3_ASAP7_75t_R rebuffer1085 (.A(_05056_),
    .Y(net1490));
 BUFx2_ASAP7_75t_R rebuffer1086 (.A(net1490),
    .Y(net1491));
 BUFx6f_ASAP7_75t_R split1087 (.A(_10759_),
    .Y(net1492));
 BUFx6f_ASAP7_75t_R rebuffer1088 (.A(_09628_),
    .Y(net1493));
 BUFx4f_ASAP7_75t_R split1089 (.A(_10365_),
    .Y(net1494));
 BUFx2_ASAP7_75t_R rebuffer1090 (.A(net1885),
    .Y(net1495));
 BUFx2_ASAP7_75t_R rebuffer1091 (.A(net1495),
    .Y(net1496));
 BUFx3_ASAP7_75t_R rebuffer1092 (.A(_10343_),
    .Y(net1497));
 BUFx2_ASAP7_75t_R rebuffer1093 (.A(net1497),
    .Y(net1498));
 BUFx2_ASAP7_75t_R rebuffer1094 (.A(net1497),
    .Y(net1499));
 BUFx2_ASAP7_75t_R rebuffer1095 (.A(net1885),
    .Y(net1500));
 BUFx6f_ASAP7_75t_R split1096 (.A(net1715),
    .Y(net1501));
 BUFx3_ASAP7_75t_R rebuffer1097 (.A(_09748_),
    .Y(net1502));
 BUFx2_ASAP7_75t_R rebuffer1098 (.A(net1502),
    .Y(net1503));
 BUFx6f_ASAP7_75t_R rebuffer1099 (.A(net1502),
    .Y(net1504));
 BUFx2_ASAP7_75t_R rebuffer1100 (.A(net1504),
    .Y(net1505));
 BUFx2_ASAP7_75t_R rebuffer1101 (.A(net1502),
    .Y(net1506));
 BUFx6f_ASAP7_75t_R rebuffer1102 (.A(_09748_),
    .Y(net1507));
 BUFx2_ASAP7_75t_R rebuffer1103 (.A(net1507),
    .Y(net1508));
 BUFx2_ASAP7_75t_R rebuffer1104 (.A(net1507),
    .Y(net1509));
 BUFx2_ASAP7_75t_R rebuffer1105 (.A(_10312_),
    .Y(net1510));
 BUFx2_ASAP7_75t_R rebuffer1106 (.A(net1510),
    .Y(net1511));
 BUFx2_ASAP7_75t_R rebuffer1107 (.A(_10312_),
    .Y(net1512));
 BUFx2_ASAP7_75t_R rebuffer1108 (.A(_10312_),
    .Y(net1513));
 BUFx2_ASAP7_75t_R rebuffer1109 (.A(net1513),
    .Y(net1514));
 BUFx6f_ASAP7_75t_R rebuffer1110 (.A(net1514),
    .Y(net1515));
 BUFx2_ASAP7_75t_R rebuffer1111 (.A(_10312_),
    .Y(net1516));
 BUFx2_ASAP7_75t_R rebuffer1112 (.A(net1516),
    .Y(net1517));
 BUFx3_ASAP7_75t_R rebuffer1113 (.A(_09738_),
    .Y(net1518));
 BUFx3_ASAP7_75t_R rebuffer1114 (.A(net1518),
    .Y(net1519));
 BUFx2_ASAP7_75t_R rebuffer1115 (.A(_05083_),
    .Y(net1520));
 BUFx2_ASAP7_75t_R rebuffer1116 (.A(_05083_),
    .Y(net1521));
 BUFx2_ASAP7_75t_R rebuffer1117 (.A(_05083_),
    .Y(net1522));
 BUFx2_ASAP7_75t_R rebuffer1118 (.A(net1522),
    .Y(net1523));
 BUFx2_ASAP7_75t_R rebuffer1119 (.A(_05083_),
    .Y(net1524));
 BUFx3_ASAP7_75t_R rebuffer1120 (.A(net1524),
    .Y(net1525));
 BUFx2_ASAP7_75t_R rebuffer1121 (.A(net1524),
    .Y(net1526));
 BUFx6f_ASAP7_75t_R split1122 (.A(_01824_),
    .Y(net1527));
 BUFx6f_ASAP7_75t_R split1123 (.A(_05561_),
    .Y(net1528));
 BUFx3_ASAP7_75t_R rebuffer1124 (.A(net2824),
    .Y(net1529));
 BUFx6f_ASAP7_75t_R rebuffer1125 (.A(_17963_),
    .Y(net1530));
 BUFx2_ASAP7_75t_R rebuffer1126 (.A(net1530),
    .Y(net1531));
 BUFx3_ASAP7_75t_R rebuffer1127 (.A(net1530),
    .Y(net1532));
 BUFx2_ASAP7_75t_R rebuffer1128 (.A(_00559_),
    .Y(net1533));
 BUFx2_ASAP7_75t_R rebuffer1129 (.A(_00559_),
    .Y(net1534));
 BUFx6f_ASAP7_75t_R rebuffer1130 (.A(_00559_),
    .Y(net1535));
 BUFx3_ASAP7_75t_R rebuffer1131 (.A(net1535),
    .Y(net1536));
 BUFx12f_ASAP7_75t_R rebuffer1132 (.A(net1535),
    .Y(net1537));
 BUFx2_ASAP7_75t_R rebuffer1133 (.A(net1537),
    .Y(net1538));
 BUFx2_ASAP7_75t_R rebuffer1134 (.A(net1535),
    .Y(net1539));
 BUFx2_ASAP7_75t_R rebuffer1135 (.A(_06118_),
    .Y(net1540));
 BUFx2_ASAP7_75t_R rebuffer1136 (.A(_06118_),
    .Y(net1541));
 BUFx2_ASAP7_75t_R rebuffer1137 (.A(_17936_),
    .Y(net1542));
 BUFx2_ASAP7_75t_R rebuffer1138 (.A(_17936_),
    .Y(net1543));
 BUFx3_ASAP7_75t_R split1139 (.A(_09636_),
    .Y(net1544));
 BUFx3_ASAP7_75t_R rebuffer1140 (.A(_00632_),
    .Y(net1545));
 BUFx2_ASAP7_75t_R rebuffer1141 (.A(net1545),
    .Y(net1546));
 BUFx2_ASAP7_75t_R rebuffer1142 (.A(net1545),
    .Y(net1547));
 BUFx2_ASAP7_75t_R rebuffer1143 (.A(net1545),
    .Y(net1548));
 BUFx2_ASAP7_75t_R rebuffer1144 (.A(net1545),
    .Y(net1549));
 BUFx12f_ASAP7_75t_R rebuffer1145 (.A(_00632_),
    .Y(net1550));
 BUFx2_ASAP7_75t_R rebuffer1146 (.A(net1550),
    .Y(net1551));
 BUFx2_ASAP7_75t_R rebuffer1147 (.A(net1550),
    .Y(net1552));
 BUFx2_ASAP7_75t_R rebuffer1148 (.A(_01788_),
    .Y(net1553));
 BUFx2_ASAP7_75t_R rebuffer1149 (.A(_01788_),
    .Y(net1554));
 BUFx2_ASAP7_75t_R rebuffer1150 (.A(net1554),
    .Y(net1555));
 BUFx12f_ASAP7_75t_R rebuffer1151 (.A(_01788_),
    .Y(net1556));
 BUFx2_ASAP7_75t_R rebuffer1152 (.A(net1556),
    .Y(net1557));
 BUFx2_ASAP7_75t_R rebuffer1153 (.A(net1556),
    .Y(net1558));
 BUFx2_ASAP7_75t_R rebuffer1154 (.A(net1558),
    .Y(net1559));
 BUFx6f_ASAP7_75t_R split1155 (.A(_05796_),
    .Y(net1560));
 BUFx3_ASAP7_75t_R rebuffer1156 (.A(_09738_),
    .Y(net1561));
 BUFx3_ASAP7_75t_R split1157 (.A(_09738_),
    .Y(net1562));
 BUFx6f_ASAP7_75t_R rebuffer1158 (.A(_18540_),
    .Y(net1563));
 BUFx2_ASAP7_75t_R rebuffer1159 (.A(net1563),
    .Y(net1564));
 BUFx4f_ASAP7_75t_R rebuffer1160 (.A(_18540_),
    .Y(net1565));
 BUFx2_ASAP7_75t_R rebuffer1161 (.A(net1565),
    .Y(net1566));
 BUFx2_ASAP7_75t_R rebuffer1162 (.A(net1566),
    .Y(net1567));
 BUFx2_ASAP7_75t_R rebuffer1163 (.A(net1565),
    .Y(net1568));
 BUFx2_ASAP7_75t_R rebuffer1164 (.A(net1568),
    .Y(net1569));
 BUFx2_ASAP7_75t_R rebuffer1165 (.A(net1568),
    .Y(net1570));
 BUFx2_ASAP7_75t_R rebuffer1166 (.A(net1565),
    .Y(net1571));
 BUFx6f_ASAP7_75t_R split1167 (.A(_01125_),
    .Y(net1572));
 BUFx2_ASAP7_75t_R rebuffer1168 (.A(_01491_),
    .Y(net1573));
 BUFx2_ASAP7_75t_R rebuffer1169 (.A(_01491_),
    .Y(net1574));
 BUFx6f_ASAP7_75t_R rebuffer1170 (.A(_01491_),
    .Y(net1575));
 BUFx2_ASAP7_75t_R rebuffer1171 (.A(net1575),
    .Y(net1576));
 BUFx4f_ASAP7_75t_R split1172 (.A(_09592_),
    .Y(net1577));
 BUFx2_ASAP7_75t_R rebuffer1173 (.A(_18268_),
    .Y(net1578));
 BUFx2_ASAP7_75t_R rebuffer1174 (.A(net2093),
    .Y(net1579));
 BUFx2_ASAP7_75t_R rebuffer1175 (.A(net2825),
    .Y(net1580));
 BUFx2_ASAP7_75t_R rebuffer1176 (.A(_00576_),
    .Y(net1581));
 BUFx12f_ASAP7_75t_R rebuffer1177 (.A(_00576_),
    .Y(net1582));
 BUFx2_ASAP7_75t_R rebuffer1178 (.A(net1582),
    .Y(net1583));
 BUFx2_ASAP7_75t_R rebuffer1179 (.A(_00576_),
    .Y(net1584));
 BUFx2_ASAP7_75t_R rebuffer1180 (.A(net1584),
    .Y(net1585));
 BUFx2_ASAP7_75t_R rebuffer1181 (.A(net1585),
    .Y(net1586));
 BUFx2_ASAP7_75t_R rebuffer1182 (.A(_09798_),
    .Y(net1587));
 BUFx2_ASAP7_75t_R rebuffer1183 (.A(_06063_),
    .Y(net1588));
 BUFx2_ASAP7_75t_R rebuffer1184 (.A(net1588),
    .Y(net1589));
 BUFx2_ASAP7_75t_R rebuffer1185 (.A(net1588),
    .Y(net1590));
 BUFx2_ASAP7_75t_R rebuffer1186 (.A(_06063_),
    .Y(net1591));
 BUFx6f_ASAP7_75t_R rebuffer1187 (.A(net1591),
    .Y(net1592));
 BUFx12f_ASAP7_75t_R rebuffer1188 (.A(_00591_),
    .Y(net1593));
 BUFx6f_ASAP7_75t_R rebuffer1189 (.A(_00591_),
    .Y(net1594));
 BUFx2_ASAP7_75t_R rebuffer1190 (.A(net1594),
    .Y(net1595));
 BUFx2_ASAP7_75t_R split1191 (.A(_09752_),
    .Y(net1596));
 BUFx6f_ASAP7_75t_R split1192 (.A(_01590_),
    .Y(net1597));
 BUFx3_ASAP7_75t_R rebuffer1193 (.A(_06034_),
    .Y(net1598));
 BUFx2_ASAP7_75t_R rebuffer1194 (.A(net1598),
    .Y(net1599));
 BUFx2_ASAP7_75t_R rebuffer1195 (.A(net1598),
    .Y(net1600));
 BUFx3_ASAP7_75t_R rebuffer1196 (.A(_06034_),
    .Y(net1601));
 BUFx2_ASAP7_75t_R rebuffer1197 (.A(net1601),
    .Y(net1602));
 BUFx6f_ASAP7_75t_R rebuffer1198 (.A(_06052_),
    .Y(net1603));
 BUFx2_ASAP7_75t_R rebuffer1199 (.A(net1603),
    .Y(net1604));
 BUFx6f_ASAP7_75t_R split1200 (.A(_02361_),
    .Y(net1605));
 BUFx6f_ASAP7_75t_R split1201 (.A(_19171_),
    .Y(net1606));
 BUFx12f_ASAP7_75t_R rebuffer1202 (.A(_17570_),
    .Y(net1607));
 BUFx2_ASAP7_75t_R rebuffer1203 (.A(net1607),
    .Y(net1608));
 BUFx3_ASAP7_75t_R rebuffer1204 (.A(net1607),
    .Y(net1609));
 BUFx2_ASAP7_75t_R rebuffer1205 (.A(net1609),
    .Y(net1610));
 BUFx2_ASAP7_75t_R rebuffer1206 (.A(net1607),
    .Y(net1611));
 BUFx6f_ASAP7_75t_R split1207 (.A(_01556_),
    .Y(net1612));
 BUFx6f_ASAP7_75t_R split1208 (.A(_01553_),
    .Y(net1613));
 BUFx6f_ASAP7_75t_R rebuffer1209 (.A(_00427_),
    .Y(net1614));
 BUFx2_ASAP7_75t_R rebuffer1210 (.A(net1614),
    .Y(net1615));
 BUFx2_ASAP7_75t_R rebuffer1211 (.A(net1615),
    .Y(net1616));
 BUFx2_ASAP7_75t_R rebuffer1212 (.A(net1616),
    .Y(net1617));
 BUFx2_ASAP7_75t_R rebuffer1213 (.A(net1614),
    .Y(net1618));
 BUFx2_ASAP7_75t_R rebuffer1214 (.A(net1614),
    .Y(net1619));
 BUFx2_ASAP7_75t_R rebuffer1215 (.A(net1614),
    .Y(net1620));
 BUFx2_ASAP7_75t_R rebuffer1216 (.A(_00427_),
    .Y(net1621));
 BUFx6f_ASAP7_75t_R rebuffer1217 (.A(_17958_),
    .Y(net1622));
 BUFx2_ASAP7_75t_R rebuffer1218 (.A(net1622),
    .Y(net1623));
 BUFx2_ASAP7_75t_R rebuffer1219 (.A(_17958_),
    .Y(net1624));
 BUFx6f_ASAP7_75t_R rebuffer1220 (.A(_00613_),
    .Y(net1625));
 BUFx2_ASAP7_75t_R rebuffer1221 (.A(net1625),
    .Y(net1626));
 BUFx6f_ASAP7_75t_R split1222 (.A(_05535_),
    .Y(net1627));
 BUFx2_ASAP7_75t_R rebuffer1223 (.A(_06137_),
    .Y(net1628));
 BUFx2_ASAP7_75t_R rebuffer1224 (.A(_21922_),
    .Y(net1629));
 BUFx3_ASAP7_75t_R rebuffer1225 (.A(_21922_),
    .Y(net1630));
 BUFx2_ASAP7_75t_R rebuffer1226 (.A(net1630),
    .Y(net1631));
 BUFx2_ASAP7_75t_R rebuffer1227 (.A(net1630),
    .Y(net1632));
 BUFx2_ASAP7_75t_R rebuffer1228 (.A(net1630),
    .Y(net1633));
 BUFx2_ASAP7_75t_R rebuffer1229 (.A(net1630),
    .Y(net1634));
 BUFx12f_ASAP7_75t_R rebuffer1230 (.A(_00639_),
    .Y(net1635));
 BUFx2_ASAP7_75t_R rebuffer1231 (.A(net1635),
    .Y(net1636));
 BUFx6f_ASAP7_75t_R rebuffer1232 (.A(net1635),
    .Y(net1637));
 BUFx2_ASAP7_75t_R rebuffer1233 (.A(net1635),
    .Y(net1638));
 BUFx2_ASAP7_75t_R rebuffer1234 (.A(net1638),
    .Y(net1639));
 BUFx2_ASAP7_75t_R rebuffer1235 (.A(net1638),
    .Y(net1640));
 BUFx2_ASAP7_75t_R rebuffer1236 (.A(net1635),
    .Y(net1641));
 BUFx2_ASAP7_75t_R rebuffer1237 (.A(_00648_),
    .Y(net1642));
 BUFx6f_ASAP7_75t_R rebuffer1238 (.A(_00648_),
    .Y(net1643));
 BUFx2_ASAP7_75t_R rebuffer1239 (.A(net1643),
    .Y(net1644));
 BUFx3_ASAP7_75t_R rebuffer1240 (.A(net1644),
    .Y(net1645));
 BUFx2_ASAP7_75t_R rebuffer1241 (.A(net1643),
    .Y(net1646));
 BUFx6f_ASAP7_75t_R rebuffer1242 (.A(_00648_),
    .Y(net1647));
 BUFx3_ASAP7_75t_R rebuffer1243 (.A(_21889_),
    .Y(net1648));
 BUFx2_ASAP7_75t_R rebuffer1244 (.A(net1648),
    .Y(net1649));
 BUFx2_ASAP7_75t_R rebuffer1245 (.A(net1649),
    .Y(net1650));
 BUFx6f_ASAP7_75t_R rebuffer1246 (.A(_21889_),
    .Y(net1651));
 BUFx2_ASAP7_75t_R rebuffer1247 (.A(net1651),
    .Y(net1652));
 BUFx2_ASAP7_75t_R rebuffer1248 (.A(_05903_),
    .Y(net1653));
 BUFx8_ASAP7_75t_R rebuffer1249 (.A(_05903_),
    .Y(net1654));
 BUFx6f_ASAP7_75t_R rebuffer1250 (.A(net1654),
    .Y(net1655));
 BUFx2_ASAP7_75t_R rebuffer1251 (.A(net1655),
    .Y(net1656));
 BUFx2_ASAP7_75t_R rebuffer1252 (.A(net1654),
    .Y(net1657));
 BUFx2_ASAP7_75t_R rebuffer1253 (.A(_05903_),
    .Y(net1658));
 BUFx6f_ASAP7_75t_R split1254 (.A(_10329_),
    .Y(net1659));
 BUFx12f_ASAP7_75t_R rebuffer1255 (.A(_09919_),
    .Y(net1660));
 BUFx6f_ASAP7_75t_R split1256 (.A(_09919_),
    .Y(net1661));
 BUFx6f_ASAP7_75t_R split1257 (.A(_05767_),
    .Y(net1662));
 BUFx2_ASAP7_75t_R rebuffer1258 (.A(_06058_),
    .Y(net1663));
 BUFx2_ASAP7_75t_R rebuffer1259 (.A(net1663),
    .Y(net1664));
 BUFx2_ASAP7_75t_R rebuffer1260 (.A(net1663),
    .Y(net1665));
 BUFx12f_ASAP7_75t_R rebuffer1261 (.A(_05560_),
    .Y(net1666));
 BUFx2_ASAP7_75t_R rebuffer1262 (.A(net1666),
    .Y(net1667));
 BUFx2_ASAP7_75t_R rebuffer1263 (.A(net1666),
    .Y(net1668));
 BUFx2_ASAP7_75t_R rebuffer1264 (.A(net1666),
    .Y(net1669));
 BUFx2_ASAP7_75t_R rebuffer1265 (.A(net1666),
    .Y(net1670));
 BUFx2_ASAP7_75t_R rebuffer1266 (.A(net1670),
    .Y(net1671));
 BUFx2_ASAP7_75t_R rebuffer1267 (.A(net1666),
    .Y(net1672));
 BUFx2_ASAP7_75t_R rebuffer1268 (.A(_05560_),
    .Y(net1673));
 BUFx2_ASAP7_75t_R rebuffer1269 (.A(net1673),
    .Y(net1674));
 BUFx6f_ASAP7_75t_R rebuffer1270 (.A(_17938_),
    .Y(net1675));
 BUFx2_ASAP7_75t_R rebuffer1271 (.A(net1675),
    .Y(net1676));
 BUFx2_ASAP7_75t_R rebuffer1272 (.A(net3000),
    .Y(net1677));
 BUFx12f_ASAP7_75t_R rebuffer1273 (.A(_00607_),
    .Y(net1678));
 BUFx2_ASAP7_75t_R rebuffer1274 (.A(net1678),
    .Y(net1679));
 BUFx3_ASAP7_75t_R rebuffer1275 (.A(_00607_),
    .Y(net1680));
 BUFx2_ASAP7_75t_R rebuffer1276 (.A(_00607_),
    .Y(net1681));
 BUFx2_ASAP7_75t_R rebuffer1277 (.A(_00592_),
    .Y(net1682));
 BUFx2_ASAP7_75t_R rebuffer1278 (.A(net1682),
    .Y(net1683));
 BUFx2_ASAP7_75t_R rebuffer1279 (.A(net1683),
    .Y(net1684));
 BUFx6f_ASAP7_75t_R rebuffer1280 (.A(net1684),
    .Y(net1685));
 BUFx12f_ASAP7_75t_R rebuffer1281 (.A(_00592_),
    .Y(net1686));
 BUFx2_ASAP7_75t_R rebuffer1282 (.A(net1686),
    .Y(net1687));
 BUFx2_ASAP7_75t_R rebuffer1283 (.A(net1686),
    .Y(net1688));
 BUFx2_ASAP7_75t_R rebuffer1284 (.A(net3307),
    .Y(net1689));
 BUFx6f_ASAP7_75t_R rebuffer1285 (.A(_17943_),
    .Y(net1690));
 BUFx2_ASAP7_75t_R rebuffer1286 (.A(net1690),
    .Y(net1691));
 BUFx2_ASAP7_75t_R rebuffer1287 (.A(net1690),
    .Y(net1692));
 BUFx2_ASAP7_75t_R rebuffer1288 (.A(_17943_),
    .Y(net1693));
 BUFx6f_ASAP7_75t_R rebuffer1289 (.A(_06449_),
    .Y(net1694));
 BUFx2_ASAP7_75t_R rebuffer1290 (.A(net1694),
    .Y(net1695));
 BUFx6f_ASAP7_75t_R rebuffer1291 (.A(_01148_),
    .Y(net1696));
 BUFx2_ASAP7_75t_R rebuffer1292 (.A(net1696),
    .Y(net1697));
 BUFx4f_ASAP7_75t_R rebuffer1293 (.A(_01148_),
    .Y(net1698));
 BUFx12f_ASAP7_75t_R rebuffer1294 (.A(_09887_),
    .Y(net1699));
 BUFx2_ASAP7_75t_R rebuffer1295 (.A(net1699),
    .Y(net1700));
 BUFx2_ASAP7_75t_R rebuffer1296 (.A(net1699),
    .Y(net1701));
 BUFx4f_ASAP7_75t_R rebuffer1297 (.A(_18254_),
    .Y(net1702));
 BUFx12f_ASAP7_75t_R rebuffer1298 (.A(_09958_),
    .Y(net1703));
 BUFx6f_ASAP7_75t_R rebuffer1299 (.A(net1703),
    .Y(net1704));
 BUFx2_ASAP7_75t_R rebuffer1300 (.A(net1704),
    .Y(net1705));
 BUFx2_ASAP7_75t_R rebuffer1301 (.A(net1703),
    .Y(net1706));
 BUFx2_ASAP7_75t_R rebuffer1302 (.A(net1703),
    .Y(net1707));
 BUFx2_ASAP7_75t_R rebuffer1303 (.A(_21873_),
    .Y(net1708));
 BUFx2_ASAP7_75t_R rebuffer1304 (.A(net1708),
    .Y(net1709));
 BUFx2_ASAP7_75t_R rebuffer1305 (.A(_21873_),
    .Y(net1710));
 BUFx2_ASAP7_75t_R rebuffer1306 (.A(_21873_),
    .Y(net1711));
 BUFx6f_ASAP7_75t_R rebuffer1307 (.A(_21873_),
    .Y(net1712));
 BUFx2_ASAP7_75t_R rebuffer1308 (.A(net1712),
    .Y(net1713));
 BUFx2_ASAP7_75t_R rebuffer1309 (.A(net1712),
    .Y(net1714));
 BUFx2_ASAP7_75t_R rebuffer1310 (.A(_00535_),
    .Y(net1715));
 BUFx12f_ASAP7_75t_R rebuffer1311 (.A(_00535_),
    .Y(net1716));
 BUFx2_ASAP7_75t_R rebuffer1312 (.A(net1716),
    .Y(net1717));
 BUFx2_ASAP7_75t_R rebuffer1313 (.A(net1716),
    .Y(net1718));
 BUFx6f_ASAP7_75t_R rebuffer1314 (.A(net1718),
    .Y(net1719));
 BUFx2_ASAP7_75t_R rebuffer1315 (.A(net1716),
    .Y(net1720));
 BUFx2_ASAP7_75t_R rebuffer1316 (.A(_00535_),
    .Y(net1721));
 BUFx3_ASAP7_75t_R rebuffer1317 (.A(_00614_),
    .Y(net1722));
 BUFx6f_ASAP7_75t_R rebuffer1318 (.A(_00614_),
    .Y(net1723));
 BUFx2_ASAP7_75t_R rebuffer1319 (.A(net1723),
    .Y(net1724));
 BUFx2_ASAP7_75t_R rebuffer1320 (.A(net1723),
    .Y(net1725));
 BUFx3_ASAP7_75t_R rebuffer1321 (.A(_18556_),
    .Y(net1726));
 BUFx2_ASAP7_75t_R rebuffer1322 (.A(net1726),
    .Y(net1727));
 BUFx6f_ASAP7_75t_R rebuffer1323 (.A(_18556_),
    .Y(net1728));
 BUFx2_ASAP7_75t_R rebuffer1324 (.A(net1728),
    .Y(net1729));
 BUFx2_ASAP7_75t_R rebuffer1325 (.A(net1728),
    .Y(net1730));
 BUFx6f_ASAP7_75t_R rebuffer1326 (.A(_00568_),
    .Y(net1731));
 BUFx2_ASAP7_75t_R rebuffer1327 (.A(net1731),
    .Y(net1732));
 BUFx2_ASAP7_75t_R rebuffer1328 (.A(net1732),
    .Y(net1733));
 BUFx2_ASAP7_75t_R rebuffer1329 (.A(net1731),
    .Y(net1734));
 BUFx6f_ASAP7_75t_R rebuffer1330 (.A(_00568_),
    .Y(net1735));
 BUFx2_ASAP7_75t_R rebuffer1331 (.A(net1735),
    .Y(net1736));
 BUFx2_ASAP7_75t_R rebuffer1332 (.A(net1735),
    .Y(net1737));
 BUFx2_ASAP7_75t_R rebuffer1333 (.A(net1735),
    .Y(net1738));
 BUFx16f_ASAP7_75t_R rebuffer1334 (.A(_09108_),
    .Y(net1739));
 BUFx6f_ASAP7_75t_R rebuffer1335 (.A(_10328_),
    .Y(net1740));
 BUFx2_ASAP7_75t_R rebuffer1336 (.A(net3035),
    .Y(net1741));
 BUFx2_ASAP7_75t_R rebuffer1337 (.A(_10328_),
    .Y(net1742));
 BUFx6f_ASAP7_75t_R split1338 (.A(_09695_),
    .Y(net1743));
 BUFx3_ASAP7_75t_R rebuffer1339 (.A(_16386_),
    .Y(net1744));
 BUFx2_ASAP7_75t_R rebuffer1340 (.A(net1744),
    .Y(net1745));
 BUFx4f_ASAP7_75t_R split1341 (.A(_17931_),
    .Y(net1746));
 BUFx2_ASAP7_75t_R rebuffer1342 (.A(net2302),
    .Y(net1747));
 BUFx2_ASAP7_75t_R rebuffer1343 (.A(net2302),
    .Y(net1748));
 BUFx3_ASAP7_75t_R rebuffer1344 (.A(net2387),
    .Y(net1749));
 BUFx2_ASAP7_75t_R rebuffer1345 (.A(net1749),
    .Y(net1750));
 BUFx6f_ASAP7_75t_R split1346 (.A(_21901_),
    .Y(net1751));
 BUFx10_ASAP7_75t_R split1347 (.A(_01146_),
    .Y(net1752));
 BUFx3_ASAP7_75t_R rebuffer1348 (.A(_18411_),
    .Y(net1753));
 BUFx2_ASAP7_75t_R rebuffer1349 (.A(net1753),
    .Y(net1754));
 BUFx2_ASAP7_75t_R rebuffer1350 (.A(net2701),
    .Y(net1755));
 BUFx2_ASAP7_75t_R rebuffer1351 (.A(_09925_),
    .Y(net1756));
 BUFx6f_ASAP7_75t_R split1352 (.A(_09925_),
    .Y(net1757));
 BUFx2_ASAP7_75t_R rebuffer1353 (.A(_06047_),
    .Y(net1758));
 BUFx2_ASAP7_75t_R rebuffer1354 (.A(net1758),
    .Y(net1759));
 BUFx6f_ASAP7_75t_R rebuffer1355 (.A(_00609_),
    .Y(net1760));
 BUFx2_ASAP7_75t_R rebuffer1356 (.A(net1760),
    .Y(net1761));
 BUFx2_ASAP7_75t_R rebuffer1357 (.A(net1761),
    .Y(net1762));
 BUFx2_ASAP7_75t_R rebuffer1358 (.A(net1760),
    .Y(net1763));
 BUFx6f_ASAP7_75t_R rebuffer1359 (.A(_05070_),
    .Y(net1764));
 BUFx2_ASAP7_75t_R rebuffer1360 (.A(net1764),
    .Y(net1765));
 BUFx3_ASAP7_75t_R rebuffer1361 (.A(net1764),
    .Y(net1766));
 BUFx6f_ASAP7_75t_R rebuffer1362 (.A(_05070_),
    .Y(net1767));
 BUFx2_ASAP7_75t_R rebuffer1363 (.A(_05156_),
    .Y(net1768));
 BUFx2_ASAP7_75t_R rebuffer1364 (.A(_14615_),
    .Y(net1769));
 BUFx2_ASAP7_75t_R rebuffer1365 (.A(_14615_),
    .Y(net1770));
 BUFx2_ASAP7_75t_R rebuffer1366 (.A(net2835),
    .Y(net1771));
 BUFx3_ASAP7_75t_R rebuffer1367 (.A(_05502_),
    .Y(net1772));
 BUFx6f_ASAP7_75t_R rebuffer1368 (.A(net1772),
    .Y(net1773));
 BUFx12f_ASAP7_75t_R rebuffer1369 (.A(_00544_),
    .Y(net1774));
 BUFx2_ASAP7_75t_R rebuffer1370 (.A(net1774),
    .Y(net1775));
 BUFx2_ASAP7_75t_R rebuffer1371 (.A(net1775),
    .Y(net1776));
 BUFx2_ASAP7_75t_R rebuffer1372 (.A(net1775),
    .Y(net1777));
 BUFx2_ASAP7_75t_R rebuffer1373 (.A(net1774),
    .Y(net1778));
 BUFx2_ASAP7_75t_R rebuffer1374 (.A(net1778),
    .Y(net1779));
 BUFx3_ASAP7_75t_R rebuffer1375 (.A(_00631_),
    .Y(net1780));
 BUFx3_ASAP7_75t_R rebuffer1376 (.A(net1780),
    .Y(net1781));
 BUFx3_ASAP7_75t_R rebuffer1377 (.A(_00631_),
    .Y(net1782));
 BUFx2_ASAP7_75t_R rebuffer1378 (.A(net1782),
    .Y(net1783));
 BUFx2_ASAP7_75t_R rebuffer1379 (.A(net1782),
    .Y(net1784));
 BUFx6f_ASAP7_75t_R rebuffer1380 (.A(_00631_),
    .Y(net1785));
 BUFx6f_ASAP7_75t_R rebuffer1381 (.A(_06449_),
    .Y(net1786));
 BUFx2_ASAP7_75t_R split1382 (.A(_06449_),
    .Y(net1787));
 BUFx2_ASAP7_75t_R rebuffer1383 (.A(_17815_),
    .Y(net1788));
 BUFx2_ASAP7_75t_R rebuffer1384 (.A(net1788),
    .Y(net1789));
 BUFx12f_ASAP7_75t_R rebuffer1385 (.A(_17934_),
    .Y(net1790));
 BUFx2_ASAP7_75t_R rebuffer1386 (.A(net3343),
    .Y(net1791));
 BUFx6f_ASAP7_75t_R split1387 (.A(_21997_),
    .Y(net1792));
 BUFx2_ASAP7_75t_R rebuffer1388 (.A(_05095_),
    .Y(net1793));
 BUFx2_ASAP7_75t_R rebuffer1389 (.A(_05095_),
    .Y(net1794));
 BUFx6f_ASAP7_75t_R split1390 (.A(_18052_),
    .Y(net1795));
 BUFx3_ASAP7_75t_R rebuffer1391 (.A(_09939_),
    .Y(net1796));
 BUFx2_ASAP7_75t_R rebuffer1392 (.A(net1796),
    .Y(net1797));
 BUFx2_ASAP7_75t_R rebuffer1393 (.A(_09939_),
    .Y(net1798));
 BUFx2_ASAP7_75t_R rebuffer1394 (.A(net1798),
    .Y(net1799));
 BUFx2_ASAP7_75t_R rebuffer1395 (.A(net1798),
    .Y(net1800));
 BUFx2_ASAP7_75t_R rebuffer1396 (.A(net1798),
    .Y(net1801));
 BUFx12f_ASAP7_75t_R rebuffer1397 (.A(_01384_),
    .Y(net1802));
 BUFx6f_ASAP7_75t_R rebuffer1398 (.A(net1802),
    .Y(net1803));
 BUFx2_ASAP7_75t_R rebuffer1399 (.A(_05772_),
    .Y(net1804));
 BUFx3_ASAP7_75t_R rebuffer1400 (.A(_05772_),
    .Y(net1805));
 BUFx6f_ASAP7_75t_R rebuffer1401 (.A(net1805),
    .Y(net1806));
 BUFx4f_ASAP7_75t_R split1402 (.A(_06429_),
    .Y(net1807));
 BUFx2_ASAP7_75t_R rebuffer1403 (.A(net3475),
    .Y(net1808));
 BUFx2_ASAP7_75t_R rebuffer1404 (.A(_05766_),
    .Y(net1809));
 BUFx2_ASAP7_75t_R rebuffer1405 (.A(_05766_),
    .Y(net1810));
 BUFx2_ASAP7_75t_R rebuffer1406 (.A(net1810),
    .Y(net1811));
 BUFx12f_ASAP7_75t_R rebuffer1407 (.A(_00629_),
    .Y(net1812));
 BUFx2_ASAP7_75t_R rebuffer1408 (.A(net1812),
    .Y(net1813));
 BUFx6f_ASAP7_75t_R rebuffer1409 (.A(net1812),
    .Y(net1814));
 BUFx3_ASAP7_75t_R split1410 (.A(_17946_),
    .Y(net1815));
 BUFx3_ASAP7_75t_R rebuffer1411 (.A(_17596_),
    .Y(net1816));
 BUFx2_ASAP7_75t_R rebuffer1412 (.A(_14622_),
    .Y(net1817));
 BUFx6f_ASAP7_75t_R rebuffer1413 (.A(_14622_),
    .Y(net1818));
 BUFx2_ASAP7_75t_R rebuffer1414 (.A(net1818),
    .Y(net1819));
 BUFx2_ASAP7_75t_R rebuffer1415 (.A(net1819),
    .Y(net1820));
 BUFx3_ASAP7_75t_R split1416 (.A(_18297_),
    .Y(net1821));
 BUFx6f_ASAP7_75t_R split1417 (.A(_05157_),
    .Y(net1822));
 BUFx2_ASAP7_75t_R rebuffer1418 (.A(_18516_),
    .Y(net1823));
 BUFx2_ASAP7_75t_R rebuffer1419 (.A(net1823),
    .Y(net1824));
 BUFx2_ASAP7_75t_R rebuffer1420 (.A(_18516_),
    .Y(net1825));
 BUFx2_ASAP7_75t_R rebuffer1421 (.A(_01292_),
    .Y(net1826));
 BUFx8_ASAP7_75t_R rebuffer1422 (.A(_01292_),
    .Y(net1827));
 BUFx2_ASAP7_75t_R rebuffer1423 (.A(net1827),
    .Y(net1828));
 BUFx4f_ASAP7_75t_R split1424 (.A(_22002_),
    .Y(net1829));
 BUFx6f_ASAP7_75t_R split1425 (.A(_14735_),
    .Y(net1830));
 BUFx6f_ASAP7_75t_R rebuffer1426 (.A(_17600_),
    .Y(net1831));
 BUFx2_ASAP7_75t_R rebuffer1427 (.A(_17600_),
    .Y(net1832));
 BUFx3_ASAP7_75t_R rebuffer1428 (.A(_21997_),
    .Y(net1833));
 BUFx2_ASAP7_75t_R rebuffer1429 (.A(_21997_),
    .Y(net1834));
 BUFx2_ASAP7_75t_R rebuffer1430 (.A(_05150_),
    .Y(net1835));
 BUFx6f_ASAP7_75t_R rebuffer1431 (.A(_05150_),
    .Y(net1836));
 BUFx2_ASAP7_75t_R rebuffer1432 (.A(net1836),
    .Y(net1837));
 BUFx2_ASAP7_75t_R rebuffer1433 (.A(net1836),
    .Y(net1838));
 BUFx2_ASAP7_75t_R split1434 (.A(_17956_),
    .Y(net1839));
 BUFx4f_ASAP7_75t_R split1435 (.A(_10578_),
    .Y(net1840));
 BUFx6f_ASAP7_75t_R rebuffer1436 (.A(_10343_),
    .Y(net1841));
 BUFx2_ASAP7_75t_R rebuffer1437 (.A(_00610_),
    .Y(net1842));
 BUFx2_ASAP7_75t_R rebuffer1438 (.A(_09583_),
    .Y(net1843));
 BUFx2_ASAP7_75t_R rebuffer1439 (.A(net1843),
    .Y(net1844));
 BUFx6f_ASAP7_75t_R rebuffer1440 (.A(_21904_),
    .Y(net1845));
 BUFx2_ASAP7_75t_R rebuffer1441 (.A(net1845),
    .Y(net1846));
 BUFx2_ASAP7_75t_R rebuffer1442 (.A(net1845),
    .Y(net1847));
 BUFx2_ASAP7_75t_R rebuffer1443 (.A(net1847),
    .Y(net1848));
 BUFx2_ASAP7_75t_R rebuffer1444 (.A(_21904_),
    .Y(net1849));
 BUFx2_ASAP7_75t_R rebuffer1445 (.A(net1849),
    .Y(net1850));
 BUFx6f_ASAP7_75t_R rebuffer1446 (.A(_21904_),
    .Y(net1851));
 BUFx2_ASAP7_75t_R rebuffer1447 (.A(net1851),
    .Y(net1852));
 BUFx2_ASAP7_75t_R rebuffer1448 (.A(net1851),
    .Y(net1853));
 BUFx10_ASAP7_75t_R split1449 (.A(_00435_),
    .Y(net1854));
 BUFx6f_ASAP7_75t_R rebuffer1450 (.A(_10451_),
    .Y(net1855));
 BUFx2_ASAP7_75t_R rebuffer1451 (.A(net1855),
    .Y(net1856));
 BUFx4f_ASAP7_75t_R rebuffer1452 (.A(_18178_),
    .Y(net1857));
 BUFx2_ASAP7_75t_R rebuffer1453 (.A(net1857),
    .Y(net1858));
 BUFx2_ASAP7_75t_R rebuffer1454 (.A(_18178_),
    .Y(net1859));
 BUFx6f_ASAP7_75t_R rebuffer1455 (.A(_08420_),
    .Y(net1860));
 BUFx2_ASAP7_75t_R rebuffer1456 (.A(net1860),
    .Y(net1861));
 BUFx6f_ASAP7_75t_R split1457 (.A(_10768_),
    .Y(net1862));
 BUFx6f_ASAP7_75t_R rebuffer1458 (.A(_18272_),
    .Y(net1863));
 BUFx6f_ASAP7_75t_R rebuffer1459 (.A(net1863),
    .Y(net1864));
 BUFx6f_ASAP7_75t_R rebuffer1460 (.A(_01252_),
    .Y(net1865));
 BUFx2_ASAP7_75t_R rebuffer1461 (.A(net1865),
    .Y(net1866));
 BUFx4f_ASAP7_75t_R split1462 (.A(_05156_),
    .Y(net1867));
 BUFx6f_ASAP7_75t_R rebuffer1463 (.A(_09718_),
    .Y(net1868));
 BUFx2_ASAP7_75t_R rebuffer1464 (.A(net1868),
    .Y(net1869));
 BUFx2_ASAP7_75t_R rebuffer1465 (.A(net1868),
    .Y(net1870));
 BUFx2_ASAP7_75t_R rebuffer1466 (.A(net1868),
    .Y(net1871));
 BUFx2_ASAP7_75t_R rebuffer1467 (.A(net1871),
    .Y(net1872));
 BUFx2_ASAP7_75t_R rebuffer1468 (.A(_14715_),
    .Y(net1873));
 BUFx2_ASAP7_75t_R rebuffer1469 (.A(net1873),
    .Y(net1874));
 BUFx2_ASAP7_75t_R rebuffer1470 (.A(net1874),
    .Y(net1875));
 BUFx3_ASAP7_75t_R split1471 (.A(_10394_),
    .Y(net1876));
 BUFx12f_ASAP7_75t_R rebuffer1472 (.A(_05337_),
    .Y(net1877));
 BUFx2_ASAP7_75t_R rebuffer1473 (.A(net1877),
    .Y(net1878));
 BUFx2_ASAP7_75t_R rebuffer1474 (.A(net1877),
    .Y(net1879));
 BUFx2_ASAP7_75t_R split1475 (.A(_05754_),
    .Y(net1880));
 BUFx6f_ASAP7_75t_R split1476 (.A(_10431_),
    .Y(net1881));
 BUFx3_ASAP7_75t_R rebuffer1477 (.A(_10121_),
    .Y(net1882));
 BUFx6f_ASAP7_75t_R rebuffer1478 (.A(_10121_),
    .Y(net1883));
 BUFx4f_ASAP7_75t_R split1479 (.A(_01252_),
    .Y(net1884));
 BUFx6f_ASAP7_75t_R split1480 (.A(_10343_),
    .Y(net1885));
 BUFx2_ASAP7_75t_R rebuffer1481 (.A(net2031),
    .Y(net1886));
 BUFx6f_ASAP7_75t_R rebuffer1482 (.A(_01589_),
    .Y(net1887));
 BUFx2_ASAP7_75t_R rebuffer1483 (.A(net1887),
    .Y(net1888));
 BUFx2_ASAP7_75t_R rebuffer1484 (.A(net1887),
    .Y(net1889));
 BUFx2_ASAP7_75t_R rebuffer1485 (.A(_10004_),
    .Y(net1890));
 BUFx2_ASAP7_75t_R rebuffer1486 (.A(net1890),
    .Y(net1891));
 BUFx2_ASAP7_75t_R rebuffer1487 (.A(net1890),
    .Y(net1892));
 BUFx2_ASAP7_75t_R rebuffer1488 (.A(_10004_),
    .Y(net1893));
 BUFx4f_ASAP7_75t_R split1489 (.A(_05073_),
    .Y(net1894));
 BUFx2_ASAP7_75t_R rebuffer1490 (.A(_00640_),
    .Y(net1895));
 BUFx12f_ASAP7_75t_R rebuffer1491 (.A(_00640_),
    .Y(net1896));
 BUFx2_ASAP7_75t_R rebuffer1492 (.A(net1896),
    .Y(net1897));
 BUFx2_ASAP7_75t_R rebuffer1493 (.A(net1896),
    .Y(net1898));
 BUFx2_ASAP7_75t_R rebuffer1494 (.A(net1896),
    .Y(net1899));
 BUFx3_ASAP7_75t_R rebuffer1495 (.A(net1896),
    .Y(net1900));
 BUFx3_ASAP7_75t_R rebuffer1496 (.A(_17676_),
    .Y(net1901));
 BUFx3_ASAP7_75t_R rebuffer1497 (.A(_05535_),
    .Y(net1902));
 BUFx2_ASAP7_75t_R rebuffer1498 (.A(net2703),
    .Y(net1903));
 BUFx2_ASAP7_75t_R rebuffer1499 (.A(_21884_),
    .Y(net1904));
 BUFx2_ASAP7_75t_R rebuffer1500 (.A(net1904),
    .Y(net1905));
 BUFx2_ASAP7_75t_R rebuffer1501 (.A(_21884_),
    .Y(net1906));
 BUFx2_ASAP7_75t_R rebuffer1502 (.A(_18065_),
    .Y(net1907));
 BUFx2_ASAP7_75t_R rebuffer1503 (.A(net1907),
    .Y(net1908));
 BUFx2_ASAP7_75t_R rebuffer1504 (.A(net1907),
    .Y(net1909));
 BUFx6f_ASAP7_75t_R rebuffer1505 (.A(_18065_),
    .Y(net1910));
 BUFx2_ASAP7_75t_R rebuffer1506 (.A(net1910),
    .Y(net1911));
 BUFx2_ASAP7_75t_R rebuffer1507 (.A(net1910),
    .Y(net1912));
 BUFx6f_ASAP7_75t_R split1508 (.A(_05943_),
    .Y(net1913));
 BUFx3_ASAP7_75t_R rebuffer1509 (.A(_01159_),
    .Y(net1914));
 BUFx2_ASAP7_75t_R rebuffer1510 (.A(net1914),
    .Y(net1915));
 BUFx2_ASAP7_75t_R rebuffer1511 (.A(net1915),
    .Y(net1916));
 BUFx2_ASAP7_75t_R rebuffer1512 (.A(_01159_),
    .Y(net1917));
 BUFx2_ASAP7_75t_R rebuffer1513 (.A(_01159_),
    .Y(net1918));
 BUFx2_ASAP7_75t_R rebuffer1514 (.A(_01159_),
    .Y(net1919));
 BUFx2_ASAP7_75t_R rebuffer1515 (.A(net1919),
    .Y(net1920));
 BUFx2_ASAP7_75t_R rebuffer1516 (.A(_05222_),
    .Y(net1921));
 BUFx2_ASAP7_75t_R rebuffer1517 (.A(_05222_),
    .Y(net1922));
 BUFx2_ASAP7_75t_R rebuffer1518 (.A(_09611_),
    .Y(net1923));
 BUFx2_ASAP7_75t_R rebuffer1519 (.A(net1923),
    .Y(net1924));
 BUFx2_ASAP7_75t_R rebuffer1520 (.A(_09611_),
    .Y(net1925));
 BUFx2_ASAP7_75t_R rebuffer1521 (.A(net2589),
    .Y(net1926));
 BUFx6f_ASAP7_75t_R rebuffer1522 (.A(_06681_),
    .Y(net1927));
 BUFx2_ASAP7_75t_R rebuffer1523 (.A(net1927),
    .Y(net1928));
 BUFx2_ASAP7_75t_R rebuffer1524 (.A(_06681_),
    .Y(net1929));
 BUFx2_ASAP7_75t_R rebuffer1525 (.A(_09603_),
    .Y(net1930));
 BUFx2_ASAP7_75t_R rebuffer1526 (.A(net1930),
    .Y(net1931));
 BUFx3_ASAP7_75t_R rebuffer1527 (.A(_09603_),
    .Y(net1932));
 BUFx12f_ASAP7_75t_R rebuffer1528 (.A(_09603_),
    .Y(net1933));
 BUFx2_ASAP7_75t_R rebuffer1529 (.A(net1933),
    .Y(net1934));
 BUFx6f_ASAP7_75t_R rebuffer1530 (.A(_06200_),
    .Y(net1935));
 BUFx6f_ASAP7_75t_R rebuffer1531 (.A(net1935),
    .Y(net1936));
 BUFx2_ASAP7_75t_R rebuffer1532 (.A(net1936),
    .Y(net1937));
 BUFx2_ASAP7_75t_R rebuffer1533 (.A(net1937),
    .Y(net1938));
 BUFx2_ASAP7_75t_R rebuffer1534 (.A(_06200_),
    .Y(net1939));
 BUFx2_ASAP7_75t_R rebuffer1535 (.A(net1939),
    .Y(net1940));
 BUFx2_ASAP7_75t_R rebuffer1536 (.A(net1940),
    .Y(net1941));
 BUFx6f_ASAP7_75t_R split1537 (.A(_09755_),
    .Y(net1942));
 BUFx4f_ASAP7_75t_R split1538 (.A(_14660_),
    .Y(net1943));
 BUFx2_ASAP7_75t_R rebuffer1539 (.A(_05135_),
    .Y(net1944));
 BUFx6f_ASAP7_75t_R rebuffer1540 (.A(_05135_),
    .Y(net1945));
 BUFx2_ASAP7_75t_R rebuffer1541 (.A(net1945),
    .Y(net1946));
 BUFx2_ASAP7_75t_R rebuffer1542 (.A(net1945),
    .Y(net1947));
 BUFx3_ASAP7_75t_R split1543 (.A(_08853_),
    .Y(net1948));
 BUFx3_ASAP7_75t_R rebuffer1544 (.A(_09943_),
    .Y(net1949));
 BUFx2_ASAP7_75t_R rebuffer1545 (.A(net1949),
    .Y(net1950));
 BUFx2_ASAP7_75t_R rebuffer1546 (.A(_09943_),
    .Y(net1951));
 BUFx2_ASAP7_75t_R rebuffer1547 (.A(net1951),
    .Y(net1952));
 BUFx2_ASAP7_75t_R rebuffer1548 (.A(net1951),
    .Y(net1953));
 BUFx6f_ASAP7_75t_R split1549 (.A(_18327_),
    .Y(net1954));
 BUFx6f_ASAP7_75t_R split1550 (.A(_17977_),
    .Y(net1955));
 BUFx6f_ASAP7_75t_R rebuffer1551 (.A(_00645_),
    .Y(net1956));
 BUFx3_ASAP7_75t_R rebuffer1552 (.A(net1956),
    .Y(net1957));
 BUFx2_ASAP7_75t_R rebuffer1553 (.A(net2093),
    .Y(net1958));
 BUFx2_ASAP7_75t_R rebuffer1554 (.A(net1958),
    .Y(net1959));
 BUFx6f_ASAP7_75t_R rebuffer1555 (.A(_00573_),
    .Y(net1960));
 BUFx3_ASAP7_75t_R rebuffer1556 (.A(_10013_),
    .Y(net1961));
 BUFx2_ASAP7_75t_R rebuffer1557 (.A(net1961),
    .Y(net1962));
 BUFx3_ASAP7_75t_R rebuffer1558 (.A(_10013_),
    .Y(net1963));
 BUFx3_ASAP7_75t_R rebuffer1559 (.A(net2402),
    .Y(net1964));
 BUFx6f_ASAP7_75t_R split1560 (.A(_18518_),
    .Y(net1965));
 BUFx6f_ASAP7_75t_R rebuffer1561 (.A(_18518_),
    .Y(net1966));
 BUFx6f_ASAP7_75t_R rebuffer1562 (.A(_01145_),
    .Y(net1967));
 BUFx2_ASAP7_75t_R rebuffer1563 (.A(net1967),
    .Y(net1968));
 BUFx2_ASAP7_75t_R rebuffer1564 (.A(net1967),
    .Y(net1969));
 BUFx2_ASAP7_75t_R rebuffer1565 (.A(_01145_),
    .Y(net1970));
 BUFx2_ASAP7_75t_R rebuffer1566 (.A(net1970),
    .Y(net1971));
 BUFx2_ASAP7_75t_R rebuffer1567 (.A(net1971),
    .Y(net1972));
 BUFx4f_ASAP7_75t_R rebuffer1568 (.A(_17557_),
    .Y(net1973));
 BUFx2_ASAP7_75t_R rebuffer1569 (.A(net1973),
    .Y(net1974));
 BUFx10_ASAP7_75t_R rebuffer1570 (.A(net1973),
    .Y(net1975));
 BUFx2_ASAP7_75t_R rebuffer1571 (.A(net1975),
    .Y(net1976));
 BUFx2_ASAP7_75t_R rebuffer1572 (.A(net1976),
    .Y(net1977));
 BUFx12f_ASAP7_75t_R rebuffer1573 (.A(_05794_),
    .Y(net1978));
 BUFx3_ASAP7_75t_R rebuffer1574 (.A(_10468_),
    .Y(net1979));
 BUFx2_ASAP7_75t_R rebuffer1575 (.A(net1979),
    .Y(net1980));
 BUFx2_ASAP7_75t_R rebuffer1576 (.A(_10468_),
    .Y(net1981));
 BUFx6f_ASAP7_75t_R split1577 (.A(_10672_),
    .Y(net1982));
 BUFx2_ASAP7_75t_R rebuffer1578 (.A(_14605_),
    .Y(net1983));
 BUFx2_ASAP7_75t_R rebuffer1579 (.A(net1983),
    .Y(net1984));
 BUFx2_ASAP7_75t_R rebuffer1580 (.A(_14605_),
    .Y(net1985));
 BUFx2_ASAP7_75t_R rebuffer1581 (.A(net1985),
    .Y(net1986));
 BUFx2_ASAP7_75t_R rebuffer1582 (.A(net1985),
    .Y(net1987));
 BUFx2_ASAP7_75t_R rebuffer1583 (.A(net1987),
    .Y(net1988));
 BUFx2_ASAP7_75t_R rebuffer1584 (.A(net1985),
    .Y(net1989));
 BUFx10_ASAP7_75t_R rebuffer1585 (.A(_10680_),
    .Y(net1990));
 BUFx6f_ASAP7_75t_R rebuffer1586 (.A(net1990),
    .Y(net1991));
 BUFx2_ASAP7_75t_R rebuffer1587 (.A(net1991),
    .Y(net1992));
 BUFx2_ASAP7_75t_R rebuffer1588 (.A(_10680_),
    .Y(net1993));
 BUFx2_ASAP7_75t_R rebuffer1589 (.A(net1993),
    .Y(net1994));
 BUFx6f_ASAP7_75t_R rebuffer1590 (.A(_10680_),
    .Y(net1995));
 BUFx2_ASAP7_75t_R rebuffer1591 (.A(net1995),
    .Y(net1996));
 BUFx2_ASAP7_75t_R rebuffer1592 (.A(net1996),
    .Y(net1997));
 BUFx2_ASAP7_75t_R rebuffer1593 (.A(_09678_),
    .Y(net1998));
 BUFx2_ASAP7_75t_R rebuffer1594 (.A(net1998),
    .Y(net1999));
 BUFx3_ASAP7_75t_R rebuffer1595 (.A(_09678_),
    .Y(net2000));
 BUFx2_ASAP7_75t_R rebuffer1596 (.A(net2000),
    .Y(net2001));
 BUFx6f_ASAP7_75t_R rebuffer1597 (.A(_09678_),
    .Y(net2002));
 BUFx6f_ASAP7_75t_R split1598 (.A(_06574_),
    .Y(net2003));
 BUFx6f_ASAP7_75t_R split1599 (.A(_18333_),
    .Y(net2004));
 BUFx6f_ASAP7_75t_R rebuffer1600 (.A(_00549_),
    .Y(net2005));
 BUFx2_ASAP7_75t_R rebuffer1601 (.A(net2005),
    .Y(net2006));
 BUFx2_ASAP7_75t_R rebuffer1602 (.A(net2005),
    .Y(net2007));
 BUFx2_ASAP7_75t_R rebuffer1603 (.A(net3246),
    .Y(net2008));
 BUFx2_ASAP7_75t_R rebuffer1604 (.A(_18253_),
    .Y(net2009));
 BUFx2_ASAP7_75t_R rebuffer1605 (.A(net2009),
    .Y(net2010));
 BUFx2_ASAP7_75t_R rebuffer1606 (.A(_18253_),
    .Y(net2011));
 BUFx6f_ASAP7_75t_R rebuffer1607 (.A(_18575_),
    .Y(net2012));
 BUFx6f_ASAP7_75t_R rebuffer1608 (.A(_17582_),
    .Y(net2013));
 BUFx3_ASAP7_75t_R rebuffer1609 (.A(net2013),
    .Y(net2014));
 BUFx3_ASAP7_75t_R rebuffer1610 (.A(_17582_),
    .Y(net2015));
 BUFx2_ASAP7_75t_R rebuffer1611 (.A(_05466_),
    .Y(net2016));
 BUFx2_ASAP7_75t_R rebuffer1612 (.A(net2016),
    .Y(net2017));
 BUFx2_ASAP7_75t_R rebuffer1613 (.A(_00641_),
    .Y(net2018));
 BUFx6f_ASAP7_75t_R rebuffer1614 (.A(_00641_),
    .Y(net2019));
 BUFx4f_ASAP7_75t_R split1615 (.A(_10454_),
    .Y(net2020));
 BUFx3_ASAP7_75t_R rebuffer1616 (.A(_10685_),
    .Y(net2021));
 BUFx2_ASAP7_75t_R rebuffer1617 (.A(net2021),
    .Y(net2022));
 BUFx3_ASAP7_75t_R rebuffer1618 (.A(net2022),
    .Y(net2023));
 BUFx2_ASAP7_75t_R rebuffer1619 (.A(_10685_),
    .Y(net2024));
 BUFx3_ASAP7_75t_R rebuffer1620 (.A(net2024),
    .Y(net2025));
 BUFx3_ASAP7_75t_R rebuffer1621 (.A(_10685_),
    .Y(net2026));
 BUFx4f_ASAP7_75t_R split1622 (.A(_05095_),
    .Y(net2027));
 BUFx6f_ASAP7_75t_R rebuffer1623 (.A(_18657_),
    .Y(net2028));
 BUFx2_ASAP7_75t_R rebuffer1624 (.A(_18657_),
    .Y(net2029));
 BUFx2_ASAP7_75t_R rebuffer1625 (.A(net2029),
    .Y(net2030));
 BUFx6f_ASAP7_75t_R split1626 (.A(_04453_),
    .Y(net2031));
 BUFx4f_ASAP7_75t_R split1627 (.A(_05530_),
    .Y(net2032));
 BUFx2_ASAP7_75t_R rebuffer1628 (.A(_05530_),
    .Y(net2033));
 BUFx2_ASAP7_75t_R rebuffer1629 (.A(net2033),
    .Y(net2034));
 BUFx3_ASAP7_75t_R rebuffer1630 (.A(_05530_),
    .Y(net2035));
 BUFx6f_ASAP7_75t_R rebuffer1631 (.A(net2035),
    .Y(net2036));
 BUFx3_ASAP7_75t_R rebuffer1632 (.A(_09890_),
    .Y(net2037));
 BUFx12f_ASAP7_75t_R rebuffer1633 (.A(_22046_),
    .Y(net2038));
 BUFx6f_ASAP7_75t_R rebuffer1634 (.A(net2038),
    .Y(net2039));
 BUFx6f_ASAP7_75t_R rebuffer1635 (.A(net2038),
    .Y(net2040));
 BUFx3_ASAP7_75t_R rebuffer1636 (.A(_02091_),
    .Y(net2041));
 BUFx2_ASAP7_75t_R rebuffer1637 (.A(_02091_),
    .Y(net2042));
 BUFx6f_ASAP7_75t_R rebuffer1638 (.A(_18314_),
    .Y(net2043));
 BUFx2_ASAP7_75t_R rebuffer1639 (.A(net2043),
    .Y(net2044));
 BUFx2_ASAP7_75t_R rebuffer1640 (.A(_18314_),
    .Y(net2045));
 BUFx2_ASAP7_75t_R rebuffer1641 (.A(_09739_),
    .Y(net2046));
 BUFx2_ASAP7_75t_R rebuffer1642 (.A(_09739_),
    .Y(net2047));
 BUFx2_ASAP7_75t_R rebuffer1643 (.A(net2047),
    .Y(net2048));
 BUFx3_ASAP7_75t_R split1644 (.A(_09889_),
    .Y(net2049));
 BUFx6f_ASAP7_75t_R rebuffer1645 (.A(_18333_),
    .Y(net2050));
 BUFx2_ASAP7_75t_R rebuffer1646 (.A(net2466),
    .Y(net2051));
 BUFx2_ASAP7_75t_R rebuffer1647 (.A(_18516_),
    .Y(net2052));
 BUFx4f_ASAP7_75t_R split1648 (.A(_10768_),
    .Y(net2053));
 BUFx3_ASAP7_75t_R rebuffer1649 (.A(_13096_),
    .Y(net2054));
 BUFx6f_ASAP7_75t_R split1650 (.A(net3390),
    .Y(net2055));
 BUFx6f_ASAP7_75t_R split1651 (.A(_05157_),
    .Y(net2056));
 BUFx2_ASAP7_75t_R rebuffer1652 (.A(_17951_),
    .Y(net2057));
 BUFx2_ASAP7_75t_R rebuffer1653 (.A(net2057),
    .Y(net2058));
 BUFx2_ASAP7_75t_R rebuffer1654 (.A(_17951_),
    .Y(net2059));
 BUFx2_ASAP7_75t_R rebuffer1655 (.A(_17951_),
    .Y(net2060));
 BUFx2_ASAP7_75t_R rebuffer1656 (.A(_10672_),
    .Y(net2061));
 BUFx12f_ASAP7_75t_R rebuffer1657 (.A(_01553_),
    .Y(net2062));
 BUFx2_ASAP7_75t_R rebuffer1658 (.A(net2062),
    .Y(net2063));
 BUFx2_ASAP7_75t_R rebuffer1659 (.A(net2062),
    .Y(net2064));
 BUFx2_ASAP7_75t_R rebuffer1660 (.A(net2062),
    .Y(net2065));
 BUFx2_ASAP7_75t_R rebuffer1661 (.A(net2062),
    .Y(net2066));
 BUFx6f_ASAP7_75t_R split1662 (.A(_18575_),
    .Y(net2067));
 BUFx12f_ASAP7_75t_R rebuffer1663 (.A(_09596_),
    .Y(net2068));
 BUFx2_ASAP7_75t_R rebuffer1664 (.A(_10482_),
    .Y(net2069));
 BUFx4f_ASAP7_75t_R rebuffer1665 (.A(_10482_),
    .Y(net2070));
 BUFx2_ASAP7_75t_R rebuffer1666 (.A(_01510_),
    .Y(net2071));
 BUFx2_ASAP7_75t_R rebuffer1667 (.A(_01510_),
    .Y(net2072));
 BUFx6f_ASAP7_75t_R rebuffer1668 (.A(_01510_),
    .Y(net2073));
 BUFx2_ASAP7_75t_R rebuffer1669 (.A(net2073),
    .Y(net2074));
 BUFx2_ASAP7_75t_R rebuffer1670 (.A(net2074),
    .Y(net2075));
 BUFx2_ASAP7_75t_R rebuffer1671 (.A(net2073),
    .Y(net2076));
 BUFx2_ASAP7_75t_R rebuffer1672 (.A(net2073),
    .Y(net2077));
 BUFx2_ASAP7_75t_R rebuffer1673 (.A(net2077),
    .Y(net2078));
 BUFx2_ASAP7_75t_R rebuffer1674 (.A(net2077),
    .Y(net2079));
 BUFx2_ASAP7_75t_R rebuffer1675 (.A(net2079),
    .Y(net2080));
 BUFx4f_ASAP7_75t_R rebuffer1676 (.A(_05747_),
    .Y(net2081));
 BUFx3_ASAP7_75t_R rebuffer1677 (.A(net2081),
    .Y(net2082));
 BUFx2_ASAP7_75t_R rebuffer1678 (.A(net2081),
    .Y(net2083));
 BUFx6f_ASAP7_75t_R rebuffer1679 (.A(_06213_),
    .Y(net2084));
 BUFx6f_ASAP7_75t_R split1680 (.A(_09770_),
    .Y(net2085));
 BUFx12f_ASAP7_75t_R rebuffer1681 (.A(_17592_),
    .Y(net2086));
 BUFx2_ASAP7_75t_R rebuffer1682 (.A(net2086),
    .Y(net2087));
 BUFx2_ASAP7_75t_R rebuffer1683 (.A(_17592_),
    .Y(net2088));
 BUFx2_ASAP7_75t_R rebuffer1684 (.A(_18600_),
    .Y(net2089));
 BUFx2_ASAP7_75t_R rebuffer1685 (.A(_05440_),
    .Y(net2090));
 BUFx2_ASAP7_75t_R rebuffer1686 (.A(_05440_),
    .Y(net2091));
 BUFx2_ASAP7_75t_R rebuffer1687 (.A(_05440_),
    .Y(net2092));
 BUFx3_ASAP7_75t_R split1688 (.A(_18268_),
    .Y(net2093));
 BUFx2_ASAP7_75t_R rebuffer1689 (.A(net2161),
    .Y(net2094));
 BUFx6f_ASAP7_75t_R rebuffer1690 (.A(_18351_),
    .Y(net2095));
 BUFx3_ASAP7_75t_R rebuffer1691 (.A(net2095),
    .Y(net2096));
 BUFx2_ASAP7_75t_R rebuffer1692 (.A(net2096),
    .Y(net2097));
 BUFx16f_ASAP7_75t_R rebuffer1693 (.A(_05943_),
    .Y(net2098));
 BUFx2_ASAP7_75t_R rebuffer1694 (.A(_18518_),
    .Y(net2099));
 BUFx2_ASAP7_75t_R rebuffer1695 (.A(_09585_),
    .Y(net2100));
 BUFx2_ASAP7_75t_R rebuffer1696 (.A(_18511_),
    .Y(net2101));
 BUFx2_ASAP7_75t_R rebuffer1697 (.A(_18511_),
    .Y(net2102));
 BUFx4f_ASAP7_75t_R rebuffer1698 (.A(_09715_),
    .Y(net2103));
 BUFx6f_ASAP7_75t_R rebuffer1699 (.A(_09715_),
    .Y(net2104));
 BUFx2_ASAP7_75t_R rebuffer1700 (.A(net2104),
    .Y(net2105));
 BUFx3_ASAP7_75t_R rebuffer1701 (.A(_18239_),
    .Y(net2106));
 BUFx2_ASAP7_75t_R rebuffer1702 (.A(_18239_),
    .Y(net2107));
 BUFx3_ASAP7_75t_R rebuffer1703 (.A(_00605_),
    .Y(net2108));
 BUFx2_ASAP7_75t_R rebuffer1704 (.A(net2108),
    .Y(net2109));
 BUFx6f_ASAP7_75t_R rebuffer1705 (.A(_00577_),
    .Y(net2110));
 BUFx2_ASAP7_75t_R rebuffer1706 (.A(net2110),
    .Y(net2111));
 BUFx2_ASAP7_75t_R rebuffer1707 (.A(net2110),
    .Y(net2112));
 BUFx2_ASAP7_75t_R rebuffer1708 (.A(net2112),
    .Y(net2113));
 BUFx3_ASAP7_75t_R rebuffer1709 (.A(_00577_),
    .Y(net2114));
 BUFx2_ASAP7_75t_R rebuffer1710 (.A(_05619_),
    .Y(net2115));
 BUFx4f_ASAP7_75t_R rebuffer1711 (.A(_05619_),
    .Y(net2116));
 BUFx6f_ASAP7_75t_R rebuffer1712 (.A(_03881_),
    .Y(net2117));
 BUFx3_ASAP7_75t_R rebuffer1713 (.A(_10669_),
    .Y(net2118));
 BUFx2_ASAP7_75t_R rebuffer1714 (.A(net2118),
    .Y(net2119));
 BUFx6f_ASAP7_75t_R rebuffer1715 (.A(_01246_),
    .Y(net2120));
 BUFx2_ASAP7_75t_R rebuffer1716 (.A(net2120),
    .Y(net2121));
 BUFx2_ASAP7_75t_R rebuffer1717 (.A(net2120),
    .Y(net2122));
 BUFx2_ASAP7_75t_R rebuffer1718 (.A(net2120),
    .Y(net2123));
 BUFx2_ASAP7_75t_R rebuffer1719 (.A(net2120),
    .Y(net2124));
 BUFx2_ASAP7_75t_R rebuffer1720 (.A(net2120),
    .Y(net2125));
 BUFx3_ASAP7_75t_R split1721 (.A(_05222_),
    .Y(net2126));
 BUFx2_ASAP7_75t_R rebuffer1722 (.A(_11600_),
    .Y(net2127));
 BUFx2_ASAP7_75t_R rebuffer1723 (.A(_00428_),
    .Y(net2128));
 BUFx2_ASAP7_75t_R rebuffer1724 (.A(_00428_),
    .Y(net2129));
 BUFx6f_ASAP7_75t_R rebuffer1725 (.A(_00428_),
    .Y(net2130));
 BUFx2_ASAP7_75t_R rebuffer1726 (.A(net2130),
    .Y(net2131));
 BUFx2_ASAP7_75t_R rebuffer1727 (.A(net2131),
    .Y(net2132));
 BUFx2_ASAP7_75t_R rebuffer1728 (.A(_00428_),
    .Y(net2133));
 BUFx6f_ASAP7_75t_R rebuffer1729 (.A(net2133),
    .Y(net2134));
 BUFx2_ASAP7_75t_R rebuffer1730 (.A(net2134),
    .Y(net2135));
 BUFx6f_ASAP7_75t_R split1731 (.A(net3535),
    .Y(net2136));
 BUFx6f_ASAP7_75t_R rebuffer1732 (.A(_05211_),
    .Y(net2137));
 BUFx2_ASAP7_75t_R rebuffer1733 (.A(net2137),
    .Y(net2138));
 BUFx3_ASAP7_75t_R rebuffer1734 (.A(net2137),
    .Y(net2139));
 BUFx4f_ASAP7_75t_R split1735 (.A(_01916_),
    .Y(net2140));
 BUFx3_ASAP7_75t_R rebuffer1736 (.A(_19961_),
    .Y(net2141));
 BUFx4f_ASAP7_75t_R split1737 (.A(_18643_),
    .Y(net2142));
 BUFx12f_ASAP7_75t_R rebuffer1738 (.A(_18230_),
    .Y(net2143));
 BUFx2_ASAP7_75t_R rebuffer1739 (.A(net2143),
    .Y(net2144));
 BUFx2_ASAP7_75t_R rebuffer1740 (.A(net2143),
    .Y(net2145));
 BUFx6f_ASAP7_75t_R split1741 (.A(_05163_),
    .Y(net2146));
 BUFx12f_ASAP7_75t_R rebuffer1742 (.A(_10650_),
    .Y(net2147));
 BUFx2_ASAP7_75t_R rebuffer1743 (.A(net2147),
    .Y(net2148));
 BUFx6f_ASAP7_75t_R rebuffer1744 (.A(_05119_),
    .Y(net2149));
 BUFx2_ASAP7_75t_R rebuffer1745 (.A(_05119_),
    .Y(net2150));
 BUFx2_ASAP7_75t_R rebuffer1746 (.A(_09591_),
    .Y(net2151));
 BUFx2_ASAP7_75t_R rebuffer1747 (.A(_09591_),
    .Y(net2152));
 BUFx3_ASAP7_75t_R split1748 (.A(_05502_),
    .Y(net2153));
 BUFx6f_ASAP7_75t_R rebuffer1749 (.A(_00646_),
    .Y(net2154));
 BUFx2_ASAP7_75t_R rebuffer1750 (.A(net2154),
    .Y(net2155));
 BUFx2_ASAP7_75t_R rebuffer1751 (.A(_06920_),
    .Y(net2156));
 BUFx2_ASAP7_75t_R rebuffer1752 (.A(_16263_),
    .Y(net2157));
 BUFx2_ASAP7_75t_R rebuffer1753 (.A(_16263_),
    .Y(net2158));
 BUFx2_ASAP7_75t_R rebuffer1754 (.A(net2158),
    .Y(net2159));
 BUFx2_ASAP7_75t_R split1755 (.A(_10013_),
    .Y(net2160));
 BUFx2_ASAP7_75t_R split1756 (.A(_05239_),
    .Y(net2161));
 BUFx6f_ASAP7_75t_R rebuffer1757 (.A(_18155_),
    .Y(net2162));
 BUFx3_ASAP7_75t_R rebuffer1758 (.A(_18155_),
    .Y(net2163));
 BUFx3_ASAP7_75t_R rebuffer1759 (.A(net2163),
    .Y(net2164));
 BUFx2_ASAP7_75t_R rebuffer1760 (.A(_18107_),
    .Y(net2165));
 BUFx2_ASAP7_75t_R rebuffer1761 (.A(net2680),
    .Y(net2166));
 BUFx6f_ASAP7_75t_R rebuffer1762 (.A(_21123_),
    .Y(net2167));
 BUFx6f_ASAP7_75t_R rebuffer1763 (.A(_21123_),
    .Y(net2168));
 BUFx12f_ASAP7_75t_R rebuffer1764 (.A(_05066_),
    .Y(net2169));
 BUFx2_ASAP7_75t_R rebuffer1765 (.A(net2169),
    .Y(net2170));
 BUFx6f_ASAP7_75t_R rebuffer1766 (.A(_05066_),
    .Y(net2171));
 BUFx2_ASAP7_75t_R rebuffer1767 (.A(net2533),
    .Y(net2172));
 BUFx6f_ASAP7_75t_R rebuffer1768 (.A(_00612_),
    .Y(net2173));
 BUFx2_ASAP7_75t_R rebuffer1769 (.A(net2173),
    .Y(net2174));
 BUFx6f_ASAP7_75t_R split1770 (.A(_01831_),
    .Y(net2175));
 BUFx6f_ASAP7_75t_R split1771 (.A(net2713),
    .Y(net2176));
 BUFx3_ASAP7_75t_R split1772 (.A(_18600_),
    .Y(net2177));
 BUFx4f_ASAP7_75t_R split1773 (.A(net3518),
    .Y(net2178));
 BUFx6f_ASAP7_75t_R split1774 (.A(_14716_),
    .Y(net2179));
 BUFx3_ASAP7_75t_R split1775 (.A(_10600_),
    .Y(net2180));
 BUFx4f_ASAP7_75t_R split1776 (.A(_18074_),
    .Y(net2181));
 BUFx3_ASAP7_75t_R rebuffer1777 (.A(_18695_),
    .Y(net2182));
 BUFx6f_ASAP7_75t_R rebuffer1778 (.A(_05741_),
    .Y(net2183));
 BUFx2_ASAP7_75t_R rebuffer1779 (.A(net2183),
    .Y(net2184));
 BUFx6f_ASAP7_75t_R rebuffer1780 (.A(net2184),
    .Y(net2185));
 BUFx2_ASAP7_75t_R rebuffer1781 (.A(net2185),
    .Y(net2186));
 BUFx2_ASAP7_75t_R rebuffer1782 (.A(_10389_),
    .Y(net2187));
 BUFx6f_ASAP7_75t_R rebuffer1783 (.A(net3010),
    .Y(net2188));
 BUFx2_ASAP7_75t_R rebuffer1784 (.A(net3010),
    .Y(net2189));
 BUFx2_ASAP7_75t_R rebuffer1785 (.A(net3010),
    .Y(net2190));
 BUFx4f_ASAP7_75t_R split1786 (.A(_05447_),
    .Y(net2191));
 BUFx6f_ASAP7_75t_R rebuffer1787 (.A(_09881_),
    .Y(net2192));
 BUFx2_ASAP7_75t_R rebuffer1788 (.A(_01936_),
    .Y(net2193));
 BUFx2_ASAP7_75t_R rebuffer1789 (.A(_01936_),
    .Y(net2194));
 BUFx2_ASAP7_75t_R rebuffer1790 (.A(net2194),
    .Y(net2195));
 BUFx2_ASAP7_75t_R rebuffer1791 (.A(_00451_),
    .Y(net2196));
 BUFx6f_ASAP7_75t_R rebuffer1792 (.A(_00451_),
    .Y(net2197));
 BUFx2_ASAP7_75t_R rebuffer1793 (.A(net2197),
    .Y(net2198));
 BUFx2_ASAP7_75t_R rebuffer1794 (.A(_00451_),
    .Y(net2199));
 BUFx3_ASAP7_75t_R rebuffer1795 (.A(net2199),
    .Y(net2200));
 BUFx2_ASAP7_75t_R rebuffer1796 (.A(_00451_),
    .Y(net2201));
 BUFx6f_ASAP7_75t_R split1797 (.A(_17687_),
    .Y(net2202));
 BUFx2_ASAP7_75t_R rebuffer1798 (.A(_00436_),
    .Y(net2203));
 BUFx2_ASAP7_75t_R rebuffer1799 (.A(_00436_),
    .Y(net2204));
 BUFx2_ASAP7_75t_R rebuffer1800 (.A(net2204),
    .Y(net2205));
 BUFx2_ASAP7_75t_R rebuffer1801 (.A(net2205),
    .Y(net2206));
 BUFx12f_ASAP7_75t_R rebuffer1802 (.A(_00436_),
    .Y(net2207));
 BUFx2_ASAP7_75t_R rebuffer1803 (.A(net2207),
    .Y(net2208));
 BUFx2_ASAP7_75t_R rebuffer1804 (.A(net2207),
    .Y(net2209));
 BUFx2_ASAP7_75t_R rebuffer1805 (.A(net2207),
    .Y(net2210));
 BUFx4f_ASAP7_75t_R split1806 (.A(_10567_),
    .Y(net2211));
 BUFx2_ASAP7_75t_R rebuffer1807 (.A(_09895_),
    .Y(net2212));
 BUFx2_ASAP7_75t_R rebuffer1808 (.A(_09895_),
    .Y(net2213));
 BUFx2_ASAP7_75t_R rebuffer1809 (.A(_09895_),
    .Y(net2214));
 BUFx4f_ASAP7_75t_R rebuffer1810 (.A(net3170),
    .Y(net2215));
 BUFx4f_ASAP7_75t_R rebuffer1811 (.A(_09717_),
    .Y(net2216));
 BUFx2_ASAP7_75t_R rebuffer1812 (.A(net2216),
    .Y(net2217));
 BUFx3_ASAP7_75t_R rebuffer1813 (.A(_01821_),
    .Y(net2218));
 BUFx2_ASAP7_75t_R rebuffer1814 (.A(net2218),
    .Y(net2219));
 BUFx3_ASAP7_75t_R rebuffer1815 (.A(_05579_),
    .Y(net2220));
 BUFx2_ASAP7_75t_R rebuffer1816 (.A(net2220),
    .Y(net2221));
 BUFx4f_ASAP7_75t_R split1817 (.A(_10097_),
    .Y(net2222));
 BUFx12f_ASAP7_75t_R rebuffer1818 (.A(_05094_),
    .Y(net2223));
 BUFx2_ASAP7_75t_R rebuffer1819 (.A(net2223),
    .Y(net2224));
 BUFx2_ASAP7_75t_R rebuffer1820 (.A(net2223),
    .Y(net2225));
 BUFx4f_ASAP7_75t_R rebuffer1821 (.A(_05094_),
    .Y(net2226));
 BUFx2_ASAP7_75t_R split1822 (.A(_10586_),
    .Y(net2227));
 BUFx4f_ASAP7_75t_R split1823 (.A(_10515_),
    .Y(net2228));
 BUFx3_ASAP7_75t_R rebuffer1824 (.A(_05796_),
    .Y(net2229));
 BUFx2_ASAP7_75t_R rebuffer1825 (.A(_05796_),
    .Y(net2230));
 BUFx6f_ASAP7_75t_R rebuffer1826 (.A(_05747_),
    .Y(net2231));
 BUFx6f_ASAP7_75t_R rebuffer1827 (.A(net2231),
    .Y(net2232));
 BUFx3_ASAP7_75t_R split1828 (.A(_10468_),
    .Y(net2233));
 BUFx6f_ASAP7_75t_R split1829 (.A(_06050_),
    .Y(net2234));
 BUFx6f_ASAP7_75t_R split1830 (.A(_09998_),
    .Y(net2235));
 BUFx4f_ASAP7_75t_R rebuffer1831 (.A(_17815_),
    .Y(net2236));
 BUFx2_ASAP7_75t_R rebuffer1832 (.A(net2236),
    .Y(net2237));
 BUFx2_ASAP7_75t_R rebuffer1833 (.A(net2236),
    .Y(net2238));
 BUFx3_ASAP7_75t_R split1834 (.A(_01797_),
    .Y(net2239));
 BUFx2_ASAP7_75t_R rebuffer1835 (.A(_10358_),
    .Y(net2240));
 BUFx2_ASAP7_75t_R rebuffer1836 (.A(_10358_),
    .Y(net2241));
 BUFx4f_ASAP7_75t_R rebuffer1837 (.A(_06153_),
    .Y(net2242));
 BUFx2_ASAP7_75t_R rebuffer1838 (.A(_05444_),
    .Y(net2243));
 BUFx2_ASAP7_75t_R rebuffer1839 (.A(_18175_),
    .Y(net2244));
 BUFx2_ASAP7_75t_R rebuffer1840 (.A(_18175_),
    .Y(net2245));
 BUFx3_ASAP7_75t_R rebuffer1841 (.A(net2245),
    .Y(net2246));
 BUFx6f_ASAP7_75t_R rebuffer1842 (.A(_10498_),
    .Y(net2247));
 BUFx2_ASAP7_75t_R rebuffer1843 (.A(net2247),
    .Y(net2248));
 BUFx6f_ASAP7_75t_R rebuffer1844 (.A(_10498_),
    .Y(net2249));
 BUFx4f_ASAP7_75t_R split1845 (.A(_19171_),
    .Y(net2250));
 BUFx2_ASAP7_75t_R split1846 (.A(_18411_),
    .Y(net2251));
 BUFx4f_ASAP7_75t_R rebuffer1847 (.A(_10070_),
    .Y(net2252));
 BUFx2_ASAP7_75t_R rebuffer1848 (.A(net2252),
    .Y(net2253));
 BUFx12f_ASAP7_75t_R rebuffer1849 (.A(_01556_),
    .Y(net2254));
 BUFx2_ASAP7_75t_R rebuffer1850 (.A(net2254),
    .Y(net2255));
 BUFx6f_ASAP7_75t_R rebuffer1851 (.A(net2254),
    .Y(net2256));
 BUFx6f_ASAP7_75t_R rebuffer1852 (.A(net2256),
    .Y(net2257));
 BUFx12f_ASAP7_75t_R rebuffer1853 (.A(_21938_),
    .Y(net2258));
 BUFx2_ASAP7_75t_R rebuffer1854 (.A(net2258),
    .Y(net2259));
 BUFx2_ASAP7_75t_R rebuffer1855 (.A(_21938_),
    .Y(net2260));
 BUFx6f_ASAP7_75t_R rebuffer1856 (.A(net2260),
    .Y(net2261));
 BUFx2_ASAP7_75t_R rebuffer1857 (.A(_01949_),
    .Y(net2262));
 BUFx2_ASAP7_75t_R rebuffer1858 (.A(_01949_),
    .Y(net2263));
 BUFx2_ASAP7_75t_R rebuffer1859 (.A(_01949_),
    .Y(net2264));
 BUFx2_ASAP7_75t_R rebuffer1860 (.A(_02259_),
    .Y(net2265));
 BUFx2_ASAP7_75t_R rebuffer1861 (.A(_02259_),
    .Y(net2266));
 BUFx2_ASAP7_75t_R rebuffer1862 (.A(_02259_),
    .Y(net2267));
 BUFx3_ASAP7_75t_R rebuffer1863 (.A(_09692_),
    .Y(net2268));
 BUFx2_ASAP7_75t_R rebuffer1864 (.A(net2268),
    .Y(net2269));
 BUFx2_ASAP7_75t_R rebuffer1865 (.A(_05819_),
    .Y(net2270));
 BUFx3_ASAP7_75t_R split1866 (.A(_05819_),
    .Y(net2271));
 BUFx2_ASAP7_75t_R rebuffer1867 (.A(_05177_),
    .Y(net2272));
 BUFx2_ASAP7_75t_R rebuffer1868 (.A(net2272),
    .Y(net2273));
 BUFx2_ASAP7_75t_R rebuffer1869 (.A(_05177_),
    .Y(net2274));
 BUFx4f_ASAP7_75t_R split1870 (.A(_01603_),
    .Y(net2275));
 BUFx6f_ASAP7_75t_R rebuffer1871 (.A(_21502_),
    .Y(net2276));
 BUFx3_ASAP7_75t_R rebuffer1872 (.A(_16321_),
    .Y(net2277));
 BUFx3_ASAP7_75t_R rebuffer1873 (.A(_16321_),
    .Y(net2278));
 BUFx2_ASAP7_75t_R rebuffer1874 (.A(net2278),
    .Y(net2279));
 BUFx2_ASAP7_75t_R rebuffer1875 (.A(net2382),
    .Y(net2280));
 BUFx2_ASAP7_75t_R rebuffer1876 (.A(_09911_),
    .Y(net2281));
 BUFx6f_ASAP7_75t_R rebuffer1877 (.A(_09911_),
    .Y(net2282));
 BUFx2_ASAP7_75t_R rebuffer1878 (.A(net2282),
    .Y(net2283));
 BUFx2_ASAP7_75t_R rebuffer1879 (.A(net2282),
    .Y(net2284));
 BUFx2_ASAP7_75t_R rebuffer1880 (.A(_09911_),
    .Y(net2285));
 BUFx4f_ASAP7_75t_R split1881 (.A(_01892_),
    .Y(net2286));
 BUFx3_ASAP7_75t_R rebuffer1882 (.A(_00610_),
    .Y(net2287));
 BUFx2_ASAP7_75t_R rebuffer1883 (.A(_05805_),
    .Y(net2288));
 BUFx2_ASAP7_75t_R rebuffer1884 (.A(net3016),
    .Y(net2289));
 BUFx2_ASAP7_75t_R rebuffer1885 (.A(_09620_),
    .Y(net2290));
 BUFx6f_ASAP7_75t_R rebuffer1886 (.A(_09620_),
    .Y(net2291));
 BUFx2_ASAP7_75t_R rebuffer1887 (.A(_18695_),
    .Y(net2292));
 BUFx3_ASAP7_75t_R rebuffer1888 (.A(_22002_),
    .Y(net2293));
 BUFx2_ASAP7_75t_R rebuffer1889 (.A(net2293),
    .Y(net2294));
 BUFx2_ASAP7_75t_R rebuffer1890 (.A(_21879_),
    .Y(net2295));
 BUFx6f_ASAP7_75t_R rebuffer1891 (.A(_22002_),
    .Y(net2296));
 BUFx2_ASAP7_75t_R rebuffer1892 (.A(net2296),
    .Y(net2297));
 BUFx6f_ASAP7_75t_R rebuffer1893 (.A(_22002_),
    .Y(net2298));
 BUFx12f_ASAP7_75t_R rebuffer1894 (.A(_01773_),
    .Y(net2299));
 BUFx2_ASAP7_75t_R rebuffer1895 (.A(net2299),
    .Y(net2300));
 BUFx2_ASAP7_75t_R rebuffer1896 (.A(net2299),
    .Y(net2301));
 BUFx3_ASAP7_75t_R split1897 (.A(_18527_),
    .Y(net2302));
 BUFx4f_ASAP7_75t_R split1898 (.A(_18054_),
    .Y(net2303));
 BUFx3_ASAP7_75t_R split1899 (.A(_18695_),
    .Y(net2304));
 BUFx6f_ASAP7_75t_R rebuffer1900 (.A(_08946_),
    .Y(net2305));
 BUFx4f_ASAP7_75t_R rebuffer1901 (.A(_01836_),
    .Y(net2306));
 BUFx6f_ASAP7_75t_R rebuffer1902 (.A(_01836_),
    .Y(net2307));
 BUFx2_ASAP7_75t_R rebuffer1903 (.A(net3209),
    .Y(net2308));
 BUFx2_ASAP7_75t_R rebuffer1904 (.A(net3210),
    .Y(net2309));
 BUFx3_ASAP7_75t_R split1905 (.A(_13696_),
    .Y(net2310));
 BUFx6f_ASAP7_75t_R rebuffer1906 (.A(_00574_),
    .Y(net2311));
 BUFx3_ASAP7_75t_R rebuffer1907 (.A(_10578_),
    .Y(net2312));
 BUFx6f_ASAP7_75t_R rebuffer1908 (.A(net2312),
    .Y(net2313));
 BUFx2_ASAP7_75t_R rebuffer1909 (.A(_05165_),
    .Y(net2314));
 BUFx3_ASAP7_75t_R rebuffer1910 (.A(_05165_),
    .Y(net2315));
 BUFx6f_ASAP7_75t_R rebuffer1911 (.A(net3321),
    .Y(net2316));
 BUFx6f_ASAP7_75t_R rebuffer1912 (.A(_18723_),
    .Y(net2317));
 BUFx2_ASAP7_75t_R rebuffer1913 (.A(_05501_),
    .Y(net2318));
 BUFx2_ASAP7_75t_R rebuffer1914 (.A(_05501_),
    .Y(net2319));
 BUFx2_ASAP7_75t_R rebuffer1915 (.A(net2319),
    .Y(net2320));
 BUFx2_ASAP7_75t_R rebuffer1916 (.A(_06145_),
    .Y(net2321));
 BUFx2_ASAP7_75t_R rebuffer1917 (.A(_06145_),
    .Y(net2322));
 BUFx6f_ASAP7_75t_R rebuffer1918 (.A(_00589_),
    .Y(net2323));
 BUFx2_ASAP7_75t_R rebuffer1919 (.A(net2323),
    .Y(net2324));
 BUFx2_ASAP7_75t_R rebuffer1920 (.A(net2323),
    .Y(net2325));
 BUFx2_ASAP7_75t_R rebuffer1921 (.A(net2323),
    .Y(net2326));
 BUFx6f_ASAP7_75t_R rebuffer1922 (.A(_09717_),
    .Y(net2327));
 BUFx2_ASAP7_75t_R rebuffer1923 (.A(net2327),
    .Y(net2328));
 BUFx2_ASAP7_75t_R rebuffer1924 (.A(_10415_),
    .Y(net2329));
 BUFx3_ASAP7_75t_R split1925 (.A(_01890_),
    .Y(net2330));
 BUFx2_ASAP7_75t_R rebuffer1926 (.A(_10333_),
    .Y(net2331));
 BUFx2_ASAP7_75t_R rebuffer1927 (.A(_10333_),
    .Y(net2332));
 BUFx6f_ASAP7_75t_R rebuffer1928 (.A(_10333_),
    .Y(net2333));
 BUFx12f_ASAP7_75t_R rebuffer1929 (.A(_01532_),
    .Y(net2334));
 BUFx2_ASAP7_75t_R rebuffer1930 (.A(net2334),
    .Y(net2335));
 BUFx2_ASAP7_75t_R rebuffer1931 (.A(net2334),
    .Y(net2336));
 BUFx2_ASAP7_75t_R rebuffer1932 (.A(_22018_),
    .Y(net2337));
 BUFx6f_ASAP7_75t_R rebuffer1933 (.A(_00542_),
    .Y(net2338));
 BUFx12f_ASAP7_75t_R rebuffer1934 (.A(_09770_),
    .Y(net2339));
 BUFx2_ASAP7_75t_R rebuffer1935 (.A(net2339),
    .Y(net2340));
 BUFx6f_ASAP7_75t_R rebuffer1936 (.A(_21723_),
    .Y(net2341));
 BUFx6f_ASAP7_75t_R rebuffer1937 (.A(_21420_),
    .Y(net2342));
 BUFx2_ASAP7_75t_R rebuffer1938 (.A(_06158_),
    .Y(net2343));
 BUFx2_ASAP7_75t_R rebuffer1939 (.A(_06158_),
    .Y(net2344));
 BUFx2_ASAP7_75t_R rebuffer1940 (.A(net2344),
    .Y(net2345));
 BUFx2_ASAP7_75t_R rebuffer1941 (.A(_06158_),
    .Y(net2346));
 BUFx2_ASAP7_75t_R rebuffer1942 (.A(_19171_),
    .Y(net2347));
 BUFx4f_ASAP7_75t_R split1943 (.A(_01586_),
    .Y(net2348));
 BUFx3_ASAP7_75t_R rebuffer1944 (.A(_07287_),
    .Y(net2349));
 BUFx6f_ASAP7_75t_R rebuffer1945 (.A(_05479_),
    .Y(net2350));
 BUFx2_ASAP7_75t_R rebuffer1946 (.A(_10098_),
    .Y(net2351));
 BUFx6f_ASAP7_75t_R split1947 (.A(_01955_),
    .Y(net2352));
 BUFx10_ASAP7_75t_R split1948 (.A(_10086_),
    .Y(net2353));
 BUFx6f_ASAP7_75t_R rebuffer1949 (.A(_10451_),
    .Y(net2354));
 BUFx2_ASAP7_75t_R rebuffer1950 (.A(_10322_),
    .Y(net2355));
 BUFx3_ASAP7_75t_R rebuffer1951 (.A(_09914_),
    .Y(net2356));
 BUFx2_ASAP7_75t_R rebuffer1952 (.A(_09914_),
    .Y(net2357));
 BUFx6f_ASAP7_75t_R split1953 (.A(_09914_),
    .Y(net2358));
 BUFx2_ASAP7_75t_R rebuffer1954 (.A(_05743_),
    .Y(net2359));
 BUFx2_ASAP7_75t_R rebuffer1955 (.A(_05743_),
    .Y(net2360));
 BUFx12f_ASAP7_75t_R rebuffer1956 (.A(_01188_),
    .Y(net2361));
 BUFx4f_ASAP7_75t_R rebuffer1957 (.A(_01094_),
    .Y(net2362));
 BUFx6f_ASAP7_75t_R rebuffer1958 (.A(_21292_),
    .Y(net2363));
 BUFx4f_ASAP7_75t_R split1959 (.A(_17968_),
    .Y(net2364));
 BUFx6f_ASAP7_75t_R split1960 (.A(_21934_),
    .Y(net2365));
 BUFx6f_ASAP7_75t_R split1961 (.A(_01607_),
    .Y(net2366));
 BUFx2_ASAP7_75t_R rebuffer1962 (.A(_01607_),
    .Y(net2367));
 BUFx6f_ASAP7_75t_R rebuffer1963 (.A(_01607_),
    .Y(net2368));
 BUFx3_ASAP7_75t_R rebuffer1964 (.A(_01837_),
    .Y(net2369));
 BUFx2_ASAP7_75t_R rebuffer1965 (.A(net2369),
    .Y(net2370));
 BUFx2_ASAP7_75t_R rebuffer1966 (.A(_01837_),
    .Y(net2371));
 BUFx2_ASAP7_75t_R rebuffer1967 (.A(net2371),
    .Y(net2372));
 BUFx2_ASAP7_75t_R rebuffer1968 (.A(net2591),
    .Y(net2373));
 BUFx6f_ASAP7_75t_R rebuffer1969 (.A(_09890_),
    .Y(net2374));
 BUFx2_ASAP7_75t_R rebuffer1970 (.A(net2374),
    .Y(net2375));
 BUFx12f_ASAP7_75t_R rebuffer1971 (.A(_01521_),
    .Y(net2376));
 BUFx2_ASAP7_75t_R rebuffer1972 (.A(net2376),
    .Y(net2377));
 BUFx2_ASAP7_75t_R rebuffer1973 (.A(net2376),
    .Y(net2378));
 BUFx2_ASAP7_75t_R rebuffer1974 (.A(_01521_),
    .Y(net2379));
 BUFx2_ASAP7_75t_R rebuffer1975 (.A(net2379),
    .Y(net2380));
 BUFx2_ASAP7_75t_R rebuffer1976 (.A(net2380),
    .Y(net2381));
 BUFx12f_ASAP7_75t_R rebuffer1977 (.A(_10122_),
    .Y(net2382));
 BUFx2_ASAP7_75t_R rebuffer1978 (.A(net2382),
    .Y(net2383));
 BUFx4f_ASAP7_75t_R rebuffer1979 (.A(net3170),
    .Y(net2384));
 BUFx6f_ASAP7_75t_R rebuffer1980 (.A(_17645_),
    .Y(net2385));
 BUFx4f_ASAP7_75t_R split1981 (.A(_18594_),
    .Y(net2386));
 BUFx6f_ASAP7_75t_R rebuffer1982 (.A(_18527_),
    .Y(net2387));
 BUFx4f_ASAP7_75t_R rebuffer1983 (.A(net2387),
    .Y(net2388));
 BUFx12f_ASAP7_75t_R rebuffer1984 (.A(_05563_),
    .Y(net2389));
 BUFx2_ASAP7_75t_R rebuffer1985 (.A(net2389),
    .Y(net2390));
 BUFx6f_ASAP7_75t_R rebuffer1986 (.A(net2408),
    .Y(net2391));
 BUFx3_ASAP7_75t_R split1987 (.A(_01480_),
    .Y(net2392));
 BUFx2_ASAP7_75t_R rebuffer1988 (.A(_01194_),
    .Y(net2393));
 BUFx6f_ASAP7_75t_R split1989 (.A(_18714_),
    .Y(net2394));
 BUFx2_ASAP7_75t_R rebuffer1990 (.A(net2563),
    .Y(net2395));
 BUFx3_ASAP7_75t_R rebuffer1991 (.A(_03618_),
    .Y(net2396));
 BUFx4f_ASAP7_75t_R split1992 (.A(_09996_),
    .Y(net2397));
 BUFx3_ASAP7_75t_R rebuffer1993 (.A(_18532_),
    .Y(net2398));
 BUFx6f_ASAP7_75t_R split1994 (.A(_06104_),
    .Y(net2399));
 BUFx3_ASAP7_75t_R split1995 (.A(_05619_),
    .Y(net2400));
 BUFx6f_ASAP7_75t_R rebuffer1996 (.A(_05451_),
    .Y(net2401));
 BUFx3_ASAP7_75t_R rebuffer1997 (.A(_08946_),
    .Y(net2402));
 BUFx3_ASAP7_75t_R rebuffer1998 (.A(_06517_),
    .Y(net2403));
 BUFx2_ASAP7_75t_R rebuffer1999 (.A(_06517_),
    .Y(net2404));
 BUFx6f_ASAP7_75t_R split2000 (.A(_18721_),
    .Y(net2405));
 BUFx2_ASAP7_75t_R rebuffer2001 (.A(_01688_),
    .Y(net2406));
 BUFx3_ASAP7_75t_R rebuffer2002 (.A(_18239_),
    .Y(net2407));
 BUFx12f_ASAP7_75t_R rebuffer2003 (.A(_09996_),
    .Y(net2408));
 BUFx6f_ASAP7_75t_R rebuffer2004 (.A(net2408),
    .Y(net2409));
 BUFx2_ASAP7_75t_R rebuffer2005 (.A(_05626_),
    .Y(net2410));
 BUFx3_ASAP7_75t_R rebuffer2006 (.A(_05626_),
    .Y(net2411));
 BUFx6f_ASAP7_75t_R split2007 (.A(_06229_),
    .Y(net2412));
 BUFx2_ASAP7_75t_R rebuffer2008 (.A(net2545),
    .Y(net2413));
 BUFx12f_ASAP7_75t_R rebuffer2009 (.A(_18611_),
    .Y(net2414));
 BUFx2_ASAP7_75t_R rebuffer2010 (.A(net2414),
    .Y(net2415));
 BUFx3_ASAP7_75t_R split2011 (.A(_05805_),
    .Y(net2416));
 BUFx2_ASAP7_75t_R rebuffer2012 (.A(_05105_),
    .Y(net2417));
 BUFx2_ASAP7_75t_R rebuffer2013 (.A(_05105_),
    .Y(net2418));
 BUFx2_ASAP7_75t_R rebuffer2014 (.A(_18327_),
    .Y(net2419));
 BUFx6f_ASAP7_75t_R split2015 (.A(_21940_),
    .Y(net2420));
 BUFx6f_ASAP7_75t_R rebuffer2016 (.A(_18559_),
    .Y(net2421));
 BUFx6f_ASAP7_75t_R rebuffer2017 (.A(net2603),
    .Y(net2422));
 BUFx4f_ASAP7_75t_R split2018 (.A(_05879_),
    .Y(net2423));
 BUFx2_ASAP7_75t_R rebuffer2019 (.A(_01078_),
    .Y(net2424));
 BUFx6f_ASAP7_75t_R rebuffer2020 (.A(_01078_),
    .Y(net2425));
 BUFx3_ASAP7_75t_R rebuffer2021 (.A(_21917_),
    .Y(net2426));
 BUFx2_ASAP7_75t_R rebuffer2022 (.A(_21917_),
    .Y(net2427));
 BUFx3_ASAP7_75t_R rebuffer2023 (.A(_21212_),
    .Y(net2428));
 BUFx2_ASAP7_75t_R rebuffer2024 (.A(_09974_),
    .Y(net2429));
 BUFx2_ASAP7_75t_R rebuffer2025 (.A(_09974_),
    .Y(net2430));
 BUFx2_ASAP7_75t_R rebuffer2026 (.A(_09974_),
    .Y(net2431));
 BUFx2_ASAP7_75t_R rebuffer2027 (.A(_18144_),
    .Y(net2432));
 BUFx6f_ASAP7_75t_R split2028 (.A(_18594_),
    .Y(net2433));
 BUFx4f_ASAP7_75t_R split2029 (.A(_09739_),
    .Y(net2434));
 BUFx2_ASAP7_75t_R rebuffer2030 (.A(net2439),
    .Y(net2435));
 BUFx2_ASAP7_75t_R rebuffer2031 (.A(net2439),
    .Y(net2436));
 BUFx6f_ASAP7_75t_R split2032 (.A(_18322_),
    .Y(net2437));
 BUFx2_ASAP7_75t_R rebuffer2033 (.A(_18322_),
    .Y(net2438));
 BUFx6f_ASAP7_75t_R rebuffer2034 (.A(_18322_),
    .Y(net2439));
 BUFx2_ASAP7_75t_R rebuffer2035 (.A(net2439),
    .Y(net2440));
 BUFx6f_ASAP7_75t_R rebuffer2036 (.A(_10396_),
    .Y(net2441));
 BUFx6f_ASAP7_75t_R rebuffer2037 (.A(net2441),
    .Y(net2442));
 BUFx6f_ASAP7_75t_R split2038 (.A(_01179_),
    .Y(net2443));
 BUFx6f_ASAP7_75t_R rebuffer2039 (.A(_09908_),
    .Y(net2444));
 BUFx3_ASAP7_75t_R rebuffer2040 (.A(_09908_),
    .Y(net2445));
 BUFx3_ASAP7_75t_R split2041 (.A(_18144_),
    .Y(net2446));
 BUFx4f_ASAP7_75t_R rebuffer2042 (.A(_05616_),
    .Y(net2447));
 BUFx2_ASAP7_75t_R rebuffer2043 (.A(_10431_),
    .Y(net2448));
 BUFx2_ASAP7_75t_R rebuffer2044 (.A(_10431_),
    .Y(net2449));
 BUFx2_ASAP7_75t_R rebuffer2045 (.A(_10431_),
    .Y(net2450));
 BUFx3_ASAP7_75t_R split2046 (.A(_17665_),
    .Y(net2451));
 BUFx6f_ASAP7_75t_R split2047 (.A(_18316_),
    .Y(net2452));
 BUFx6f_ASAP7_75t_R split2048 (.A(_09717_),
    .Y(net2453));
 BUFx6f_ASAP7_75t_R rebuffer2049 (.A(_10385_),
    .Y(net2454));
 BUFx2_ASAP7_75t_R rebuffer2050 (.A(net2454),
    .Y(net2455));
 BUFx6f_ASAP7_75t_R rebuffer2051 (.A(_10385_),
    .Y(net2456));
 BUFx3_ASAP7_75t_R rebuffer2052 (.A(net2713),
    .Y(net2457));
 BUFx4f_ASAP7_75t_R rebuffer2053 (.A(_01894_),
    .Y(net2458));
 BUFx2_ASAP7_75t_R rebuffer2054 (.A(net2458),
    .Y(net2459));
 BUFx4f_ASAP7_75t_R split2055 (.A(_01322_),
    .Y(net2460));
 BUFx3_ASAP7_75t_R rebuffer2056 (.A(_05634_),
    .Y(net2461));
 BUFx6f_ASAP7_75t_R rebuffer2057 (.A(net2461),
    .Y(net2462));
 BUFx4f_ASAP7_75t_R split2058 (.A(_10449_),
    .Y(net2463));
 BUFx4f_ASAP7_75t_R rebuffer2059 (.A(_10454_),
    .Y(net2464));
 BUFx2_ASAP7_75t_R rebuffer2060 (.A(net2464),
    .Y(net2465));
 BUFx3_ASAP7_75t_R rebuffer2061 (.A(net2713),
    .Y(net2466));
 BUFx2_ASAP7_75t_R rebuffer2062 (.A(_00621_),
    .Y(net2467));
 BUFx6f_ASAP7_75t_R rebuffer2063 (.A(_00621_),
    .Y(net2468));
 BUFx2_ASAP7_75t_R rebuffer2064 (.A(net2468),
    .Y(net2469));
 BUFx6f_ASAP7_75t_R rebuffer2065 (.A(_09889_),
    .Y(net2470));
 BUFx2_ASAP7_75t_R rebuffer2066 (.A(_08771_),
    .Y(net2471));
 BUFx2_ASAP7_75t_R rebuffer2067 (.A(net2471),
    .Y(net2472));
 BUFx6f_ASAP7_75t_R split2068 (.A(_18283_),
    .Y(net2473));
 BUFx6f_ASAP7_75t_R rebuffer2069 (.A(_00607_),
    .Y(net2474));
 BUFx2_ASAP7_75t_R rebuffer2070 (.A(_00607_),
    .Y(net2475));
 BUFx2_ASAP7_75t_R rebuffer2071 (.A(_18283_),
    .Y(net2476));
 BUFx3_ASAP7_75t_R rebuffer2072 (.A(_05486_),
    .Y(net2477));
 BUFx2_ASAP7_75t_R rebuffer2073 (.A(net2477),
    .Y(net2478));
 BUFx6f_ASAP7_75t_R split2074 (.A(_18545_),
    .Y(net2479));
 BUFx2_ASAP7_75t_R split2075 (.A(_06153_),
    .Y(net2480));
 BUFx3_ASAP7_75t_R rebuffer2076 (.A(_09585_),
    .Y(net2481));
 BUFx3_ASAP7_75t_R split2077 (.A(_06213_),
    .Y(net2482));
 BUFx3_ASAP7_75t_R rebuffer2078 (.A(_05985_),
    .Y(net2483));
 BUFx6f_ASAP7_75t_R split2079 (.A(_17641_),
    .Y(net2484));
 BUFx6f_ASAP7_75t_R split2080 (.A(_05860_),
    .Y(net2485));
 BUFx6f_ASAP7_75t_R rebuffer2081 (.A(_00597_),
    .Y(net2486));
 BUFx2_ASAP7_75t_R rebuffer2082 (.A(net2486),
    .Y(net2487));
 BUFx3_ASAP7_75t_R rebuffer2083 (.A(net2894),
    .Y(net2488));
 BUFx4f_ASAP7_75t_R rebuffer2084 (.A(_05746_),
    .Y(net2489));
 BUFx2_ASAP7_75t_R rebuffer2085 (.A(_05746_),
    .Y(net2490));
 BUFx4f_ASAP7_75t_R rebuffer2086 (.A(_10430_),
    .Y(net2491));
 BUFx2_ASAP7_75t_R rebuffer2087 (.A(_16560_),
    .Y(net2492));
 BUFx4f_ASAP7_75t_R split2088 (.A(_05079_),
    .Y(net2493));
 BUFx3_ASAP7_75t_R split2089 (.A(_01863_),
    .Y(net2494));
 BUFx3_ASAP7_75t_R rebuffer2090 (.A(_21893_),
    .Y(net2495));
 BUFx2_ASAP7_75t_R rebuffer2091 (.A(net2495),
    .Y(net2496));
 BUFx2_ASAP7_75t_R rebuffer2092 (.A(_21893_),
    .Y(net2497));
 BUFx12f_ASAP7_75t_R rebuffer2093 (.A(_18290_),
    .Y(net2498));
 BUFx2_ASAP7_75t_R rebuffer2094 (.A(net2498),
    .Y(net2499));
 BUFx2_ASAP7_75t_R rebuffer2095 (.A(net2498),
    .Y(net2500));
 BUFx6f_ASAP7_75t_R rebuffer2096 (.A(_09655_),
    .Y(net2501));
 BUFx3_ASAP7_75t_R rebuffer2097 (.A(_09655_),
    .Y(net2502));
 BUFx2_ASAP7_75t_R split2098 (.A(_09611_),
    .Y(net2503));
 BUFx2_ASAP7_75t_R split2099 (.A(_18643_),
    .Y(net2504));
 BUFx6f_ASAP7_75t_R rebuffer2100 (.A(_19171_),
    .Y(net2505));
 BUFx2_ASAP7_75t_R rebuffer2101 (.A(net2505),
    .Y(net2506));
 BUFx12f_ASAP7_75t_R rebuffer2102 (.A(_06049_),
    .Y(net2507));
 BUFx2_ASAP7_75t_R rebuffer2103 (.A(net2507),
    .Y(net2508));
 BUFx6f_ASAP7_75t_R split2104 (.A(_05497_),
    .Y(net2509));
 BUFx4f_ASAP7_75t_R split2105 (.A(_22018_),
    .Y(net2510));
 BUFx2_ASAP7_75t_R rebuffer2106 (.A(net2661),
    .Y(net2511));
 BUFx3_ASAP7_75t_R rebuffer2107 (.A(_22015_),
    .Y(net2512));
 BUFx3_ASAP7_75t_R rebuffer2108 (.A(net2512),
    .Y(net2513));
 BUFx3_ASAP7_75t_R rebuffer2109 (.A(_10877_),
    .Y(net2514));
 BUFx2_ASAP7_75t_R rebuffer2110 (.A(_10877_),
    .Y(net2515));
 BUFx2_ASAP7_75t_R rebuffer2111 (.A(net2515),
    .Y(net2516));
 BUFx2_ASAP7_75t_R rebuffer2112 (.A(_05758_),
    .Y(net2517));
 BUFx2_ASAP7_75t_R rebuffer2113 (.A(_05758_),
    .Y(net2518));
 BUFx2_ASAP7_75t_R rebuffer2114 (.A(_05758_),
    .Y(net2519));
 BUFx2_ASAP7_75t_R rebuffer2115 (.A(_05938_),
    .Y(net2520));
 BUFx2_ASAP7_75t_R rebuffer2116 (.A(_05938_),
    .Y(net2521));
 BUFx6f_ASAP7_75t_R split2117 (.A(_01146_),
    .Y(net2522));
 BUFx6f_ASAP7_75t_R split2118 (.A(_02692_),
    .Y(net2523));
 BUFx6f_ASAP7_75t_R split2119 (.A(_01670_),
    .Y(net2524));
 BUFx6f_ASAP7_75t_R split2120 (.A(_05993_),
    .Y(net2525));
 BUFx3_ASAP7_75t_R split2121 (.A(_10600_),
    .Y(net2526));
 BUFx2_ASAP7_75t_R rebuffer2122 (.A(_18581_),
    .Y(net2527));
 BUFx3_ASAP7_75t_R rebuffer2123 (.A(_21467_),
    .Y(net2528));
 BUFx4f_ASAP7_75t_R split2124 (.A(_05174_),
    .Y(net2529));
 BUFx3_ASAP7_75t_R rebuffer2125 (.A(_06072_),
    .Y(net2530));
 BUFx2_ASAP7_75t_R rebuffer2126 (.A(net2530),
    .Y(net2531));
 BUFx4f_ASAP7_75t_R split2127 (.A(_17593_),
    .Y(net2532));
 BUFx3_ASAP7_75t_R split2128 (.A(_18281_),
    .Y(net2533));
 BUFx6f_ASAP7_75t_R rebuffer2129 (.A(_00606_),
    .Y(net2534));
 BUFx4f_ASAP7_75t_R split2130 (.A(_10098_),
    .Y(net2535));
 BUFx2_ASAP7_75t_R split2131 (.A(_10415_),
    .Y(net2536));
 BUFx4f_ASAP7_75t_R split2132 (.A(_20170_),
    .Y(net2537));
 BUFx3_ASAP7_75t_R rebuffer2133 (.A(_02363_),
    .Y(net2538));
 BUFx3_ASAP7_75t_R rebuffer2134 (.A(net2538),
    .Y(net2539));
 BUFx12f_ASAP7_75t_R rebuffer2135 (.A(_05775_),
    .Y(net2540));
 BUFx2_ASAP7_75t_R rebuffer2136 (.A(net2540),
    .Y(net2541));
 BUFx6f_ASAP7_75t_R rebuffer2137 (.A(net2540),
    .Y(net2542));
 BUFx2_ASAP7_75t_R rebuffer2138 (.A(net2542),
    .Y(net2543));
 BUFx6f_ASAP7_75t_R rebuffer2139 (.A(_01172_),
    .Y(net2544));
 BUFx6f_ASAP7_75t_R rebuffer2140 (.A(_18682_),
    .Y(net2545));
 BUFx2_ASAP7_75t_R rebuffer2141 (.A(net2545),
    .Y(net2546));
 BUFx4f_ASAP7_75t_R split2142 (.A(_09692_),
    .Y(net2547));
 BUFx12f_ASAP7_75t_R rebuffer2143 (.A(_05490_),
    .Y(net2548));
 BUFx3_ASAP7_75t_R split2144 (.A(_01926_),
    .Y(net2549));
 BUFx2_ASAP7_75t_R rebuffer2145 (.A(_09574_),
    .Y(net2550));
 BUFx2_ASAP7_75t_R rebuffer2146 (.A(net2550),
    .Y(net2551));
 BUFx6f_ASAP7_75t_R rebuffer2147 (.A(_09574_),
    .Y(net2552));
 BUFx2_ASAP7_75t_R rebuffer2148 (.A(net2552),
    .Y(net2553));
 BUFx2_ASAP7_75t_R rebuffer2149 (.A(net2553),
    .Y(net2554));
 BUFx4f_ASAP7_75t_R split2150 (.A(_18565_),
    .Y(net2555));
 BUFx3_ASAP7_75t_R split2151 (.A(_22028_),
    .Y(net2556));
 BUFx6f_ASAP7_75t_R rebuffer2152 (.A(_17974_),
    .Y(net2557));
 BUFx3_ASAP7_75t_R rebuffer2153 (.A(_09717_),
    .Y(net2558));
 BUFx2_ASAP7_75t_R rebuffer2154 (.A(_09922_),
    .Y(net2559));
 BUFx6f_ASAP7_75t_R split2155 (.A(_01965_),
    .Y(net2560));
 BUFx4f_ASAP7_75t_R rebuffer2156 (.A(_10365_),
    .Y(net2561));
 BUFx2_ASAP7_75t_R rebuffer2157 (.A(net2561),
    .Y(net2562));
 BUFx6f_ASAP7_75t_R split2158 (.A(_01819_),
    .Y(net2563));
 BUFx4f_ASAP7_75t_R rebuffer2159 (.A(_00653_),
    .Y(net2564));
 BUFx2_ASAP7_75t_R rebuffer2160 (.A(net2564),
    .Y(net2565));
 BUFx4f_ASAP7_75t_R split2161 (.A(_10339_),
    .Y(net2566));
 BUFx2_ASAP7_75t_R rebuffer2162 (.A(_05579_),
    .Y(net2567));
 BUFx2_ASAP7_75t_R rebuffer2163 (.A(_05579_),
    .Y(net2568));
 BUFx6f_ASAP7_75t_R rebuffer2164 (.A(_05754_),
    .Y(net2569));
 BUFx6f_ASAP7_75t_R rebuffer2165 (.A(net2572),
    .Y(net2570));
 BUFx2_ASAP7_75t_R rebuffer2166 (.A(net2570),
    .Y(net2571));
 BUFx12f_ASAP7_75t_R rebuffer2167 (.A(_01577_),
    .Y(net2572));
 BUFx2_ASAP7_75t_R rebuffer2168 (.A(_02467_),
    .Y(net2573));
 BUFx2_ASAP7_75t_R rebuffer2169 (.A(_02467_),
    .Y(net2574));
 BUFx3_ASAP7_75t_R rebuffer2170 (.A(_11566_),
    .Y(net2575));
 BUFx2_ASAP7_75t_R rebuffer2171 (.A(net2575),
    .Y(net2576));
 BUFx6f_ASAP7_75t_R rebuffer2172 (.A(_01194_),
    .Y(net2577));
 BUFx2_ASAP7_75t_R rebuffer2173 (.A(_18604_),
    .Y(net2578));
 BUFx2_ASAP7_75t_R rebuffer2174 (.A(net2578),
    .Y(net2579));
 BUFx4f_ASAP7_75t_R rebuffer2175 (.A(_18604_),
    .Y(net2580));
 BUFx2_ASAP7_75t_R rebuffer2176 (.A(_12126_),
    .Y(net2581));
 BUFx3_ASAP7_75t_R split2177 (.A(_07287_),
    .Y(net2582));
 BUFx6f_ASAP7_75t_R rebuffer2178 (.A(_10097_),
    .Y(net2583));
 BUFx6f_ASAP7_75t_R rebuffer2179 (.A(_09971_),
    .Y(net2584));
 BUFx2_ASAP7_75t_R rebuffer2180 (.A(_01589_),
    .Y(net2585));
 BUFx3_ASAP7_75t_R split2181 (.A(_06046_),
    .Y(net2586));
 BUFx4f_ASAP7_75t_R rebuffer2182 (.A(_16275_),
    .Y(net2587));
 BUFx2_ASAP7_75t_R rebuffer2183 (.A(net2587),
    .Y(net2588));
 BUFx2_ASAP7_75t_R split2184 (.A(_21919_),
    .Y(net2589));
 BUFx4f_ASAP7_75t_R split2185 (.A(_06182_),
    .Y(net2590));
 BUFx3_ASAP7_75t_R split2186 (.A(_09893_),
    .Y(net2591));
 BUFx2_ASAP7_75t_R rebuffer2187 (.A(_13842_),
    .Y(net2592));
 BUFx2_ASAP7_75t_R rebuffer2188 (.A(net2592),
    .Y(net2593));
 BUFx2_ASAP7_75t_R rebuffer2189 (.A(net2592),
    .Y(net2594));
 BUFx4f_ASAP7_75t_R split2190 (.A(_18490_),
    .Y(net2595));
 BUFx2_ASAP7_75t_R rebuffer2191 (.A(net3287),
    .Y(net2596));
 BUFx2_ASAP7_75t_R rebuffer2192 (.A(_17687_),
    .Y(net2597));
 BUFx6f_ASAP7_75t_R rebuffer2193 (.A(_17687_),
    .Y(net2598));
 BUFx4f_ASAP7_75t_R rebuffer2194 (.A(net2598),
    .Y(net2599));
 BUFx2_ASAP7_75t_R rebuffer2195 (.A(net2598),
    .Y(net2600));
 BUFx2_ASAP7_75t_R rebuffer2196 (.A(_18281_),
    .Y(net2601));
 BUFx6f_ASAP7_75t_R rebuffer2197 (.A(_18281_),
    .Y(net2602));
 BUFx12f_ASAP7_75t_R rebuffer2198 (.A(_05879_),
    .Y(net2603));
 BUFx2_ASAP7_75t_R rebuffer2199 (.A(net2603),
    .Y(net2604));
 BUFx6f_ASAP7_75t_R rebuffer2200 (.A(_09801_),
    .Y(net2605));
 BUFx2_ASAP7_75t_R rebuffer2201 (.A(net2605),
    .Y(net2606));
 BUFx2_ASAP7_75t_R rebuffer2202 (.A(net2605),
    .Y(net2607));
 BUFx2_ASAP7_75t_R rebuffer2203 (.A(_21937_),
    .Y(net2608));
 BUFx4f_ASAP7_75t_R split2204 (.A(_06375_),
    .Y(net2609));
 BUFx3_ASAP7_75t_R split2205 (.A(net1084),
    .Y(net2610));
 BUFx6f_ASAP7_75t_R rebuffer2206 (.A(_05532_),
    .Y(net2611));
 BUFx2_ASAP7_75t_R rebuffer2207 (.A(net2611),
    .Y(net2612));
 BUFx2_ASAP7_75t_R rebuffer2208 (.A(net2611),
    .Y(net2613));
 BUFx6f_ASAP7_75t_R rebuffer2209 (.A(_06182_),
    .Y(net2614));
 BUFx2_ASAP7_75t_R split2210 (.A(_18604_),
    .Y(net2615));
 BUFx12f_ASAP7_75t_R rebuffer2211 (.A(_05640_),
    .Y(net2616));
 BUFx6f_ASAP7_75t_R rebuffer2212 (.A(net2616),
    .Y(net2617));
 BUFx4f_ASAP7_75t_R rebuffer2213 (.A(_05640_),
    .Y(net2618));
 BUFx6f_ASAP7_75t_R split2214 (.A(_01778_),
    .Y(net2619));
 BUFx2_ASAP7_75t_R rebuffer2215 (.A(_18641_),
    .Y(net2620));
 BUFx3_ASAP7_75t_R split2216 (.A(_05107_),
    .Y(net2621));
 BUFx2_ASAP7_75t_R rebuffer2217 (.A(_16318_),
    .Y(net2622));
 BUFx6f_ASAP7_75t_R rebuffer2218 (.A(_00637_),
    .Y(net2623));
 BUFx2_ASAP7_75t_R rebuffer2219 (.A(net2623),
    .Y(net2624));
 BUFx2_ASAP7_75t_R rebuffer2220 (.A(net2623),
    .Y(net2625));
 BUFx2_ASAP7_75t_R split2221 (.A(_18723_),
    .Y(net2626));
 BUFx3_ASAP7_75t_R split2222 (.A(_10161_),
    .Y(net2627));
 BUFx2_ASAP7_75t_R rebuffer2223 (.A(_10106_),
    .Y(net2628));
 BUFx2_ASAP7_75t_R rebuffer2224 (.A(_10106_),
    .Y(net2629));
 BUFx6f_ASAP7_75t_R split2225 (.A(_17551_),
    .Y(net2630));
 BUFx4f_ASAP7_75t_R split2226 (.A(_18581_),
    .Y(net2631));
 BUFx2_ASAP7_75t_R rebuffer2227 (.A(_18569_),
    .Y(net2632));
 BUFx6f_ASAP7_75t_R split2228 (.A(_18685_),
    .Y(net2633));
 BUFx4f_ASAP7_75t_R split2229 (.A(_18357_),
    .Y(net2634));
 BUFx4f_ASAP7_75t_R rebuffer2230 (.A(_18357_),
    .Y(net2635));
 BUFx6f_ASAP7_75t_R split2231 (.A(_05966_),
    .Y(net2636));
 BUFx2_ASAP7_75t_R rebuffer2232 (.A(_21925_),
    .Y(net2637));
 BUFx6f_ASAP7_75t_R split2233 (.A(_18383_),
    .Y(net2638));
 BUFx6f_ASAP7_75t_R split2234 (.A(_06131_),
    .Y(net2639));
 BUFx6f_ASAP7_75t_R rebuffer2235 (.A(_17616_),
    .Y(net2640));
 BUFx3_ASAP7_75t_R rebuffer2236 (.A(net2640),
    .Y(net2641));
 BUFx2_ASAP7_75t_R rebuffer2237 (.A(net2640),
    .Y(net2642));
 BUFx6f_ASAP7_75t_R rebuffer2238 (.A(_05131_),
    .Y(net2643));
 BUFx6f_ASAP7_75t_R rebuffer2239 (.A(net2643),
    .Y(net2644));
 BUFx3_ASAP7_75t_R rebuffer2240 (.A(_05131_),
    .Y(net2645));
 BUFx6f_ASAP7_75t_R rebuffer2241 (.A(_03618_),
    .Y(net2646));
 BUFx6f_ASAP7_75t_R rebuffer2242 (.A(_00590_),
    .Y(net2647));
 BUFx6f_ASAP7_75t_R rebuffer2243 (.A(net2647),
    .Y(net2648));
 BUFx2_ASAP7_75t_R rebuffer2244 (.A(net2648),
    .Y(net2649));
 BUFx2_ASAP7_75t_R rebuffer2245 (.A(_00590_),
    .Y(net2650));
 BUFx10_ASAP7_75t_R rebuffer2246 (.A(_01115_),
    .Y(net2651));
 BUFx6f_ASAP7_75t_R rebuffer2247 (.A(net2651),
    .Y(net2652));
 BUFx6f_ASAP7_75t_R rebuffer2248 (.A(_01916_),
    .Y(net2653));
 BUFx2_ASAP7_75t_R rebuffer2249 (.A(_02544_),
    .Y(net2654));
 BUFx2_ASAP7_75t_R rebuffer2250 (.A(net2654),
    .Y(net2655));
 BUFx4f_ASAP7_75t_R rebuffer2251 (.A(_09594_),
    .Y(net2656));
 BUFx2_ASAP7_75t_R rebuffer2252 (.A(net3113),
    .Y(net2657));
 BUFx4f_ASAP7_75t_R split2253 (.A(_05508_),
    .Y(net2658));
 BUFx2_ASAP7_75t_R rebuffer2254 (.A(_05503_),
    .Y(net2659));
 BUFx4f_ASAP7_75t_R split2255 (.A(_09922_),
    .Y(net2660));
 BUFx6f_ASAP7_75t_R split2256 (.A(_05514_),
    .Y(net2661));
 BUFx6f_ASAP7_75t_R split2257 (.A(_10040_),
    .Y(net2662));
 BUFx3_ASAP7_75t_R split2258 (.A(_05451_),
    .Y(net2663));
 BUFx2_ASAP7_75t_R rebuffer2259 (.A(net3493),
    .Y(net2664));
 BUFx2_ASAP7_75t_R rebuffer2260 (.A(net3493),
    .Y(net2665));
 BUFx2_ASAP7_75t_R rebuffer2261 (.A(net3493),
    .Y(net2666));
 BUFx2_ASAP7_75t_R rebuffer2262 (.A(_09945_),
    .Y(net2667));
 BUFx2_ASAP7_75t_R rebuffer2263 (.A(_18270_),
    .Y(net2668));
 BUFx2_ASAP7_75t_R rebuffer2264 (.A(_18270_),
    .Y(net2669));
 BUFx3_ASAP7_75t_R rebuffer2265 (.A(_05485_),
    .Y(net2670));
 BUFx3_ASAP7_75t_R split2266 (.A(_18239_),
    .Y(net2671));
 BUFx3_ASAP7_75t_R rebuffer2267 (.A(_03001_),
    .Y(net2672));
 BUFx2_ASAP7_75t_R rebuffer2268 (.A(net2672),
    .Y(net2673));
 BUFx2_ASAP7_75t_R rebuffer2269 (.A(net2672),
    .Y(net2674));
 BUFx2_ASAP7_75t_R rebuffer2270 (.A(net2674),
    .Y(net2675));
 BUFx3_ASAP7_75t_R rebuffer2271 (.A(_00565_),
    .Y(net2676));
 BUFx3_ASAP7_75t_R rebuffer2272 (.A(_00565_),
    .Y(net2677));
 BUFx2_ASAP7_75t_R rebuffer2273 (.A(_00565_),
    .Y(net2678));
 BUFx4f_ASAP7_75t_R split2274 (.A(_05854_),
    .Y(net2679));
 BUFx3_ASAP7_75t_R split2275 (.A(_18107_),
    .Y(net2680));
 BUFx12f_ASAP7_75t_R rebuffer2276 (.A(_10300_),
    .Y(net2681));
 BUFx2_ASAP7_75t_R rebuffer2277 (.A(net2681),
    .Y(net2682));
 BUFx2_ASAP7_75t_R rebuffer2278 (.A(net2681),
    .Y(net2683));
 BUFx2_ASAP7_75t_R rebuffer2279 (.A(_01807_),
    .Y(net2684));
 BUFx2_ASAP7_75t_R rebuffer2280 (.A(_01807_),
    .Y(net2685));
 BUFx2_ASAP7_75t_R rebuffer2281 (.A(_09612_),
    .Y(net2686));
 BUFx2_ASAP7_75t_R rebuffer2282 (.A(_09612_),
    .Y(net2687));
 BUFx3_ASAP7_75t_R rebuffer2283 (.A(net2687),
    .Y(net2688));
 BUFx6f_ASAP7_75t_R rebuffer2284 (.A(_01360_),
    .Y(net2689));
 BUFx3_ASAP7_75t_R split2285 (.A(_18524_),
    .Y(net2690));
 BUFx3_ASAP7_75t_R rebuffer2286 (.A(_09695_),
    .Y(net2691));
 BUFx2_ASAP7_75t_R rebuffer2287 (.A(_09695_),
    .Y(net2692));
 BUFx2_ASAP7_75t_R rebuffer2288 (.A(_18729_),
    .Y(net2693));
 BUFx6f_ASAP7_75t_R rebuffer2289 (.A(_18729_),
    .Y(net2694));
 BUFx3_ASAP7_75t_R rebuffer2290 (.A(_10420_),
    .Y(net2695));
 BUFx6f_ASAP7_75t_R rebuffer2291 (.A(_00561_),
    .Y(net2696));
 BUFx2_ASAP7_75t_R rebuffer2292 (.A(net2696),
    .Y(net2697));
 BUFx6f_ASAP7_75t_R rebuffer2293 (.A(_05447_),
    .Y(net2698));
 BUFx6f_ASAP7_75t_R split2294 (.A(_18357_),
    .Y(net2699));
 BUFx4f_ASAP7_75t_R split2295 (.A(_03193_),
    .Y(net2700));
 BUFx4f_ASAP7_75t_R rebuffer2296 (.A(_18411_),
    .Y(net2701));
 BUFx3_ASAP7_75t_R rebuffer2297 (.A(_05656_),
    .Y(net2702));
 BUFx3_ASAP7_75t_R rebuffer2298 (.A(_05535_),
    .Y(net2703));
 BUFx2_ASAP7_75t_R rebuffer2299 (.A(_00541_),
    .Y(net2704));
 BUFx2_ASAP7_75t_R rebuffer2300 (.A(_00541_),
    .Y(net2705));
 BUFx3_ASAP7_75t_R rebuffer2301 (.A(net2705),
    .Y(net2706));
 BUFx6f_ASAP7_75t_R rebuffer2302 (.A(_01797_),
    .Y(net2707));
 BUFx2_ASAP7_75t_R rebuffer2303 (.A(net2707),
    .Y(net2708));
 BUFx2_ASAP7_75t_R rebuffer2304 (.A(net2707),
    .Y(net2709));
 BUFx4f_ASAP7_75t_R rebuffer2305 (.A(_01987_),
    .Y(net2710));
 BUFx6f_ASAP7_75t_R rebuffer2306 (.A(_00582_),
    .Y(net2711));
 BUFx2_ASAP7_75t_R rebuffer2307 (.A(net2711),
    .Y(net2712));
 BUFx6f_ASAP7_75t_R rebuffer2308 (.A(_18283_),
    .Y(net2713));
 BUFx2_ASAP7_75t_R rebuffer2309 (.A(_10350_),
    .Y(net2714));
 BUFx3_ASAP7_75t_R rebuffer2310 (.A(_10350_),
    .Y(net2715));
 BUFx2_ASAP7_75t_R rebuffer2311 (.A(net2715),
    .Y(net2716));
 BUFx2_ASAP7_75t_R rebuffer2312 (.A(_01172_),
    .Y(net2717));
 BUFx2_ASAP7_75t_R rebuffer2313 (.A(_18036_),
    .Y(net2718));
 BUFx3_ASAP7_75t_R rebuffer2314 (.A(_18036_),
    .Y(net2719));
 BUFx2_ASAP7_75t_R rebuffer2315 (.A(net2719),
    .Y(net2720));
 BUFx2_ASAP7_75t_R rebuffer2316 (.A(_14630_),
    .Y(net2721));
 BUFx2_ASAP7_75t_R rebuffer2317 (.A(_14630_),
    .Y(net2722));
 BUFx4f_ASAP7_75t_R split2318 (.A(_01172_),
    .Y(net2723));
 BUFx2_ASAP7_75t_R rebuffer2319 (.A(_09684_),
    .Y(net2724));
 BUFx2_ASAP7_75t_R rebuffer2320 (.A(_17955_),
    .Y(net2725));
 BUFx6f_ASAP7_75t_R rebuffer2321 (.A(_00581_),
    .Y(net2726));
 BUFx6f_ASAP7_75t_R rebuffer2322 (.A(_00569_),
    .Y(net2727));
 BUFx2_ASAP7_75t_R rebuffer2323 (.A(_01496_),
    .Y(net2728));
 BUFx2_ASAP7_75t_R rebuffer2324 (.A(net2728),
    .Y(net2729));
 BUFx2_ASAP7_75t_R rebuffer2325 (.A(net3092),
    .Y(net2730));
 BUFx3_ASAP7_75t_R rebuffer2326 (.A(_01318_),
    .Y(net2731));
 BUFx4f_ASAP7_75t_R split2327 (.A(_09714_),
    .Y(net2732));
 BUFx4f_ASAP7_75t_R split2328 (.A(_01675_),
    .Y(net2733));
 BUFx2_ASAP7_75t_R rebuffer2329 (.A(_09928_),
    .Y(net2734));
 BUFx2_ASAP7_75t_R rebuffer2330 (.A(_19057_),
    .Y(net2735));
 BUFx3_ASAP7_75t_R rebuffer2331 (.A(_05887_),
    .Y(net2736));
 BUFx2_ASAP7_75t_R rebuffer2332 (.A(_05887_),
    .Y(net2737));
 BUFx2_ASAP7_75t_R rebuffer2333 (.A(net2737),
    .Y(net2738));
 BUFx6f_ASAP7_75t_R rebuffer2334 (.A(_05737_),
    .Y(net2739));
 BUFx2_ASAP7_75t_R rebuffer2335 (.A(_05528_),
    .Y(net2740));
 BUFx6f_ASAP7_75t_R rebuffer2336 (.A(_00572_),
    .Y(net2741));
 BUFx2_ASAP7_75t_R rebuffer2337 (.A(net2741),
    .Y(net2742));
 BUFx6f_ASAP7_75t_R split2338 (.A(_05857_),
    .Y(net2743));
 BUFx6f_ASAP7_75t_R split2339 (.A(_06071_),
    .Y(net2744));
 BUFx3_ASAP7_75t_R rebuffer2340 (.A(_10328_),
    .Y(net2745));
 BUFx4f_ASAP7_75t_R split2341 (.A(_01636_),
    .Y(net2746));
 BUFx2_ASAP7_75t_R rebuffer2342 (.A(_18305_),
    .Y(net2747));
 BUFx6f_ASAP7_75t_R rebuffer2343 (.A(_18305_),
    .Y(net2748));
 BUFx2_ASAP7_75t_R rebuffer2344 (.A(_00642_),
    .Y(net2749));
 BUFx2_ASAP7_75t_R rebuffer2345 (.A(_00642_),
    .Y(net2750));
 BUFx2_ASAP7_75t_R rebuffer2346 (.A(_00642_),
    .Y(net2751));
 BUFx4f_ASAP7_75t_R split2347 (.A(_21967_),
    .Y(net2752));
 BUFx3_ASAP7_75t_R rebuffer2348 (.A(_18357_),
    .Y(net2753));
 BUFx2_ASAP7_75t_R rebuffer2349 (.A(_18254_),
    .Y(net2754));
 BUFx3_ASAP7_75t_R split2350 (.A(_05528_),
    .Y(net2755));
 BUFx2_ASAP7_75t_R rebuffer2351 (.A(_07297_),
    .Y(net2756));
 BUFx6f_ASAP7_75t_R split2352 (.A(_18081_),
    .Y(net2757));
 BUFx3_ASAP7_75t_R rebuffer2353 (.A(_17770_),
    .Y(net2758));
 BUFx2_ASAP7_75t_R rebuffer2354 (.A(net2758),
    .Y(net2759));
 BUFx3_ASAP7_75t_R split2355 (.A(_18532_),
    .Y(net2760));
 BUFx2_ASAP7_75t_R rebuffer2356 (.A(_05803_),
    .Y(net2761));
 BUFx2_ASAP7_75t_R rebuffer2357 (.A(_21919_),
    .Y(net2762));
 BUFx2_ASAP7_75t_R rebuffer2358 (.A(_21919_),
    .Y(net2763));
 BUFx4f_ASAP7_75t_R split2359 (.A(_06081_),
    .Y(net2764));
 BUFx2_ASAP7_75t_R rebuffer2360 (.A(_16304_),
    .Y(net2765));
 BUFx2_ASAP7_75t_R rebuffer2361 (.A(_16304_),
    .Y(net2766));
 BUFx2_ASAP7_75t_R rebuffer2362 (.A(net2766),
    .Y(net2767));
 BUFx2_ASAP7_75t_R rebuffer2363 (.A(net2766),
    .Y(net2768));
 BUFx2_ASAP7_75t_R rebuffer2364 (.A(net2766),
    .Y(net2769));
 BUFx4f_ASAP7_75t_R split2365 (.A(net1184),
    .Y(net2770));
 BUFx6f_ASAP7_75t_R rebuffer2366 (.A(_09636_),
    .Y(net2771));
 BUFx2_ASAP7_75t_R rebuffer2367 (.A(_10169_),
    .Y(net2772));
 BUFx2_ASAP7_75t_R rebuffer2368 (.A(_15504_),
    .Y(net2773));
 BUFx6f_ASAP7_75t_R rebuffer2369 (.A(_08338_),
    .Y(net2774));
 BUFx2_ASAP7_75t_R rebuffer2370 (.A(_09672_),
    .Y(net2775));
 BUFx2_ASAP7_75t_R rebuffer2371 (.A(_19108_),
    .Y(net2776));
 BUFx6f_ASAP7_75t_R rebuffer2372 (.A(_00633_),
    .Y(net2777));
 BUFx2_ASAP7_75t_R rebuffer2373 (.A(net2777),
    .Y(net2778));
 BUFx2_ASAP7_75t_R rebuffer2374 (.A(net2778),
    .Y(net2779));
 BUFx2_ASAP7_75t_R rebuffer2375 (.A(net2779),
    .Y(net2780));
 BUFx3_ASAP7_75t_R rebuffer2376 (.A(_10768_),
    .Y(net2781));
 BUFx2_ASAP7_75t_R rebuffer2377 (.A(_00622_),
    .Y(net2782));
 BUFx2_ASAP7_75t_R rebuffer2378 (.A(net2782),
    .Y(net2783));
 BUFx2_ASAP7_75t_R rebuffer2379 (.A(_05069_),
    .Y(net2784));
 BUFx2_ASAP7_75t_R rebuffer2380 (.A(_22015_),
    .Y(net2785));
 BUFx12f_ASAP7_75t_R rebuffer2381 (.A(_06044_),
    .Y(net2786));
 BUFx2_ASAP7_75t_R rebuffer2382 (.A(net2786),
    .Y(net2787));
 BUFx2_ASAP7_75t_R rebuffer2383 (.A(_18242_),
    .Y(net2788));
 BUFx3_ASAP7_75t_R rebuffer2384 (.A(_21914_),
    .Y(net2789));
 BUFx2_ASAP7_75t_R rebuffer2385 (.A(net2789),
    .Y(net2790));
 BUFx2_ASAP7_75t_R rebuffer2386 (.A(_21914_),
    .Y(net2791));
 BUFx3_ASAP7_75t_R rebuffer2387 (.A(_18131_),
    .Y(net2792));
 BUFx4f_ASAP7_75t_R split2388 (.A(_03090_),
    .Y(net2793));
 BUFx2_ASAP7_75t_R split2389 (.A(_01586_),
    .Y(net2794));
 BUFx4f_ASAP7_75t_R rebuffer2390 (.A(_01496_),
    .Y(net2795));
 BUFx2_ASAP7_75t_R rebuffer2391 (.A(net3186),
    .Y(net2796));
 BUFx6f_ASAP7_75t_R rebuffer2392 (.A(_00643_),
    .Y(net2797));
 BUFx4f_ASAP7_75t_R rebuffer2393 (.A(_09607_),
    .Y(net2798));
 BUFx2_ASAP7_75t_R rebuffer2394 (.A(net2798),
    .Y(net2799));
 BUFx6f_ASAP7_75t_R rebuffer2395 (.A(_20818_),
    .Y(net2800));
 BUFx2_ASAP7_75t_R rebuffer2396 (.A(_21927_),
    .Y(net2801));
 BUFx12f_ASAP7_75t_R split2397 (.A(net2038),
    .Y(net2802));
 BUFx2_ASAP7_75t_R rebuffer2398 (.A(_03617_),
    .Y(net2803));
 BUFx12f_ASAP7_75t_R rebuffer2399 (.A(_10144_),
    .Y(net2804));
 BUFx6f_ASAP7_75t_R rebuffer2400 (.A(net2804),
    .Y(net2805));
 BUFx6f_ASAP7_75t_R rebuffer2401 (.A(_10383_),
    .Y(net2806));
 BUFx2_ASAP7_75t_R rebuffer2402 (.A(_10383_),
    .Y(net2807));
 BUFx6f_ASAP7_75t_R rebuffer2403 (.A(_09906_),
    .Y(net2808));
 BUFx2_ASAP7_75t_R rebuffer2404 (.A(_05520_),
    .Y(net2809));
 BUFx2_ASAP7_75t_R rebuffer2405 (.A(_05520_),
    .Y(net2810));
 BUFx2_ASAP7_75t_R rebuffer2406 (.A(_18575_),
    .Y(net2811));
 BUFx6f_ASAP7_75t_R rebuffer2407 (.A(_20267_),
    .Y(net2812));
 BUFx4f_ASAP7_75t_R rebuffer2408 (.A(_06142_),
    .Y(net2813));
 BUFx10_ASAP7_75t_R split2409 (.A(net3121),
    .Y(net2814));
 BUFx6f_ASAP7_75t_R rebuffer2410 (.A(_05497_),
    .Y(net2815));
 BUFx6f_ASAP7_75t_R rebuffer2411 (.A(net2815),
    .Y(net2816));
 BUFx6f_ASAP7_75t_R rebuffer2412 (.A(_09662_),
    .Y(net2817));
 BUFx6f_ASAP7_75t_R rebuffer2413 (.A(_02361_),
    .Y(net2818));
 BUFx2_ASAP7_75t_R rebuffer2414 (.A(net2818),
    .Y(net2819));
 BUFx6f_ASAP7_75t_R rebuffer2415 (.A(_18971_),
    .Y(net2820));
 BUFx6f_ASAP7_75t_R rebuffer2416 (.A(net3186),
    .Y(net2821));
 BUFx6f_ASAP7_75t_R rebuffer2417 (.A(_21603_),
    .Y(net2822));
 BUFx2_ASAP7_75t_R rebuffer2418 (.A(_17957_),
    .Y(net2823));
 BUFx6f_ASAP7_75t_R rebuffer2419 (.A(_17963_),
    .Y(net2824));
 BUFx3_ASAP7_75t_R rebuffer2420 (.A(_18268_),
    .Y(net2825));
 BUFx2_ASAP7_75t_R rebuffer2421 (.A(_17561_),
    .Y(net2826));
 BUFx2_ASAP7_75t_R rebuffer2422 (.A(_03711_),
    .Y(net2827));
 BUFx4f_ASAP7_75t_R rebuffer2423 (.A(_09711_),
    .Y(net2828));
 BUFx3_ASAP7_75t_R rebuffer2424 (.A(_18532_),
    .Y(net2829));
 BUFx6f_ASAP7_75t_R rebuffer2425 (.A(_00650_),
    .Y(net2830));
 BUFx2_ASAP7_75t_R rebuffer2426 (.A(net2830),
    .Y(net2831));
 BUFx2_ASAP7_75t_R rebuffer2427 (.A(net2830),
    .Y(net2832));
 BUFx6f_ASAP7_75t_R split2428 (.A(_05579_),
    .Y(net2833));
 BUFx3_ASAP7_75t_R split2429 (.A(_05642_),
    .Y(net2834));
 BUFx3_ASAP7_75t_R rebuffer2430 (.A(_05502_),
    .Y(net2835));
 BUFx2_ASAP7_75t_R rebuffer2431 (.A(net2835),
    .Y(net2836));
 BUFx2_ASAP7_75t_R rebuffer2432 (.A(_00654_),
    .Y(net2837));
 BUFx2_ASAP7_75t_R rebuffer2433 (.A(_00654_),
    .Y(net2838));
 BUFx2_ASAP7_75t_R rebuffer2434 (.A(net3361),
    .Y(net2839));
 BUFx2_ASAP7_75t_R rebuffer2435 (.A(_16295_),
    .Y(net2840));
 BUFx3_ASAP7_75t_R split2436 (.A(_10329_),
    .Y(net2841));
 BUFx2_ASAP7_75t_R rebuffer2437 (.A(_18048_),
    .Y(net2842));
 BUFx6f_ASAP7_75t_R rebuffer2438 (.A(_18048_),
    .Y(net2843));
 BUFx3_ASAP7_75t_R rebuffer2439 (.A(net2843),
    .Y(net2844));
 BUFx2_ASAP7_75t_R rebuffer2440 (.A(_05860_),
    .Y(net2845));
 BUFx3_ASAP7_75t_R rebuffer2441 (.A(_05860_),
    .Y(net2846));
 BUFx4f_ASAP7_75t_R split2442 (.A(_17657_),
    .Y(net2847));
 BUFx2_ASAP7_75t_R rebuffer2443 (.A(_17954_),
    .Y(net2848));
 BUFx3_ASAP7_75t_R rebuffer2444 (.A(_18259_),
    .Y(net2849));
 BUFx4_ASAP7_75t_R rebuffer2445 (.A(_12290_),
    .Y(net2850));
 BUFx3_ASAP7_75t_R split2446 (.A(_10370_),
    .Y(net2851));
 BUFx2_ASAP7_75t_R rebuffer2447 (.A(net3009),
    .Y(net2852));
 BUFx2_ASAP7_75t_R rebuffer2448 (.A(_17942_),
    .Y(net2853));
 BUFx2_ASAP7_75t_R rebuffer2449 (.A(_10485_),
    .Y(net2854));
 BUFx2_ASAP7_75t_R rebuffer2450 (.A(_06188_),
    .Y(net2855));
 BUFx6f_ASAP7_75t_R rebuffer2451 (.A(_06188_),
    .Y(net2856));
 BUFx2_ASAP7_75t_R rebuffer2452 (.A(net2856),
    .Y(net2857));
 BUFx12f_ASAP7_75t_R rebuffer2453 (.A(_05859_),
    .Y(net2858));
 BUFx2_ASAP7_75t_R rebuffer2454 (.A(net2858),
    .Y(net2859));
 BUFx3_ASAP7_75t_R rebuffer2455 (.A(_09867_),
    .Y(net2860));
 BUFx2_ASAP7_75t_R rebuffer2456 (.A(_09710_),
    .Y(net2861));
 BUFx6f_ASAP7_75t_R split2457 (.A(net2907),
    .Y(net2862));
 BUFx6f_ASAP7_75t_R rebuffer2458 (.A(_05485_),
    .Y(net2863));
 BUFx2_ASAP7_75t_R rebuffer2459 (.A(net2863),
    .Y(net2864));
 BUFx2_ASAP7_75t_R rebuffer2460 (.A(_05485_),
    .Y(net2865));
 BUFx2_ASAP7_75t_R rebuffer2461 (.A(_09936_),
    .Y(net2866));
 BUFx2_ASAP7_75t_R rebuffer2462 (.A(_09936_),
    .Y(net2867));
 BUFx2_ASAP7_75t_R rebuffer2463 (.A(_10326_),
    .Y(net2868));
 BUFx2_ASAP7_75t_R rebuffer2464 (.A(_00562_),
    .Y(net2869));
 BUFx4f_ASAP7_75t_R split2465 (.A(_05508_),
    .Y(net2870));
 BUFx2_ASAP7_75t_R rebuffer2466 (.A(_17536_),
    .Y(net2871));
 BUFx6f_ASAP7_75t_R split2467 (.A(net3142),
    .Y(net2872));
 BUFx6f_ASAP7_75t_R rebuffer2468 (.A(_00630_),
    .Y(net2873));
 BUFx2_ASAP7_75t_R rebuffer2469 (.A(net2873),
    .Y(net2874));
 BUFx3_ASAP7_75t_R rebuffer2470 (.A(_05767_),
    .Y(net2875));
 BUFx6f_ASAP7_75t_R rebuffer2471 (.A(_05767_),
    .Y(net2876));
 BUFx3_ASAP7_75t_R rebuffer2472 (.A(_18901_),
    .Y(net2877));
 BUFx2_ASAP7_75t_R rebuffer2473 (.A(net2877),
    .Y(net2878));
 BUFx6f_ASAP7_75t_R split2474 (.A(_17533_),
    .Y(net2879));
 BUFx2_ASAP7_75t_R rebuffer2475 (.A(_17550_),
    .Y(net2880));
 BUFx6f_ASAP7_75t_R rebuffer2476 (.A(_17712_),
    .Y(net2881));
 BUFx2_ASAP7_75t_R rebuffer2477 (.A(_17712_),
    .Y(net2882));
 BUFx2_ASAP7_75t_R rebuffer2478 (.A(net2882),
    .Y(net2883));
 BUFx6f_ASAP7_75t_R rebuffer2479 (.A(_17712_),
    .Y(net2884));
 BUFx3_ASAP7_75t_R split2480 (.A(_19143_),
    .Y(net2885));
 BUFx2_ASAP7_75t_R rebuffer2481 (.A(_00563_),
    .Y(net2886));
 BUFx2_ASAP7_75t_R rebuffer2482 (.A(net2886),
    .Y(net2887));
 BUFx4f_ASAP7_75t_R rebuffer2483 (.A(_19145_),
    .Y(net2888));
 BUFx12f_ASAP7_75t_R rebuffer2484 (.A(_17670_),
    .Y(net2889));
 BUFx2_ASAP7_75t_R rebuffer2485 (.A(net2889),
    .Y(net2890));
 BUFx4f_ASAP7_75t_R split2486 (.A(_17533_),
    .Y(net2891));
 BUFx3_ASAP7_75t_R split2487 (.A(_17596_),
    .Y(net2892));
 BUFx4f_ASAP7_75t_R split2488 (.A(net1098),
    .Y(net2893));
 BUFx3_ASAP7_75t_R rebuffer2489 (.A(_17593_),
    .Y(net2894));
 BUFx6f_ASAP7_75t_R rebuffer2490 (.A(_17593_),
    .Y(net2895));
 BUFx3_ASAP7_75t_R rebuffer2491 (.A(_17656_),
    .Y(net2896));
 BUFx3_ASAP7_75t_R rebuffer2492 (.A(_17622_),
    .Y(net2897));
 BUFx2_ASAP7_75t_R rebuffer2493 (.A(_18229_),
    .Y(net2898));
 BUFx4f_ASAP7_75t_R split2494 (.A(_17624_),
    .Y(net2899));
 BUFx2_ASAP7_75t_R rebuffer2495 (.A(_17624_),
    .Y(net2900));
 BUFx4f_ASAP7_75t_R rebuffer2496 (.A(_17624_),
    .Y(net2901));
 BUFx12f_ASAP7_75t_R rebuffer2497 (.A(_17530_),
    .Y(net2902));
 BUFx2_ASAP7_75t_R rebuffer2498 (.A(net2902),
    .Y(net2903));
 BUFx2_ASAP7_75t_R rebuffer2499 (.A(net2902),
    .Y(net2904));
 BUFx2_ASAP7_75t_R rebuffer2500 (.A(net2902),
    .Y(net2905));
 BUFx6f_ASAP7_75t_R rebuffer2501 (.A(_17535_),
    .Y(net2906));
 BUFx4f_ASAP7_75t_R split2502 (.A(_17580_),
    .Y(net2907));
 BUFx6f_ASAP7_75t_R split2503 (.A(_17993_),
    .Y(net2908));
 BUFx3_ASAP7_75t_R split2504 (.A(_17770_),
    .Y(net2909));
 BUFx2_ASAP7_75t_R rebuffer2505 (.A(_00558_),
    .Y(net2910));
 BUFx6f_ASAP7_75t_R rebuffer2506 (.A(_09801_),
    .Y(net2911));
 BUFx2_ASAP7_75t_R rebuffer2507 (.A(_09730_),
    .Y(net2912));
 BUFx2_ASAP7_75t_R rebuffer2508 (.A(net2912),
    .Y(net2913));
 BUFx3_ASAP7_75t_R split2509 (.A(_09695_),
    .Y(net2914));
 BUFx2_ASAP7_75t_R rebuffer2510 (.A(_09629_),
    .Y(net2915));
 BUFx2_ASAP7_75t_R rebuffer2511 (.A(_09672_),
    .Y(net2916));
 BUFx3_ASAP7_75t_R split2512 (.A(_09594_),
    .Y(net2917));
 BUFx2_ASAP7_75t_R rebuffer2513 (.A(_09580_),
    .Y(net2918));
 BUFx6f_ASAP7_75t_R rebuffer2514 (.A(_09580_),
    .Y(net2919));
 BUFx2_ASAP7_75t_R rebuffer2515 (.A(net2919),
    .Y(net2920));
 BUFx3_ASAP7_75t_R rebuffer2516 (.A(_09642_),
    .Y(net2921));
 BUFx12f_ASAP7_75t_R rebuffer2517 (.A(_09755_),
    .Y(net2922));
 BUFx2_ASAP7_75t_R rebuffer2518 (.A(net2922),
    .Y(net2923));
 BUFx2_ASAP7_75t_R rebuffer2519 (.A(net2922),
    .Y(net2924));
 BUFx4f_ASAP7_75t_R split2520 (.A(_10106_),
    .Y(net2925));
 BUFx2_ASAP7_75t_R rebuffer2521 (.A(_11141_),
    .Y(net2926));
 BUFx12f_ASAP7_75t_R rebuffer2522 (.A(_09586_),
    .Y(net2927));
 BUFx2_ASAP7_75t_R rebuffer2523 (.A(net2927),
    .Y(net2928));
 BUFx2_ASAP7_75t_R rebuffer2524 (.A(_00611_),
    .Y(net2929));
 BUFx2_ASAP7_75t_R rebuffer2525 (.A(net2929),
    .Y(net2930));
 BUFx2_ASAP7_75t_R rebuffer2526 (.A(_09625_),
    .Y(net2931));
 BUFx3_ASAP7_75t_R rebuffer2527 (.A(_10884_),
    .Y(net2932));
 BUFx6f_ASAP7_75t_R rebuffer2528 (.A(_00533_),
    .Y(net2933));
 BUFx2_ASAP7_75t_R rebuffer2529 (.A(net2933),
    .Y(net2934));
 BUFx2_ASAP7_75t_R rebuffer2530 (.A(net2933),
    .Y(net2935));
 BUFx6f_ASAP7_75t_R rebuffer2531 (.A(_09919_),
    .Y(net2936));
 BUFx6f_ASAP7_75t_R rebuffer2532 (.A(_09854_),
    .Y(net2937));
 BUFx2_ASAP7_75t_R rebuffer2533 (.A(net2937),
    .Y(net2938));
 BUFx3_ASAP7_75t_R rebuffer2534 (.A(net2937),
    .Y(net2939));
 BUFx3_ASAP7_75t_R split2535 (.A(_09592_),
    .Y(net2940));
 BUFx4f_ASAP7_75t_R split2536 (.A(_09822_),
    .Y(net2941));
 BUFx2_ASAP7_75t_R rebuffer2537 (.A(_09649_),
    .Y(net2942));
 BUFx2_ASAP7_75t_R rebuffer2538 (.A(_09649_),
    .Y(net2943));
 BUFx6f_ASAP7_75t_R rebuffer2539 (.A(_17956_),
    .Y(net2944));
 BUFx2_ASAP7_75t_R split2540 (.A(_18316_),
    .Y(net2945));
 BUFx3_ASAP7_75t_R rebuffer2541 (.A(_18144_),
    .Y(net2946));
 BUFx3_ASAP7_75t_R split2546 (.A(_10419_),
    .Y(net2951));
 BUFx2_ASAP7_75t_R rebuffer2547 (.A(_11364_),
    .Y(net2952));
 BUFx2_ASAP7_75t_R rebuffer2548 (.A(net2952),
    .Y(net2953));
 BUFx3_ASAP7_75t_R rebuffer2549 (.A(_10408_),
    .Y(net2954));
 BUFx2_ASAP7_75t_R rebuffer2550 (.A(net2954),
    .Y(net2955));
 BUFx4f_ASAP7_75t_R split2551 (.A(_09809_),
    .Y(net2956));
 BUFx6f_ASAP7_75t_R split2552 (.A(_10485_),
    .Y(net2957));
 BUFx4f_ASAP7_75t_R rebuffer2553 (.A(_09998_),
    .Y(net2958));
 BUFx4f_ASAP7_75t_R rebuffer2554 (.A(_09718_),
    .Y(net2959));
 BUFx3_ASAP7_75t_R rebuffer2555 (.A(net2959),
    .Y(net2960));
 BUFx2_ASAP7_75t_R rebuffer2556 (.A(net2959),
    .Y(net2961));
 BUFx2_ASAP7_75t_R split2557 (.A(_10384_),
    .Y(net2962));
 BUFx6f_ASAP7_75t_R split2558 (.A(_18305_),
    .Y(net2963));
 BUFx6f_ASAP7_75t_R rebuffer2559 (.A(_18316_),
    .Y(net2964));
 BUFx6f_ASAP7_75t_R rebuffer2560 (.A(_18453_),
    .Y(net2965));
 BUFx2_ASAP7_75t_R rebuffer2561 (.A(net2965),
    .Y(net2966));
 BUFx2_ASAP7_75t_R rebuffer2562 (.A(net2965),
    .Y(net2967));
 BUFx2_ASAP7_75t_R rebuffer2563 (.A(_18238_),
    .Y(net2968));
 BUFx2_ASAP7_75t_R rebuffer2564 (.A(_18305_),
    .Y(net2969));
 BUFx4f_ASAP7_75t_R split2565 (.A(_18300_),
    .Y(net2970));
 BUFx2_ASAP7_75t_R rebuffer2566 (.A(_18256_),
    .Y(net2971));
 BUFx2_ASAP7_75t_R rebuffer2567 (.A(net2971),
    .Y(net2972));
 BUFx2_ASAP7_75t_R rebuffer2568 (.A(_18366_),
    .Y(net2973));
 BUFx2_ASAP7_75t_R rebuffer2569 (.A(net2973),
    .Y(net2974));
 BUFx2_ASAP7_75t_R rebuffer2570 (.A(_18366_),
    .Y(net2975));
 BUFx2_ASAP7_75t_R rebuffer2571 (.A(net2975),
    .Y(net2976));
 BUFx2_ASAP7_75t_R rebuffer2572 (.A(_18366_),
    .Y(net2977));
 BUFx2_ASAP7_75t_R rebuffer2573 (.A(net2977),
    .Y(net2978));
 BUFx3_ASAP7_75t_R split2574 (.A(_18650_),
    .Y(net2979));
 BUFx2_ASAP7_75t_R rebuffer2575 (.A(_18252_),
    .Y(net2980));
 BUFx4f_ASAP7_75t_R split2576 (.A(_18377_),
    .Y(net2981));
 BUFx6f_ASAP7_75t_R rebuffer2577 (.A(_18287_),
    .Y(net2982));
 BUFx2_ASAP7_75t_R rebuffer2578 (.A(net2982),
    .Y(net2983));
 BUFx3_ASAP7_75t_R rebuffer2579 (.A(_00568_),
    .Y(net2984));
 BUFx2_ASAP7_75t_R split2580 (.A(_18287_),
    .Y(net2985));
 BUFx6f_ASAP7_75t_R rebuffer2581 (.A(_20049_),
    .Y(net2986));
 BUFx2_ASAP7_75t_R rebuffer2582 (.A(net2986),
    .Y(net2987));
 BUFx6f_ASAP7_75t_R rebuffer2583 (.A(_00566_),
    .Y(net2988));
 BUFx4f_ASAP7_75t_R split2584 (.A(_18439_),
    .Y(net2989));
 BUFx2_ASAP7_75t_R split2585 (.A(net1393),
    .Y(net2990));
 BUFx2_ASAP7_75t_R rebuffer2586 (.A(_18690_),
    .Y(net2991));
 BUFx2_ASAP7_75t_R rebuffer2587 (.A(_18690_),
    .Y(net2992));
 BUFx2_ASAP7_75t_R rebuffer2588 (.A(_18523_),
    .Y(net2993));
 BUFx3_ASAP7_75t_R split2589 (.A(_18490_),
    .Y(net2994));
 BUFx2_ASAP7_75t_R rebuffer2590 (.A(_18235_),
    .Y(net2995));
 BUFx6f_ASAP7_75t_R rebuffer2591 (.A(_00601_),
    .Y(net2996));
 BUFx2_ASAP7_75t_R rebuffer2592 (.A(net2996),
    .Y(net2997));
 BUFx2_ASAP7_75t_R rebuffer2593 (.A(net2996),
    .Y(net2998));
 BUFx6f_ASAP7_75t_R split2594 (.A(_18240_),
    .Y(net2999));
 BUFx3_ASAP7_75t_R rebuffer2595 (.A(_00607_),
    .Y(net3000));
 BUFx2_ASAP7_75t_R rebuffer2596 (.A(_18272_),
    .Y(net3001));
 BUFx3_ASAP7_75t_R rebuffer2597 (.A(_18281_),
    .Y(net3002));
 BUFx3_ASAP7_75t_R split2598 (.A(_18442_),
    .Y(net3003));
 BUFx6f_ASAP7_75t_R rebuffer2599 (.A(_18517_),
    .Y(net3004));
 BUFx3_ASAP7_75t_R split2600 (.A(_18240_),
    .Y(net3005));
 BUFx2_ASAP7_75t_R rebuffer2601 (.A(_18655_),
    .Y(net3006));
 BUFx2_ASAP7_75t_R rebuffer2602 (.A(_00565_),
    .Y(net3007));
 BUFx3_ASAP7_75t_R rebuffer2603 (.A(_00565_),
    .Y(net3008));
 BUFx3_ASAP7_75t_R rebuffer2604 (.A(_00565_),
    .Y(net3009));
 BUFx3_ASAP7_75t_R rebuffer2605 (.A(_10389_),
    .Y(net3010));
 BUFx2_ASAP7_75t_R rebuffer2606 (.A(_10389_),
    .Y(net3011));
 BUFx2_ASAP7_75t_R rebuffer2607 (.A(net3011),
    .Y(net3012));
 BUFx2_ASAP7_75t_R rebuffer2608 (.A(net3011),
    .Y(net3013));
 BUFx2_ASAP7_75t_R rebuffer2609 (.A(_11954_),
    .Y(net3014));
 BUFx6f_ASAP7_75t_R split2610 (.A(_09888_),
    .Y(net3015));
 BUFx3_ASAP7_75t_R split2611 (.A(_09620_),
    .Y(net3016));
 BUFx6f_ASAP7_75t_R rebuffer2612 (.A(_09888_),
    .Y(net3017));
 BUFx6f_ASAP7_75t_R rebuffer2613 (.A(_10318_),
    .Y(net3018));
 BUFx2_ASAP7_75t_R rebuffer2614 (.A(_10318_),
    .Y(net3019));
 BUFx6f_ASAP7_75t_R split2615 (.A(_10624_),
    .Y(net3020));
 BUFx4f_ASAP7_75t_R split2616 (.A(_10664_),
    .Y(net3021));
 BUFx4f_ASAP7_75t_R rebuffer2617 (.A(_10744_),
    .Y(net3022));
 BUFx2_ASAP7_75t_R rebuffer2618 (.A(net3022),
    .Y(net3023));
 BUFx2_ASAP7_75t_R rebuffer2619 (.A(_00534_),
    .Y(net3024));
 BUFx3_ASAP7_75t_R rebuffer2620 (.A(_00534_),
    .Y(net3025));
 BUFx2_ASAP7_75t_R rebuffer2621 (.A(net3025),
    .Y(net3026));
 BUFx2_ASAP7_75t_R rebuffer2622 (.A(net3026),
    .Y(net3027));
 BUFx3_ASAP7_75t_R rebuffer2623 (.A(_00534_),
    .Y(net3028));
 BUFx2_ASAP7_75t_R rebuffer2624 (.A(_10826_),
    .Y(net3029));
 BUFx6f_ASAP7_75t_R rebuffer2625 (.A(_10826_),
    .Y(net3030));
 BUFx3_ASAP7_75t_R rebuffer2626 (.A(_10826_),
    .Y(net3031));
 BUFx6f_ASAP7_75t_R rebuffer2627 (.A(_10339_),
    .Y(net3032));
 BUFx4f_ASAP7_75t_R split2628 (.A(_10851_),
    .Y(net3033));
 BUFx3_ASAP7_75t_R split2629 (.A(_10551_),
    .Y(net3034));
 BUFx6f_ASAP7_75t_R rebuffer2630 (.A(_10328_),
    .Y(net3035));
 BUFx2_ASAP7_75t_R rebuffer2631 (.A(_10380_),
    .Y(net3036));
 BUFx3_ASAP7_75t_R rebuffer2632 (.A(_10394_),
    .Y(net3037));
 BUFx6f_ASAP7_75t_R rebuffer2633 (.A(_10369_),
    .Y(net3038));
 BUFx2_ASAP7_75t_R rebuffer2634 (.A(net3038),
    .Y(net3039));
 BUFx12f_ASAP7_75t_R rebuffer2635 (.A(_10769_),
    .Y(net3040));
 BUFx2_ASAP7_75t_R rebuffer2636 (.A(net3040),
    .Y(net3041));
 BUFx2_ASAP7_75t_R rebuffer2637 (.A(net3040),
    .Y(net3042));
 BUFx12f_ASAP7_75t_R rebuffer2638 (.A(_10546_),
    .Y(net3043));
 BUFx2_ASAP7_75t_R rebuffer2639 (.A(_10637_),
    .Y(net3044));
 BUFx2_ASAP7_75t_R rebuffer2640 (.A(_10637_),
    .Y(net3045));
 BUFx2_ASAP7_75t_R rebuffer2641 (.A(_10628_),
    .Y(net3046));
 BUFx2_ASAP7_75t_R rebuffer2642 (.A(_10628_),
    .Y(net3047));
 BUFx3_ASAP7_75t_R split2643 (.A(_10628_),
    .Y(net3048));
 BUFx4f_ASAP7_75t_R split2644 (.A(_10660_),
    .Y(net3049));
 BUFx2_ASAP7_75t_R rebuffer2645 (.A(_13869_),
    .Y(net3050));
 BUFx4f_ASAP7_75t_R split2646 (.A(_10375_),
    .Y(net3051));
 BUFx6f_ASAP7_75t_R split2647 (.A(_10449_),
    .Y(net3052));
 BUFx6f_ASAP7_75t_R split2648 (.A(_10751_),
    .Y(net3053));
 BUFx4f_ASAP7_75t_R split2649 (.A(_10864_),
    .Y(net3054));
 BUFx2_ASAP7_75t_R rebuffer2650 (.A(_10585_),
    .Y(net3055));
 BUFx4f_ASAP7_75t_R split2651 (.A(_10816_),
    .Y(net3056));
 BUFx4f_ASAP7_75t_R split2652 (.A(_10744_),
    .Y(net3057));
 BUFx6f_ASAP7_75t_R split2653 (.A(_10645_),
    .Y(net3058));
 BUFx6f_ASAP7_75t_R rebuffer2654 (.A(_09925_),
    .Y(net3059));
 BUFx3_ASAP7_75t_R rebuffer2655 (.A(_00610_),
    .Y(net3060));
 BUFx2_ASAP7_75t_R split2656 (.A(_10711_),
    .Y(net3061));
 BUFx3_ASAP7_75t_R rebuffer2657 (.A(_10106_),
    .Y(net3062));
 BUFx3_ASAP7_75t_R rebuffer2658 (.A(net3062),
    .Y(net3063));
 BUFx2_ASAP7_75t_R rebuffer2659 (.A(_10106_),
    .Y(net3064));
 BUFx3_ASAP7_75t_R split2660 (.A(_10751_),
    .Y(net3065));
 BUFx3_ASAP7_75t_R split2661 (.A(net1476),
    .Y(net3066));
 BUFx4f_ASAP7_75t_R split2662 (.A(_09689_),
    .Y(net3067));
 BUFx2_ASAP7_75t_R rebuffer2663 (.A(_10782_),
    .Y(net3068));
 BUFx4f_ASAP7_75t_R split2664 (.A(_09642_),
    .Y(net3069));
 BUFx4f_ASAP7_75t_R rebuffer2669 (.A(_00653_),
    .Y(net3074));
 BUFx3_ASAP7_75t_R split2670 (.A(_22015_),
    .Y(net3075));
 BUFx3_ASAP7_75t_R rebuffer2671 (.A(_21927_),
    .Y(net3076));
 BUFx2_ASAP7_75t_R rebuffer2672 (.A(net3076),
    .Y(net3077));
 BUFx6f_ASAP7_75t_R rebuffer2673 (.A(_21975_),
    .Y(net3078));
 BUFx2_ASAP7_75t_R rebuffer2674 (.A(_21975_),
    .Y(net3079));
 BUFx2_ASAP7_75t_R rebuffer2675 (.A(_22100_),
    .Y(net3080));
 BUFx6f_ASAP7_75t_R rebuffer2676 (.A(_22100_),
    .Y(net3081));
 BUFx3_ASAP7_75t_R rebuffer2677 (.A(net3081),
    .Y(net3082));
 BUFx6f_ASAP7_75t_R rebuffer2678 (.A(_22075_),
    .Y(net3083));
 BUFx3_ASAP7_75t_R split2679 (.A(net1374),
    .Y(net3084));
 BUFx2_ASAP7_75t_R rebuffer2680 (.A(_17700_),
    .Y(net3085));
 BUFx3_ASAP7_75t_R split2681 (.A(_17700_),
    .Y(net3086));
 BUFx2_ASAP7_75t_R rebuffer2682 (.A(_18295_),
    .Y(net3087));
 BUFx2_ASAP7_75t_R rebuffer2683 (.A(_17691_),
    .Y(net3088));
 BUFx2_ASAP7_75t_R rebuffer2684 (.A(_17691_),
    .Y(net3089));
 BUFx4f_ASAP7_75t_R split2685 (.A(_18530_),
    .Y(net3090));
 BUFx4f_ASAP7_75t_R split2686 (.A(_18900_),
    .Y(net3091));
 BUFx4f_ASAP7_75t_R split2687 (.A(_18020_),
    .Y(net3092));
 BUFx3_ASAP7_75t_R split2688 (.A(_10098_),
    .Y(net3093));
 BUFx2_ASAP7_75t_R rebuffer2689 (.A(_00621_),
    .Y(net3094));
 BUFx4f_ASAP7_75t_R split2690 (.A(_05240_),
    .Y(net3095));
 BUFx6f_ASAP7_75t_R rebuffer2691 (.A(_05337_),
    .Y(net3096));
 BUFx2_ASAP7_75t_R rebuffer2692 (.A(_05072_),
    .Y(net3097));
 BUFx6f_ASAP7_75t_R split2693 (.A(_05500_),
    .Y(net3098));
 BUFx6f_ASAP7_75t_R rebuffer2694 (.A(_00622_),
    .Y(net3099));
 BUFx2_ASAP7_75t_R rebuffer2695 (.A(_05069_),
    .Y(net3100));
 BUFx3_ASAP7_75t_R rebuffer2696 (.A(_05225_),
    .Y(net3101));
 BUFx3_ASAP7_75t_R rebuffer2697 (.A(_05225_),
    .Y(net3102));
 BUFx6f_ASAP7_75t_R rebuffer2698 (.A(_05086_),
    .Y(net3103));
 BUFx6f_ASAP7_75t_R rebuffer2699 (.A(net3103),
    .Y(net3104));
 BUFx2_ASAP7_75t_R rebuffer2700 (.A(_05165_),
    .Y(net3105));
 BUFx6f_ASAP7_75t_R split2701 (.A(_05664_),
    .Y(net3106));
 BUFx3_ASAP7_75t_R rebuffer2702 (.A(_05079_),
    .Y(net3107));
 BUFx3_ASAP7_75t_R rebuffer2703 (.A(_05079_),
    .Y(net3108));
 BUFx2_ASAP7_75t_R rebuffer2704 (.A(_05513_),
    .Y(net3109));
 BUFx4f_ASAP7_75t_R split2705 (.A(_05443_),
    .Y(net3110));
 BUFx3_ASAP7_75t_R split2706 (.A(_05500_),
    .Y(net3111));
 BUFx6f_ASAP7_75t_R rebuffer2707 (.A(_00580_),
    .Y(net3112));
 BUFx6f_ASAP7_75t_R rebuffer2708 (.A(_05451_),
    .Y(net3113));
 BUFx6f_ASAP7_75t_R rebuffer2709 (.A(_05427_),
    .Y(net3114));
 BUFx3_ASAP7_75t_R split2710 (.A(_05580_),
    .Y(net3115));
 BUFx2_ASAP7_75t_R rebuffer2711 (.A(_05434_),
    .Y(net3116));
 BUFx2_ASAP7_75t_R rebuffer2712 (.A(_05434_),
    .Y(net3117));
 BUFx6f_ASAP7_75t_R rebuffer2713 (.A(_05528_),
    .Y(net3118));
 BUFx6f_ASAP7_75t_R rebuffer2714 (.A(_09109_),
    .Y(net3119));
 BUFx2_ASAP7_75t_R rebuffer2715 (.A(net3447),
    .Y(net3120));
 BUFx4f_ASAP7_75t_R split2716 (.A(_05443_),
    .Y(net3121));
 BUFx2_ASAP7_75t_R rebuffer2717 (.A(_00579_),
    .Y(net3122));
 BUFx2_ASAP7_75t_R rebuffer2718 (.A(_18012_),
    .Y(net3123));
 BUFx4f_ASAP7_75t_R split2719 (.A(_17953_),
    .Y(net3124));
 BUFx3_ASAP7_75t_R split2720 (.A(_01949_),
    .Y(net3125));
 BUFx2_ASAP7_75t_R rebuffer2721 (.A(_01539_),
    .Y(net3126));
 BUFx2_ASAP7_75t_R rebuffer2722 (.A(_01539_),
    .Y(net3127));
 BUFx2_ASAP7_75t_R split2723 (.A(_01894_),
    .Y(net3128));
 BUFx6f_ASAP7_75t_R rebuffer2724 (.A(_00638_),
    .Y(net3129));
 BUFx2_ASAP7_75t_R rebuffer2725 (.A(net3129),
    .Y(net3130));
 BUFx2_ASAP7_75t_R rebuffer2726 (.A(_01815_),
    .Y(net3131));
 BUFx3_ASAP7_75t_R rebuffer2727 (.A(_01815_),
    .Y(net3132));
 BUFx6f_ASAP7_75t_R rebuffer2728 (.A(_00598_),
    .Y(net3133));
 BUFx2_ASAP7_75t_R rebuffer2729 (.A(net3133),
    .Y(net3134));
 BUFx6f_ASAP7_75t_R rebuffer2730 (.A(_01670_),
    .Y(net3135));
 BUFx2_ASAP7_75t_R rebuffer2731 (.A(net3135),
    .Y(net3136));
 BUFx2_ASAP7_75t_R rebuffer2732 (.A(net3135),
    .Y(net3137));
 BUFx4f_ASAP7_75t_R split2733 (.A(_01125_),
    .Y(net3138));
 BUFx6f_ASAP7_75t_R rebuffer2734 (.A(_04358_),
    .Y(net3139));
 BUFx3_ASAP7_75t_R rebuffer2735 (.A(net3139),
    .Y(net3140));
 BUFx2_ASAP7_75t_R rebuffer2736 (.A(net3140),
    .Y(net3141));
 BUFx4f_ASAP7_75t_R split2737 (.A(_01136_),
    .Y(net3142));
 BUFx2_ASAP7_75t_R rebuffer2738 (.A(_01078_),
    .Y(net3143));
 BUFx6f_ASAP7_75t_R split2739 (.A(_01191_),
    .Y(net3144));
 BUFx6f_ASAP7_75t_R split2740 (.A(_01287_),
    .Y(net3145));
 BUFx2_ASAP7_75t_R rebuffer2741 (.A(_01552_),
    .Y(net3146));
 BUFx2_ASAP7_75t_R rebuffer2742 (.A(net3146),
    .Y(net3147));
 BUFx2_ASAP7_75t_R rebuffer2743 (.A(_22004_),
    .Y(net3148));
 BUFx3_ASAP7_75t_R split2744 (.A(_01612_),
    .Y(net3149));
 BUFx2_ASAP7_75t_R rebuffer2745 (.A(_03466_),
    .Y(net3150));
 BUFx3_ASAP7_75t_R split2746 (.A(_21992_),
    .Y(net3151));
 BUFx3_ASAP7_75t_R split2747 (.A(_01078_),
    .Y(net3152));
 BUFx2_ASAP7_75t_R rebuffer2748 (.A(net3416),
    .Y(net3153));
 BUFx6f_ASAP7_75t_R split2749 (.A(_01202_),
    .Y(net3154));
 BUFx6f_ASAP7_75t_R split2750 (.A(_21934_),
    .Y(net3155));
 BUFx6f_ASAP7_75t_R rebuffer2751 (.A(_22028_),
    .Y(net3156));
 BUFx3_ASAP7_75t_R rebuffer2752 (.A(_10421_),
    .Y(net3157));
 BUFx2_ASAP7_75t_R rebuffer2753 (.A(net3157),
    .Y(net3158));
 BUFx2_ASAP7_75t_R rebuffer2754 (.A(_00651_),
    .Y(net3159));
 BUFx2_ASAP7_75t_R rebuffer2755 (.A(net3159),
    .Y(net3160));
 BUFx4f_ASAP7_75t_R split2756 (.A(net1114),
    .Y(net3161));
 BUFx2_ASAP7_75t_R rebuffer2759 (.A(net3373),
    .Y(net3164));
 BUFx6f_ASAP7_75t_R rebuffer2760 (.A(_07049_),
    .Y(net3165));
 BUFx6f_ASAP7_75t_R rebuffer2762 (.A(_22083_),
    .Y(net3167));
 BUFx3_ASAP7_75t_R rebuffer2763 (.A(_01892_),
    .Y(net3168));
 BUFx2_ASAP7_75t_R rebuffer2764 (.A(_01892_),
    .Y(net3169));
 BUFx6f_ASAP7_75t_R rebuffer2765 (.A(_01926_),
    .Y(net3170));
 BUFx2_ASAP7_75t_R rebuffer2766 (.A(net3170),
    .Y(net3171));
 BUFx12f_ASAP7_75t_R rebuffer2767 (.A(_21920_),
    .Y(net3172));
 BUFx2_ASAP7_75t_R rebuffer2768 (.A(_21920_),
    .Y(net3173));
 BUFx6f_ASAP7_75t_R rebuffer2769 (.A(_00567_),
    .Y(net3174));
 BUFx4f_ASAP7_75t_R split2770 (.A(_01728_),
    .Y(net3175));
 BUFx3_ASAP7_75t_R split2771 (.A(_03291_),
    .Y(net3176));
 BUFx4f_ASAP7_75t_R rebuffer2772 (.A(_09822_),
    .Y(net3177));
 BUFx4f_ASAP7_75t_R split2773 (.A(_18354_),
    .Y(net3178));
 BUFx6f_ASAP7_75t_R rebuffer2774 (.A(_00644_),
    .Y(net3179));
 BUFx2_ASAP7_75t_R rebuffer2775 (.A(_19846_),
    .Y(net3180));
 BUFx2_ASAP7_75t_R rebuffer2776 (.A(_18333_),
    .Y(net3181));
 BUFx4f_ASAP7_75t_R rebuffer2777 (.A(_18383_),
    .Y(net3182));
 BUFx2_ASAP7_75t_R rebuffer2778 (.A(_18383_),
    .Y(net3183));
 BUFx2_ASAP7_75t_R rebuffer2779 (.A(net3199),
    .Y(net3184));
 BUFx2_ASAP7_75t_R rebuffer2780 (.A(net3188),
    .Y(net3185));
 BUFx12f_ASAP7_75t_R rebuffer2781 (.A(_17993_),
    .Y(net3186));
 BUFx2_ASAP7_75t_R rebuffer2782 (.A(net3186),
    .Y(net3187));
 BUFx2_ASAP7_75t_R split2783 (.A(_18052_),
    .Y(net3188));
 BUFx2_ASAP7_75t_R rebuffer2784 (.A(_18014_),
    .Y(net3189));
 BUFx2_ASAP7_75t_R rebuffer2785 (.A(net3189),
    .Y(net3190));
 BUFx2_ASAP7_75t_R split2786 (.A(_18014_),
    .Y(net3191));
 BUFx3_ASAP7_75t_R split2787 (.A(_18155_),
    .Y(net3192));
 BUFx12f_ASAP7_75t_R split2788 (.A(net1030),
    .Y(net3193));
 BUFx6f_ASAP7_75t_R rebuffer2789 (.A(_17551_),
    .Y(net3194));
 BUFx6f_ASAP7_75t_R rebuffer2790 (.A(_17551_),
    .Y(net3195));
 BUFx6f_ASAP7_75t_R rebuffer2791 (.A(_18020_),
    .Y(net3196));
 BUFx3_ASAP7_75t_R rebuffer2792 (.A(_17955_),
    .Y(net3197));
 BUFx2_ASAP7_75t_R rebuffer2793 (.A(_17955_),
    .Y(net3198));
 BUFx3_ASAP7_75t_R rebuffer2794 (.A(_18052_),
    .Y(net3199));
 BUFx3_ASAP7_75t_R rebuffer2795 (.A(_18074_),
    .Y(net3200));
 BUFx6f_ASAP7_75t_R split2796 (.A(net3366),
    .Y(net3201));
 BUFx2_ASAP7_75t_R rebuffer2797 (.A(_18131_),
    .Y(net3202));
 BUFx3_ASAP7_75t_R rebuffer2798 (.A(_18014_),
    .Y(net3203));
 BUFx3_ASAP7_75t_R split2799 (.A(net1058),
    .Y(net3204));
 BUFx3_ASAP7_75t_R split2800 (.A(_17977_),
    .Y(net3205));
 BUFx3_ASAP7_75t_R rebuffer2801 (.A(_17957_),
    .Y(net3206));
 BUFx6f_ASAP7_75t_R split2802 (.A(_18131_),
    .Y(net3207));
 BUFx6f_ASAP7_75t_R rebuffer2803 (.A(_18535_),
    .Y(net3208));
 BUFx3_ASAP7_75t_R rebuffer2804 (.A(_18535_),
    .Y(net3209));
 BUFx3_ASAP7_75t_R rebuffer2805 (.A(_18535_),
    .Y(net3210));
 BUFx6f_ASAP7_75t_R rebuffer2806 (.A(_00564_),
    .Y(net3211));
 BUFx2_ASAP7_75t_R rebuffer2807 (.A(_18881_),
    .Y(net3212));
 BUFx2_ASAP7_75t_R rebuffer2808 (.A(_18881_),
    .Y(net3213));
 BUFx2_ASAP7_75t_R rebuffer2809 (.A(net3213),
    .Y(net3214));
 BUFx3_ASAP7_75t_R split2810 (.A(_18685_),
    .Y(net3215));
 BUFx4f_ASAP7_75t_R split2811 (.A(_18012_),
    .Y(net3216));
 BUFx2_ASAP7_75t_R rebuffer2812 (.A(_18081_),
    .Y(net3217));
 BUFx6f_ASAP7_75t_R rebuffer2813 (.A(_18047_),
    .Y(net3218));
 BUFx2_ASAP7_75t_R rebuffer2814 (.A(net3218),
    .Y(net3219));
 BUFx2_ASAP7_75t_R rebuffer2815 (.A(net3218),
    .Y(net3220));
 BUFx2_ASAP7_75t_R rebuffer2816 (.A(_18108_),
    .Y(net3221));
 BUFx2_ASAP7_75t_R rebuffer2817 (.A(_18108_),
    .Y(net3222));
 BUFx4f_ASAP7_75t_R rebuffer2818 (.A(_18116_),
    .Y(net3223));
 BUFx2_ASAP7_75t_R rebuffer2819 (.A(_17980_),
    .Y(net3224));
 BUFx3_ASAP7_75t_R rebuffer2820 (.A(_21983_),
    .Y(net3225));
 BUFx3_ASAP7_75t_R rebuffer2825 (.A(_06039_),
    .Y(net3230));
 BUFx4f_ASAP7_75t_R split2826 (.A(_06084_),
    .Y(net3231));
 BUFx6f_ASAP7_75t_R rebuffer2827 (.A(_00625_),
    .Y(net3232));
 BUFx2_ASAP7_75t_R rebuffer2828 (.A(net3232),
    .Y(net3233));
 BUFx3_ASAP7_75t_R rebuffer2829 (.A(net3232),
    .Y(net3234));
 BUFx6f_ASAP7_75t_R split2830 (.A(_06210_),
    .Y(net3235));
 BUFx6f_ASAP7_75t_R rebuffer2831 (.A(_21934_),
    .Y(net3236));
 BUFx6f_ASAP7_75t_R rebuffer2832 (.A(_04201_),
    .Y(net3237));
 BUFx2_ASAP7_75t_R rebuffer2833 (.A(_20436_),
    .Y(net3238));
 BUFx6f_ASAP7_75t_R rebuffer2834 (.A(_18969_),
    .Y(net3239));
 BUFx6f_ASAP7_75t_R split2835 (.A(_01345_),
    .Y(net3240));
 BUFx3_ASAP7_75t_R split2836 (.A(_09655_),
    .Y(net3241));
 BUFx6f_ASAP7_75t_R rebuffer2837 (.A(_11730_),
    .Y(net3242));
 BUFx2_ASAP7_75t_R rebuffer2838 (.A(_09798_),
    .Y(net3243));
 BUFx3_ASAP7_75t_R split2839 (.A(_10086_),
    .Y(net3244));
 BUFx2_ASAP7_75t_R rebuffer2840 (.A(_09882_),
    .Y(net3245));
 BUFx3_ASAP7_75t_R split2841 (.A(_18253_),
    .Y(net3246));
 BUFx3_ASAP7_75t_R rebuffer2842 (.A(_18297_),
    .Y(net3247));
 BUFx2_ASAP7_75t_R rebuffer2843 (.A(_18297_),
    .Y(net3248));
 BUFx3_ASAP7_75t_R rebuffer2844 (.A(_05508_),
    .Y(net3249));
 BUFx2_ASAP7_75t_R rebuffer2845 (.A(_05508_),
    .Y(net3250));
 BUFx3_ASAP7_75t_R rebuffer2848 (.A(_01965_),
    .Y(net3253));
 BUFx2_ASAP7_75t_R rebuffer2849 (.A(_01965_),
    .Y(net3254));
 BUFx2_ASAP7_75t_R rebuffer2850 (.A(_01592_),
    .Y(net3255));
 BUFx3_ASAP7_75t_R split2851 (.A(_01707_),
    .Y(net3256));
 BUFx3_ASAP7_75t_R split2852 (.A(_01635_),
    .Y(net3257));
 BUFx3_ASAP7_75t_R rebuffer2853 (.A(_01786_),
    .Y(net3258));
 BUFx2_ASAP7_75t_R rebuffer2854 (.A(net3258),
    .Y(net3259));
 BUFx4f_ASAP7_75t_R split2855 (.A(_04606_),
    .Y(net3260));
 BUFx4f_ASAP7_75t_R split2856 (.A(_01641_),
    .Y(net3261));
 BUFx6f_ASAP7_75t_R rebuffer2857 (.A(_00593_),
    .Y(net3262));
 BUFx2_ASAP7_75t_R rebuffer2858 (.A(net3262),
    .Y(net3263));
 BUFx2_ASAP7_75t_R rebuffer2859 (.A(_01543_),
    .Y(net3264));
 BUFx2_ASAP7_75t_R rebuffer2860 (.A(_02361_),
    .Y(net3265));
 BUFx2_ASAP7_75t_R rebuffer2861 (.A(_02361_),
    .Y(net3266));
 BUFx2_ASAP7_75t_R rebuffer2862 (.A(_01607_),
    .Y(net3267));
 BUFx3_ASAP7_75t_R rebuffer2863 (.A(_02888_),
    .Y(net3268));
 BUFx12f_ASAP7_75t_R split2864 (.A(_04747_),
    .Y(net3269));
 BUFx6f_ASAP7_75t_R rebuffer2865 (.A(_04683_),
    .Y(net3270));
 BUFx3_ASAP7_75t_R rebuffer2866 (.A(_01769_),
    .Y(net3271));
 BUFx2_ASAP7_75t_R rebuffer2867 (.A(net3271),
    .Y(net3272));
 BUFx6f_ASAP7_75t_R rebuffer2868 (.A(_00595_),
    .Y(net3273));
 BUFx3_ASAP7_75t_R split2869 (.A(_02117_),
    .Y(net3274));
 BUFx12f_ASAP7_75t_R rebuffer2870 (.A(_01778_),
    .Y(net3275));
 BUFx4f_ASAP7_75t_R split2871 (.A(_01831_),
    .Y(net3276));
 BUFx2_ASAP7_75t_R rebuffer2872 (.A(_01824_),
    .Y(net3277));
 BUFx6f_ASAP7_75t_R rebuffer2873 (.A(_00545_),
    .Y(net3278));
 BUFx2_ASAP7_75t_R rebuffer2874 (.A(net3278),
    .Y(net3279));
 BUFx4f_ASAP7_75t_R split2875 (.A(_21927_),
    .Y(net3280));
 BUFx2_ASAP7_75t_R rebuffer2876 (.A(_18269_),
    .Y(net3281));
 BUFx3_ASAP7_75t_R split2877 (.A(_18479_),
    .Y(net3282));
 BUFx6f_ASAP7_75t_R rebuffer2878 (.A(_18445_),
    .Y(net3283));
 BUFx6f_ASAP7_75t_R split2879 (.A(net3285),
    .Y(net3284));
 BUFx4f_ASAP7_75t_R split2880 (.A(_17947_),
    .Y(net3285));
 BUFx2_ASAP7_75t_R rebuffer2881 (.A(_20112_),
    .Y(net3286));
 BUFx6f_ASAP7_75t_R split2882 (.A(_03809_),
    .Y(net3287));
 BUFx2_ASAP7_75t_R rebuffer2883 (.A(_03013_),
    .Y(net3288));
 BUFx6f_ASAP7_75t_R split2884 (.A(_01096_),
    .Y(net3289));
 BUFx6f_ASAP7_75t_R rebuffer2885 (.A(_10349_),
    .Y(net3290));
 BUFx2_ASAP7_75t_R rebuffer2886 (.A(net3290),
    .Y(net3291));
 BUFx4f_ASAP7_75t_R split2887 (.A(_10471_),
    .Y(net3292));
 BUFx3_ASAP7_75t_R rebuffer2888 (.A(_10343_),
    .Y(net3293));
 BUFx2_ASAP7_75t_R rebuffer2889 (.A(_13021_),
    .Y(net3294));
 BUFx3_ASAP7_75t_R rebuffer2890 (.A(_14154_),
    .Y(net3295));
 BUFx2_ASAP7_75t_R rebuffer2891 (.A(_10317_),
    .Y(net3296));
 BUFx3_ASAP7_75t_R rebuffer2892 (.A(_10505_),
    .Y(net3297));
 BUFx2_ASAP7_75t_R rebuffer2893 (.A(net3297),
    .Y(net3298));
 BUFx3_ASAP7_75t_R rebuffer2894 (.A(_18165_),
    .Y(net3299));
 BUFx3_ASAP7_75t_R rebuffer2895 (.A(_18028_),
    .Y(net3300));
 BUFx2_ASAP7_75t_R rebuffer2896 (.A(net3300),
    .Y(net3301));
 BUFx2_ASAP7_75t_R rebuffer2897 (.A(_18028_),
    .Y(net3302));
 BUFx2_ASAP7_75t_R rebuffer2898 (.A(_18039_),
    .Y(net3303));
 BUFx6f_ASAP7_75t_R rebuffer2899 (.A(_18039_),
    .Y(net3304));
 BUFx2_ASAP7_75t_R rebuffer2900 (.A(net3304),
    .Y(net3305));
 BUFx4f_ASAP7_75t_R split2901 (.A(_17980_),
    .Y(net3306));
 BUFx3_ASAP7_75t_R rebuffer2902 (.A(_17943_),
    .Y(net3307));
 BUFx3_ASAP7_75t_R split2903 (.A(_17953_),
    .Y(net3308));
 BUFx6f_ASAP7_75t_R split2904 (.A(_09892_),
    .Y(net3309));
 BUFx2_ASAP7_75t_R rebuffer2905 (.A(_18464_),
    .Y(net3310));
 BUFx2_ASAP7_75t_R rebuffer2906 (.A(_17529_),
    .Y(net3311));
 BUFx3_ASAP7_75t_R split2907 (.A(_18464_),
    .Y(net3312));
 BUFx3_ASAP7_75t_R rebuffer2908 (.A(_17670_),
    .Y(net3313));
 BUFx6f_ASAP7_75t_R rebuffer2909 (.A(_04917_),
    .Y(net3314));
 BUFx16f_ASAP7_75t_R rebuffer2910 (.A(_01256_),
    .Y(net3315));
 BUFx2_ASAP7_75t_R rebuffer2911 (.A(net3315),
    .Y(net3316));
 BUFx6f_ASAP7_75t_R split2912 (.A(_19356_),
    .Y(net3317));
 BUFx4f_ASAP7_75t_R split2913 (.A(net1414),
    .Y(net3318));
 BUFx2_ASAP7_75t_R rebuffer2914 (.A(_10311_),
    .Y(net3319));
 BUFx4f_ASAP7_75t_R split2915 (.A(net1752),
    .Y(net3320));
 BUFx6f_ASAP7_75t_R rebuffer2916 (.A(_01146_),
    .Y(net3321));
 BUFx2_ASAP7_75t_R rebuffer2917 (.A(net3321),
    .Y(net3322));
 BUFx6f_ASAP7_75t_R rebuffer2918 (.A(_17534_),
    .Y(net3323));
 BUFx3_ASAP7_75t_R rebuffer2919 (.A(_18712_),
    .Y(net3324));
 BUFx3_ASAP7_75t_R rebuffer2920 (.A(_18712_),
    .Y(net3325));
 BUFx6f_ASAP7_75t_R rebuffer2921 (.A(_18295_),
    .Y(net3326));
 BUFx3_ASAP7_75t_R split2922 (.A(_06142_),
    .Y(net3327));
 BUFx6f_ASAP7_75t_R split2923 (.A(_06129_),
    .Y(net3328));
 BUFx3_ASAP7_75t_R split2924 (.A(_06141_),
    .Y(net3329));
 BUFx6f_ASAP7_75t_R split2925 (.A(_06107_),
    .Y(net3330));
 BUFx2_ASAP7_75t_R rebuffer2926 (.A(_06089_),
    .Y(net3331));
 BUFx3_ASAP7_75t_R rebuffer2927 (.A(_01815_),
    .Y(net3332));
 BUFx3_ASAP7_75t_R rebuffer2928 (.A(_10578_),
    .Y(net3333));
 BUFx6f_ASAP7_75t_R rebuffer2929 (.A(_13906_),
    .Y(net3334));
 BUFx3_ASAP7_75t_R split2930 (.A(net1855),
    .Y(net3335));
 BUFx6f_ASAP7_75t_R rebuffer2931 (.A(_11426_),
    .Y(net3336));
 BUFx2_ASAP7_75t_R rebuffer2932 (.A(net3336),
    .Y(net3337));
 BUFx6f_ASAP7_75t_R split2933 (.A(_10316_),
    .Y(net3338));
 BUFx4f_ASAP7_75t_R split2935 (.A(_04525_),
    .Y(net3340));
 BUFx6f_ASAP7_75t_R rebuffer2936 (.A(_01128_),
    .Y(net3341));
 BUFx3_ASAP7_75t_R rebuffer2937 (.A(_19451_),
    .Y(net3342));
 BUFx3_ASAP7_75t_R split2938 (.A(net1790),
    .Y(net3343));
 BUFx6f_ASAP7_75t_R rebuffer2941 (.A(_19356_),
    .Y(net3346));
 BUFx3_ASAP7_75t_R rebuffer2942 (.A(_08850_),
    .Y(net3347));
 BUFx3_ASAP7_75t_R split2943 (.A(_05845_),
    .Y(net3348));
 BUFx4f_ASAP7_75t_R split2944 (.A(_05462_),
    .Y(net3349));
 BUFx3_ASAP7_75t_R split2945 (.A(_05643_),
    .Y(net3350));
 BUFx4f_ASAP7_75t_R split2946 (.A(_05821_),
    .Y(net3351));
 BUFx12f_ASAP7_75t_R rebuffer2947 (.A(_05951_),
    .Y(net3352));
 BUFx2_ASAP7_75t_R rebuffer2948 (.A(_05717_),
    .Y(net3353));
 BUFx2_ASAP7_75t_R rebuffer2949 (.A(_05717_),
    .Y(net3354));
 BUFx2_ASAP7_75t_R rebuffer2950 (.A(_05887_),
    .Y(net3355));
 BUFx6f_ASAP7_75t_R rebuffer2951 (.A(_05643_),
    .Y(net3356));
 BUFx3_ASAP7_75t_R split2952 (.A(_05857_),
    .Y(net3357));
 BUFx2_ASAP7_75t_R rebuffer2953 (.A(_00540_),
    .Y(net3358));
 BUFx6f_ASAP7_75t_R rebuffer2954 (.A(_00540_),
    .Y(net3359));
 BUFx2_ASAP7_75t_R rebuffer2955 (.A(net3359),
    .Y(net3360));
 BUFx6f_ASAP7_75t_R rebuffer2956 (.A(_00571_),
    .Y(net3361));
 BUFx2_ASAP7_75t_R rebuffer2957 (.A(net3361),
    .Y(net3362));
 BUFx3_ASAP7_75t_R rebuffer2958 (.A(_14093_),
    .Y(net3363));
 BUFx6f_ASAP7_75t_R rebuffer2959 (.A(_14090_),
    .Y(net3364));
 BUFx4f_ASAP7_75t_R split2961 (.A(_17941_),
    .Y(net3366));
 BUFx3_ASAP7_75t_R rebuffer2962 (.A(_18130_),
    .Y(net3367));
 BUFx4f_ASAP7_75t_R split2963 (.A(_05728_),
    .Y(net3368));
 BUFx6f_ASAP7_75t_R split2964 (.A(_05156_),
    .Y(net3369));
 BUFx12f_ASAP7_75t_R rebuffer2965 (.A(_05825_),
    .Y(net3370));
 BUFx2_ASAP7_75t_R rebuffer2966 (.A(net3370),
    .Y(net3371));
 BUFx4f_ASAP7_75t_R rebuffer2967 (.A(net3370),
    .Y(net3372));
 BUFx12f_ASAP7_75t_R rebuffer2968 (.A(_05510_),
    .Y(net3373));
 BUFx2_ASAP7_75t_R rebuffer2969 (.A(net3373),
    .Y(net3374));
 BUFx4f_ASAP7_75t_R split2970 (.A(net980),
    .Y(net3375));
 BUFx4f_ASAP7_75t_R split2971 (.A(_18559_),
    .Y(net3376));
 BUFx6f_ASAP7_75t_R rebuffer2972 (.A(_18559_),
    .Y(net3377));
 BUFx4f_ASAP7_75t_R rebuffer2973 (.A(_18528_),
    .Y(net3378));
 BUFx2_ASAP7_75t_R rebuffer2974 (.A(net3378),
    .Y(net3379));
 BUFx4f_ASAP7_75t_R split2975 (.A(_18554_),
    .Y(net3380));
 BUFx3_ASAP7_75t_R split2976 (.A(_18721_),
    .Y(net3381));
 BUFx6f_ASAP7_75t_R rebuffer2977 (.A(_07499_),
    .Y(net3382));
 BUFx2_ASAP7_75t_R rebuffer2978 (.A(net3382),
    .Y(net3383));
 BUFx2_ASAP7_75t_R rebuffer2979 (.A(_00578_),
    .Y(net3384));
 BUFx2_ASAP7_75t_R rebuffer2980 (.A(_00421_),
    .Y(net3385));
 BUFx2_ASAP7_75t_R rebuffer2981 (.A(_00421_),
    .Y(net3386));
 BUFx2_ASAP7_75t_R rebuffer2982 (.A(_00421_),
    .Y(net3387));
 BUFx2_ASAP7_75t_R rebuffer2983 (.A(_05870_),
    .Y(net3388));
 BUFx2_ASAP7_75t_R rebuffer2984 (.A(_05870_),
    .Y(net3389));
 BUFx2_ASAP7_75t_R rebuffer2985 (.A(_06123_),
    .Y(net3390));
 BUFx2_ASAP7_75t_R rebuffer2986 (.A(net3390),
    .Y(net3391));
 BUFx4f_ASAP7_75t_R split2987 (.A(_05958_),
    .Y(net3392));
 BUFx2_ASAP7_75t_R rebuffer2988 (.A(_06277_),
    .Y(net3393));
 BUFx2_ASAP7_75t_R rebuffer2989 (.A(net3393),
    .Y(net3394));
 BUFx12f_ASAP7_75t_R rebuffer2990 (.A(_00426_),
    .Y(net3395));
 BUFx2_ASAP7_75t_R rebuffer2991 (.A(net3395),
    .Y(net3396));
 BUFx2_ASAP7_75t_R rebuffer2992 (.A(_00426_),
    .Y(net3397));
 BUFx3_ASAP7_75t_R split2993 (.A(_05958_),
    .Y(net3398));
 BUFx6f_ASAP7_75t_R rebuffer2994 (.A(_00425_),
    .Y(net3399));
 BUFx2_ASAP7_75t_R rebuffer2995 (.A(net3399),
    .Y(net3400));
 BUFx2_ASAP7_75t_R rebuffer2996 (.A(net3400),
    .Y(net3401));
 BUFx2_ASAP7_75t_R rebuffer2997 (.A(net3399),
    .Y(net3402));
 BUFx3_ASAP7_75t_R split2998 (.A(_06277_),
    .Y(net3403));
 BUFx3_ASAP7_75t_R rebuffer3004 (.A(_05191_),
    .Y(net3409));
 BUFx2_ASAP7_75t_R rebuffer3005 (.A(_05126_),
    .Y(net3410));
 BUFx3_ASAP7_75t_R rebuffer3006 (.A(net3410),
    .Y(net3411));
 BUFx6f_ASAP7_75t_R rebuffer3007 (.A(_05126_),
    .Y(net3412));
 BUFx2_ASAP7_75t_R rebuffer3010 (.A(_01496_),
    .Y(net3415));
 BUFx6f_ASAP7_75t_R rebuffer3011 (.A(_01495_),
    .Y(net3416));
 BUFx6f_ASAP7_75t_R split3012 (.A(_01276_),
    .Y(net3417));
 BUFx2_ASAP7_75t_R rebuffer3013 (.A(_07593_),
    .Y(net3418));
 BUFx4f_ASAP7_75t_R split3014 (.A(_06420_),
    .Y(net3419));
 BUFx6f_ASAP7_75t_R rebuffer3015 (.A(_07159_),
    .Y(net3420));
 BUFx2_ASAP7_75t_R rebuffer3016 (.A(_06097_),
    .Y(net3421));
 BUFx2_ASAP7_75t_R rebuffer3017 (.A(_06097_),
    .Y(net3422));
 BUFx2_ASAP7_75t_R rebuffer3018 (.A(_06097_),
    .Y(net3423));
 BUFx6f_ASAP7_75t_R rebuffer3019 (.A(_06097_),
    .Y(net3424));
 BUFx2_ASAP7_75t_R rebuffer3020 (.A(net3424),
    .Y(net3425));
 BUFx6f_ASAP7_75t_R split3021 (.A(net1822),
    .Y(net3426));
 BUFx3_ASAP7_75t_R rebuffer3022 (.A(_05157_),
    .Y(net3427));
 BUFx2_ASAP7_75t_R rebuffer3023 (.A(_05329_),
    .Y(net3428));
 BUFx4f_ASAP7_75t_R rebuffer3024 (.A(_06071_),
    .Y(net3429));
 BUFx2_ASAP7_75t_R rebuffer3025 (.A(_06109_),
    .Y(net3430));
 BUFx2_ASAP7_75t_R rebuffer3026 (.A(_06765_),
    .Y(net3431));
 BUFx2_ASAP7_75t_R rebuffer3027 (.A(_06765_),
    .Y(net3432));
 BUFx3_ASAP7_75t_R split3028 (.A(_06063_),
    .Y(net3433));
 BUFx2_ASAP7_75t_R rebuffer3029 (.A(_06131_),
    .Y(net3434));
 BUFx6f_ASAP7_75t_R rebuffer3030 (.A(_06420_),
    .Y(net3435));
 BUFx4f_ASAP7_75t_R split3031 (.A(net3439),
    .Y(net3436));
 BUFx2_ASAP7_75t_R rebuffer3032 (.A(_06363_),
    .Y(net3437));
 BUFx4f_ASAP7_75t_R split3033 (.A(net1319),
    .Y(net3438));
 BUFx3_ASAP7_75t_R split3034 (.A(_05103_),
    .Y(net3439));
 BUFx4f_ASAP7_75t_R split3035 (.A(_05163_),
    .Y(net3440));
 BUFx2_ASAP7_75t_R rebuffer3036 (.A(_06889_),
    .Y(net3441));
 BUFx4f_ASAP7_75t_R split3037 (.A(_05068_),
    .Y(net3442));
 BUFx3_ASAP7_75t_R rebuffer3038 (.A(_05104_),
    .Y(net3443));
 BUFx3_ASAP7_75t_R rebuffer3039 (.A(_05118_),
    .Y(net3444));
 BUFx2_ASAP7_75t_R rebuffer3040 (.A(_05190_),
    .Y(net3445));
 BUFx6f_ASAP7_75t_R split3041 (.A(_05225_),
    .Y(net3446));
 BUFx2_ASAP7_75t_R rebuffer3042 (.A(_05449_),
    .Y(net3447));
 BUFx6f_ASAP7_75t_R rebuffer3043 (.A(_08853_),
    .Y(net3448));
 BUFx6f_ASAP7_75t_R rebuffer3044 (.A(_05156_),
    .Y(net3449));
 BUFx2_ASAP7_75t_R rebuffer3045 (.A(_05561_),
    .Y(net3450));
 BUFx3_ASAP7_75t_R rebuffer3046 (.A(_05185_),
    .Y(net3451));
 BUFx2_ASAP7_75t_R rebuffer3047 (.A(net3451),
    .Y(net3452));
 BUFx2_ASAP7_75t_R rebuffer3048 (.A(net3451),
    .Y(net3453));
 BUFx2_ASAP7_75t_R rebuffer3049 (.A(_05185_),
    .Y(net3454));
 BUFx3_ASAP7_75t_R split3050 (.A(_05174_),
    .Y(net3455));
 BUFx6f_ASAP7_75t_R rebuffer3051 (.A(_05104_),
    .Y(net3456));
 BUFx2_ASAP7_75t_R rebuffer3052 (.A(net3456),
    .Y(net3457));
 BUFx2_ASAP7_75t_R rebuffer3053 (.A(_05515_),
    .Y(net3458));
 BUFx2_ASAP7_75t_R rebuffer3054 (.A(_05515_),
    .Y(net3459));
 BUFx2_ASAP7_75t_R rebuffer3055 (.A(net3459),
    .Y(net3460));
 BUFx6f_ASAP7_75t_R split3056 (.A(net2548),
    .Y(net3461));
 BUFx3_ASAP7_75t_R rebuffer3057 (.A(_05535_),
    .Y(net3462));
 BUFx3_ASAP7_75t_R rebuffer3058 (.A(_05466_),
    .Y(net3463));
 BUFx2_ASAP7_75t_R rebuffer3061 (.A(_06429_),
    .Y(net3466));
 BUFx3_ASAP7_75t_R rebuffer3062 (.A(_05833_),
    .Y(net3467));
 BUFx2_ASAP7_75t_R rebuffer3063 (.A(net3467),
    .Y(net3468));
 BUFx2_ASAP7_75t_R rebuffer3064 (.A(net3467),
    .Y(net3469));
 BUFx2_ASAP7_75t_R rebuffer3065 (.A(net3467),
    .Y(net3470));
 BUFx3_ASAP7_75t_R rebuffer3066 (.A(_06429_),
    .Y(net3471));
 BUFx6f_ASAP7_75t_R rebuffer3067 (.A(_06158_),
    .Y(net3472));
 BUFx3_ASAP7_75t_R rebuffer3068 (.A(_06799_),
    .Y(net3473));
 BUFx2_ASAP7_75t_R rebuffer3069 (.A(_05766_),
    .Y(net3474));
 BUFx6f_ASAP7_75t_R rebuffer3070 (.A(_05766_),
    .Y(net3475));
 BUFx2_ASAP7_75t_R rebuffer3071 (.A(net3475),
    .Y(net3476));
 BUFx3_ASAP7_75t_R rebuffer3072 (.A(_00435_),
    .Y(net3477));
 BUFx2_ASAP7_75t_R rebuffer3073 (.A(net3477),
    .Y(net3478));
 BUFx12f_ASAP7_75t_R rebuffer3074 (.A(_00435_),
    .Y(net3479));
 BUFx2_ASAP7_75t_R rebuffer3075 (.A(net3479),
    .Y(net3480));
 BUFx2_ASAP7_75t_R rebuffer3076 (.A(net3480),
    .Y(net3481));
 BUFx2_ASAP7_75t_R rebuffer3077 (.A(_00435_),
    .Y(net3482));
 BUFx2_ASAP7_75t_R rebuffer3078 (.A(_00434_),
    .Y(net3483));
 BUFx3_ASAP7_75t_R rebuffer3079 (.A(_00434_),
    .Y(net3484));
 BUFx2_ASAP7_75t_R rebuffer3080 (.A(net3484),
    .Y(net3485));
 BUFx6f_ASAP7_75t_R rebuffer3081 (.A(net3485),
    .Y(net3486));
 BUFx2_ASAP7_75t_R rebuffer3082 (.A(_00433_),
    .Y(net3487));
 BUFx2_ASAP7_75t_R rebuffer3083 (.A(net3487),
    .Y(net3488));
 BUFx6f_ASAP7_75t_R rebuffer3084 (.A(_00433_),
    .Y(net3489));
 BUFx2_ASAP7_75t_R rebuffer3085 (.A(net3489),
    .Y(net3490));
 BUFx2_ASAP7_75t_R rebuffer3086 (.A(net3489),
    .Y(net3491));
 BUFx2_ASAP7_75t_R rebuffer3087 (.A(_00433_),
    .Y(net3492));
 BUFx2_ASAP7_75t_R split3088 (.A(_16277_),
    .Y(net3493));
 BUFx6f_ASAP7_75t_R rebuffer3089 (.A(_00431_),
    .Y(net3494));
 BUFx2_ASAP7_75t_R rebuffer3090 (.A(net3494),
    .Y(net3495));
 BUFx2_ASAP7_75t_R rebuffer3091 (.A(net3495),
    .Y(net3496));
 BUFx2_ASAP7_75t_R rebuffer3092 (.A(net3494),
    .Y(net3497));
 BUFx2_ASAP7_75t_R rebuffer3093 (.A(_16267_),
    .Y(net3498));
 BUFx4f_ASAP7_75t_R split3094 (.A(_16542_),
    .Y(net3499));
 BUFx2_ASAP7_75t_R rebuffer3095 (.A(_00432_),
    .Y(net3500));
 BUFx2_ASAP7_75t_R rebuffer3096 (.A(_00432_),
    .Y(net3501));
 BUFx2_ASAP7_75t_R rebuffer3097 (.A(net3501),
    .Y(net3502));
 BUFx2_ASAP7_75t_R rebuffer3098 (.A(_16293_),
    .Y(net3503));
 BUFx2_ASAP7_75t_R rebuffer3099 (.A(net3503),
    .Y(net3504));
 BUFx2_ASAP7_75t_R rebuffer3100 (.A(_14633_),
    .Y(net3505));
 BUFx6f_ASAP7_75t_R rebuffer3101 (.A(_14625_),
    .Y(net3506));
 BUFx3_ASAP7_75t_R rebuffer3102 (.A(net3506),
    .Y(net3507));
 BUFx2_ASAP7_75t_R rebuffer3103 (.A(net3507),
    .Y(net3508));
 BUFx6f_ASAP7_75t_R split3104 (.A(_14764_),
    .Y(net3509));
 BUFx6f_ASAP7_75t_R rebuffer3105 (.A(_14692_),
    .Y(net3510));
 BUFx2_ASAP7_75t_R rebuffer3106 (.A(net3510),
    .Y(net3511));
 BUFx2_ASAP7_75t_R rebuffer3107 (.A(_00452_),
    .Y(net3512));
 BUFx6f_ASAP7_75t_R rebuffer3108 (.A(_00452_),
    .Y(net3513));
 BUFx2_ASAP7_75t_R rebuffer3109 (.A(net3513),
    .Y(net3514));
 BUFx6f_ASAP7_75t_R rebuffer3110 (.A(net3513),
    .Y(net3515));
 BUFx2_ASAP7_75t_R rebuffer3111 (.A(_00452_),
    .Y(net3516));
 BUFx2_ASAP7_75t_R rebuffer3112 (.A(net3516),
    .Y(net3517));
 BUFx3_ASAP7_75t_R rebuffer3113 (.A(_14617_),
    .Y(net3518));
 BUFx2_ASAP7_75t_R rebuffer3114 (.A(net3518),
    .Y(net3519));
 BUFx2_ASAP7_75t_R rebuffer3115 (.A(net3518),
    .Y(net3520));
 BUFx2_ASAP7_75t_R rebuffer3116 (.A(_14660_),
    .Y(net3521));
 BUFx2_ASAP7_75t_R rebuffer3117 (.A(net3521),
    .Y(net3522));
 BUFx2_ASAP7_75t_R rebuffer3118 (.A(_14635_),
    .Y(net3523));
 BUFx2_ASAP7_75t_R split3119 (.A(_14622_),
    .Y(net3524));
 BUFx2_ASAP7_75t_R rebuffer3120 (.A(_14614_),
    .Y(net3525));
 BUFx12f_ASAP7_75t_R rebuffer3121 (.A(_00450_),
    .Y(net3526));
 BUFx2_ASAP7_75t_R rebuffer3122 (.A(net3526),
    .Y(net3527));
 BUFx2_ASAP7_75t_R rebuffer3123 (.A(net3526),
    .Y(net3528));
 BUFx2_ASAP7_75t_R rebuffer3124 (.A(net3526),
    .Y(net3529));
 BUFx2_ASAP7_75t_R rebuffer3125 (.A(net3526),
    .Y(net3530));
 BUFx2_ASAP7_75t_R rebuffer3126 (.A(_00449_),
    .Y(net3531));
 BUFx2_ASAP7_75t_R rebuffer3127 (.A(_00449_),
    .Y(net3532));
 BUFx2_ASAP7_75t_R rebuffer3128 (.A(net3532),
    .Y(net3533));
 BUFx2_ASAP7_75t_R rebuffer3129 (.A(_00449_),
    .Y(net3534));
 BUFx6f_ASAP7_75t_R rebuffer3130 (.A(_14766_),
    .Y(net3535));
 BUFx2_ASAP7_75t_R rebuffer3131 (.A(net3535),
    .Y(net3536));
 BUFx3_ASAP7_75t_R rebuffer3132 (.A(net3535),
    .Y(net3537));
 BUFx2_ASAP7_75t_R rebuffer3133 (.A(net3535),
    .Y(net3538));
 BUFx2_ASAP7_75t_R rebuffer3134 (.A(_14735_),
    .Y(net3539));
 BUFx3_ASAP7_75t_R split3135 (.A(_15504_),
    .Y(net3540));
 BUFx4f_ASAP7_75t_R split3136 (.A(_15496_),
    .Y(net3541));
 BUFx2_ASAP7_75t_R split3137 (.A(_15694_),
    .Y(net3542));
 BUFx2_ASAP7_75t_R rebuffer3138 (.A(_00443_),
    .Y(net3543));
 BUFx12f_ASAP7_75t_R rebuffer3139 (.A(_00443_),
    .Y(net3544));
 BUFx2_ASAP7_75t_R rebuffer3140 (.A(net3544),
    .Y(net3545));
 BUFx2_ASAP7_75t_R rebuffer3141 (.A(_00443_),
    .Y(net3546));
 BUFx2_ASAP7_75t_R rebuffer3142 (.A(_00444_),
    .Y(net3547));
 BUFx6f_ASAP7_75t_R rebuffer3143 (.A(_00444_),
    .Y(net3548));
 BUFx2_ASAP7_75t_R rebuffer3144 (.A(net3548),
    .Y(net3549));
 BUFx2_ASAP7_75t_R rebuffer3145 (.A(net3549),
    .Y(net3550));
 BUFx2_ASAP7_75t_R rebuffer3146 (.A(_00444_),
    .Y(net3551));
 BUFx2_ASAP7_75t_R rebuffer3147 (.A(_00444_),
    .Y(net3552));
 BUFx12f_ASAP7_75t_R rebuffer3148 (.A(_15434_),
    .Y(net3553));
 BUFx6f_ASAP7_75t_R rebuffer3149 (.A(net3553),
    .Y(net3554));
 BUFx2_ASAP7_75t_R rebuffer3150 (.A(net3553),
    .Y(net3555));
 BUFx2_ASAP7_75t_R rebuffer3151 (.A(_15428_),
    .Y(net3556));
 BUFx2_ASAP7_75t_R rebuffer3152 (.A(net3556),
    .Y(net3557));
 BUFx2_ASAP7_75t_R rebuffer3153 (.A(_15428_),
    .Y(net3558));
 BUFx2_ASAP7_75t_R rebuffer3154 (.A(_15428_),
    .Y(net3559));
 BUFx2_ASAP7_75t_R rebuffer3155 (.A(net3561),
    .Y(net3560));
 BUFx3_ASAP7_75t_R split3156 (.A(_15415_),
    .Y(net3561));
 BUFx4f_ASAP7_75t_R split3157 (.A(_15409_),
    .Y(net3562));
 BUFx2_ASAP7_75t_R rebuffer3158 (.A(_15409_),
    .Y(net3563));
 BUFx2_ASAP7_75t_R hold3159 (.A(net4212),
    .Y(net3564));
 BUFx2_ASAP7_75t_R hold3160 (.A(net247),
    .Y(net3565));
 BUFx2_ASAP7_75t_R hold3161 (.A(_00938_),
    .Y(net3566));
 BUFx2_ASAP7_75t_R hold3162 (.A(net4213),
    .Y(net3567));
 BUFx2_ASAP7_75t_R hold3163 (.A(net139),
    .Y(net3568));
 BUFx2_ASAP7_75t_R hold3164 (.A(_01037_),
    .Y(net3569));
 BUFx2_ASAP7_75t_R hold3165 (.A(net4214),
    .Y(net3570));
 BUFx2_ASAP7_75t_R hold3166 (.A(net225),
    .Y(net3571));
 BUFx2_ASAP7_75t_R hold3167 (.A(_00936_),
    .Y(net3572));
 BUFx2_ASAP7_75t_R hold3168 (.A(net4215),
    .Y(net3573));
 BUFx2_ASAP7_75t_R hold3169 (.A(net258),
    .Y(net3574));
 BUFx2_ASAP7_75t_R hold3170 (.A(_00939_),
    .Y(net3575));
 BUFx2_ASAP7_75t_R hold3171 (.A(net4216),
    .Y(net3576));
 BUFx2_ASAP7_75t_R hold3172 (.A(net173),
    .Y(net3577));
 BUFx2_ASAP7_75t_R hold3173 (.A(_00952_),
    .Y(net3578));
 BUFx2_ASAP7_75t_R hold3174 (.A(net4220),
    .Y(net3579));
 BUFx2_ASAP7_75t_R hold3175 (.A(net209),
    .Y(net3580));
 BUFx2_ASAP7_75t_R hold3176 (.A(_00985_),
    .Y(net3581));
 BUFx2_ASAP7_75t_R hold3177 (.A(net4217),
    .Y(net3582));
 BUFx2_ASAP7_75t_R hold3178 (.A(net219),
    .Y(net3583));
 BUFx2_ASAP7_75t_R hold3179 (.A(_00994_),
    .Y(net3584));
 BUFx2_ASAP7_75t_R hold3180 (.A(net4219),
    .Y(net3585));
 BUFx2_ASAP7_75t_R hold3181 (.A(net142),
    .Y(net3586));
 BUFx2_ASAP7_75t_R hold3182 (.A(_00940_),
    .Y(net3587));
 BUFx2_ASAP7_75t_R hold3183 (.A(net4218),
    .Y(net3588));
 BUFx2_ASAP7_75t_R hold3184 (.A(net246),
    .Y(net3589));
 BUFx2_ASAP7_75t_R hold3185 (.A(_01019_),
    .Y(net3590));
 BUFx2_ASAP7_75t_R hold3186 (.A(net4207),
    .Y(net3591));
 BUFx2_ASAP7_75t_R hold3187 (.A(net17),
    .Y(net3592));
 BUFx2_ASAP7_75t_R hold3188 (.A(net4222),
    .Y(net3593));
 BUFx2_ASAP7_75t_R hold3189 (.A(net207),
    .Y(net3594));
 BUFx2_ASAP7_75t_R hold3190 (.A(_00983_),
    .Y(net3595));
 BUFx2_ASAP7_75t_R hold3191 (.A(net4224),
    .Y(net3596));
 BUFx2_ASAP7_75t_R hold3192 (.A(net241),
    .Y(net3597));
 BUFx2_ASAP7_75t_R hold3193 (.A(_01014_),
    .Y(net3598));
 BUFx2_ASAP7_75t_R hold3194 (.A(net4223),
    .Y(net3599));
 BUFx2_ASAP7_75t_R hold3195 (.A(net251),
    .Y(net3600));
 BUFx2_ASAP7_75t_R hold3196 (.A(_01023_),
    .Y(net3601));
 BUFx2_ASAP7_75t_R hold3197 (.A(net4225),
    .Y(net3602));
 BUFx2_ASAP7_75t_R hold3198 (.A(net253),
    .Y(net3603));
 BUFx2_ASAP7_75t_R hold3199 (.A(_01025_),
    .Y(net3604));
 BUFx2_ASAP7_75t_R hold3200 (.A(net4233),
    .Y(net3605));
 BUFx2_ASAP7_75t_R hold3201 (.A(net233),
    .Y(net3606));
 BUFx2_ASAP7_75t_R hold3202 (.A(_01007_),
    .Y(net3607));
 BUFx2_ASAP7_75t_R hold3203 (.A(net4231),
    .Y(net3608));
 BUFx2_ASAP7_75t_R hold3204 (.A(net204),
    .Y(net3609));
 BUFx2_ASAP7_75t_R hold3205 (.A(_00980_),
    .Y(net3610));
 BUFx2_ASAP7_75t_R hold3206 (.A(text_in[83]),
    .Y(net3611));
 BUFx2_ASAP7_75t_R hold3207 (.A(net240),
    .Y(net3612));
 BUFx2_ASAP7_75t_R hold3208 (.A(_01013_),
    .Y(net3613));
 BUFx2_ASAP7_75t_R hold3209 (.A(net4227),
    .Y(net3614));
 BUFx2_ASAP7_75t_R hold3210 (.A(net220),
    .Y(net3615));
 BUFx2_ASAP7_75t_R hold3211 (.A(_00995_),
    .Y(net3616));
 BUFx2_ASAP7_75t_R hold3212 (.A(net4229),
    .Y(net3617));
 BUFx2_ASAP7_75t_R hold3213 (.A(net215),
    .Y(net3618));
 BUFx2_ASAP7_75t_R hold3214 (.A(_00990_),
    .Y(net3619));
 BUFx2_ASAP7_75t_R hold3215 (.A(net4226),
    .Y(net3620));
 BUFx2_ASAP7_75t_R hold3216 (.A(net236),
    .Y(net3621));
 BUFx2_ASAP7_75t_R hold3217 (.A(_00937_),
    .Y(net3622));
 BUFx2_ASAP7_75t_R hold3218 (.A(net4234),
    .Y(net3623));
 BUFx2_ASAP7_75t_R hold3219 (.A(net198),
    .Y(net3624));
 BUFx2_ASAP7_75t_R hold3220 (.A(_00975_),
    .Y(net3625));
 BUFx2_ASAP7_75t_R hold3221 (.A(net4230),
    .Y(net3626));
 BUFx2_ASAP7_75t_R hold3222 (.A(net245),
    .Y(net3627));
 BUFx2_ASAP7_75t_R hold3223 (.A(_01018_),
    .Y(net3628));
 BUFx2_ASAP7_75t_R hold3224 (.A(net4228),
    .Y(net3629));
 BUFx2_ASAP7_75t_R hold3225 (.A(net237),
    .Y(net3630));
 BUFx2_ASAP7_75t_R hold3226 (.A(_01010_),
    .Y(net3631));
 BUFx2_ASAP7_75t_R hold3227 (.A(text_in[54]),
    .Y(net3632));
 BUFx2_ASAP7_75t_R hold3228 (.A(net208),
    .Y(net3633));
 BUFx2_ASAP7_75t_R hold3229 (.A(_00984_),
    .Y(net3634));
 BUFx2_ASAP7_75t_R hold3230 (.A(text_in[44]),
    .Y(net3635));
 BUFx2_ASAP7_75t_R hold3231 (.A(net197),
    .Y(net3636));
 BUFx2_ASAP7_75t_R hold3232 (.A(_00974_),
    .Y(net3637));
 BUFx2_ASAP7_75t_R hold3233 (.A(text_in[35]),
    .Y(net3638));
 BUFx2_ASAP7_75t_R hold3234 (.A(net187),
    .Y(net3639));
 BUFx2_ASAP7_75t_R hold3235 (.A(_00965_),
    .Y(net3640));
 BUFx2_ASAP7_75t_R hold3236 (.A(net4232),
    .Y(net3641));
 BUFx2_ASAP7_75t_R hold3237 (.A(net203),
    .Y(net3642));
 BUFx2_ASAP7_75t_R hold3238 (.A(_00934_),
    .Y(net3643));
 BUFx2_ASAP7_75t_R hold3239 (.A(text_in[43]),
    .Y(net3644));
 BUFx2_ASAP7_75t_R hold3240 (.A(net196),
    .Y(net3645));
 BUFx2_ASAP7_75t_R hold3241 (.A(_00973_),
    .Y(net3646));
 BUFx2_ASAP7_75t_R hold3242 (.A(text_in[58]),
    .Y(net3647));
 BUFx2_ASAP7_75t_R hold3243 (.A(net212),
    .Y(net3648));
 BUFx2_ASAP7_75t_R hold3244 (.A(_00988_),
    .Y(net3649));
 BUFx2_ASAP7_75t_R hold3245 (.A(net4209),
    .Y(net3650));
 BUFx2_ASAP7_75t_R hold3246 (.A(net74),
    .Y(net3651));
 BUFx2_ASAP7_75t_R hold3247 (.A(text_in[81]),
    .Y(net3652));
 BUFx2_ASAP7_75t_R hold3248 (.A(net238),
    .Y(net3653));
 BUFx2_ASAP7_75t_R hold3249 (.A(_01011_),
    .Y(net3654));
 BUFx2_ASAP7_75t_R hold3250 (.A(text_in[63]),
    .Y(net3655));
 BUFx2_ASAP7_75t_R hold3251 (.A(net218),
    .Y(net3656));
 BUFx2_ASAP7_75t_R hold3252 (.A(_00993_),
    .Y(net3657));
 BUFx2_ASAP7_75t_R hold3253 (.A(key[21]),
    .Y(net3658));
 BUFx2_ASAP7_75t_R hold3254 (.A(net42),
    .Y(net3659));
 BUFx2_ASAP7_75t_R hold3255 (.A(_16056_),
    .Y(net3660));
 BUFx2_ASAP7_75t_R hold3256 (.A(text_in[72]),
    .Y(net3661));
 BUFx2_ASAP7_75t_R hold3257 (.A(net228),
    .Y(net3662));
 BUFx2_ASAP7_75t_R hold3258 (.A(_01002_),
    .Y(net3663));
 BUFx2_ASAP7_75t_R hold3259 (.A(text_in[17]),
    .Y(net3664));
 BUFx2_ASAP7_75t_R hold3260 (.A(net167),
    .Y(net3665));
 BUFx2_ASAP7_75t_R hold3261 (.A(_00947_),
    .Y(net3666));
 BUFx2_ASAP7_75t_R hold3262 (.A(text_in[49]),
    .Y(net3667));
 BUFx2_ASAP7_75t_R hold3263 (.A(net202),
    .Y(net3668));
 BUFx2_ASAP7_75t_R hold3264 (.A(_00979_),
    .Y(net3669));
 BUFx2_ASAP7_75t_R hold3265 (.A(text_in[66]),
    .Y(net3670));
 BUFx2_ASAP7_75t_R hold3266 (.A(net221),
    .Y(net3671));
 BUFx2_ASAP7_75t_R hold3267 (.A(_00996_),
    .Y(net3672));
 BUFx2_ASAP7_75t_R hold3268 (.A(text_in[90]),
    .Y(net3673));
 BUFx2_ASAP7_75t_R hold3269 (.A(net248),
    .Y(net3674));
 BUFx2_ASAP7_75t_R hold3270 (.A(_01020_),
    .Y(net3675));
 BUFx2_ASAP7_75t_R hold3271 (.A(text_in[92]),
    .Y(net3676));
 BUFx2_ASAP7_75t_R hold3272 (.A(net250),
    .Y(net3677));
 BUFx2_ASAP7_75t_R hold3273 (.A(_01022_),
    .Y(net3678));
 BUFx2_ASAP7_75t_R hold3274 (.A(text_in[41]),
    .Y(net3679));
 BUFx2_ASAP7_75t_R hold3275 (.A(net194),
    .Y(net3680));
 BUFx2_ASAP7_75t_R hold3276 (.A(_00971_),
    .Y(net3681));
 BUFx2_ASAP7_75t_R hold3277 (.A(text_in[48]),
    .Y(net3682));
 BUFx2_ASAP7_75t_R hold3278 (.A(net201),
    .Y(net3683));
 BUFx2_ASAP7_75t_R hold3279 (.A(_00978_),
    .Y(net3684));
 BUFx2_ASAP7_75t_R hold3280 (.A(text_in[23]),
    .Y(net3685));
 BUFx2_ASAP7_75t_R hold3281 (.A(net174),
    .Y(net3686));
 BUFx2_ASAP7_75t_R hold3282 (.A(_00953_),
    .Y(net3687));
 BUFx2_ASAP7_75t_R hold3283 (.A(text_in[62]),
    .Y(net3688));
 BUFx2_ASAP7_75t_R hold3284 (.A(net217),
    .Y(net3689));
 BUFx2_ASAP7_75t_R hold3285 (.A(_00992_),
    .Y(net3690));
 BUFx2_ASAP7_75t_R hold3286 (.A(text_in[40]),
    .Y(net3691));
 BUFx2_ASAP7_75t_R hold3287 (.A(net193),
    .Y(net3692));
 BUFx2_ASAP7_75t_R hold3288 (.A(_00970_),
    .Y(net3693));
 BUFx2_ASAP7_75t_R hold3289 (.A(text_in[51]),
    .Y(net3694));
 BUFx2_ASAP7_75t_R hold3290 (.A(net205),
    .Y(net3695));
 BUFx2_ASAP7_75t_R hold3291 (.A(_00981_),
    .Y(net3696));
 BUFx2_ASAP7_75t_R hold3292 (.A(text_in[42]),
    .Y(net3697));
 BUFx2_ASAP7_75t_R hold3293 (.A(net195),
    .Y(net3698));
 BUFx2_ASAP7_75t_R hold3294 (.A(_00972_),
    .Y(net3699));
 BUFx2_ASAP7_75t_R hold3295 (.A(text_in[12]),
    .Y(net3700));
 BUFx2_ASAP7_75t_R hold3296 (.A(net162),
    .Y(net3701));
 BUFx2_ASAP7_75t_R hold3297 (.A(_00942_),
    .Y(net3702));
 BUFx2_ASAP7_75t_R hold3298 (.A(text_in[59]),
    .Y(net3703));
 BUFx2_ASAP7_75t_R hold3299 (.A(net213),
    .Y(net3704));
 BUFx2_ASAP7_75t_R hold3300 (.A(_00989_),
    .Y(net3705));
 BUFx2_ASAP7_75t_R hold3301 (.A(text_in[57]),
    .Y(net3706));
 BUFx2_ASAP7_75t_R hold3302 (.A(net211),
    .Y(net3707));
 BUFx2_ASAP7_75t_R hold3303 (.A(_00987_),
    .Y(net3708));
 BUFx2_ASAP7_75t_R hold3304 (.A(text_in[21]),
    .Y(net3709));
 BUFx2_ASAP7_75t_R hold3305 (.A(net172),
    .Y(net3710));
 BUFx2_ASAP7_75t_R hold3306 (.A(_00951_),
    .Y(net3711));
 BUFx2_ASAP7_75t_R hold3307 (.A(text_in[16]),
    .Y(net3712));
 BUFx2_ASAP7_75t_R hold3308 (.A(net166),
    .Y(net3713));
 BUFx2_ASAP7_75t_R hold3309 (.A(_00946_),
    .Y(net3714));
 BUFx2_ASAP7_75t_R hold3310 (.A(text_in[33]),
    .Y(net3715));
 BUFx2_ASAP7_75t_R hold3311 (.A(net185),
    .Y(net3716));
 BUFx2_ASAP7_75t_R hold3312 (.A(_00963_),
    .Y(net3717));
 BUFx2_ASAP7_75t_R hold3313 (.A(text_in[39]),
    .Y(net3718));
 BUFx2_ASAP7_75t_R hold3314 (.A(net191),
    .Y(net3719));
 BUFx2_ASAP7_75t_R hold3315 (.A(_00969_),
    .Y(net3720));
 BUFx2_ASAP7_75t_R hold3316 (.A(text_in[20]),
    .Y(net3721));
 BUFx2_ASAP7_75t_R hold3317 (.A(net171),
    .Y(net3722));
 BUFx2_ASAP7_75t_R hold3318 (.A(_00950_),
    .Y(net3723));
 BUFx2_ASAP7_75t_R hold3319 (.A(text_in[15]),
    .Y(net3724));
 BUFx2_ASAP7_75t_R hold3320 (.A(net165),
    .Y(net3725));
 BUFx2_ASAP7_75t_R hold3321 (.A(_00945_),
    .Y(net3726));
 BUFx2_ASAP7_75t_R hold3322 (.A(text_in[76]),
    .Y(net3727));
 BUFx2_ASAP7_75t_R hold3323 (.A(net232),
    .Y(net3728));
 BUFx2_ASAP7_75t_R hold3324 (.A(_01006_),
    .Y(net3729));
 BUFx2_ASAP7_75t_R hold3325 (.A(text_in[18]),
    .Y(net3730));
 BUFx2_ASAP7_75t_R hold3326 (.A(net168),
    .Y(net3731));
 BUFx2_ASAP7_75t_R hold3327 (.A(_00948_),
    .Y(net3732));
 BUFx2_ASAP7_75t_R hold3328 (.A(text_in[34]),
    .Y(net3733));
 BUFx2_ASAP7_75t_R hold3329 (.A(net186),
    .Y(net3734));
 BUFx2_ASAP7_75t_R hold3330 (.A(_00964_),
    .Y(net3735));
 BUFx2_ASAP7_75t_R hold3331 (.A(text_in[14]),
    .Y(net3736));
 BUFx2_ASAP7_75t_R hold3332 (.A(net164),
    .Y(net3737));
 BUFx2_ASAP7_75t_R hold3333 (.A(_00944_),
    .Y(net3738));
 BUFx2_ASAP7_75t_R hold3334 (.A(text_in[38]),
    .Y(net3739));
 BUFx2_ASAP7_75t_R hold3335 (.A(net190),
    .Y(net3740));
 BUFx2_ASAP7_75t_R hold3336 (.A(_00968_),
    .Y(net3741));
 BUFx2_ASAP7_75t_R hold3337 (.A(text_in[75]),
    .Y(net3742));
 BUFx2_ASAP7_75t_R hold3338 (.A(net231),
    .Y(net3743));
 BUFx2_ASAP7_75t_R hold3339 (.A(_01005_),
    .Y(net3744));
 BUFx2_ASAP7_75t_R hold3340 (.A(text_in[56]),
    .Y(net3745));
 BUFx2_ASAP7_75t_R hold3341 (.A(net210),
    .Y(net3746));
 BUFx2_ASAP7_75t_R hold3342 (.A(_00986_),
    .Y(net3747));
 BUFx2_ASAP7_75t_R hold3343 (.A(text_in[32]),
    .Y(net3748));
 BUFx2_ASAP7_75t_R hold3344 (.A(net184),
    .Y(net3749));
 BUFx2_ASAP7_75t_R hold3345 (.A(_00962_),
    .Y(net3750));
 BUFx2_ASAP7_75t_R hold3346 (.A(text_in[19]),
    .Y(net3751));
 BUFx2_ASAP7_75t_R hold3347 (.A(net169),
    .Y(net3752));
 BUFx2_ASAP7_75t_R hold3348 (.A(_00949_),
    .Y(net3753));
 BUFx2_ASAP7_75t_R hold3349 (.A(text_in[13]),
    .Y(net3754));
 BUFx2_ASAP7_75t_R hold3350 (.A(net163),
    .Y(net3755));
 BUFx2_ASAP7_75t_R hold3351 (.A(_00943_),
    .Y(net3756));
 BUFx2_ASAP7_75t_R hold3352 (.A(text_in[2]),
    .Y(net3757));
 BUFx2_ASAP7_75t_R hold3353 (.A(net181),
    .Y(net3758));
 BUFx2_ASAP7_75t_R hold3354 (.A(_00932_),
    .Y(net3759));
 BUFx2_ASAP7_75t_R hold3355 (.A(text_in[122]),
    .Y(net3760));
 BUFx2_ASAP7_75t_R hold3356 (.A(net156),
    .Y(net3761));
 BUFx2_ASAP7_75t_R hold3357 (.A(_01052_),
    .Y(net3762));
 BUFx2_ASAP7_75t_R hold3358 (.A(text_in[11]),
    .Y(net3763));
 BUFx2_ASAP7_75t_R hold3359 (.A(net153),
    .Y(net3764));
 BUFx2_ASAP7_75t_R hold3360 (.A(_00941_),
    .Y(net3765));
 BUFx2_ASAP7_75t_R hold3361 (.A(text_in[26]),
    .Y(net3766));
 BUFx2_ASAP7_75t_R hold3362 (.A(net177),
    .Y(net3767));
 BUFx2_ASAP7_75t_R hold3363 (.A(_00956_),
    .Y(net3768));
 BUFx2_ASAP7_75t_R hold3364 (.A(key[82]),
    .Y(net3769));
 BUFx2_ASAP7_75t_R hold3365 (.A(net109),
    .Y(net3770));
 BUFx2_ASAP7_75t_R hold3366 (.A(_17371_),
    .Y(net3771));
 BUFx2_ASAP7_75t_R hold3367 (.A(text_in[31]),
    .Y(net3772));
 BUFx2_ASAP7_75t_R hold3368 (.A(net183),
    .Y(net3773));
 BUFx2_ASAP7_75t_R hold3369 (.A(_00961_),
    .Y(net3774));
 BUFx2_ASAP7_75t_R hold3370 (.A(text_in[79]),
    .Y(net3775));
 BUFx2_ASAP7_75t_R hold3371 (.A(net235),
    .Y(net3776));
 BUFx2_ASAP7_75t_R hold3372 (.A(_01009_),
    .Y(net3777));
 BUFx2_ASAP7_75t_R hold3373 (.A(text_in[30]),
    .Y(net3778));
 BUFx2_ASAP7_75t_R hold3374 (.A(net182),
    .Y(net3779));
 BUFx2_ASAP7_75t_R hold3375 (.A(_00960_),
    .Y(net3780));
 BUFx2_ASAP7_75t_R hold3376 (.A(text_in[112]),
    .Y(net3781));
 BUFx2_ASAP7_75t_R hold3377 (.A(net145),
    .Y(net3782));
 BUFx2_ASAP7_75t_R hold3378 (.A(_01042_),
    .Y(net3783));
 BUFx2_ASAP7_75t_R hold3379 (.A(text_in[124]),
    .Y(net3784));
 BUFx2_ASAP7_75t_R hold3380 (.A(net158),
    .Y(net3785));
 BUFx2_ASAP7_75t_R hold3381 (.A(_01054_),
    .Y(net3786));
 BUFx2_ASAP7_75t_R hold3382 (.A(text_in[69]),
    .Y(net3787));
 BUFx2_ASAP7_75t_R hold3383 (.A(net224),
    .Y(net3788));
 BUFx2_ASAP7_75t_R hold3384 (.A(_00999_),
    .Y(net3789));
 BUFx2_ASAP7_75t_R hold3385 (.A(text_in[97]),
    .Y(net3790));
 BUFx2_ASAP7_75t_R hold3386 (.A(net255),
    .Y(net3791));
 BUFx2_ASAP7_75t_R hold3387 (.A(_01027_),
    .Y(net3792));
 BUFx2_ASAP7_75t_R hold3388 (.A(key[17]),
    .Y(net3793));
 BUFx2_ASAP7_75t_R hold3389 (.A(net37),
    .Y(net3794));
 BUFx2_ASAP7_75t_R hold3390 (.A(_15667_),
    .Y(net3795));
 BUFx2_ASAP7_75t_R hold3391 (.A(text_in[85]),
    .Y(net3796));
 BUFx2_ASAP7_75t_R hold3392 (.A(net242),
    .Y(net3797));
 BUFx2_ASAP7_75t_R hold3393 (.A(_01015_),
    .Y(net3798));
 BUFx2_ASAP7_75t_R hold3394 (.A(text_in[28]),
    .Y(net3799));
 BUFx2_ASAP7_75t_R hold3395 (.A(net179),
    .Y(net3800));
 BUFx2_ASAP7_75t_R hold3396 (.A(_00958_),
    .Y(net3801));
 BUFx2_ASAP7_75t_R hold3397 (.A(text_in[113]),
    .Y(net3802));
 BUFx2_ASAP7_75t_R hold3398 (.A(net146),
    .Y(net3803));
 BUFx2_ASAP7_75t_R hold3399 (.A(_01043_),
    .Y(net3804));
 BUFx2_ASAP7_75t_R hold3400 (.A(text_in[70]),
    .Y(net3805));
 BUFx2_ASAP7_75t_R hold3401 (.A(net226),
    .Y(net3806));
 BUFx2_ASAP7_75t_R hold3402 (.A(_01000_),
    .Y(net3807));
 BUFx2_ASAP7_75t_R hold3403 (.A(text_in[111]),
    .Y(net3808));
 BUFx2_ASAP7_75t_R hold3404 (.A(net144),
    .Y(net3809));
 BUFx2_ASAP7_75t_R hold3405 (.A(_01041_),
    .Y(net3810));
 BUFx2_ASAP7_75t_R hold3406 (.A(text_in[78]),
    .Y(net3811));
 BUFx2_ASAP7_75t_R hold3407 (.A(net234),
    .Y(net3812));
 BUFx2_ASAP7_75t_R hold3408 (.A(_01008_),
    .Y(net3813));
 BUFx2_ASAP7_75t_R hold3409 (.A(net3847),
    .Y(net3814));
 BUFx2_ASAP7_75t_R hold3410 (.A(net130),
    .Y(net3815));
 BUFx2_ASAP7_75t_R hold3411 (.A(_01059_),
    .Y(net3816));
 BUFx2_ASAP7_75t_R hold3412 (.A(text_in[96]),
    .Y(net3817));
 BUFx2_ASAP7_75t_R hold3413 (.A(net254),
    .Y(net3818));
 BUFx2_ASAP7_75t_R hold3414 (.A(_01026_),
    .Y(net3819));
 BUFx2_ASAP7_75t_R hold3415 (.A(text_in[123]),
    .Y(net3820));
 BUFx2_ASAP7_75t_R hold3416 (.A(net157),
    .Y(net3821));
 BUFx2_ASAP7_75t_R hold3417 (.A(_01053_),
    .Y(net3822));
 BUFx2_ASAP7_75t_R hold3418 (.A(text_in[127]),
    .Y(net3823));
 BUFx2_ASAP7_75t_R hold3419 (.A(net161),
    .Y(net3824));
 BUFx2_ASAP7_75t_R hold3420 (.A(_01057_),
    .Y(net3825));
 BUFx2_ASAP7_75t_R hold3421 (.A(text_in[82]),
    .Y(net3826));
 BUFx2_ASAP7_75t_R hold3422 (.A(net239),
    .Y(net3827));
 BUFx2_ASAP7_75t_R hold3423 (.A(_01012_),
    .Y(net3828));
 BUFx2_ASAP7_75t_R hold3424 (.A(text_in[126]),
    .Y(net3829));
 BUFx2_ASAP7_75t_R hold3425 (.A(net160),
    .Y(net3830));
 BUFx2_ASAP7_75t_R hold3426 (.A(_01056_),
    .Y(net3831));
 BUFx2_ASAP7_75t_R hold3427 (.A(text_in[105]),
    .Y(net3832));
 BUFx2_ASAP7_75t_R hold3428 (.A(net137),
    .Y(net3833));
 BUFx2_ASAP7_75t_R hold3429 (.A(_01035_),
    .Y(net3834));
 BUFx2_ASAP7_75t_R hold3430 (.A(text_in[68]),
    .Y(net3835));
 BUFx2_ASAP7_75t_R hold3431 (.A(net223),
    .Y(net3836));
 BUFx2_ASAP7_75t_R hold3432 (.A(_00998_),
    .Y(net3837));
 BUFx2_ASAP7_75t_R hold3433 (.A(ld),
    .Y(net3838));
 BUFx2_ASAP7_75t_R hold3434 (.A(net129),
    .Y(net3839));
 BUFx2_ASAP7_75t_R hold3435 (.A(_01058_),
    .Y(net3840));
 BUFx2_ASAP7_75t_R hold3436 (.A(text_in[87]),
    .Y(net3841));
 BUFx2_ASAP7_75t_R hold3437 (.A(net244),
    .Y(net3842));
 BUFx2_ASAP7_75t_R hold3438 (.A(_01017_),
    .Y(net3843));
 BUFx2_ASAP7_75t_R hold3439 (.A(text_in[73]),
    .Y(net3844));
 BUFx2_ASAP7_75t_R hold3440 (.A(net229),
    .Y(net3845));
 BUFx2_ASAP7_75t_R hold3441 (.A(_01003_),
    .Y(net3846));
 BUFx2_ASAP7_75t_R hold3442 (.A(rst),
    .Y(net3847));
 BUFx2_ASAP7_75t_R hold3443 (.A(text_in[67]),
    .Y(net3848));
 BUFx2_ASAP7_75t_R hold3444 (.A(net222),
    .Y(net3849));
 BUFx2_ASAP7_75t_R hold3445 (.A(_00997_),
    .Y(net3850));
 BUFx2_ASAP7_75t_R hold3446 (.A(text_in[121]),
    .Y(net3851));
 BUFx2_ASAP7_75t_R hold3447 (.A(net155),
    .Y(net3852));
 BUFx2_ASAP7_75t_R hold3448 (.A(_01051_),
    .Y(net3853));
 BUFx2_ASAP7_75t_R hold3449 (.A(key[90]),
    .Y(net3854));
 BUFx2_ASAP7_75t_R hold3450 (.A(net118),
    .Y(net3855));
 BUFx2_ASAP7_75t_R hold3451 (.A(_17397_),
    .Y(net3856));
 BUFx2_ASAP7_75t_R hold3452 (.A(text_in[94]),
    .Y(net3857));
 BUFx2_ASAP7_75t_R hold3453 (.A(net252),
    .Y(net3858));
 BUFx2_ASAP7_75t_R hold3454 (.A(_01024_),
    .Y(net3859));
 BUFx2_ASAP7_75t_R hold3455 (.A(key[58]),
    .Y(net3860));
 BUFx2_ASAP7_75t_R hold3456 (.A(net82),
    .Y(net3861));
 BUFx2_ASAP7_75t_R hold3457 (.A(_17273_),
    .Y(net3862));
 BUFx2_ASAP7_75t_R hold3458 (.A(key[26]),
    .Y(net3863));
 BUFx2_ASAP7_75t_R hold3459 (.A(net47),
    .Y(net3864));
 BUFx2_ASAP7_75t_R hold3460 (.A(_00371_),
    .Y(net3865));
 BUFx2_ASAP7_75t_R hold3461 (.A(text_in[1]),
    .Y(net3866));
 BUFx2_ASAP7_75t_R hold3462 (.A(net170),
    .Y(net3867));
 BUFx2_ASAP7_75t_R hold3463 (.A(_00931_),
    .Y(net3868));
 BUFx2_ASAP7_75t_R hold3464 (.A(text_in[24]),
    .Y(net3869));
 BUFx2_ASAP7_75t_R hold3465 (.A(net175),
    .Y(net3870));
 BUFx2_ASAP7_75t_R hold3466 (.A(_00954_),
    .Y(net3871));
 BUFx2_ASAP7_75t_R hold3467 (.A(key[20]),
    .Y(net3872));
 BUFx2_ASAP7_75t_R hold3468 (.A(net41),
    .Y(net3873));
 BUFx2_ASAP7_75t_R hold3469 (.A(_16055_),
    .Y(net3874));
 BUFx2_ASAP7_75t_R hold3470 (.A(net4210),
    .Y(net3875));
 BUFx2_ASAP7_75t_R hold3471 (.A(net26),
    .Y(net3876));
 BUFx2_ASAP7_75t_R hold3472 (.A(text_in[86]),
    .Y(net3877));
 BUFx2_ASAP7_75t_R hold3473 (.A(net243),
    .Y(net3878));
 BUFx2_ASAP7_75t_R hold3474 (.A(_01016_),
    .Y(net3879));
 BUFx2_ASAP7_75t_R hold3475 (.A(key[29]),
    .Y(net3880));
 BUFx2_ASAP7_75t_R hold3476 (.A(net50),
    .Y(net3881));
 BUFx2_ASAP7_75t_R hold3477 (.A(_16992_),
    .Y(net3882));
 BUFx2_ASAP7_75t_R hold3478 (.A(text_in[109]),
    .Y(net3883));
 BUFx2_ASAP7_75t_R hold3479 (.A(net141),
    .Y(net3884));
 BUFx2_ASAP7_75t_R hold3480 (.A(_01039_),
    .Y(net3885));
 BUFx2_ASAP7_75t_R hold3481 (.A(text_in[120]),
    .Y(net3886));
 BUFx2_ASAP7_75t_R hold3482 (.A(net154),
    .Y(net3887));
 BUFx2_ASAP7_75t_R hold3483 (.A(_01050_),
    .Y(net3888));
 BUFx2_ASAP7_75t_R hold3484 (.A(key[44]),
    .Y(net3889));
 BUFx2_ASAP7_75t_R hold3485 (.A(net67),
    .Y(net3890));
 BUFx2_ASAP7_75t_R hold3486 (.A(_17198_),
    .Y(net3891));
 BUFx2_ASAP7_75t_R hold3487 (.A(key[112]),
    .Y(net3892));
 BUFx2_ASAP7_75t_R hold3488 (.A(net15),
    .Y(net3893));
 BUFx2_ASAP7_75t_R hold3489 (.A(_17477_),
    .Y(net3894));
 BUFx2_ASAP7_75t_R hold3490 (.A(text_in[104]),
    .Y(net3895));
 BUFx2_ASAP7_75t_R hold3491 (.A(net136),
    .Y(net3896));
 BUFx2_ASAP7_75t_R hold3492 (.A(_01034_),
    .Y(net3897));
 BUFx2_ASAP7_75t_R hold3493 (.A(text_in[71]),
    .Y(net3898));
 BUFx2_ASAP7_75t_R hold3494 (.A(net227),
    .Y(net3899));
 BUFx2_ASAP7_75t_R hold3495 (.A(_01001_),
    .Y(net3900));
 BUFx2_ASAP7_75t_R hold3496 (.A(text_in[46]),
    .Y(net3901));
 BUFx2_ASAP7_75t_R hold3497 (.A(net199),
    .Y(net3902));
 BUFx2_ASAP7_75t_R hold3498 (.A(_00976_),
    .Y(net3903));
 BUFx2_ASAP7_75t_R hold3499 (.A(text_in[91]),
    .Y(net3904));
 BUFx2_ASAP7_75t_R hold3500 (.A(net249),
    .Y(net3905));
 BUFx2_ASAP7_75t_R hold3501 (.A(_01021_),
    .Y(net3906));
 BUFx2_ASAP7_75t_R hold3502 (.A(net4211),
    .Y(net3907));
 BUFx2_ASAP7_75t_R hold3503 (.A(net28),
    .Y(net3908));
 BUFx2_ASAP7_75t_R hold3504 (.A(text_in[125]),
    .Y(net3909));
 BUFx2_ASAP7_75t_R hold3505 (.A(net159),
    .Y(net3910));
 BUFx2_ASAP7_75t_R hold3506 (.A(_01055_),
    .Y(net3911));
 BUFx2_ASAP7_75t_R hold3507 (.A(text_in[74]),
    .Y(net3912));
 BUFx2_ASAP7_75t_R hold3508 (.A(net230),
    .Y(net3913));
 BUFx2_ASAP7_75t_R hold3509 (.A(_01004_),
    .Y(net3914));
 BUFx2_ASAP7_75t_R hold3510 (.A(key[113]),
    .Y(net3915));
 BUFx2_ASAP7_75t_R hold3511 (.A(net16),
    .Y(net3916));
 BUFx2_ASAP7_75t_R hold3512 (.A(_17480_),
    .Y(net3917));
 BUFx2_ASAP7_75t_R hold3513 (.A(text_in[99]),
    .Y(net3918));
 BUFx2_ASAP7_75t_R hold3514 (.A(net257),
    .Y(net3919));
 BUFx2_ASAP7_75t_R hold3515 (.A(_01029_),
    .Y(net3920));
 BUFx2_ASAP7_75t_R hold3516 (.A(text_in[106]),
    .Y(net3921));
 BUFx2_ASAP7_75t_R hold3517 (.A(net138),
    .Y(net3922));
 BUFx2_ASAP7_75t_R hold3518 (.A(_01036_),
    .Y(net3923));
 BUFx2_ASAP7_75t_R hold3519 (.A(text_in[102]),
    .Y(net3924));
 BUFx2_ASAP7_75t_R hold3520 (.A(net134),
    .Y(net3925));
 BUFx2_ASAP7_75t_R hold3521 (.A(_01032_),
    .Y(net3926));
 BUFx2_ASAP7_75t_R hold3522 (.A(text_in[27]),
    .Y(net3927));
 BUFx2_ASAP7_75t_R hold3523 (.A(net178),
    .Y(net3928));
 BUFx2_ASAP7_75t_R hold3524 (.A(_00957_),
    .Y(net3929));
 BUFx2_ASAP7_75t_R hold3525 (.A(text_in[114]),
    .Y(net3930));
 BUFx2_ASAP7_75t_R hold3526 (.A(net147),
    .Y(net3931));
 BUFx2_ASAP7_75t_R hold3527 (.A(_01044_),
    .Y(net3932));
 BUFx2_ASAP7_75t_R hold3528 (.A(text_in[29]),
    .Y(net3933));
 BUFx2_ASAP7_75t_R hold3529 (.A(net180),
    .Y(net3934));
 BUFx2_ASAP7_75t_R hold3530 (.A(_00959_),
    .Y(net3935));
 BUFx2_ASAP7_75t_R hold3531 (.A(text_in[108]),
    .Y(net3936));
 BUFx2_ASAP7_75t_R hold3532 (.A(net140),
    .Y(net3937));
 BUFx2_ASAP7_75t_R hold3533 (.A(_01038_),
    .Y(net3938));
 BUFx2_ASAP7_75t_R hold3534 (.A(key[51]),
    .Y(net3939));
 BUFx2_ASAP7_75t_R hold3535 (.A(net75),
    .Y(net3940));
 BUFx2_ASAP7_75t_R hold3536 (.A(_00331_),
    .Y(net3941));
 BUFx2_ASAP7_75t_R hold3537 (.A(text_in[52]),
    .Y(net3942));
 BUFx2_ASAP7_75t_R hold3538 (.A(net206),
    .Y(net3943));
 BUFx2_ASAP7_75t_R hold3539 (.A(_00982_),
    .Y(net3944));
 BUFx2_ASAP7_75t_R hold3540 (.A(text_in[115]),
    .Y(net3945));
 BUFx2_ASAP7_75t_R hold3541 (.A(net148),
    .Y(net3946));
 BUFx2_ASAP7_75t_R hold3542 (.A(_01045_),
    .Y(net3947));
 BUFx2_ASAP7_75t_R hold3543 (.A(text_in[98]),
    .Y(net3948));
 BUFx2_ASAP7_75t_R hold3544 (.A(net256),
    .Y(net3949));
 BUFx2_ASAP7_75t_R hold3545 (.A(_01028_),
    .Y(net3950));
 BUFx2_ASAP7_75t_R hold3546 (.A(text_in[25]),
    .Y(net3951));
 BUFx2_ASAP7_75t_R hold3547 (.A(net176),
    .Y(net3952));
 BUFx2_ASAP7_75t_R hold3548 (.A(_00955_),
    .Y(net3953));
 BUFx2_ASAP7_75t_R hold3549 (.A(text_in[61]),
    .Y(net3954));
 BUFx2_ASAP7_75t_R hold3550 (.A(net216),
    .Y(net3955));
 BUFx2_ASAP7_75t_R hold3551 (.A(_00991_),
    .Y(net3956));
 BUFx2_ASAP7_75t_R hold3552 (.A(text_in[100]),
    .Y(net3957));
 BUFx2_ASAP7_75t_R hold3553 (.A(net132),
    .Y(net3958));
 BUFx2_ASAP7_75t_R hold3554 (.A(_01030_),
    .Y(net3959));
 BUFx2_ASAP7_75t_R hold3555 (.A(text_in[101]),
    .Y(net3960));
 BUFx2_ASAP7_75t_R hold3556 (.A(net133),
    .Y(net3961));
 BUFx2_ASAP7_75t_R hold3557 (.A(_01031_),
    .Y(net3962));
 BUFx2_ASAP7_75t_R hold3558 (.A(text_in[0]),
    .Y(net3963));
 BUFx2_ASAP7_75t_R hold3559 (.A(net131),
    .Y(net3964));
 BUFx2_ASAP7_75t_R hold3560 (.A(_00930_),
    .Y(net3965));
 BUFx2_ASAP7_75t_R hold3561 (.A(key[16]),
    .Y(net3966));
 BUFx2_ASAP7_75t_R hold3562 (.A(net36),
    .Y(net3967));
 BUFx2_ASAP7_75t_R hold3563 (.A(_15396_),
    .Y(net3968));
 BUFx2_ASAP7_75t_R hold3564 (.A(key[22]),
    .Y(net3969));
 BUFx2_ASAP7_75t_R hold3565 (.A(net43),
    .Y(net3970));
 BUFx2_ASAP7_75t_R hold3566 (.A(_16127_),
    .Y(net3971));
 BUFx2_ASAP7_75t_R hold3567 (.A(text_in[117]),
    .Y(net3972));
 BUFx2_ASAP7_75t_R hold3568 (.A(net150),
    .Y(net3973));
 BUFx2_ASAP7_75t_R hold3569 (.A(_01047_),
    .Y(net3974));
 BUFx2_ASAP7_75t_R hold3570 (.A(text_in[36]),
    .Y(net3975));
 BUFx2_ASAP7_75t_R hold3571 (.A(net188),
    .Y(net3976));
 BUFx2_ASAP7_75t_R hold3572 (.A(_00966_),
    .Y(net3977));
 BUFx2_ASAP7_75t_R hold3573 (.A(text_in[119]),
    .Y(net3978));
 BUFx2_ASAP7_75t_R hold3574 (.A(net152),
    .Y(net3979));
 BUFx2_ASAP7_75t_R hold3575 (.A(_01049_),
    .Y(net3980));
 BUFx2_ASAP7_75t_R hold3576 (.A(key[47]),
    .Y(net3981));
 BUFx2_ASAP7_75t_R hold3577 (.A(net70),
    .Y(net3982));
 BUFx2_ASAP7_75t_R hold3578 (.A(_17219_),
    .Y(net3983));
 BUFx2_ASAP7_75t_R hold3579 (.A(text_in[110]),
    .Y(net3984));
 BUFx2_ASAP7_75t_R hold3580 (.A(net143),
    .Y(net3985));
 BUFx2_ASAP7_75t_R hold3581 (.A(_01040_),
    .Y(net3986));
 BUFx2_ASAP7_75t_R hold3582 (.A(text_in[103]),
    .Y(net3987));
 BUFx2_ASAP7_75t_R hold3583 (.A(net135),
    .Y(net3988));
 BUFx2_ASAP7_75t_R hold3584 (.A(_01033_),
    .Y(net3989));
 BUFx2_ASAP7_75t_R hold3585 (.A(net4221),
    .Y(net3990));
 BUFx2_ASAP7_75t_R hold3586 (.A(net27),
    .Y(net3991));
 BUFx2_ASAP7_75t_R hold3587 (.A(text_in[3]),
    .Y(net3992));
 BUFx2_ASAP7_75t_R hold3588 (.A(net192),
    .Y(net3993));
 BUFx2_ASAP7_75t_R hold3589 (.A(_00933_),
    .Y(net3994));
 BUFx2_ASAP7_75t_R hold3590 (.A(text_in[116]),
    .Y(net3995));
 BUFx2_ASAP7_75t_R hold3591 (.A(net149),
    .Y(net3996));
 BUFx2_ASAP7_75t_R hold3592 (.A(_01046_),
    .Y(net3997));
 BUFx2_ASAP7_75t_R hold3593 (.A(key[43]),
    .Y(net3998));
 BUFx2_ASAP7_75t_R hold3594 (.A(net66),
    .Y(net3999));
 BUFx2_ASAP7_75t_R hold3595 (.A(_17193_),
    .Y(net4000));
 BUFx2_ASAP7_75t_R hold3596 (.A(text_in[47]),
    .Y(net4001));
 BUFx2_ASAP7_75t_R hold3597 (.A(net200),
    .Y(net4002));
 BUFx2_ASAP7_75t_R hold3598 (.A(_00977_),
    .Y(net4003));
 BUFx2_ASAP7_75t_R hold3599 (.A(key[109]),
    .Y(net4004));
 BUFx2_ASAP7_75t_R hold3600 (.A(net11),
    .Y(net4005));
 BUFx2_ASAP7_75t_R hold3601 (.A(_17468_),
    .Y(net4006));
 BUFx2_ASAP7_75t_R hold3602 (.A(key[74]),
    .Y(net4007));
 BUFx2_ASAP7_75t_R hold3603 (.A(net100),
    .Y(net4008));
 BUFx2_ASAP7_75t_R hold3604 (.A(_17347_),
    .Y(net4009));
 BUFx2_ASAP7_75t_R hold3605 (.A(key[97]),
    .Y(net4010));
 BUFx2_ASAP7_75t_R hold3606 (.A(net125),
    .Y(net4011));
 BUFx2_ASAP7_75t_R hold3607 (.A(_17437_),
    .Y(net4012));
 BUFx2_ASAP7_75t_R hold3608 (.A(key[96]),
    .Y(net4013));
 BUFx2_ASAP7_75t_R hold3609 (.A(net124),
    .Y(net4014));
 BUFx2_ASAP7_75t_R hold3610 (.A(_17434_),
    .Y(net4015));
 BUFx2_ASAP7_75t_R hold3611 (.A(key[1]),
    .Y(net4016));
 BUFx2_ASAP7_75t_R hold3612 (.A(net40),
    .Y(net4017));
 BUFx2_ASAP7_75t_R hold3613 (.A(key[48]),
    .Y(net4018));
 BUFx2_ASAP7_75t_R hold3614 (.A(net71),
    .Y(net4019));
 BUFx2_ASAP7_75t_R hold3615 (.A(_17229_),
    .Y(net4020));
 BUFx2_ASAP7_75t_R hold3616 (.A(key[127]),
    .Y(net4021));
 BUFx2_ASAP7_75t_R hold3617 (.A(net31),
    .Y(net4022));
 BUFx2_ASAP7_75t_R hold3618 (.A(key[80]),
    .Y(net4023));
 BUFx2_ASAP7_75t_R hold3619 (.A(net107),
    .Y(net4024));
 BUFx2_ASAP7_75t_R hold3620 (.A(_17365_),
    .Y(net4025));
 BUFx2_ASAP7_75t_R hold3621 (.A(text_in[5]),
    .Y(net4026));
 BUFx2_ASAP7_75t_R hold3622 (.A(net214),
    .Y(net4027));
 BUFx2_ASAP7_75t_R hold3623 (.A(text_in[37]),
    .Y(net4028));
 BUFx2_ASAP7_75t_R hold3624 (.A(net189),
    .Y(net4029));
 BUFx2_ASAP7_75t_R hold3625 (.A(key[81]),
    .Y(net4030));
 BUFx2_ASAP7_75t_R hold3626 (.A(net108),
    .Y(net4031));
 BUFx2_ASAP7_75t_R hold3627 (.A(_17367_),
    .Y(net4032));
 BUFx2_ASAP7_75t_R hold3628 (.A(key[95]),
    .Y(net4033));
 BUFx2_ASAP7_75t_R hold3629 (.A(net123),
    .Y(net4034));
 BUFx2_ASAP7_75t_R hold3630 (.A(key[13]),
    .Y(net4035));
 BUFx2_ASAP7_75t_R hold3631 (.A(net33),
    .Y(net4036));
 BUFx2_ASAP7_75t_R hold3632 (.A(key[49]),
    .Y(net4037));
 BUFx2_ASAP7_75t_R hold3633 (.A(net72),
    .Y(net4038));
 BUFx2_ASAP7_75t_R hold3634 (.A(key[84]),
    .Y(net4039));
 BUFx2_ASAP7_75t_R hold3635 (.A(net111),
    .Y(net4040));
 BUFx2_ASAP7_75t_R hold3636 (.A(key[40]),
    .Y(net4041));
 BUFx2_ASAP7_75t_R hold3637 (.A(net63),
    .Y(net4042));
 BUFx2_ASAP7_75t_R hold3638 (.A(key[5]),
    .Y(net4043));
 BUFx2_ASAP7_75t_R hold3639 (.A(net84),
    .Y(net4044));
 BUFx2_ASAP7_75t_R hold3640 (.A(key[56]),
    .Y(net4045));
 BUFx2_ASAP7_75t_R hold3641 (.A(net80),
    .Y(net4046));
 BUFx2_ASAP7_75t_R hold3642 (.A(key[121]),
    .Y(net4047));
 BUFx2_ASAP7_75t_R hold3643 (.A(net25),
    .Y(net4048));
 BUFx2_ASAP7_75t_R hold3644 (.A(key[46]),
    .Y(net4049));
 BUFx2_ASAP7_75t_R hold3645 (.A(net69),
    .Y(net4050));
 BUFx2_ASAP7_75t_R hold3646 (.A(key[12]),
    .Y(net4051));
 BUFx2_ASAP7_75t_R hold3647 (.A(net32),
    .Y(net4052));
 BUFx2_ASAP7_75t_R hold3648 (.A(key[89]),
    .Y(net4053));
 BUFx2_ASAP7_75t_R hold3649 (.A(net116),
    .Y(net4054));
 BUFx2_ASAP7_75t_R hold3650 (.A(key[6]),
    .Y(net4055));
 BUFx2_ASAP7_75t_R hold3651 (.A(net95),
    .Y(net4056));
 BUFx2_ASAP7_75t_R hold3652 (.A(key[41]),
    .Y(net4057));
 BUFx2_ASAP7_75t_R hold3653 (.A(net64),
    .Y(net4058));
 BUFx2_ASAP7_75t_R hold3654 (.A(key[52]),
    .Y(net4059));
 BUFx2_ASAP7_75t_R hold3655 (.A(net76),
    .Y(net4060));
 BUFx2_ASAP7_75t_R hold3656 (.A(key[115]),
    .Y(net4061));
 BUFx2_ASAP7_75t_R hold3657 (.A(net18),
    .Y(net4062));
 BUFx2_ASAP7_75t_R hold3658 (.A(key[45]),
    .Y(net4063));
 BUFx2_ASAP7_75t_R hold3659 (.A(net68),
    .Y(net4064));
 BUFx2_ASAP7_75t_R hold3660 (.A(key[34]),
    .Y(net4065));
 BUFx2_ASAP7_75t_R hold3661 (.A(net56),
    .Y(net4066));
 BUFx2_ASAP7_75t_R hold3662 (.A(key[77]),
    .Y(net4067));
 BUFx2_ASAP7_75t_R hold3663 (.A(net103),
    .Y(net4068));
 BUFx2_ASAP7_75t_R hold3664 (.A(key[83]),
    .Y(net4069));
 BUFx2_ASAP7_75t_R hold3665 (.A(net110),
    .Y(net4070));
 BUFx2_ASAP7_75t_R hold3666 (.A(key[57]),
    .Y(net4071));
 BUFx2_ASAP7_75t_R hold3667 (.A(net81),
    .Y(net4072));
 BUFx2_ASAP7_75t_R hold3668 (.A(key[8]),
    .Y(net4073));
 BUFx2_ASAP7_75t_R hold3669 (.A(net117),
    .Y(net4074));
 BUFx2_ASAP7_75t_R hold3670 (.A(key[101]),
    .Y(net4075));
 BUFx2_ASAP7_75t_R hold3671 (.A(net3),
    .Y(net4076));
 BUFx2_ASAP7_75t_R hold3672 (.A(key[65]),
    .Y(net4077));
 BUFx2_ASAP7_75t_R hold3673 (.A(net90),
    .Y(net4078));
 BUFx2_ASAP7_75t_R hold3674 (.A(key[91]),
    .Y(net4079));
 BUFx2_ASAP7_75t_R hold3675 (.A(net119),
    .Y(net4080));
 BUFx2_ASAP7_75t_R hold3676 (.A(key[53]),
    .Y(net4081));
 BUFx2_ASAP7_75t_R hold3677 (.A(net77),
    .Y(net4082));
 BUFx2_ASAP7_75t_R hold3678 (.A(key[35]),
    .Y(net4083));
 BUFx2_ASAP7_75t_R hold3679 (.A(net57),
    .Y(net4084));
 BUFx2_ASAP7_75t_R hold3680 (.A(key[92]),
    .Y(net4085));
 BUFx2_ASAP7_75t_R hold3681 (.A(net120),
    .Y(net4086));
 BUFx2_ASAP7_75t_R hold3682 (.A(key[60]),
    .Y(net4087));
 BUFx2_ASAP7_75t_R hold3683 (.A(net85),
    .Y(net4088));
 BUFx2_ASAP7_75t_R hold3684 (.A(key[59]),
    .Y(net4089));
 BUFx2_ASAP7_75t_R hold3685 (.A(net83),
    .Y(net4090));
 BUFx2_ASAP7_75t_R hold3686 (.A(key[36]),
    .Y(net4091));
 BUFx2_ASAP7_75t_R hold3687 (.A(net58),
    .Y(net4092));
 BUFx2_ASAP7_75t_R hold3688 (.A(text_in[118]),
    .Y(net4093));
 BUFx2_ASAP7_75t_R hold3689 (.A(net151),
    .Y(net4094));
 BUFx2_ASAP7_75t_R hold3690 (.A(key[64]),
    .Y(net4095));
 BUFx2_ASAP7_75t_R hold3691 (.A(net89),
    .Y(net4096));
 BUFx2_ASAP7_75t_R hold3692 (.A(key[72]),
    .Y(net4097));
 BUFx2_ASAP7_75t_R hold3693 (.A(net98),
    .Y(net4098));
 BUFx2_ASAP7_75t_R hold3694 (.A(key[42]),
    .Y(net4099));
 BUFx2_ASAP7_75t_R hold3695 (.A(net65),
    .Y(net4100));
 BUFx2_ASAP7_75t_R hold3696 (.A(key[33]),
    .Y(net4101));
 BUFx2_ASAP7_75t_R hold3697 (.A(net55),
    .Y(net4102));
 BUFx2_ASAP7_75t_R hold3698 (.A(key[32]),
    .Y(net4103));
 BUFx2_ASAP7_75t_R hold3699 (.A(net54),
    .Y(net4104));
 BUFx2_ASAP7_75t_R hold3700 (.A(key[75]),
    .Y(net4105));
 BUFx2_ASAP7_75t_R hold3701 (.A(net101),
    .Y(net4106));
 BUFx2_ASAP7_75t_R hold3702 (.A(key[107]),
    .Y(net4107));
 BUFx2_ASAP7_75t_R hold3703 (.A(net9),
    .Y(net4108));
 BUFx2_ASAP7_75t_R hold3704 (.A(key[37]),
    .Y(net4109));
 BUFx2_ASAP7_75t_R hold3705 (.A(net59),
    .Y(net4110));
 BUFx2_ASAP7_75t_R hold3706 (.A(key[55]),
    .Y(net4111));
 BUFx2_ASAP7_75t_R hold3707 (.A(net79),
    .Y(net4112));
 BUFx2_ASAP7_75t_R hold3708 (.A(key[87]),
    .Y(net4113));
 BUFx2_ASAP7_75t_R hold3709 (.A(net114),
    .Y(net4114));
 BUFx2_ASAP7_75t_R hold3710 (.A(key[39]),
    .Y(net4115));
 BUFx2_ASAP7_75t_R hold3711 (.A(net61),
    .Y(net4116));
 BUFx2_ASAP7_75t_R hold3712 (.A(key[119]),
    .Y(net4117));
 BUFx2_ASAP7_75t_R hold3713 (.A(net22),
    .Y(net4118));
 BUFx2_ASAP7_75t_R hold3714 (.A(key[11]),
    .Y(net4119));
 BUFx2_ASAP7_75t_R hold3715 (.A(net23),
    .Y(net4120));
 BUFx2_ASAP7_75t_R hold3716 (.A(key[23]),
    .Y(net4121));
 BUFx2_ASAP7_75t_R hold3717 (.A(net44),
    .Y(net4122));
 BUFx2_ASAP7_75t_R hold3718 (.A(key[63]),
    .Y(net4123));
 BUFx2_ASAP7_75t_R hold3719 (.A(net88),
    .Y(net4124));
 BUFx2_ASAP7_75t_R hold3720 (.A(key[76]),
    .Y(net4125));
 BUFx2_ASAP7_75t_R hold3721 (.A(net102),
    .Y(net4126));
 BUFx2_ASAP7_75t_R hold3722 (.A(key[79]),
    .Y(net4127));
 BUFx2_ASAP7_75t_R hold3723 (.A(net105),
    .Y(net4128));
 BUFx2_ASAP7_75t_R hold3724 (.A(key[3]),
    .Y(net4129));
 BUFx2_ASAP7_75t_R hold3725 (.A(net62),
    .Y(net4130));
 BUFx2_ASAP7_75t_R hold3726 (.A(key[66]),
    .Y(net4131));
 BUFx2_ASAP7_75t_R hold3727 (.A(net91),
    .Y(net4132));
 BUFx2_ASAP7_75t_R hold3728 (.A(key[88]),
    .Y(net4133));
 BUFx2_ASAP7_75t_R hold3729 (.A(net115),
    .Y(net4134));
 BUFx2_ASAP7_75t_R hold3730 (.A(key[98]),
    .Y(net4135));
 BUFx2_ASAP7_75t_R hold3731 (.A(net126),
    .Y(net4136));
 BUFx2_ASAP7_75t_R hold3732 (.A(key[67]),
    .Y(net4137));
 BUFx2_ASAP7_75t_R hold3733 (.A(net92),
    .Y(net4138));
 BUFx2_ASAP7_75t_R hold3734 (.A(key[117]),
    .Y(net4139));
 BUFx2_ASAP7_75t_R hold3735 (.A(net20),
    .Y(net4140));
 BUFx2_ASAP7_75t_R hold3736 (.A(key[24]),
    .Y(net4141));
 BUFx2_ASAP7_75t_R hold3737 (.A(net45),
    .Y(net4142));
 BUFx2_ASAP7_75t_R hold3738 (.A(key[18]),
    .Y(net4143));
 BUFx2_ASAP7_75t_R hold3739 (.A(net38),
    .Y(net4144));
 BUFx2_ASAP7_75t_R hold3740 (.A(key[126]),
    .Y(net4145));
 BUFx2_ASAP7_75t_R hold3741 (.A(net30),
    .Y(net4146));
 BUFx2_ASAP7_75t_R hold3742 (.A(key[85]),
    .Y(net4147));
 BUFx2_ASAP7_75t_R hold3743 (.A(net112),
    .Y(net4148));
 BUFx2_ASAP7_75t_R hold3744 (.A(key[61]),
    .Y(net4149));
 BUFx2_ASAP7_75t_R hold3745 (.A(net86),
    .Y(net4150));
 BUFx2_ASAP7_75t_R hold3746 (.A(key[30]),
    .Y(net4151));
 BUFx2_ASAP7_75t_R hold3747 (.A(net52),
    .Y(net4152));
 BUFx2_ASAP7_75t_R hold3748 (.A(key[19]),
    .Y(net4153));
 BUFx2_ASAP7_75t_R hold3749 (.A(net39),
    .Y(net4154));
 BUFx2_ASAP7_75t_R hold3750 (.A(key[15]),
    .Y(net4155));
 BUFx2_ASAP7_75t_R hold3751 (.A(net35),
    .Y(net4156));
 BUFx2_ASAP7_75t_R hold3752 (.A(key[110]),
    .Y(net4157));
 BUFx2_ASAP7_75t_R hold3753 (.A(net13),
    .Y(net4158));
 BUFx2_ASAP7_75t_R hold3754 (.A(key[25]),
    .Y(net4159));
 BUFx2_ASAP7_75t_R hold3755 (.A(net46),
    .Y(net4160));
 BUFx2_ASAP7_75t_R hold3756 (.A(key[93]),
    .Y(net4161));
 BUFx2_ASAP7_75t_R hold3757 (.A(net121),
    .Y(net4162));
 BUFx2_ASAP7_75t_R hold3758 (.A(key[2]),
    .Y(net4163));
 BUFx2_ASAP7_75t_R hold3759 (.A(net51),
    .Y(net4164));
 BUFx2_ASAP7_75t_R hold3760 (.A(key[125]),
    .Y(net4165));
 BUFx2_ASAP7_75t_R hold3761 (.A(net29),
    .Y(net4166));
 BUFx2_ASAP7_75t_R hold3762 (.A(key[78]),
    .Y(net4167));
 BUFx2_ASAP7_75t_R hold3763 (.A(net104),
    .Y(net4168));
 BUFx2_ASAP7_75t_R hold3764 (.A(key[14]),
    .Y(net4169));
 BUFx2_ASAP7_75t_R hold3765 (.A(net34),
    .Y(net4170));
 BUFx2_ASAP7_75t_R hold3766 (.A(key[105]),
    .Y(net4171));
 BUFx2_ASAP7_75t_R hold3767 (.A(net7),
    .Y(net4172));
 BUFx2_ASAP7_75t_R hold3768 (.A(key[116]),
    .Y(net4173));
 BUFx2_ASAP7_75t_R hold3769 (.A(net19),
    .Y(net4174));
 BUFx2_ASAP7_75t_R hold3770 (.A(key[108]),
    .Y(net4175));
 BUFx2_ASAP7_75t_R hold3771 (.A(net10),
    .Y(net4176));
 BUFx2_ASAP7_75t_R hold3772 (.A(key[86]),
    .Y(net4177));
 BUFx2_ASAP7_75t_R hold3773 (.A(net113),
    .Y(net4178));
 BUFx2_ASAP7_75t_R hold3774 (.A(key[120]),
    .Y(net4179));
 BUFx2_ASAP7_75t_R hold3775 (.A(net24),
    .Y(net4180));
 BUFx2_ASAP7_75t_R hold3776 (.A(key[111]),
    .Y(net4181));
 BUFx2_ASAP7_75t_R hold3777 (.A(net14),
    .Y(net4182));
 BUFx2_ASAP7_75t_R hold3778 (.A(key[62]),
    .Y(net4183));
 BUFx2_ASAP7_75t_R hold3779 (.A(key[94]),
    .Y(net4184));
 BUFx2_ASAP7_75t_R hold3780 (.A(key[27]),
    .Y(net4185));
 BUFx2_ASAP7_75t_R hold3781 (.A(key[4]),
    .Y(net4186));
 BUFx2_ASAP7_75t_R hold3782 (.A(key[7]),
    .Y(net4187));
 BUFx2_ASAP7_75t_R hold3783 (.A(key[0]),
    .Y(net4188));
 BUFx2_ASAP7_75t_R hold3784 (.A(key[118]),
    .Y(net4189));
 BUFx2_ASAP7_75t_R hold3785 (.A(key[103]),
    .Y(net4190));
 BUFx2_ASAP7_75t_R hold3786 (.A(key[69]),
    .Y(net4191));
 BUFx2_ASAP7_75t_R hold3787 (.A(key[71]),
    .Y(net4192));
 BUFx2_ASAP7_75t_R hold3788 (.A(key[28]),
    .Y(net4193));
 BUFx2_ASAP7_75t_R hold3789 (.A(key[70]),
    .Y(net4194));
 BUFx2_ASAP7_75t_R hold3790 (.A(key[54]),
    .Y(net4195));
 BUFx2_ASAP7_75t_R hold3791 (.A(key[31]),
    .Y(net4196));
 BUFx2_ASAP7_75t_R hold3792 (.A(key[100]),
    .Y(net4197));
 BUFx2_ASAP7_75t_R hold3793 (.A(key[99]),
    .Y(net4198));
 BUFx2_ASAP7_75t_R hold3794 (.A(key[68]),
    .Y(net4199));
 BUFx2_ASAP7_75t_R hold3795 (.A(key[38]),
    .Y(net4200));
 BUFx2_ASAP7_75t_R hold3796 (.A(key[102]),
    .Y(net4201));
 BUFx2_ASAP7_75t_R hold3797 (.A(key[73]),
    .Y(net4202));
 BUFx2_ASAP7_75t_R hold3798 (.A(key[10]),
    .Y(net4203));
 BUFx2_ASAP7_75t_R hold3799 (.A(key[9]),
    .Y(net4204));
 BUFx2_ASAP7_75t_R hold3800 (.A(key[106]),
    .Y(net4205));
 BUFx2_ASAP7_75t_R hold3801 (.A(key[104]),
    .Y(net4206));
 BUFx2_ASAP7_75t_R hold3802 (.A(key[114]),
    .Y(net4207));
 BUFx2_ASAP7_75t_R hold3803 (.A(net3591),
    .Y(net4208));
 BUFx2_ASAP7_75t_R hold3804 (.A(key[50]),
    .Y(net4209));
 BUFx2_ASAP7_75t_R hold3805 (.A(key[122]),
    .Y(net4210));
 BUFx2_ASAP7_75t_R hold3806 (.A(key[124]),
    .Y(net4211));
 BUFx2_ASAP7_75t_R hold3807 (.A(text_in[8]),
    .Y(net4212));
 BUFx2_ASAP7_75t_R hold3808 (.A(text_in[107]),
    .Y(net4213));
 BUFx2_ASAP7_75t_R hold3809 (.A(text_in[6]),
    .Y(net4214));
 BUFx2_ASAP7_75t_R hold3810 (.A(text_in[9]),
    .Y(net4215));
 BUFx2_ASAP7_75t_R hold3811 (.A(text_in[22]),
    .Y(net4216));
 BUFx2_ASAP7_75t_R hold3812 (.A(text_in[64]),
    .Y(net4217));
 BUFx2_ASAP7_75t_R hold3813 (.A(text_in[89]),
    .Y(net4218));
 BUFx2_ASAP7_75t_R hold3814 (.A(text_in[10]),
    .Y(net4219));
 BUFx2_ASAP7_75t_R hold3815 (.A(text_in[55]),
    .Y(net4220));
 BUFx2_ASAP7_75t_R hold3816 (.A(key[123]),
    .Y(net4221));
 BUFx2_ASAP7_75t_R hold3817 (.A(text_in[53]),
    .Y(net4222));
 BUFx2_ASAP7_75t_R hold3818 (.A(text_in[93]),
    .Y(net4223));
 BUFx2_ASAP7_75t_R hold3819 (.A(text_in[84]),
    .Y(net4224));
 BUFx2_ASAP7_75t_R hold3820 (.A(text_in[95]),
    .Y(net4225));
 BUFx2_ASAP7_75t_R hold3821 (.A(text_in[7]),
    .Y(net4226));
 BUFx2_ASAP7_75t_R hold3822 (.A(text_in[65]),
    .Y(net4227));
 BUFx2_ASAP7_75t_R hold3823 (.A(text_in[80]),
    .Y(net4228));
 BUFx2_ASAP7_75t_R hold3824 (.A(text_in[60]),
    .Y(net4229));
 BUFx2_ASAP7_75t_R hold3825 (.A(text_in[88]),
    .Y(net4230));
 BUFx2_ASAP7_75t_R hold3826 (.A(text_in[50]),
    .Y(net4231));
 BUFx2_ASAP7_75t_R hold3827 (.A(text_in[4]),
    .Y(net4232));
 BUFx2_ASAP7_75t_R hold3828 (.A(text_in[77]),
    .Y(net4233));
 BUFx2_ASAP7_75t_R hold3829 (.A(text_in[45]),
    .Y(net4234));
 DECAPx10_ASAP7_75t_R FILLER_0_0_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_354 ();
 DECAPx2_ASAP7_75t_R FILLER_0_0_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_432 ();
 DECAPx2_ASAP7_75t_R FILLER_0_0_454 ();
 FILLER_ASAP7_75t_R FILLER_0_0_460 ();
 FILLER_ASAP7_75t_R FILLER_0_0_464 ();
 DECAPx4_ASAP7_75t_R FILLER_0_0_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_481 ();
 FILLER_ASAP7_75t_R FILLER_0_0_487 ();
 FILLER_ASAP7_75t_R FILLER_0_0_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_496 ();
 FILLER_ASAP7_75t_R FILLER_0_0_502 ();
 FILLER_ASAP7_75t_R FILLER_0_0_509 ();
 FILLER_ASAP7_75t_R FILLER_0_0_516 ();
 FILLER_ASAP7_75t_R FILLER_0_0_523 ();
 FILLER_ASAP7_75t_R FILLER_0_0_530 ();
 FILLER_ASAP7_75t_R FILLER_0_0_537 ();
 FILLER_ASAP7_75t_R FILLER_0_0_544 ();
 FILLER_ASAP7_75t_R FILLER_0_0_551 ();
 FILLER_ASAP7_75t_R FILLER_0_0_558 ();
 FILLER_ASAP7_75t_R FILLER_0_0_565 ();
 FILLER_ASAP7_75t_R FILLER_0_0_572 ();
 FILLER_ASAP7_75t_R FILLER_0_0_579 ();
 FILLER_ASAP7_75t_R FILLER_0_0_586 ();
 FILLER_ASAP7_75t_R FILLER_0_0_593 ();
 FILLER_ASAP7_75t_R FILLER_0_0_600 ();
 FILLER_ASAP7_75t_R FILLER_0_0_607 ();
 FILLER_ASAP7_75t_R FILLER_0_0_614 ();
 FILLER_ASAP7_75t_R FILLER_0_0_621 ();
 FILLER_ASAP7_75t_R FILLER_0_0_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_631 ();
 FILLER_ASAP7_75t_R FILLER_0_0_637 ();
 FILLER_ASAP7_75t_R FILLER_0_0_644 ();
 FILLER_ASAP7_75t_R FILLER_0_0_651 ();
 FILLER_ASAP7_75t_R FILLER_0_0_658 ();
 FILLER_ASAP7_75t_R FILLER_0_0_665 ();
 FILLER_ASAP7_75t_R FILLER_0_0_672 ();
 FILLER_ASAP7_75t_R FILLER_0_0_679 ();
 FILLER_ASAP7_75t_R FILLER_0_0_686 ();
 FILLER_ASAP7_75t_R FILLER_0_0_693 ();
 FILLER_ASAP7_75t_R FILLER_0_0_700 ();
 FILLER_ASAP7_75t_R FILLER_0_0_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_710 ();
 FILLER_ASAP7_75t_R FILLER_0_0_716 ();
 FILLER_ASAP7_75t_R FILLER_0_0_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_725 ();
 FILLER_ASAP7_75t_R FILLER_0_0_736 ();
 FILLER_ASAP7_75t_R FILLER_0_0_744 ();
 FILLER_ASAP7_75t_R FILLER_0_0_751 ();
 FILLER_ASAP7_75t_R FILLER_0_0_758 ();
 FILLER_ASAP7_75t_R FILLER_0_0_765 ();
 FILLER_ASAP7_75t_R FILLER_0_0_772 ();
 FILLER_ASAP7_75t_R FILLER_0_0_779 ();
 FILLER_ASAP7_75t_R FILLER_0_0_787 ();
 FILLER_ASAP7_75t_R FILLER_0_0_794 ();
 FILLER_ASAP7_75t_R FILLER_0_0_801 ();
 FILLER_ASAP7_75t_R FILLER_0_0_808 ();
 DECAPx2_ASAP7_75t_R FILLER_0_0_815 ();
 FILLER_ASAP7_75t_R FILLER_0_0_831 ();
 FILLER_ASAP7_75t_R FILLER_0_0_838 ();
 FILLER_ASAP7_75t_R FILLER_0_0_845 ();
 FILLER_ASAP7_75t_R FILLER_0_0_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_854 ();
 FILLER_ASAP7_75t_R FILLER_0_0_865 ();
 FILLER_ASAP7_75t_R FILLER_0_0_872 ();
 FILLER_ASAP7_75t_R FILLER_0_0_879 ();
 FILLER_ASAP7_75t_R FILLER_0_0_886 ();
 FILLER_ASAP7_75t_R FILLER_0_0_893 ();
 FILLER_ASAP7_75t_R FILLER_0_0_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_902 ();
 FILLER_ASAP7_75t_R FILLER_0_0_909 ();
 FILLER_ASAP7_75t_R FILLER_0_0_917 ();
 FILLER_ASAP7_75t_R FILLER_0_0_922 ();
 FILLER_ASAP7_75t_R FILLER_0_0_926 ();
 FILLER_ASAP7_75t_R FILLER_0_0_935 ();
 DECAPx2_ASAP7_75t_R FILLER_0_0_942 ();
 FILLER_ASAP7_75t_R FILLER_0_0_954 ();
 FILLER_ASAP7_75t_R FILLER_0_0_966 ();
 DECAPx1_ASAP7_75t_R FILLER_0_0_973 ();
 FILLER_ASAP7_75t_R FILLER_0_0_987 ();
 FILLER_ASAP7_75t_R FILLER_0_0_994 ();
 FILLER_ASAP7_75t_R FILLER_0_0_1001 ();
 FILLER_ASAP7_75t_R FILLER_0_0_1008 ();
 FILLER_ASAP7_75t_R FILLER_0_0_1015 ();
 FILLER_ASAP7_75t_R FILLER_0_0_1022 ();
 FILLER_ASAP7_75t_R FILLER_0_0_1029 ();
 FILLER_ASAP7_75t_R FILLER_0_0_1036 ();
 FILLER_ASAP7_75t_R FILLER_0_0_1044 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1056 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1100 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1166 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1254 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1276 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1298 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1342 ();
 DECAPx6_ASAP7_75t_R FILLER_0_0_1364 ();
 DECAPx1_ASAP7_75t_R FILLER_0_0_1378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_332 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1_354 ();
 FILLER_ASAP7_75t_R FILLER_0_1_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_370 ();
 FILLER_ASAP7_75t_R FILLER_0_1_392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_400 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_422 ();
 FILLER_ASAP7_75t_R FILLER_0_1_431 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_436 ();
 FILLER_ASAP7_75t_R FILLER_0_1_443 ();
 FILLER_ASAP7_75t_R FILLER_0_1_451 ();
 FILLER_ASAP7_75t_R FILLER_0_1_459 ();
 FILLER_ASAP7_75t_R FILLER_0_1_467 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_475 ();
 FILLER_ASAP7_75t_R FILLER_0_1_481 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_505 ();
 FILLER_ASAP7_75t_R FILLER_0_1_514 ();
 FILLER_ASAP7_75t_R FILLER_0_1_521 ();
 FILLER_ASAP7_75t_R FILLER_0_1_528 ();
 FILLER_ASAP7_75t_R FILLER_0_1_535 ();
 FILLER_ASAP7_75t_R FILLER_0_1_542 ();
 FILLER_ASAP7_75t_R FILLER_0_1_549 ();
 FILLER_ASAP7_75t_R FILLER_0_1_556 ();
 FILLER_ASAP7_75t_R FILLER_0_1_564 ();
 FILLER_ASAP7_75t_R FILLER_0_1_572 ();
 FILLER_ASAP7_75t_R FILLER_0_1_579 ();
 FILLER_ASAP7_75t_R FILLER_0_1_586 ();
 FILLER_ASAP7_75t_R FILLER_0_1_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_596 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_603 ();
 FILLER_ASAP7_75t_R FILLER_0_1_612 ();
 FILLER_ASAP7_75t_R FILLER_0_1_619 ();
 FILLER_ASAP7_75t_R FILLER_0_1_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_645 ();
 FILLER_ASAP7_75t_R FILLER_0_1_649 ();
 FILLER_ASAP7_75t_R FILLER_0_1_656 ();
 FILLER_ASAP7_75t_R FILLER_0_1_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_666 ();
 FILLER_ASAP7_75t_R FILLER_0_1_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_691 ();
 FILLER_ASAP7_75t_R FILLER_0_1_697 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_709 ();
 FILLER_ASAP7_75t_R FILLER_0_1_718 ();
 FILLER_ASAP7_75t_R FILLER_0_1_723 ();
 FILLER_ASAP7_75t_R FILLER_0_1_746 ();
 FILLER_ASAP7_75t_R FILLER_0_1_753 ();
 FILLER_ASAP7_75t_R FILLER_0_1_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_760 ();
 FILLER_ASAP7_75t_R FILLER_0_1_782 ();
 FILLER_ASAP7_75t_R FILLER_0_1_790 ();
 FILLER_ASAP7_75t_R FILLER_0_1_798 ();
 FILLER_ASAP7_75t_R FILLER_0_1_805 ();
 FILLER_ASAP7_75t_R FILLER_0_1_810 ();
 FILLER_ASAP7_75t_R FILLER_0_1_818 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_829 ();
 FILLER_ASAP7_75t_R FILLER_0_1_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_853 ();
 FILLER_ASAP7_75t_R FILLER_0_1_860 ();
 FILLER_ASAP7_75t_R FILLER_0_1_865 ();
 FILLER_ASAP7_75t_R FILLER_0_1_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_891 ();
 FILLER_ASAP7_75t_R FILLER_0_1_913 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_924 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_931 ();
 FILLER_ASAP7_75t_R FILLER_0_1_952 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_974 ();
 FILLER_ASAP7_75t_R FILLER_0_1_984 ();
 FILLER_ASAP7_75t_R FILLER_0_1_991 ();
 FILLER_ASAP7_75t_R FILLER_0_1_998 ();
 FILLER_ASAP7_75t_R FILLER_0_1_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_1007 ();
 FILLER_ASAP7_75t_R FILLER_0_1_1019 ();
 FILLER_ASAP7_75t_R FILLER_0_1_1027 ();
 FILLER_ASAP7_75t_R FILLER_0_1_1034 ();
 FILLER_ASAP7_75t_R FILLER_0_1_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_1043 ();
 FILLER_ASAP7_75t_R FILLER_0_1_1050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1057 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1079 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1101 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1123 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1145 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1167 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1189 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1255 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1277 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1299 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1321 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1343 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1_1365 ();
 FILLER_ASAP7_75t_R FILLER_0_1_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_354 ();
 DECAPx6_ASAP7_75t_R FILLER_0_2_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_393 ();
 FILLER_ASAP7_75t_R FILLER_0_2_419 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_433 ();
 FILLER_ASAP7_75t_R FILLER_0_2_443 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_453 ();
 FILLER_ASAP7_75t_R FILLER_0_2_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_461 ();
 FILLER_ASAP7_75t_R FILLER_0_2_464 ();
 DECAPx4_ASAP7_75t_R FILLER_0_2_472 ();
 FILLER_ASAP7_75t_R FILLER_0_2_488 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_493 ();
 FILLER_ASAP7_75t_R FILLER_0_2_499 ();
 DECAPx6_ASAP7_75t_R FILLER_0_2_504 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_518 ();
 FILLER_ASAP7_75t_R FILLER_0_2_527 ();
 FILLER_ASAP7_75t_R FILLER_0_2_535 ();
 FILLER_ASAP7_75t_R FILLER_0_2_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_545 ();
 FILLER_ASAP7_75t_R FILLER_0_2_551 ();
 FILLER_ASAP7_75t_R FILLER_0_2_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_576 ();
 FILLER_ASAP7_75t_R FILLER_0_2_582 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_594 ();
 FILLER_ASAP7_75t_R FILLER_0_2_603 ();
 FILLER_ASAP7_75t_R FILLER_0_2_610 ();
 FILLER_ASAP7_75t_R FILLER_0_2_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_635 ();
 FILLER_ASAP7_75t_R FILLER_0_2_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_660 ();
 FILLER_ASAP7_75t_R FILLER_0_2_667 ();
 FILLER_ASAP7_75t_R FILLER_0_2_674 ();
 FILLER_ASAP7_75t_R FILLER_0_2_698 ();
 FILLER_ASAP7_75t_R FILLER_0_2_705 ();
 FILLER_ASAP7_75t_R FILLER_0_2_712 ();
 FILLER_ASAP7_75t_R FILLER_0_2_719 ();
 FILLER_ASAP7_75t_R FILLER_0_2_726 ();
 FILLER_ASAP7_75t_R FILLER_0_2_734 ();
 FILLER_ASAP7_75t_R FILLER_0_2_742 ();
 FILLER_ASAP7_75t_R FILLER_0_2_749 ();
 FILLER_ASAP7_75t_R FILLER_0_2_756 ();
 FILLER_ASAP7_75t_R FILLER_0_2_763 ();
 FILLER_ASAP7_75t_R FILLER_0_2_770 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_781 ();
 FILLER_ASAP7_75t_R FILLER_0_2_788 ();
 FILLER_ASAP7_75t_R FILLER_0_2_795 ();
 FILLER_ASAP7_75t_R FILLER_0_2_802 ();
 FILLER_ASAP7_75t_R FILLER_0_2_826 ();
 FILLER_ASAP7_75t_R FILLER_0_2_831 ();
 FILLER_ASAP7_75t_R FILLER_0_2_839 ();
 FILLER_ASAP7_75t_R FILLER_0_2_847 ();
 FILLER_ASAP7_75t_R FILLER_0_2_871 ();
 FILLER_ASAP7_75t_R FILLER_0_2_878 ();
 FILLER_ASAP7_75t_R FILLER_0_2_885 ();
 FILLER_ASAP7_75t_R FILLER_0_2_892 ();
 FILLER_ASAP7_75t_R FILLER_0_2_899 ();
 FILLER_ASAP7_75t_R FILLER_0_2_906 ();
 FILLER_ASAP7_75t_R FILLER_0_2_913 ();
 FILLER_ASAP7_75t_R FILLER_0_2_918 ();
 FILLER_ASAP7_75t_R FILLER_0_2_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_942 ();
 FILLER_ASAP7_75t_R FILLER_0_2_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_955 ();
 FILLER_ASAP7_75t_R FILLER_0_2_966 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_974 ();
 FILLER_ASAP7_75t_R FILLER_0_2_988 ();
 FILLER_ASAP7_75t_R FILLER_0_2_996 ();
 FILLER_ASAP7_75t_R FILLER_0_2_1004 ();
 FILLER_ASAP7_75t_R FILLER_0_2_1012 ();
 FILLER_ASAP7_75t_R FILLER_0_2_1020 ();
 FILLER_ASAP7_75t_R FILLER_0_2_1028 ();
 FILLER_ASAP7_75t_R FILLER_0_2_1036 ();
 FILLER_ASAP7_75t_R FILLER_0_2_1043 ();
 FILLER_ASAP7_75t_R FILLER_0_2_1048 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_1057 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1063 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1085 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1107 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1129 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1151 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1173 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1305 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1327 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1349 ();
 DECAPx4_ASAP7_75t_R FILLER_0_2_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_354 ();
 DECAPx6_ASAP7_75t_R FILLER_0_3_376 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_390 ();
 FILLER_ASAP7_75t_R FILLER_0_3_402 ();
 DECAPx4_ASAP7_75t_R FILLER_0_3_410 ();
 FILLER_ASAP7_75t_R FILLER_0_3_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_422 ();
 DECAPx6_ASAP7_75t_R FILLER_0_3_429 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_447 ();
 DECAPx4_ASAP7_75t_R FILLER_0_3_451 ();
 FILLER_ASAP7_75t_R FILLER_0_3_461 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_473 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_477 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_499 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_521 ();
 FILLER_ASAP7_75t_R FILLER_0_3_532 ();
 FILLER_ASAP7_75t_R FILLER_0_3_539 ();
 FILLER_ASAP7_75t_R FILLER_0_3_546 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_558 ();
 FILLER_ASAP7_75t_R FILLER_0_3_567 ();
 FILLER_ASAP7_75t_R FILLER_0_3_575 ();
 FILLER_ASAP7_75t_R FILLER_0_3_599 ();
 FILLER_ASAP7_75t_R FILLER_0_3_604 ();
 FILLER_ASAP7_75t_R FILLER_0_3_611 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_618 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_632 ();
 FILLER_ASAP7_75t_R FILLER_0_3_638 ();
 FILLER_ASAP7_75t_R FILLER_0_3_645 ();
 FILLER_ASAP7_75t_R FILLER_0_3_652 ();
 FILLER_ASAP7_75t_R FILLER_0_3_675 ();
 FILLER_ASAP7_75t_R FILLER_0_3_680 ();
 FILLER_ASAP7_75t_R FILLER_0_3_687 ();
 FILLER_ASAP7_75t_R FILLER_0_3_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_696 ();
 FILLER_ASAP7_75t_R FILLER_0_3_702 ();
 FILLER_ASAP7_75t_R FILLER_0_3_709 ();
 FILLER_ASAP7_75t_R FILLER_0_3_716 ();
 FILLER_ASAP7_75t_R FILLER_0_3_724 ();
 FILLER_ASAP7_75t_R FILLER_0_3_748 ();
 FILLER_ASAP7_75t_R FILLER_0_3_756 ();
 FILLER_ASAP7_75t_R FILLER_0_3_763 ();
 FILLER_ASAP7_75t_R FILLER_0_3_770 ();
 FILLER_ASAP7_75t_R FILLER_0_3_777 ();
 FILLER_ASAP7_75t_R FILLER_0_3_784 ();
 FILLER_ASAP7_75t_R FILLER_0_3_808 ();
 FILLER_ASAP7_75t_R FILLER_0_3_815 ();
 FILLER_ASAP7_75t_R FILLER_0_3_822 ();
 FILLER_ASAP7_75t_R FILLER_0_3_829 ();
 FILLER_ASAP7_75t_R FILLER_0_3_836 ();
 FILLER_ASAP7_75t_R FILLER_0_3_841 ();
 FILLER_ASAP7_75t_R FILLER_0_3_865 ();
 FILLER_ASAP7_75t_R FILLER_0_3_872 ();
 FILLER_ASAP7_75t_R FILLER_0_3_879 ();
 FILLER_ASAP7_75t_R FILLER_0_3_886 ();
 FILLER_ASAP7_75t_R FILLER_0_3_893 ();
 FILLER_ASAP7_75t_R FILLER_0_3_900 ();
 FILLER_ASAP7_75t_R FILLER_0_3_912 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_919 ();
 FILLER_ASAP7_75t_R FILLER_0_3_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_929 ();
 FILLER_ASAP7_75t_R FILLER_0_3_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_942 ();
 FILLER_ASAP7_75t_R FILLER_0_3_953 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_963 ();
 FILLER_ASAP7_75t_R FILLER_0_3_976 ();
 FILLER_ASAP7_75t_R FILLER_0_3_983 ();
 FILLER_ASAP7_75t_R FILLER_0_3_995 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_1006 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_1021 ();
 FILLER_ASAP7_75t_R FILLER_0_3_1032 ();
 FILLER_ASAP7_75t_R FILLER_0_3_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_1039 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_1046 ();
 FILLER_ASAP7_75t_R FILLER_0_3_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_1054 ();
 FILLER_ASAP7_75t_R FILLER_0_3_1065 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_1078 ();
 DECAPx4_ASAP7_75t_R FILLER_0_3_1085 ();
 FILLER_ASAP7_75t_R FILLER_0_3_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1117 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1139 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1161 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1293 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1315 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1337 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1359 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_310 ();
 FILLER_ASAP7_75t_R FILLER_0_4_332 ();
 FILLER_ASAP7_75t_R FILLER_0_4_340 ();
 FILLER_ASAP7_75t_R FILLER_0_4_349 ();
 DECAPx2_ASAP7_75t_R FILLER_0_4_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_4_363 ();
 FILLER_ASAP7_75t_R FILLER_0_4_367 ();
 DECAPx1_ASAP7_75t_R FILLER_0_4_375 ();
 FILLER_ASAP7_75t_R FILLER_0_4_385 ();
 FILLER_ASAP7_75t_R FILLER_0_4_397 ();
 FILLER_ASAP7_75t_R FILLER_0_4_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_4_407 ();
 FILLER_ASAP7_75t_R FILLER_0_4_419 ();
 FILLER_ASAP7_75t_R FILLER_0_4_427 ();
 DECAPx6_ASAP7_75t_R FILLER_0_4_435 ();
 DECAPx1_ASAP7_75t_R FILLER_0_4_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_4_453 ();
 FILLER_ASAP7_75t_R FILLER_0_4_460 ();
 DECAPx1_ASAP7_75t_R FILLER_0_4_464 ();
 DECAPx6_ASAP7_75t_R FILLER_0_4_474 ();
 FILLER_ASAP7_75t_R FILLER_0_4_494 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_499 ();
 DECAPx6_ASAP7_75t_R FILLER_0_4_521 ();
 DECAPx2_ASAP7_75t_R FILLER_0_4_540 ();
 FILLER_ASAP7_75t_R FILLER_0_4_552 ();
 FILLER_ASAP7_75t_R FILLER_0_4_557 ();
 FILLER_ASAP7_75t_R FILLER_0_4_564 ();
 FILLER_ASAP7_75t_R FILLER_0_4_572 ();
 FILLER_ASAP7_75t_R FILLER_0_4_579 ();
 FILLER_ASAP7_75t_R FILLER_0_4_586 ();
 FILLER_ASAP7_75t_R FILLER_0_4_593 ();
 FILLER_ASAP7_75t_R FILLER_0_4_600 ();
 FILLER_ASAP7_75t_R FILLER_0_4_608 ();
 DECAPx2_ASAP7_75t_R FILLER_0_4_615 ();
 FILLER_ASAP7_75t_R FILLER_0_4_626 ();
 DECAPx1_ASAP7_75t_R FILLER_0_4_633 ();
 FILLER_ASAP7_75t_R FILLER_0_4_642 ();
 DECAPx2_ASAP7_75t_R FILLER_0_4_650 ();
 FILLER_ASAP7_75t_R FILLER_0_4_661 ();
 DECAPx2_ASAP7_75t_R FILLER_0_4_685 ();
 DECAPx1_ASAP7_75t_R FILLER_0_4_696 ();
 DECAPx1_ASAP7_75t_R FILLER_0_4_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_4_724 ();
 FILLER_ASAP7_75t_R FILLER_0_4_730 ();
 FILLER_ASAP7_75t_R FILLER_0_4_737 ();
 DECAPx2_ASAP7_75t_R FILLER_0_4_760 ();
 FILLER_ASAP7_75t_R FILLER_0_4_788 ();
 FILLER_ASAP7_75t_R FILLER_0_4_795 ();
 FILLER_ASAP7_75t_R FILLER_0_4_802 ();
 FILLER_ASAP7_75t_R FILLER_0_4_809 ();
 DECAPx1_ASAP7_75t_R FILLER_0_4_816 ();
 FILLER_ASAP7_75t_R FILLER_0_4_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_4_828 ();
 FILLER_ASAP7_75t_R FILLER_0_4_835 ();
 FILLER_ASAP7_75t_R FILLER_0_4_858 ();
 FILLER_ASAP7_75t_R FILLER_0_4_865 ();
 FILLER_ASAP7_75t_R FILLER_0_4_872 ();
 FILLER_ASAP7_75t_R FILLER_0_4_879 ();
 FILLER_ASAP7_75t_R FILLER_0_4_886 ();
 FILLER_ASAP7_75t_R FILLER_0_4_893 ();
 FILLER_ASAP7_75t_R FILLER_0_4_900 ();
 FILLER_ASAP7_75t_R FILLER_0_4_907 ();
 FILLER_ASAP7_75t_R FILLER_0_4_912 ();
 FILLER_ASAP7_75t_R FILLER_0_4_920 ();
 FILLER_ASAP7_75t_R FILLER_0_4_928 ();
 FILLER_ASAP7_75t_R FILLER_0_4_935 ();
 FILLER_ASAP7_75t_R FILLER_0_4_943 ();
 FILLER_ASAP7_75t_R FILLER_0_4_955 ();
 FILLER_ASAP7_75t_R FILLER_0_4_967 ();
 FILLER_ASAP7_75t_R FILLER_0_4_975 ();
 FILLER_ASAP7_75t_R FILLER_0_4_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_4_982 ();
 DECAPx1_ASAP7_75t_R FILLER_0_4_993 ();
 FILLER_ASAP7_75t_R FILLER_0_4_1007 ();
 FILLER_ASAP7_75t_R FILLER_0_4_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_4_1021 ();
 FILLER_ASAP7_75t_R FILLER_0_4_1032 ();
 FILLER_ASAP7_75t_R FILLER_0_4_1040 ();
 FILLER_ASAP7_75t_R FILLER_0_4_1048 ();
 DECAPx2_ASAP7_75t_R FILLER_0_4_1056 ();
 FILLER_ASAP7_75t_R FILLER_0_4_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_4_1069 ();
 DECAPx1_ASAP7_75t_R FILLER_0_4_1078 ();
 FILLER_ASAP7_75t_R FILLER_0_4_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_4_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1166 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1210 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1254 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1276 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1298 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1342 ();
 DECAPx6_ASAP7_75t_R FILLER_0_4_1364 ();
 DECAPx1_ASAP7_75t_R FILLER_0_4_1378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_310 ();
 DECAPx4_ASAP7_75t_R FILLER_0_5_332 ();
 FILLER_ASAP7_75t_R FILLER_0_5_342 ();
 DECAPx1_ASAP7_75t_R FILLER_0_5_350 ();
 FILLER_ASAP7_75t_R FILLER_0_5_357 ();
 FILLER_ASAP7_75t_R FILLER_0_5_365 ();
 DECAPx4_ASAP7_75t_R FILLER_0_5_373 ();
 DECAPx2_ASAP7_75t_R FILLER_0_5_389 ();
 FILLER_ASAP7_75t_R FILLER_0_5_395 ();
 DECAPx4_ASAP7_75t_R FILLER_0_5_403 ();
 FILLER_ASAP7_75t_R FILLER_0_5_413 ();
 FILLER_ASAP7_75t_R FILLER_0_5_421 ();
 FILLER_ASAP7_75t_R FILLER_0_5_429 ();
 DECAPx6_ASAP7_75t_R FILLER_0_5_437 ();
 DECAPx2_ASAP7_75t_R FILLER_0_5_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_457 ();
 FILLER_ASAP7_75t_R FILLER_0_5_464 ();
 FILLER_ASAP7_75t_R FILLER_0_5_472 ();
 FILLER_ASAP7_75t_R FILLER_0_5_480 ();
 FILLER_ASAP7_75t_R FILLER_0_5_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_490 ();
 FILLER_ASAP7_75t_R FILLER_0_5_501 ();
 DECAPx1_ASAP7_75t_R FILLER_0_5_509 ();
 FILLER_ASAP7_75t_R FILLER_0_5_519 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_521 ();
 DECAPx6_ASAP7_75t_R FILLER_0_5_528 ();
 DECAPx1_ASAP7_75t_R FILLER_0_5_542 ();
 FILLER_ASAP7_75t_R FILLER_0_5_549 ();
 FILLER_ASAP7_75t_R FILLER_0_5_556 ();
 FILLER_ASAP7_75t_R FILLER_0_5_579 ();
 FILLER_ASAP7_75t_R FILLER_0_5_586 ();
 DECAPx2_ASAP7_75t_R FILLER_0_5_593 ();
 FILLER_ASAP7_75t_R FILLER_0_5_620 ();
 FILLER_ASAP7_75t_R FILLER_0_5_628 ();
 FILLER_ASAP7_75t_R FILLER_0_5_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_653 ();
 FILLER_ASAP7_75t_R FILLER_0_5_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_676 ();
 DECAPx1_ASAP7_75t_R FILLER_0_5_683 ();
 DECAPx1_ASAP7_75t_R FILLER_0_5_690 ();
 FILLER_ASAP7_75t_R FILLER_0_5_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_701 ();
 FILLER_ASAP7_75t_R FILLER_0_5_705 ();
 FILLER_ASAP7_75t_R FILLER_0_5_710 ();
 FILLER_ASAP7_75t_R FILLER_0_5_718 ();
 FILLER_ASAP7_75t_R FILLER_0_5_726 ();
 DECAPx4_ASAP7_75t_R FILLER_0_5_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_741 ();
 FILLER_ASAP7_75t_R FILLER_0_5_745 ();
 FILLER_ASAP7_75t_R FILLER_0_5_753 ();
 FILLER_ASAP7_75t_R FILLER_0_5_760 ();
 FILLER_ASAP7_75t_R FILLER_0_5_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_769 ();
 FILLER_ASAP7_75t_R FILLER_0_5_775 ();
 FILLER_ASAP7_75t_R FILLER_0_5_782 ();
 FILLER_ASAP7_75t_R FILLER_0_5_787 ();
 FILLER_ASAP7_75t_R FILLER_0_5_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_796 ();
 FILLER_ASAP7_75t_R FILLER_0_5_819 ();
 FILLER_ASAP7_75t_R FILLER_0_5_826 ();
 DECAPx1_ASAP7_75t_R FILLER_0_5_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_837 ();
 FILLER_ASAP7_75t_R FILLER_0_5_844 ();
 FILLER_ASAP7_75t_R FILLER_0_5_852 ();
 FILLER_ASAP7_75t_R FILLER_0_5_859 ();
 FILLER_ASAP7_75t_R FILLER_0_5_866 ();
 FILLER_ASAP7_75t_R FILLER_0_5_873 ();
 FILLER_ASAP7_75t_R FILLER_0_5_880 ();
 DECAPx1_ASAP7_75t_R FILLER_0_5_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_892 ();
 DECAPx1_ASAP7_75t_R FILLER_0_5_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_903 ();
 FILLER_ASAP7_75t_R FILLER_0_5_914 ();
 DECAPx1_ASAP7_75t_R FILLER_0_5_921 ();
 FILLER_ASAP7_75t_R FILLER_0_5_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_929 ();
 FILLER_ASAP7_75t_R FILLER_0_5_940 ();
 DECAPx1_ASAP7_75t_R FILLER_0_5_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_956 ();
 FILLER_ASAP7_75t_R FILLER_0_5_967 ();
 FILLER_ASAP7_75t_R FILLER_0_5_975 ();
 FILLER_ASAP7_75t_R FILLER_0_5_982 ();
 FILLER_ASAP7_75t_R FILLER_0_5_994 ();
 DECAPx1_ASAP7_75t_R FILLER_0_5_1006 ();
 DECAPx1_ASAP7_75t_R FILLER_0_5_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_1024 ();
 DECAPx1_ASAP7_75t_R FILLER_0_5_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_1036 ();
 DECAPx2_ASAP7_75t_R FILLER_0_5_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_1049 ();
 FILLER_ASAP7_75t_R FILLER_0_5_1057 ();
 FILLER_ASAP7_75t_R FILLER_0_5_1069 ();
 FILLER_ASAP7_75t_R FILLER_0_5_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_1079 ();
 FILLER_ASAP7_75t_R FILLER_0_5_1090 ();
 FILLER_ASAP7_75t_R FILLER_0_5_1097 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_1099 ();
 FILLER_ASAP7_75t_R FILLER_0_5_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1358 ();
 FILLER_ASAP7_75t_R FILLER_0_5_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_310 ();
 DECAPx6_ASAP7_75t_R FILLER_0_6_332 ();
 DECAPx2_ASAP7_75t_R FILLER_0_6_346 ();
 FILLER_ASAP7_75t_R FILLER_0_6_358 ();
 FILLER_ASAP7_75t_R FILLER_0_6_366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_6_374 ();
 FILLER_ASAP7_75t_R FILLER_0_6_380 ();
 DECAPx1_ASAP7_75t_R FILLER_0_6_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_394 ();
 FILLER_ASAP7_75t_R FILLER_0_6_401 ();
 DECAPx4_ASAP7_75t_R FILLER_0_6_409 ();
 FILLER_ASAP7_75t_R FILLER_0_6_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_421 ();
 FILLER_ASAP7_75t_R FILLER_0_6_428 ();
 FILLER_ASAP7_75t_R FILLER_0_6_438 ();
 FILLER_ASAP7_75t_R FILLER_0_6_450 ();
 FILLER_ASAP7_75t_R FILLER_0_6_460 ();
 DECAPx2_ASAP7_75t_R FILLER_0_6_464 ();
 FILLER_ASAP7_75t_R FILLER_0_6_470 ();
 FILLER_ASAP7_75t_R FILLER_0_6_478 ();
 FILLER_ASAP7_75t_R FILLER_0_6_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_489 ();
 FILLER_ASAP7_75t_R FILLER_0_6_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_498 ();
 FILLER_ASAP7_75t_R FILLER_0_6_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_507 ();
 DECAPx1_ASAP7_75t_R FILLER_0_6_511 ();
 FILLER_ASAP7_75t_R FILLER_0_6_521 ();
 DECAPx6_ASAP7_75t_R FILLER_0_6_529 ();
 DECAPx1_ASAP7_75t_R FILLER_0_6_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_547 ();
 FILLER_ASAP7_75t_R FILLER_0_6_554 ();
 DECAPx2_ASAP7_75t_R FILLER_0_6_561 ();
 DECAPx1_ASAP7_75t_R FILLER_0_6_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_576 ();
 DECAPx2_ASAP7_75t_R FILLER_0_6_582 ();
 DECAPx2_ASAP7_75t_R FILLER_0_6_593 ();
 FILLER_ASAP7_75t_R FILLER_0_6_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_606 ();
 FILLER_ASAP7_75t_R FILLER_0_6_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_615 ();
 FILLER_ASAP7_75t_R FILLER_0_6_619 ();
 FILLER_ASAP7_75t_R FILLER_0_6_624 ();
 FILLER_ASAP7_75t_R FILLER_0_6_629 ();
 FILLER_ASAP7_75t_R FILLER_0_6_634 ();
 FILLER_ASAP7_75t_R FILLER_0_6_639 ();
 DECAPx1_ASAP7_75t_R FILLER_0_6_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_667 ();
 FILLER_ASAP7_75t_R FILLER_0_6_673 ();
 FILLER_ASAP7_75t_R FILLER_0_6_681 ();
 FILLER_ASAP7_75t_R FILLER_0_6_688 ();
 DECAPx1_ASAP7_75t_R FILLER_0_6_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_697 ();
 DECAPx1_ASAP7_75t_R FILLER_0_6_719 ();
 FILLER_ASAP7_75t_R FILLER_0_6_729 ();
 DECAPx1_ASAP7_75t_R FILLER_0_6_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_741 ();
 FILLER_ASAP7_75t_R FILLER_0_6_745 ();
 FILLER_ASAP7_75t_R FILLER_0_6_750 ();
 FILLER_ASAP7_75t_R FILLER_0_6_755 ();
 FILLER_ASAP7_75t_R FILLER_0_6_760 ();
 FILLER_ASAP7_75t_R FILLER_0_6_784 ();
 DECAPx1_ASAP7_75t_R FILLER_0_6_792 ();
 FILLER_ASAP7_75t_R FILLER_0_6_802 ();
 FILLER_ASAP7_75t_R FILLER_0_6_809 ();
 FILLER_ASAP7_75t_R FILLER_0_6_816 ();
 FILLER_ASAP7_75t_R FILLER_0_6_823 ();
 FILLER_ASAP7_75t_R FILLER_0_6_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_830 ();
 FILLER_ASAP7_75t_R FILLER_0_6_852 ();
 FILLER_ASAP7_75t_R FILLER_0_6_859 ();
 FILLER_ASAP7_75t_R FILLER_0_6_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_868 ();
 FILLER_ASAP7_75t_R FILLER_0_6_879 ();
 FILLER_ASAP7_75t_R FILLER_0_6_887 ();
 DECAPx1_ASAP7_75t_R FILLER_0_6_899 ();
 FILLER_ASAP7_75t_R FILLER_0_6_913 ();
 DECAPx1_ASAP7_75t_R FILLER_0_6_921 ();
 FILLER_ASAP7_75t_R FILLER_0_6_931 ();
 DECAPx1_ASAP7_75t_R FILLER_0_6_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_946 ();
 DECAPx1_ASAP7_75t_R FILLER_0_6_965 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_969 ();
 DECAPx2_ASAP7_75t_R FILLER_0_6_982 ();
 FILLER_ASAP7_75t_R FILLER_0_6_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_1000 ();
 FILLER_ASAP7_75t_R FILLER_0_6_1009 ();
 FILLER_ASAP7_75t_R FILLER_0_6_1016 ();
 FILLER_ASAP7_75t_R FILLER_0_6_1024 ();
 FILLER_ASAP7_75t_R FILLER_0_6_1032 ();
 FILLER_ASAP7_75t_R FILLER_0_6_1039 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_1041 ();
 FILLER_ASAP7_75t_R FILLER_0_6_1048 ();
 FILLER_ASAP7_75t_R FILLER_0_6_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_1058 ();
 DECAPx1_ASAP7_75t_R FILLER_0_6_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_1071 ();
 FILLER_ASAP7_75t_R FILLER_0_6_1082 ();
 FILLER_ASAP7_75t_R FILLER_0_6_1122 ();
 FILLER_ASAP7_75t_R FILLER_0_6_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1141 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1251 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1273 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1295 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1317 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1339 ();
 DECAPx6_ASAP7_75t_R FILLER_0_6_1361 ();
 DECAPx2_ASAP7_75t_R FILLER_0_6_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_310 ();
 DECAPx4_ASAP7_75t_R FILLER_0_7_332 ();
 FILLER_ASAP7_75t_R FILLER_0_7_342 ();
 DECAPx6_ASAP7_75t_R FILLER_0_7_360 ();
 DECAPx2_ASAP7_75t_R FILLER_0_7_374 ();
 DECAPx6_ASAP7_75t_R FILLER_0_7_386 ();
 DECAPx1_ASAP7_75t_R FILLER_0_7_400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_415 ();
 DECAPx4_ASAP7_75t_R FILLER_0_7_437 ();
 FILLER_ASAP7_75t_R FILLER_0_7_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7_449 ();
 FILLER_ASAP7_75t_R FILLER_0_7_456 ();
 FILLER_ASAP7_75t_R FILLER_0_7_478 ();
 DECAPx2_ASAP7_75t_R FILLER_0_7_486 ();
 FILLER_ASAP7_75t_R FILLER_0_7_492 ();
 FILLER_ASAP7_75t_R FILLER_0_7_500 ();
 DECAPx4_ASAP7_75t_R FILLER_0_7_509 ();
 DECAPx1_ASAP7_75t_R FILLER_0_7_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7_528 ();
 DECAPx4_ASAP7_75t_R FILLER_0_7_535 ();
 FILLER_ASAP7_75t_R FILLER_0_7_551 ();
 FILLER_ASAP7_75t_R FILLER_0_7_559 ();
 DECAPx1_ASAP7_75t_R FILLER_0_7_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7_568 ();
 FILLER_ASAP7_75t_R FILLER_0_7_572 ();
 FILLER_ASAP7_75t_R FILLER_0_7_580 ();
 DECAPx1_ASAP7_75t_R FILLER_0_7_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7_591 ();
 FILLER_ASAP7_75t_R FILLER_0_7_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7_600 ();
 DECAPx1_ASAP7_75t_R FILLER_0_7_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7_610 ();
 FILLER_ASAP7_75t_R FILLER_0_7_614 ();
 FILLER_ASAP7_75t_R FILLER_0_7_638 ();
 FILLER_ASAP7_75t_R FILLER_0_7_643 ();
 DECAPx1_ASAP7_75t_R FILLER_0_7_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7_655 ();
 DECAPx1_ASAP7_75t_R FILLER_0_7_659 ();
 FILLER_ASAP7_75t_R FILLER_0_7_666 ();
 FILLER_ASAP7_75t_R FILLER_0_7_689 ();
 FILLER_ASAP7_75t_R FILLER_0_7_713 ();
 DECAPx1_ASAP7_75t_R FILLER_0_7_720 ();
 DECAPx2_ASAP7_75t_R FILLER_0_7_745 ();
 FILLER_ASAP7_75t_R FILLER_0_7_751 ();
 DECAPx1_ASAP7_75t_R FILLER_0_7_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7_763 ();
 FILLER_ASAP7_75t_R FILLER_0_7_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7_769 ();
 DECAPx2_ASAP7_75t_R FILLER_0_7_776 ();
 FILLER_ASAP7_75t_R FILLER_0_7_803 ();
 DECAPx1_ASAP7_75t_R FILLER_0_7_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7_815 ();
 FILLER_ASAP7_75t_R FILLER_0_7_821 ();
 FILLER_ASAP7_75t_R FILLER_0_7_829 ();
 FILLER_ASAP7_75t_R FILLER_0_7_837 ();
 FILLER_ASAP7_75t_R FILLER_0_7_844 ();
 FILLER_ASAP7_75t_R FILLER_0_7_851 ();
 FILLER_ASAP7_75t_R FILLER_0_7_858 ();
 FILLER_ASAP7_75t_R FILLER_0_7_863 ();
 FILLER_ASAP7_75t_R FILLER_0_7_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7_888 ();
 FILLER_ASAP7_75t_R FILLER_0_7_913 ();
 DECAPx1_ASAP7_75t_R FILLER_0_7_921 ();
 FILLER_ASAP7_75t_R FILLER_0_7_927 ();
 FILLER_ASAP7_75t_R FILLER_0_7_932 ();
 DECAPx2_ASAP7_75t_R FILLER_0_7_942 ();
 FILLER_ASAP7_75t_R FILLER_0_7_958 ();
 FILLER_ASAP7_75t_R FILLER_0_7_966 ();
 FILLER_ASAP7_75t_R FILLER_0_7_974 ();
 FILLER_ASAP7_75t_R FILLER_0_7_981 ();
 FILLER_ASAP7_75t_R FILLER_0_7_1001 ();
 DECAPx1_ASAP7_75t_R FILLER_0_7_1009 ();
 DECAPx1_ASAP7_75t_R FILLER_0_7_1023 ();
 DECAPx1_ASAP7_75t_R FILLER_0_7_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7_1036 ();
 FILLER_ASAP7_75t_R FILLER_0_7_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7_1049 ();
 FILLER_ASAP7_75t_R FILLER_0_7_1057 ();
 FILLER_ASAP7_75t_R FILLER_0_7_1067 ();
 FILLER_ASAP7_75t_R FILLER_0_7_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7_1078 ();
 FILLER_ASAP7_75t_R FILLER_0_7_1085 ();
 FILLER_ASAP7_75t_R FILLER_0_7_1117 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1129 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1151 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1173 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1305 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1327 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1349 ();
 DECAPx4_ASAP7_75t_R FILLER_0_7_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_310 ();
 DECAPx4_ASAP7_75t_R FILLER_0_8_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8_342 ();
 DECAPx1_ASAP7_75t_R FILLER_0_8_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8_350 ();
 DECAPx6_ASAP7_75t_R FILLER_0_8_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_383 ();
 DECAPx6_ASAP7_75t_R FILLER_0_8_405 ();
 FILLER_ASAP7_75t_R FILLER_0_8_425 ();
 DECAPx1_ASAP7_75t_R FILLER_0_8_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8_447 ();
 DECAPx2_ASAP7_75t_R FILLER_0_8_454 ();
 FILLER_ASAP7_75t_R FILLER_0_8_460 ();
 FILLER_ASAP7_75t_R FILLER_0_8_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8_498 ();
 DECAPx6_ASAP7_75t_R FILLER_0_8_505 ();
 FILLER_ASAP7_75t_R FILLER_0_8_525 ();
 FILLER_ASAP7_75t_R FILLER_0_8_530 ();
 DECAPx4_ASAP7_75t_R FILLER_0_8_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8_554 ();
 DECAPx4_ASAP7_75t_R FILLER_0_8_561 ();
 FILLER_ASAP7_75t_R FILLER_0_8_592 ();
 FILLER_ASAP7_75t_R FILLER_0_8_616 ();
 FILLER_ASAP7_75t_R FILLER_0_8_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8_623 ();
 FILLER_ASAP7_75t_R FILLER_0_8_646 ();
 FILLER_ASAP7_75t_R FILLER_0_8_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8_653 ();
 FILLER_ASAP7_75t_R FILLER_0_8_657 ();
 FILLER_ASAP7_75t_R FILLER_0_8_662 ();
 DECAPx6_ASAP7_75t_R FILLER_0_8_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8_681 ();
 FILLER_ASAP7_75t_R FILLER_0_8_685 ();
 FILLER_ASAP7_75t_R FILLER_0_8_690 ();
 FILLER_ASAP7_75t_R FILLER_0_8_698 ();
 DECAPx4_ASAP7_75t_R FILLER_0_8_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8_713 ();
 FILLER_ASAP7_75t_R FILLER_0_8_717 ();
 FILLER_ASAP7_75t_R FILLER_0_8_722 ();
 FILLER_ASAP7_75t_R FILLER_0_8_729 ();
 FILLER_ASAP7_75t_R FILLER_0_8_752 ();
 FILLER_ASAP7_75t_R FILLER_0_8_775 ();
 FILLER_ASAP7_75t_R FILLER_0_8_780 ();
 FILLER_ASAP7_75t_R FILLER_0_8_787 ();
 FILLER_ASAP7_75t_R FILLER_0_8_810 ();
 FILLER_ASAP7_75t_R FILLER_0_8_833 ();
 FILLER_ASAP7_75t_R FILLER_0_8_840 ();
 DECAPx1_ASAP7_75t_R FILLER_0_8_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8_851 ();
 FILLER_ASAP7_75t_R FILLER_0_8_873 ();
 DECAPx1_ASAP7_75t_R FILLER_0_8_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8_884 ();
 FILLER_ASAP7_75t_R FILLER_0_8_891 ();
 FILLER_ASAP7_75t_R FILLER_0_8_901 ();
 FILLER_ASAP7_75t_R FILLER_0_8_908 ();
 FILLER_ASAP7_75t_R FILLER_0_8_916 ();
 DECAPx1_ASAP7_75t_R FILLER_0_8_928 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8_932 ();
 DECAPx1_ASAP7_75t_R FILLER_0_8_939 ();
 FILLER_ASAP7_75t_R FILLER_0_8_951 ();
 FILLER_ASAP7_75t_R FILLER_0_8_963 ();
 FILLER_ASAP7_75t_R FILLER_0_8_971 ();
 DECAPx2_ASAP7_75t_R FILLER_0_8_979 ();
 DECAPx2_ASAP7_75t_R FILLER_0_8_995 ();
 FILLER_ASAP7_75t_R FILLER_0_8_1007 ();
 DECAPx1_ASAP7_75t_R FILLER_0_8_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8_1018 ();
 DECAPx2_ASAP7_75t_R FILLER_0_8_1025 ();
 FILLER_ASAP7_75t_R FILLER_0_8_1031 ();
 DECAPx2_ASAP7_75t_R FILLER_0_8_1039 ();
 DECAPx2_ASAP7_75t_R FILLER_0_8_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8_1061 ();
 FILLER_ASAP7_75t_R FILLER_0_8_1072 ();
 DECAPx1_ASAP7_75t_R FILLER_0_8_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8_1088 ();
 FILLER_ASAP7_75t_R FILLER_0_8_1094 ();
 FILLER_ASAP7_75t_R FILLER_0_8_1106 ();
 FILLER_ASAP7_75t_R FILLER_0_8_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1147 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1169 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1257 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1301 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1323 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1345 ();
 DECAPx6_ASAP7_75t_R FILLER_0_8_1367 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_310 ();
 DECAPx6_ASAP7_75t_R FILLER_0_9_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_346 ();
 FILLER_ASAP7_75t_R FILLER_0_9_353 ();
 FILLER_ASAP7_75t_R FILLER_0_9_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_363 ();
 FILLER_ASAP7_75t_R FILLER_0_9_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_372 ();
 FILLER_ASAP7_75t_R FILLER_0_9_385 ();
 DECAPx1_ASAP7_75t_R FILLER_0_9_393 ();
 DECAPx1_ASAP7_75t_R FILLER_0_9_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_407 ();
 DECAPx4_ASAP7_75t_R FILLER_0_9_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_424 ();
 DECAPx6_ASAP7_75t_R FILLER_0_9_431 ();
 FILLER_ASAP7_75t_R FILLER_0_9_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_447 ();
 DECAPx6_ASAP7_75t_R FILLER_0_9_454 ();
 DECAPx2_ASAP7_75t_R FILLER_0_9_468 ();
 FILLER_ASAP7_75t_R FILLER_0_9_480 ();
 DECAPx2_ASAP7_75t_R FILLER_0_9_485 ();
 FILLER_ASAP7_75t_R FILLER_0_9_491 ();
 FILLER_ASAP7_75t_R FILLER_0_9_499 ();
 DECAPx1_ASAP7_75t_R FILLER_0_9_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_511 ();
 FILLER_ASAP7_75t_R FILLER_0_9_517 ();
 FILLER_ASAP7_75t_R FILLER_0_9_539 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_547 ();
 FILLER_ASAP7_75t_R FILLER_0_9_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_571 ();
 FILLER_ASAP7_75t_R FILLER_0_9_575 ();
 DECAPx2_ASAP7_75t_R FILLER_0_9_583 ();
 FILLER_ASAP7_75t_R FILLER_0_9_589 ();
 FILLER_ASAP7_75t_R FILLER_0_9_594 ();
 FILLER_ASAP7_75t_R FILLER_0_9_599 ();
 DECAPx2_ASAP7_75t_R FILLER_0_9_604 ();
 FILLER_ASAP7_75t_R FILLER_0_9_613 ();
 FILLER_ASAP7_75t_R FILLER_0_9_618 ();
 FILLER_ASAP7_75t_R FILLER_0_9_626 ();
 DECAPx4_ASAP7_75t_R FILLER_0_9_631 ();
 FILLER_ASAP7_75t_R FILLER_0_9_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_643 ();
 DECAPx6_ASAP7_75t_R FILLER_0_9_654 ();
 DECAPx1_ASAP7_75t_R FILLER_0_9_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_672 ();
 DECAPx2_ASAP7_75t_R FILLER_0_9_683 ();
 FILLER_ASAP7_75t_R FILLER_0_9_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_691 ();
 DECAPx4_ASAP7_75t_R FILLER_0_9_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_708 ();
 FILLER_ASAP7_75t_R FILLER_0_9_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_717 ();
 FILLER_ASAP7_75t_R FILLER_0_9_740 ();
 DECAPx2_ASAP7_75t_R FILLER_0_9_745 ();
 FILLER_ASAP7_75t_R FILLER_0_9_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_753 ();
 FILLER_ASAP7_75t_R FILLER_0_9_757 ();
 DECAPx1_ASAP7_75t_R FILLER_0_9_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_768 ();
 FILLER_ASAP7_75t_R FILLER_0_9_775 ();
 DECAPx2_ASAP7_75t_R FILLER_0_9_787 ();
 DECAPx2_ASAP7_75t_R FILLER_0_9_799 ();
 FILLER_ASAP7_75t_R FILLER_0_9_811 ();
 FILLER_ASAP7_75t_R FILLER_0_9_818 ();
 DECAPx1_ASAP7_75t_R FILLER_0_9_825 ();
 FILLER_ASAP7_75t_R FILLER_0_9_839 ();
 FILLER_ASAP7_75t_R FILLER_0_9_847 ();
 FILLER_ASAP7_75t_R FILLER_0_9_855 ();
 FILLER_ASAP7_75t_R FILLER_0_9_862 ();
 FILLER_ASAP7_75t_R FILLER_0_9_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_871 ();
 DECAPx2_ASAP7_75t_R FILLER_0_9_878 ();
 FILLER_ASAP7_75t_R FILLER_0_9_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_893 ();
 FILLER_ASAP7_75t_R FILLER_0_9_904 ();
 FILLER_ASAP7_75t_R FILLER_0_9_914 ();
 DECAPx1_ASAP7_75t_R FILLER_0_9_921 ();
 FILLER_ASAP7_75t_R FILLER_0_9_927 ();
 FILLER_ASAP7_75t_R FILLER_0_9_934 ();
 FILLER_ASAP7_75t_R FILLER_0_9_939 ();
 FILLER_ASAP7_75t_R FILLER_0_9_947 ();
 DECAPx1_ASAP7_75t_R FILLER_0_9_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_959 ();
 FILLER_ASAP7_75t_R FILLER_0_9_970 ();
 FILLER_ASAP7_75t_R FILLER_0_9_978 ();
 FILLER_ASAP7_75t_R FILLER_0_9_983 ();
 FILLER_ASAP7_75t_R FILLER_0_9_991 ();
 FILLER_ASAP7_75t_R FILLER_0_9_998 ();
 FILLER_ASAP7_75t_R FILLER_0_9_1005 ();
 FILLER_ASAP7_75t_R FILLER_0_9_1012 ();
 FILLER_ASAP7_75t_R FILLER_0_9_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_1023 ();
 FILLER_ASAP7_75t_R FILLER_0_9_1034 ();
 DECAPx2_ASAP7_75t_R FILLER_0_9_1042 ();
 FILLER_ASAP7_75t_R FILLER_0_9_1048 ();
 DECAPx1_ASAP7_75t_R FILLER_0_9_1068 ();
 FILLER_ASAP7_75t_R FILLER_0_9_1078 ();
 FILLER_ASAP7_75t_R FILLER_0_9_1090 ();
 FILLER_ASAP7_75t_R FILLER_0_9_1102 ();
 FILLER_ASAP7_75t_R FILLER_0_9_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1120 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1142 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1164 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1252 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1274 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1296 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1318 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1340 ();
 DECAPx6_ASAP7_75t_R FILLER_0_9_1362 ();
 DECAPx2_ASAP7_75t_R FILLER_0_9_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_112 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_168 ();
 DECAPx6_ASAP7_75t_R FILLER_0_10_190 ();
 DECAPx1_ASAP7_75t_R FILLER_0_10_204 ();
 FILLER_ASAP7_75t_R FILLER_0_10_214 ();
 FILLER_ASAP7_75t_R FILLER_0_10_222 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_230 ();
 DECAPx1_ASAP7_75t_R FILLER_0_10_242 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_252 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_274 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_296 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_318 ();
 FILLER_ASAP7_75t_R FILLER_0_10_346 ();
 DECAPx6_ASAP7_75t_R FILLER_0_10_358 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_372 ();
 DECAPx1_ASAP7_75t_R FILLER_0_10_384 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_400 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_407 ();
 DECAPx1_ASAP7_75t_R FILLER_0_10_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_424 ();
 DECAPx4_ASAP7_75t_R FILLER_0_10_431 ();
 FILLER_ASAP7_75t_R FILLER_0_10_441 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_454 ();
 FILLER_ASAP7_75t_R FILLER_0_10_460 ();
 FILLER_ASAP7_75t_R FILLER_0_10_464 ();
 FILLER_ASAP7_75t_R FILLER_0_10_474 ();
 DECAPx1_ASAP7_75t_R FILLER_0_10_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_493 ();
 DECAPx4_ASAP7_75t_R FILLER_0_10_515 ();
 DECAPx1_ASAP7_75t_R FILLER_0_10_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_537 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_541 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_569 ();
 FILLER_ASAP7_75t_R FILLER_0_10_576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_584 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_606 ();
 FILLER_ASAP7_75t_R FILLER_0_10_612 ();
 DECAPx1_ASAP7_75t_R FILLER_0_10_617 ();
 DECAPx1_ASAP7_75t_R FILLER_0_10_642 ();
 FILLER_ASAP7_75t_R FILLER_0_10_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_670 ();
 FILLER_ASAP7_75t_R FILLER_0_10_677 ();
 FILLER_ASAP7_75t_R FILLER_0_10_682 ();
 FILLER_ASAP7_75t_R FILLER_0_10_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_707 ();
 FILLER_ASAP7_75t_R FILLER_0_10_715 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_723 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_739 ();
 FILLER_ASAP7_75t_R FILLER_0_10_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_763 ();
 DECAPx6_ASAP7_75t_R FILLER_0_10_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_781 ();
 FILLER_ASAP7_75t_R FILLER_0_10_787 ();
 FILLER_ASAP7_75t_R FILLER_0_10_795 ();
 FILLER_ASAP7_75t_R FILLER_0_10_800 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_807 ();
 FILLER_ASAP7_75t_R FILLER_0_10_818 ();
 FILLER_ASAP7_75t_R FILLER_0_10_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_827 ();
 FILLER_ASAP7_75t_R FILLER_0_10_833 ();
 FILLER_ASAP7_75t_R FILLER_0_10_840 ();
 FILLER_ASAP7_75t_R FILLER_0_10_850 ();
 FILLER_ASAP7_75t_R FILLER_0_10_855 ();
 FILLER_ASAP7_75t_R FILLER_0_10_869 ();
 FILLER_ASAP7_75t_R FILLER_0_10_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_878 ();
 FILLER_ASAP7_75t_R FILLER_0_10_884 ();
 FILLER_ASAP7_75t_R FILLER_0_10_891 ();
 DECAPx1_ASAP7_75t_R FILLER_0_10_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_907 ();
 FILLER_ASAP7_75t_R FILLER_0_10_915 ();
 FILLER_ASAP7_75t_R FILLER_0_10_923 ();
 FILLER_ASAP7_75t_R FILLER_0_10_928 ();
 FILLER_ASAP7_75t_R FILLER_0_10_938 ();
 FILLER_ASAP7_75t_R FILLER_0_10_949 ();
 FILLER_ASAP7_75t_R FILLER_0_10_961 ();
 FILLER_ASAP7_75t_R FILLER_0_10_969 ();
 FILLER_ASAP7_75t_R FILLER_0_10_977 ();
 FILLER_ASAP7_75t_R FILLER_0_10_984 ();
 FILLER_ASAP7_75t_R FILLER_0_10_996 ();
 DECAPx4_ASAP7_75t_R FILLER_0_10_1004 ();
 FILLER_ASAP7_75t_R FILLER_0_10_1014 ();
 DECAPx6_ASAP7_75t_R FILLER_0_10_1022 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_1042 ();
 FILLER_ASAP7_75t_R FILLER_0_10_1048 ();
 FILLER_ASAP7_75t_R FILLER_0_10_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_1062 ();
 FILLER_ASAP7_75t_R FILLER_0_10_1069 ();
 FILLER_ASAP7_75t_R FILLER_0_10_1077 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_1089 ();
 FILLER_ASAP7_75t_R FILLER_0_10_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1153 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1263 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1285 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1307 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1351 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_10_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_90 ();
 DECAPx6_ASAP7_75t_R FILLER_0_11_112 ();
 DECAPx2_ASAP7_75t_R FILLER_0_11_126 ();
 FILLER_ASAP7_75t_R FILLER_0_11_137 ();
 DECAPx4_ASAP7_75t_R FILLER_0_11_159 ();
 DECAPx1_ASAP7_75t_R FILLER_0_11_175 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_185 ();
 DECAPx2_ASAP7_75t_R FILLER_0_11_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_213 ();
 FILLER_ASAP7_75t_R FILLER_0_11_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_224 ();
 DECAPx2_ASAP7_75t_R FILLER_0_11_233 ();
 FILLER_ASAP7_75t_R FILLER_0_11_239 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_252 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_274 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_296 ();
 DECAPx4_ASAP7_75t_R FILLER_0_11_318 ();
 FILLER_ASAP7_75t_R FILLER_0_11_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_330 ();
 DECAPx1_ASAP7_75t_R FILLER_0_11_337 ();
 DECAPx1_ASAP7_75t_R FILLER_0_11_346 ();
 FILLER_ASAP7_75t_R FILLER_0_11_366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_374 ();
 FILLER_ASAP7_75t_R FILLER_0_11_396 ();
 FILLER_ASAP7_75t_R FILLER_0_11_404 ();
 FILLER_ASAP7_75t_R FILLER_0_11_426 ();
 DECAPx2_ASAP7_75t_R FILLER_0_11_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_440 ();
 FILLER_ASAP7_75t_R FILLER_0_11_447 ();
 DECAPx4_ASAP7_75t_R FILLER_0_11_455 ();
 FILLER_ASAP7_75t_R FILLER_0_11_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_467 ();
 DECAPx6_ASAP7_75t_R FILLER_0_11_471 ();
 FILLER_ASAP7_75t_R FILLER_0_11_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_487 ();
 DECAPx6_ASAP7_75t_R FILLER_0_11_491 ();
 FILLER_ASAP7_75t_R FILLER_0_11_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_507 ();
 DECAPx2_ASAP7_75t_R FILLER_0_11_514 ();
 FILLER_ASAP7_75t_R FILLER_0_11_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_522 ();
 FILLER_ASAP7_75t_R FILLER_0_11_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_535 ();
 DECAPx4_ASAP7_75t_R FILLER_0_11_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_552 ();
 DECAPx4_ASAP7_75t_R FILLER_0_11_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_569 ();
 DECAPx2_ASAP7_75t_R FILLER_0_11_591 ();
 FILLER_ASAP7_75t_R FILLER_0_11_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_599 ();
 DECAPx2_ASAP7_75t_R FILLER_0_11_606 ();
 FILLER_ASAP7_75t_R FILLER_0_11_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_614 ();
 DECAPx1_ASAP7_75t_R FILLER_0_11_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_625 ();
 FILLER_ASAP7_75t_R FILLER_0_11_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_633 ();
 DECAPx1_ASAP7_75t_R FILLER_0_11_640 ();
 FILLER_ASAP7_75t_R FILLER_0_11_647 ();
 FILLER_ASAP7_75t_R FILLER_0_11_655 ();
 DECAPx6_ASAP7_75t_R FILLER_0_11_679 ();
 FILLER_ASAP7_75t_R FILLER_0_11_698 ();
 FILLER_ASAP7_75t_R FILLER_0_11_703 ();
 DECAPx1_ASAP7_75t_R FILLER_0_11_716 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_723 ();
 FILLER_ASAP7_75t_R FILLER_0_11_767 ();
 FILLER_ASAP7_75t_R FILLER_0_11_790 ();
 FILLER_ASAP7_75t_R FILLER_0_11_798 ();
 FILLER_ASAP7_75t_R FILLER_0_11_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_812 ();
 FILLER_ASAP7_75t_R FILLER_0_11_816 ();
 FILLER_ASAP7_75t_R FILLER_0_11_821 ();
 FILLER_ASAP7_75t_R FILLER_0_11_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_833 ();
 FILLER_ASAP7_75t_R FILLER_0_11_840 ();
 FILLER_ASAP7_75t_R FILLER_0_11_850 ();
 FILLER_ASAP7_75t_R FILLER_0_11_857 ();
 FILLER_ASAP7_75t_R FILLER_0_11_864 ();
 FILLER_ASAP7_75t_R FILLER_0_11_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_873 ();
 FILLER_ASAP7_75t_R FILLER_0_11_879 ();
 FILLER_ASAP7_75t_R FILLER_0_11_891 ();
 FILLER_ASAP7_75t_R FILLER_0_11_903 ();
 FILLER_ASAP7_75t_R FILLER_0_11_915 ();
 FILLER_ASAP7_75t_R FILLER_0_11_923 ();
 DECAPx1_ASAP7_75t_R FILLER_0_11_927 ();
 DECAPx1_ASAP7_75t_R FILLER_0_11_941 ();
 FILLER_ASAP7_75t_R FILLER_0_11_955 ();
 FILLER_ASAP7_75t_R FILLER_0_11_962 ();
 FILLER_ASAP7_75t_R FILLER_0_11_969 ();
 FILLER_ASAP7_75t_R FILLER_0_11_974 ();
 FILLER_ASAP7_75t_R FILLER_0_11_986 ();
 FILLER_ASAP7_75t_R FILLER_0_11_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_993 ();
 DECAPx2_ASAP7_75t_R FILLER_0_11_1014 ();
 FILLER_ASAP7_75t_R FILLER_0_11_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_1022 ();
 DECAPx2_ASAP7_75t_R FILLER_0_11_1029 ();
 DECAPx1_ASAP7_75t_R FILLER_0_11_1041 ();
 FILLER_ASAP7_75t_R FILLER_0_11_1051 ();
 DECAPx2_ASAP7_75t_R FILLER_0_11_1062 ();
 FILLER_ASAP7_75t_R FILLER_0_11_1068 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_1070 ();
 DECAPx2_ASAP7_75t_R FILLER_0_11_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_1083 ();
 DECAPx6_ASAP7_75t_R FILLER_0_11_1094 ();
 FILLER_ASAP7_75t_R FILLER_0_11_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1143 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1319 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1341 ();
 DECAPx6_ASAP7_75t_R FILLER_0_11_1363 ();
 DECAPx1_ASAP7_75t_R FILLER_0_11_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_90 ();
 DECAPx4_ASAP7_75t_R FILLER_0_12_112 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_130 ();
 FILLER_ASAP7_75t_R FILLER_0_12_146 ();
 DECAPx1_ASAP7_75t_R FILLER_0_12_158 ();
 FILLER_ASAP7_75t_R FILLER_0_12_168 ();
 FILLER_ASAP7_75t_R FILLER_0_12_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_180 ();
 FILLER_ASAP7_75t_R FILLER_0_12_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_191 ();
 DECAPx1_ASAP7_75t_R FILLER_0_12_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_202 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_209 ();
 FILLER_ASAP7_75t_R FILLER_0_12_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_223 ();
 DECAPx1_ASAP7_75t_R FILLER_0_12_244 ();
 FILLER_ASAP7_75t_R FILLER_0_12_254 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_262 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_284 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_306 ();
 DECAPx1_ASAP7_75t_R FILLER_0_12_328 ();
 FILLER_ASAP7_75t_R FILLER_0_12_338 ();
 FILLER_ASAP7_75t_R FILLER_0_12_346 ();
 FILLER_ASAP7_75t_R FILLER_0_12_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_353 ();
 FILLER_ASAP7_75t_R FILLER_0_12_360 ();
 FILLER_ASAP7_75t_R FILLER_0_12_368 ();
 DECAPx4_ASAP7_75t_R FILLER_0_12_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_386 ();
 FILLER_ASAP7_75t_R FILLER_0_12_393 ();
 DECAPx1_ASAP7_75t_R FILLER_0_12_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_405 ();
 FILLER_ASAP7_75t_R FILLER_0_12_416 ();
 FILLER_ASAP7_75t_R FILLER_0_12_424 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_433 ();
 FILLER_ASAP7_75t_R FILLER_0_12_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_441 ();
 FILLER_ASAP7_75t_R FILLER_0_12_448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_456 ();
 FILLER_ASAP7_75t_R FILLER_0_12_464 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_474 ();
 FILLER_ASAP7_75t_R FILLER_0_12_480 ();
 DECAPx1_ASAP7_75t_R FILLER_0_12_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_497 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_514 ();
 FILLER_ASAP7_75t_R FILLER_0_12_526 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_531 ();
 FILLER_ASAP7_75t_R FILLER_0_12_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_539 ();
 FILLER_ASAP7_75t_R FILLER_0_12_543 ();
 FILLER_ASAP7_75t_R FILLER_0_12_551 ();
 DECAPx4_ASAP7_75t_R FILLER_0_12_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_569 ();
 FILLER_ASAP7_75t_R FILLER_0_12_573 ();
 DECAPx6_ASAP7_75t_R FILLER_0_12_580 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_600 ();
 FILLER_ASAP7_75t_R FILLER_0_12_622 ();
 FILLER_ASAP7_75t_R FILLER_0_12_630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_635 ();
 FILLER_ASAP7_75t_R FILLER_0_12_657 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_662 ();
 FILLER_ASAP7_75t_R FILLER_0_12_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_670 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_677 ();
 FILLER_ASAP7_75t_R FILLER_0_12_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_685 ();
 DECAPx6_ASAP7_75t_R FILLER_0_12_692 ();
 DECAPx1_ASAP7_75t_R FILLER_0_12_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_710 ();
 FILLER_ASAP7_75t_R FILLER_0_12_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_725 ();
 DECAPx4_ASAP7_75t_R FILLER_0_12_737 ();
 DECAPx6_ASAP7_75t_R FILLER_0_12_750 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_770 ();
 DECAPx4_ASAP7_75t_R FILLER_0_12_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_784 ();
 FILLER_ASAP7_75t_R FILLER_0_12_805 ();
 DECAPx1_ASAP7_75t_R FILLER_0_12_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_814 ();
 FILLER_ASAP7_75t_R FILLER_0_12_823 ();
 DECAPx1_ASAP7_75t_R FILLER_0_12_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_837 ();
 FILLER_ASAP7_75t_R FILLER_0_12_843 ();
 FILLER_ASAP7_75t_R FILLER_0_12_850 ();
 FILLER_ASAP7_75t_R FILLER_0_12_857 ();
 FILLER_ASAP7_75t_R FILLER_0_12_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_866 ();
 FILLER_ASAP7_75t_R FILLER_0_12_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_874 ();
 FILLER_ASAP7_75t_R FILLER_0_12_885 ();
 FILLER_ASAP7_75t_R FILLER_0_12_890 ();
 FILLER_ASAP7_75t_R FILLER_0_12_910 ();
 FILLER_ASAP7_75t_R FILLER_0_12_922 ();
 FILLER_ASAP7_75t_R FILLER_0_12_934 ();
 FILLER_ASAP7_75t_R FILLER_0_12_946 ();
 FILLER_ASAP7_75t_R FILLER_0_12_954 ();
 DECAPx1_ASAP7_75t_R FILLER_0_12_962 ();
 FILLER_ASAP7_75t_R FILLER_0_12_972 ();
 FILLER_ASAP7_75t_R FILLER_0_12_980 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_987 ();
 FILLER_ASAP7_75t_R FILLER_0_12_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_995 ();
 DECAPx4_ASAP7_75t_R FILLER_0_12_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_1013 ();
 FILLER_ASAP7_75t_R FILLER_0_12_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_1022 ();
 FILLER_ASAP7_75t_R FILLER_0_12_1033 ();
 FILLER_ASAP7_75t_R FILLER_0_12_1043 ();
 DECAPx1_ASAP7_75t_R FILLER_0_12_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_1057 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_1068 ();
 FILLER_ASAP7_75t_R FILLER_0_12_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_12_1214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_1228 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_1240 ();
 FILLER_ASAP7_75t_R FILLER_0_12_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1254 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1276 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1298 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1342 ();
 DECAPx6_ASAP7_75t_R FILLER_0_12_1364 ();
 DECAPx1_ASAP7_75t_R FILLER_0_12_1378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_90 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_118 ();
 FILLER_ASAP7_75t_R FILLER_0_13_130 ();
 DECAPx1_ASAP7_75t_R FILLER_0_13_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_142 ();
 FILLER_ASAP7_75t_R FILLER_0_13_163 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_171 ();
 FILLER_ASAP7_75t_R FILLER_0_13_177 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_185 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_199 ();
 FILLER_ASAP7_75t_R FILLER_0_13_205 ();
 FILLER_ASAP7_75t_R FILLER_0_13_212 ();
 FILLER_ASAP7_75t_R FILLER_0_13_220 ();
 FILLER_ASAP7_75t_R FILLER_0_13_229 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_236 ();
 FILLER_ASAP7_75t_R FILLER_0_13_242 ();
 FILLER_ASAP7_75t_R FILLER_0_13_252 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_264 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_286 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_330 ();
 DECAPx1_ASAP7_75t_R FILLER_0_13_337 ();
 FILLER_ASAP7_75t_R FILLER_0_13_347 ();
 FILLER_ASAP7_75t_R FILLER_0_13_355 ();
 DECAPx6_ASAP7_75t_R FILLER_0_13_364 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_390 ();
 FILLER_ASAP7_75t_R FILLER_0_13_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_403 ();
 FILLER_ASAP7_75t_R FILLER_0_13_410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_418 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_452 ();
 FILLER_ASAP7_75t_R FILLER_0_13_459 ();
 DECAPx4_ASAP7_75t_R FILLER_0_13_471 ();
 FILLER_ASAP7_75t_R FILLER_0_13_481 ();
 FILLER_ASAP7_75t_R FILLER_0_13_495 ();
 FILLER_ASAP7_75t_R FILLER_0_13_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_505 ();
 DECAPx4_ASAP7_75t_R FILLER_0_13_516 ();
 FILLER_ASAP7_75t_R FILLER_0_13_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_528 ();
 FILLER_ASAP7_75t_R FILLER_0_13_535 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_544 ();
 FILLER_ASAP7_75t_R FILLER_0_13_550 ();
 FILLER_ASAP7_75t_R FILLER_0_13_558 ();
 DECAPx4_ASAP7_75t_R FILLER_0_13_571 ();
 FILLER_ASAP7_75t_R FILLER_0_13_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_583 ();
 FILLER_ASAP7_75t_R FILLER_0_13_590 ();
 FILLER_ASAP7_75t_R FILLER_0_13_604 ();
 FILLER_ASAP7_75t_R FILLER_0_13_611 ();
 DECAPx4_ASAP7_75t_R FILLER_0_13_616 ();
 FILLER_ASAP7_75t_R FILLER_0_13_626 ();
 DECAPx6_ASAP7_75t_R FILLER_0_13_634 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_666 ();
 FILLER_ASAP7_75t_R FILLER_0_13_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_673 ();
 FILLER_ASAP7_75t_R FILLER_0_13_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_684 ();
 DECAPx1_ASAP7_75t_R FILLER_0_13_689 ();
 FILLER_ASAP7_75t_R FILLER_0_13_699 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_709 ();
 FILLER_ASAP7_75t_R FILLER_0_13_715 ();
 DECAPx1_ASAP7_75t_R FILLER_0_13_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_729 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_736 ();
 FILLER_ASAP7_75t_R FILLER_0_13_742 ();
 FILLER_ASAP7_75t_R FILLER_0_13_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_785 ();
 FILLER_ASAP7_75t_R FILLER_0_13_792 ();
 DECAPx6_ASAP7_75t_R FILLER_0_13_797 ();
 DECAPx1_ASAP7_75t_R FILLER_0_13_811 ();
 FILLER_ASAP7_75t_R FILLER_0_13_823 ();
 DECAPx4_ASAP7_75t_R FILLER_0_13_831 ();
 FILLER_ASAP7_75t_R FILLER_0_13_851 ();
 DECAPx1_ASAP7_75t_R FILLER_0_13_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_862 ();
 FILLER_ASAP7_75t_R FILLER_0_13_869 ();
 DECAPx1_ASAP7_75t_R FILLER_0_13_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_885 ();
 DECAPx1_ASAP7_75t_R FILLER_0_13_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_900 ();
 FILLER_ASAP7_75t_R FILLER_0_13_913 ();
 DECAPx1_ASAP7_75t_R FILLER_0_13_921 ();
 FILLER_ASAP7_75t_R FILLER_0_13_927 ();
 FILLER_ASAP7_75t_R FILLER_0_13_939 ();
 FILLER_ASAP7_75t_R FILLER_0_13_947 ();
 FILLER_ASAP7_75t_R FILLER_0_13_955 ();
 FILLER_ASAP7_75t_R FILLER_0_13_963 ();
 FILLER_ASAP7_75t_R FILLER_0_13_968 ();
 FILLER_ASAP7_75t_R FILLER_0_13_973 ();
 DECAPx6_ASAP7_75t_R FILLER_0_13_981 ();
 DECAPx4_ASAP7_75t_R FILLER_0_13_1005 ();
 DECAPx6_ASAP7_75t_R FILLER_0_13_1021 ();
 FILLER_ASAP7_75t_R FILLER_0_13_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_1043 ();
 FILLER_ASAP7_75t_R FILLER_0_13_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_1056 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_1073 ();
 FILLER_ASAP7_75t_R FILLER_0_13_1084 ();
 FILLER_ASAP7_75t_R FILLER_0_13_1092 ();
 DECAPx1_ASAP7_75t_R FILLER_0_13_1099 ();
 FILLER_ASAP7_75t_R FILLER_0_13_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_1111 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1162 ();
 DECAPx4_ASAP7_75t_R FILLER_0_13_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_1194 ();
 DECAPx4_ASAP7_75t_R FILLER_0_13_1198 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_1214 ();
 FILLER_ASAP7_75t_R FILLER_0_13_1220 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_1222 ();
 FILLER_ASAP7_75t_R FILLER_0_13_1233 ();
 DECAPx4_ASAP7_75t_R FILLER_0_13_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_1248 ();
 FILLER_ASAP7_75t_R FILLER_0_13_1255 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1260 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_1282 ();
 FILLER_ASAP7_75t_R FILLER_0_13_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_1290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_1301 ();
 FILLER_ASAP7_75t_R FILLER_0_13_1307 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1356 ();
 DECAPx1_ASAP7_75t_R FILLER_0_13_1378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_68 ();
 DECAPx6_ASAP7_75t_R FILLER_0_14_90 ();
 FILLER_ASAP7_75t_R FILLER_0_14_110 ();
 FILLER_ASAP7_75t_R FILLER_0_14_120 ();
 DECAPx1_ASAP7_75t_R FILLER_0_14_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_136 ();
 FILLER_ASAP7_75t_R FILLER_0_14_143 ();
 DECAPx1_ASAP7_75t_R FILLER_0_14_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_157 ();
 FILLER_ASAP7_75t_R FILLER_0_14_165 ();
 DECAPx2_ASAP7_75t_R FILLER_0_14_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_179 ();
 FILLER_ASAP7_75t_R FILLER_0_14_186 ();
 DECAPx6_ASAP7_75t_R FILLER_0_14_194 ();
 FILLER_ASAP7_75t_R FILLER_0_14_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_210 ();
 FILLER_ASAP7_75t_R FILLER_0_14_217 ();
 FILLER_ASAP7_75t_R FILLER_0_14_222 ();
 DECAPx1_ASAP7_75t_R FILLER_0_14_230 ();
 DECAPx1_ASAP7_75t_R FILLER_0_14_242 ();
 FILLER_ASAP7_75t_R FILLER_0_14_252 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_264 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_286 ();
 DECAPx2_ASAP7_75t_R FILLER_0_14_308 ();
 FILLER_ASAP7_75t_R FILLER_0_14_314 ();
 FILLER_ASAP7_75t_R FILLER_0_14_328 ();
 DECAPx2_ASAP7_75t_R FILLER_0_14_342 ();
 FILLER_ASAP7_75t_R FILLER_0_14_348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_392 ();
 FILLER_ASAP7_75t_R FILLER_0_14_398 ();
 DECAPx2_ASAP7_75t_R FILLER_0_14_408 ();
 FILLER_ASAP7_75t_R FILLER_0_14_414 ();
 FILLER_ASAP7_75t_R FILLER_0_14_426 ();
 DECAPx4_ASAP7_75t_R FILLER_0_14_434 ();
 FILLER_ASAP7_75t_R FILLER_0_14_444 ();
 FILLER_ASAP7_75t_R FILLER_0_14_449 ();
 FILLER_ASAP7_75t_R FILLER_0_14_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_486 ();
 DECAPx4_ASAP7_75t_R FILLER_0_14_499 ();
 DECAPx2_ASAP7_75t_R FILLER_0_14_515 ();
 FILLER_ASAP7_75t_R FILLER_0_14_521 ();
 FILLER_ASAP7_75t_R FILLER_0_14_529 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_537 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_559 ();
 DECAPx4_ASAP7_75t_R FILLER_0_14_581 ();
 FILLER_ASAP7_75t_R FILLER_0_14_591 ();
 FILLER_ASAP7_75t_R FILLER_0_14_601 ();
 DECAPx2_ASAP7_75t_R FILLER_0_14_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_639 ();
 DECAPx1_ASAP7_75t_R FILLER_0_14_661 ();
 FILLER_ASAP7_75t_R FILLER_0_14_673 ();
 FILLER_ASAP7_75t_R FILLER_0_14_683 ();
 FILLER_ASAP7_75t_R FILLER_0_14_691 ();
 DECAPx1_ASAP7_75t_R FILLER_0_14_699 ();
 DECAPx1_ASAP7_75t_R FILLER_0_14_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_715 ();
 DECAPx1_ASAP7_75t_R FILLER_0_14_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_728 ();
 DECAPx1_ASAP7_75t_R FILLER_0_14_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_741 ();
 FILLER_ASAP7_75t_R FILLER_0_14_753 ();
 FILLER_ASAP7_75t_R FILLER_0_14_776 ();
 DECAPx6_ASAP7_75t_R FILLER_0_14_790 ();
 FILLER_ASAP7_75t_R FILLER_0_14_804 ();
 FILLER_ASAP7_75t_R FILLER_0_14_817 ();
 FILLER_ASAP7_75t_R FILLER_0_14_825 ();
 DECAPx2_ASAP7_75t_R FILLER_0_14_830 ();
 FILLER_ASAP7_75t_R FILLER_0_14_836 ();
 FILLER_ASAP7_75t_R FILLER_0_14_842 ();
 FILLER_ASAP7_75t_R FILLER_0_14_854 ();
 DECAPx2_ASAP7_75t_R FILLER_0_14_866 ();
 DECAPx1_ASAP7_75t_R FILLER_0_14_882 ();
 FILLER_ASAP7_75t_R FILLER_0_14_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_898 ();
 DECAPx1_ASAP7_75t_R FILLER_0_14_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_913 ();
 FILLER_ASAP7_75t_R FILLER_0_14_920 ();
 FILLER_ASAP7_75t_R FILLER_0_14_928 ();
 FILLER_ASAP7_75t_R FILLER_0_14_937 ();
 FILLER_ASAP7_75t_R FILLER_0_14_945 ();
 FILLER_ASAP7_75t_R FILLER_0_14_953 ();
 FILLER_ASAP7_75t_R FILLER_0_14_963 ();
 FILLER_ASAP7_75t_R FILLER_0_14_973 ();
 DECAPx2_ASAP7_75t_R FILLER_0_14_981 ();
 FILLER_ASAP7_75t_R FILLER_0_14_993 ();
 FILLER_ASAP7_75t_R FILLER_0_14_1001 ();
 DECAPx1_ASAP7_75t_R FILLER_0_14_1009 ();
 FILLER_ASAP7_75t_R FILLER_0_14_1019 ();
 FILLER_ASAP7_75t_R FILLER_0_14_1028 ();
 FILLER_ASAP7_75t_R FILLER_0_14_1038 ();
 FILLER_ASAP7_75t_R FILLER_0_14_1050 ();
 FILLER_ASAP7_75t_R FILLER_0_14_1062 ();
 FILLER_ASAP7_75t_R FILLER_0_14_1070 ();
 FILLER_ASAP7_75t_R FILLER_0_14_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_0_14_1092 ();
 FILLER_ASAP7_75t_R FILLER_0_14_1104 ();
 FILLER_ASAP7_75t_R FILLER_0_14_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_1147 ();
 DECAPx6_ASAP7_75t_R FILLER_0_14_1169 ();
 FILLER_ASAP7_75t_R FILLER_0_14_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_1185 ();
 DECAPx1_ASAP7_75t_R FILLER_0_14_1192 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_1196 ();
 FILLER_ASAP7_75t_R FILLER_0_14_1203 ();
 DECAPx2_ASAP7_75t_R FILLER_0_14_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_1221 ();
 DECAPx4_ASAP7_75t_R FILLER_0_14_1228 ();
 FILLER_ASAP7_75t_R FILLER_0_14_1244 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_1258 ();
 DECAPx6_ASAP7_75t_R FILLER_0_14_1280 ();
 DECAPx1_ASAP7_75t_R FILLER_0_14_1294 ();
 FILLER_ASAP7_75t_R FILLER_0_14_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_1338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_1360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_68 ();
 DECAPx4_ASAP7_75t_R FILLER_0_15_90 ();
 FILLER_ASAP7_75t_R FILLER_0_15_100 ();
 FILLER_ASAP7_75t_R FILLER_0_15_108 ();
 FILLER_ASAP7_75t_R FILLER_0_15_116 ();
 FILLER_ASAP7_75t_R FILLER_0_15_124 ();
 FILLER_ASAP7_75t_R FILLER_0_15_136 ();
 DECAPx2_ASAP7_75t_R FILLER_0_15_148 ();
 FILLER_ASAP7_75t_R FILLER_0_15_164 ();
 FILLER_ASAP7_75t_R FILLER_0_15_172 ();
 FILLER_ASAP7_75t_R FILLER_0_15_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_182 ();
 FILLER_ASAP7_75t_R FILLER_0_15_189 ();
 DECAPx2_ASAP7_75t_R FILLER_0_15_196 ();
 FILLER_ASAP7_75t_R FILLER_0_15_202 ();
 FILLER_ASAP7_75t_R FILLER_0_15_214 ();
 FILLER_ASAP7_75t_R FILLER_0_15_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_225 ();
 FILLER_ASAP7_75t_R FILLER_0_15_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_239 ();
 FILLER_ASAP7_75t_R FILLER_0_15_260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_274 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_296 ();
 DECAPx4_ASAP7_75t_R FILLER_0_15_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_328 ();
 DECAPx6_ASAP7_75t_R FILLER_0_15_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_355 ();
 DECAPx4_ASAP7_75t_R FILLER_0_15_366 ();
 DECAPx4_ASAP7_75t_R FILLER_0_15_382 ();
 FILLER_ASAP7_75t_R FILLER_0_15_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_394 ();
 FILLER_ASAP7_75t_R FILLER_0_15_405 ();
 FILLER_ASAP7_75t_R FILLER_0_15_415 ();
 FILLER_ASAP7_75t_R FILLER_0_15_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_433 ();
 DECAPx2_ASAP7_75t_R FILLER_0_15_465 ();
 FILLER_ASAP7_75t_R FILLER_0_15_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_473 ();
 DECAPx6_ASAP7_75t_R FILLER_0_15_486 ();
 FILLER_ASAP7_75t_R FILLER_0_15_500 ();
 FILLER_ASAP7_75t_R FILLER_0_15_508 ();
 DECAPx4_ASAP7_75t_R FILLER_0_15_516 ();
 FILLER_ASAP7_75t_R FILLER_0_15_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_528 ();
 DECAPx6_ASAP7_75t_R FILLER_0_15_536 ();
 FILLER_ASAP7_75t_R FILLER_0_15_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_552 ();
 FILLER_ASAP7_75t_R FILLER_0_15_559 ();
 DECAPx1_ASAP7_75t_R FILLER_0_15_567 ();
 DECAPx2_ASAP7_75t_R FILLER_0_15_581 ();
 FILLER_ASAP7_75t_R FILLER_0_15_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_589 ();
 FILLER_ASAP7_75t_R FILLER_0_15_598 ();
 FILLER_ASAP7_75t_R FILLER_0_15_603 ();
 DECAPx1_ASAP7_75t_R FILLER_0_15_611 ();
 DECAPx1_ASAP7_75t_R FILLER_0_15_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_631 ();
 DECAPx6_ASAP7_75t_R FILLER_0_15_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_649 ();
 FILLER_ASAP7_75t_R FILLER_0_15_662 ();
 FILLER_ASAP7_75t_R FILLER_0_15_672 ();
 FILLER_ASAP7_75t_R FILLER_0_15_680 ();
 DECAPx4_ASAP7_75t_R FILLER_0_15_692 ();
 DECAPx1_ASAP7_75t_R FILLER_0_15_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_716 ();
 DECAPx1_ASAP7_75t_R FILLER_0_15_725 ();
 FILLER_ASAP7_75t_R FILLER_0_15_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_739 ();
 DECAPx2_ASAP7_75t_R FILLER_0_15_750 ();
 FILLER_ASAP7_75t_R FILLER_0_15_762 ();
 DECAPx6_ASAP7_75t_R FILLER_0_15_767 ();
 DECAPx4_ASAP7_75t_R FILLER_0_15_802 ();
 DECAPx6_ASAP7_75t_R FILLER_0_15_822 ();
 FILLER_ASAP7_75t_R FILLER_0_15_836 ();
 DECAPx1_ASAP7_75t_R FILLER_0_15_843 ();
 FILLER_ASAP7_75t_R FILLER_0_15_852 ();
 FILLER_ASAP7_75t_R FILLER_0_15_864 ();
 FILLER_ASAP7_75t_R FILLER_0_15_872 ();
 FILLER_ASAP7_75t_R FILLER_0_15_877 ();
 FILLER_ASAP7_75t_R FILLER_0_15_889 ();
 FILLER_ASAP7_75t_R FILLER_0_15_901 ();
 FILLER_ASAP7_75t_R FILLER_0_15_913 ();
 DECAPx1_ASAP7_75t_R FILLER_0_15_921 ();
 DECAPx1_ASAP7_75t_R FILLER_0_15_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_931 ();
 FILLER_ASAP7_75t_R FILLER_0_15_944 ();
 FILLER_ASAP7_75t_R FILLER_0_15_956 ();
 FILLER_ASAP7_75t_R FILLER_0_15_964 ();
 DECAPx1_ASAP7_75t_R FILLER_0_15_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_977 ();
 FILLER_ASAP7_75t_R FILLER_0_15_986 ();
 FILLER_ASAP7_75t_R FILLER_0_15_994 ();
 DECAPx4_ASAP7_75t_R FILLER_0_15_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_1012 ();
 FILLER_ASAP7_75t_R FILLER_0_15_1020 ();
 DECAPx1_ASAP7_75t_R FILLER_0_15_1032 ();
 FILLER_ASAP7_75t_R FILLER_0_15_1041 ();
 FILLER_ASAP7_75t_R FILLER_0_15_1048 ();
 DECAPx1_ASAP7_75t_R FILLER_0_15_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_1059 ();
 FILLER_ASAP7_75t_R FILLER_0_15_1070 ();
 DECAPx1_ASAP7_75t_R FILLER_0_15_1082 ();
 DECAPx1_ASAP7_75t_R FILLER_0_15_1098 ();
 FILLER_ASAP7_75t_R FILLER_0_15_1108 ();
 FILLER_ASAP7_75t_R FILLER_0_15_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_1143 ();
 DECAPx2_ASAP7_75t_R FILLER_0_15_1165 ();
 FILLER_ASAP7_75t_R FILLER_0_15_1177 ();
 FILLER_ASAP7_75t_R FILLER_0_15_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_1198 ();
 DECAPx1_ASAP7_75t_R FILLER_0_15_1220 ();
 FILLER_ASAP7_75t_R FILLER_0_15_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_1237 ();
 DECAPx6_ASAP7_75t_R FILLER_0_15_1259 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_1273 ();
 DECAPx6_ASAP7_75t_R FILLER_0_15_1280 ();
 DECAPx1_ASAP7_75t_R FILLER_0_15_1294 ();
 DECAPx1_ASAP7_75t_R FILLER_0_15_1301 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_1311 ();
 DECAPx6_ASAP7_75t_R FILLER_0_15_1333 ();
 FILLER_ASAP7_75t_R FILLER_0_15_1347 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_1349 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_1353 ();
 DECAPx2_ASAP7_75t_R FILLER_0_15_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_68 ();
 FILLER_ASAP7_75t_R FILLER_0_16_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_92 ();
 FILLER_ASAP7_75t_R FILLER_0_16_98 ();
 DECAPx1_ASAP7_75t_R FILLER_0_16_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_114 ();
 FILLER_ASAP7_75t_R FILLER_0_16_126 ();
 FILLER_ASAP7_75t_R FILLER_0_16_146 ();
 FILLER_ASAP7_75t_R FILLER_0_16_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_157 ();
 FILLER_ASAP7_75t_R FILLER_0_16_164 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_176 ();
 DECAPx6_ASAP7_75t_R FILLER_0_16_188 ();
 DECAPx1_ASAP7_75t_R FILLER_0_16_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_206 ();
 DECAPx1_ASAP7_75t_R FILLER_0_16_227 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_241 ();
 DECAPx4_ASAP7_75t_R FILLER_0_16_253 ();
 FILLER_ASAP7_75t_R FILLER_0_16_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_265 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_294 ();
 DECAPx4_ASAP7_75t_R FILLER_0_16_316 ();
 FILLER_ASAP7_75t_R FILLER_0_16_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_328 ();
 DECAPx1_ASAP7_75t_R FILLER_0_16_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_353 ();
 DECAPx6_ASAP7_75t_R FILLER_0_16_360 ();
 DECAPx1_ASAP7_75t_R FILLER_0_16_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_384 ();
 FILLER_ASAP7_75t_R FILLER_0_16_405 ();
 DECAPx4_ASAP7_75t_R FILLER_0_16_415 ();
 FILLER_ASAP7_75t_R FILLER_0_16_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_427 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_453 ();
 FILLER_ASAP7_75t_R FILLER_0_16_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_461 ();
 FILLER_ASAP7_75t_R FILLER_0_16_464 ();
 DECAPx1_ASAP7_75t_R FILLER_0_16_472 ();
 DECAPx6_ASAP7_75t_R FILLER_0_16_483 ();
 DECAPx1_ASAP7_75t_R FILLER_0_16_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_501 ();
 DECAPx6_ASAP7_75t_R FILLER_0_16_508 ();
 DECAPx1_ASAP7_75t_R FILLER_0_16_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_526 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_533 ();
 FILLER_ASAP7_75t_R FILLER_0_16_545 ();
 FILLER_ASAP7_75t_R FILLER_0_16_553 ();
 DECAPx1_ASAP7_75t_R FILLER_0_16_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_565 ();
 DECAPx4_ASAP7_75t_R FILLER_0_16_572 ();
 FILLER_ASAP7_75t_R FILLER_0_16_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_584 ();
 FILLER_ASAP7_75t_R FILLER_0_16_591 ();
 FILLER_ASAP7_75t_R FILLER_0_16_599 ();
 DECAPx6_ASAP7_75t_R FILLER_0_16_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_618 ();
 FILLER_ASAP7_75t_R FILLER_0_16_624 ();
 FILLER_ASAP7_75t_R FILLER_0_16_634 ();
 FILLER_ASAP7_75t_R FILLER_0_16_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_644 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_667 ();
 FILLER_ASAP7_75t_R FILLER_0_16_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_675 ();
 FILLER_ASAP7_75t_R FILLER_0_16_688 ();
 DECAPx6_ASAP7_75t_R FILLER_0_16_700 ();
 FILLER_ASAP7_75t_R FILLER_0_16_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_716 ();
 FILLER_ASAP7_75t_R FILLER_0_16_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_727 ();
 FILLER_ASAP7_75t_R FILLER_0_16_738 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_750 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_763 ();
 FILLER_ASAP7_75t_R FILLER_0_16_781 ();
 FILLER_ASAP7_75t_R FILLER_0_16_789 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_800 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_813 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_820 ();
 FILLER_ASAP7_75t_R FILLER_0_16_848 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_866 ();
 FILLER_ASAP7_75t_R FILLER_0_16_877 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_884 ();
 FILLER_ASAP7_75t_R FILLER_0_16_908 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_916 ();
 DECAPx1_ASAP7_75t_R FILLER_0_16_930 ();
 FILLER_ASAP7_75t_R FILLER_0_16_952 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_966 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_977 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_999 ();
 FILLER_ASAP7_75t_R FILLER_0_16_1005 ();
 FILLER_ASAP7_75t_R FILLER_0_16_1013 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_1021 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_1033 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_1039 ();
 FILLER_ASAP7_75t_R FILLER_0_16_1046 ();
 FILLER_ASAP7_75t_R FILLER_0_16_1055 ();
 FILLER_ASAP7_75t_R FILLER_0_16_1067 ();
 FILLER_ASAP7_75t_R FILLER_0_16_1079 ();
 FILLER_ASAP7_75t_R FILLER_0_16_1091 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_1099 ();
 FILLER_ASAP7_75t_R FILLER_0_16_1111 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_1119 ();
 DECAPx6_ASAP7_75t_R FILLER_0_16_1141 ();
 FILLER_ASAP7_75t_R FILLER_0_16_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_1157 ();
 FILLER_ASAP7_75t_R FILLER_0_16_1166 ();
 FILLER_ASAP7_75t_R FILLER_0_16_1174 ();
 FILLER_ASAP7_75t_R FILLER_0_16_1182 ();
 FILLER_ASAP7_75t_R FILLER_0_16_1190 ();
 FILLER_ASAP7_75t_R FILLER_0_16_1198 ();
 DECAPx1_ASAP7_75t_R FILLER_0_16_1206 ();
 FILLER_ASAP7_75t_R FILLER_0_16_1218 ();
 FILLER_ASAP7_75t_R FILLER_0_16_1228 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_1236 ();
 FILLER_ASAP7_75t_R FILLER_0_16_1248 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_1256 ();
 FILLER_ASAP7_75t_R FILLER_0_16_1262 ();
 FILLER_ASAP7_75t_R FILLER_0_16_1270 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_1278 ();
 FILLER_ASAP7_75t_R FILLER_0_16_1284 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_1292 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_1298 ();
 FILLER_ASAP7_75t_R FILLER_0_16_1319 ();
 FILLER_ASAP7_75t_R FILLER_0_16_1324 ();
 DECAPx4_ASAP7_75t_R FILLER_0_16_1332 ();
 FILLER_ASAP7_75t_R FILLER_0_16_1348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_1356 ();
 DECAPx1_ASAP7_75t_R FILLER_0_16_1378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_68 ();
 DECAPx2_ASAP7_75t_R FILLER_0_17_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_104 ();
 DECAPx1_ASAP7_75t_R FILLER_0_17_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_119 ();
 FILLER_ASAP7_75t_R FILLER_0_17_128 ();
 DECAPx2_ASAP7_75t_R FILLER_0_17_136 ();
 FILLER_ASAP7_75t_R FILLER_0_17_142 ();
 FILLER_ASAP7_75t_R FILLER_0_17_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_152 ();
 DECAPx2_ASAP7_75t_R FILLER_0_17_160 ();
 FILLER_ASAP7_75t_R FILLER_0_17_166 ();
 FILLER_ASAP7_75t_R FILLER_0_17_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_177 ();
 FILLER_ASAP7_75t_R FILLER_0_17_184 ();
 DECAPx2_ASAP7_75t_R FILLER_0_17_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_198 ();
 FILLER_ASAP7_75t_R FILLER_0_17_209 ();
 FILLER_ASAP7_75t_R FILLER_0_17_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_216 ();
 FILLER_ASAP7_75t_R FILLER_0_17_232 ();
 FILLER_ASAP7_75t_R FILLER_0_17_240 ();
 FILLER_ASAP7_75t_R FILLER_0_17_248 ();
 DECAPx2_ASAP7_75t_R FILLER_0_17_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_263 ();
 FILLER_ASAP7_75t_R FILLER_0_17_270 ();
 DECAPx1_ASAP7_75t_R FILLER_0_17_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_289 ();
 DECAPx4_ASAP7_75t_R FILLER_0_17_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_321 ();
 DECAPx6_ASAP7_75t_R FILLER_0_17_334 ();
 DECAPx1_ASAP7_75t_R FILLER_0_17_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_352 ();
 FILLER_ASAP7_75t_R FILLER_0_17_359 ();
 FILLER_ASAP7_75t_R FILLER_0_17_367 ();
 FILLER_ASAP7_75t_R FILLER_0_17_375 ();
 FILLER_ASAP7_75t_R FILLER_0_17_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_385 ();
 FILLER_ASAP7_75t_R FILLER_0_17_396 ();
 FILLER_ASAP7_75t_R FILLER_0_17_404 ();
 DECAPx6_ASAP7_75t_R FILLER_0_17_414 ();
 FILLER_ASAP7_75t_R FILLER_0_17_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_430 ();
 DECAPx2_ASAP7_75t_R FILLER_0_17_437 ();
 FILLER_ASAP7_75t_R FILLER_0_17_443 ();
 DECAPx4_ASAP7_75t_R FILLER_0_17_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_461 ();
 FILLER_ASAP7_75t_R FILLER_0_17_472 ();
 DECAPx4_ASAP7_75t_R FILLER_0_17_481 ();
 FILLER_ASAP7_75t_R FILLER_0_17_498 ();
 DECAPx2_ASAP7_75t_R FILLER_0_17_510 ();
 FILLER_ASAP7_75t_R FILLER_0_17_516 ();
 DECAPx1_ASAP7_75t_R FILLER_0_17_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_528 ();
 FILLER_ASAP7_75t_R FILLER_0_17_535 ();
 FILLER_ASAP7_75t_R FILLER_0_17_547 ();
 FILLER_ASAP7_75t_R FILLER_0_17_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_569 ();
 FILLER_ASAP7_75t_R FILLER_0_17_591 ();
 DECAPx2_ASAP7_75t_R FILLER_0_17_599 ();
 FILLER_ASAP7_75t_R FILLER_0_17_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_607 ();
 FILLER_ASAP7_75t_R FILLER_0_17_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_615 ();
 FILLER_ASAP7_75t_R FILLER_0_17_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_629 ();
 FILLER_ASAP7_75t_R FILLER_0_17_638 ();
 FILLER_ASAP7_75t_R FILLER_0_17_647 ();
 DECAPx2_ASAP7_75t_R FILLER_0_17_652 ();
 FILLER_ASAP7_75t_R FILLER_0_17_664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_684 ();
 DECAPx4_ASAP7_75t_R FILLER_0_17_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_722 ();
 DECAPx6_ASAP7_75t_R FILLER_0_17_744 ();
 DECAPx1_ASAP7_75t_R FILLER_0_17_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_762 ();
 FILLER_ASAP7_75t_R FILLER_0_17_766 ();
 DECAPx6_ASAP7_75t_R FILLER_0_17_780 ();
 FILLER_ASAP7_75t_R FILLER_0_17_794 ();
 DECAPx2_ASAP7_75t_R FILLER_0_17_804 ();
 FILLER_ASAP7_75t_R FILLER_0_17_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_812 ();
 DECAPx6_ASAP7_75t_R FILLER_0_17_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_839 ();
 DECAPx1_ASAP7_75t_R FILLER_0_17_850 ();
 DECAPx1_ASAP7_75t_R FILLER_0_17_864 ();
 FILLER_ASAP7_75t_R FILLER_0_17_878 ();
 FILLER_ASAP7_75t_R FILLER_0_17_890 ();
 FILLER_ASAP7_75t_R FILLER_0_17_900 ();
 FILLER_ASAP7_75t_R FILLER_0_17_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_909 ();
 DECAPx1_ASAP7_75t_R FILLER_0_17_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_924 ();
 FILLER_ASAP7_75t_R FILLER_0_17_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_929 ();
 FILLER_ASAP7_75t_R FILLER_0_17_938 ();
 DECAPx2_ASAP7_75t_R FILLER_0_17_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_951 ();
 FILLER_ASAP7_75t_R FILLER_0_17_958 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_990 ();
 DECAPx1_ASAP7_75t_R FILLER_0_17_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_1015 ();
 DECAPx4_ASAP7_75t_R FILLER_0_17_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_1029 ();
 FILLER_ASAP7_75t_R FILLER_0_17_1036 ();
 FILLER_ASAP7_75t_R FILLER_0_17_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_1046 ();
 DECAPx1_ASAP7_75t_R FILLER_0_17_1053 ();
 DECAPx1_ASAP7_75t_R FILLER_0_17_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_1071 ();
 FILLER_ASAP7_75t_R FILLER_0_17_1090 ();
 FILLER_ASAP7_75t_R FILLER_0_17_1102 ();
 FILLER_ASAP7_75t_R FILLER_0_17_1114 ();
 FILLER_ASAP7_75t_R FILLER_0_17_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_1132 ();
 DECAPx4_ASAP7_75t_R FILLER_0_17_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_1164 ();
 DECAPx2_ASAP7_75t_R FILLER_0_17_1173 ();
 FILLER_ASAP7_75t_R FILLER_0_17_1185 ();
 FILLER_ASAP7_75t_R FILLER_0_17_1193 ();
 FILLER_ASAP7_75t_R FILLER_0_17_1203 ();
 DECAPx2_ASAP7_75t_R FILLER_0_17_1210 ();
 FILLER_ASAP7_75t_R FILLER_0_17_1232 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_1234 ();
 FILLER_ASAP7_75t_R FILLER_0_17_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_1249 ();
 FILLER_ASAP7_75t_R FILLER_0_17_1277 ();
 FILLER_ASAP7_75t_R FILLER_0_17_1285 ();
 DECAPx6_ASAP7_75t_R FILLER_0_17_1298 ();
 FILLER_ASAP7_75t_R FILLER_0_17_1312 ();
 DECAPx1_ASAP7_75t_R FILLER_0_17_1322 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_1326 ();
 DECAPx1_ASAP7_75t_R FILLER_0_17_1335 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_1339 ();
 FILLER_ASAP7_75t_R FILLER_0_17_1346 ();
 DECAPx2_ASAP7_75t_R FILLER_0_17_1354 ();
 DECAPx6_ASAP7_75t_R FILLER_0_17_1366 ();
 FILLER_ASAP7_75t_R FILLER_0_17_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_46 ();
 DECAPx4_ASAP7_75t_R FILLER_0_18_68 ();
 FILLER_ASAP7_75t_R FILLER_0_18_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_80 ();
 FILLER_ASAP7_75t_R FILLER_0_18_89 ();
 FILLER_ASAP7_75t_R FILLER_0_18_96 ();
 FILLER_ASAP7_75t_R FILLER_0_18_108 ();
 FILLER_ASAP7_75t_R FILLER_0_18_118 ();
 DECAPx1_ASAP7_75t_R FILLER_0_18_126 ();
 FILLER_ASAP7_75t_R FILLER_0_18_136 ();
 FILLER_ASAP7_75t_R FILLER_0_18_144 ();
 FILLER_ASAP7_75t_R FILLER_0_18_152 ();
 DECAPx1_ASAP7_75t_R FILLER_0_18_160 ();
 FILLER_ASAP7_75t_R FILLER_0_18_170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_179 ();
 DECAPx6_ASAP7_75t_R FILLER_0_18_201 ();
 DECAPx2_ASAP7_75t_R FILLER_0_18_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_221 ();
 DECAPx4_ASAP7_75t_R FILLER_0_18_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_242 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_249 ();
 DECAPx4_ASAP7_75t_R FILLER_0_18_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_281 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_292 ();
 DECAPx2_ASAP7_75t_R FILLER_0_18_314 ();
 FILLER_ASAP7_75t_R FILLER_0_18_326 ();
 FILLER_ASAP7_75t_R FILLER_0_18_338 ();
 DECAPx4_ASAP7_75t_R FILLER_0_18_346 ();
 FILLER_ASAP7_75t_R FILLER_0_18_356 ();
 FILLER_ASAP7_75t_R FILLER_0_18_364 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_372 ();
 DECAPx6_ASAP7_75t_R FILLER_0_18_394 ();
 FILLER_ASAP7_75t_R FILLER_0_18_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_410 ();
 FILLER_ASAP7_75t_R FILLER_0_18_421 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_431 ();
 DECAPx2_ASAP7_75t_R FILLER_0_18_453 ();
 FILLER_ASAP7_75t_R FILLER_0_18_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_461 ();
 DECAPx2_ASAP7_75t_R FILLER_0_18_464 ();
 FILLER_ASAP7_75t_R FILLER_0_18_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_472 ();
 DECAPx2_ASAP7_75t_R FILLER_0_18_485 ();
 FILLER_ASAP7_75t_R FILLER_0_18_491 ();
 DECAPx6_ASAP7_75t_R FILLER_0_18_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_519 ();
 DECAPx6_ASAP7_75t_R FILLER_0_18_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_540 ();
 DECAPx6_ASAP7_75t_R FILLER_0_18_563 ();
 FILLER_ASAP7_75t_R FILLER_0_18_577 ();
 FILLER_ASAP7_75t_R FILLER_0_18_600 ();
 DECAPx1_ASAP7_75t_R FILLER_0_18_613 ();
 DECAPx1_ASAP7_75t_R FILLER_0_18_629 ();
 FILLER_ASAP7_75t_R FILLER_0_18_641 ();
 FILLER_ASAP7_75t_R FILLER_0_18_649 ();
 DECAPx6_ASAP7_75t_R FILLER_0_18_661 ();
 DECAPx2_ASAP7_75t_R FILLER_0_18_687 ();
 FILLER_ASAP7_75t_R FILLER_0_18_693 ();
 DECAPx4_ASAP7_75t_R FILLER_0_18_703 ();
 FILLER_ASAP7_75t_R FILLER_0_18_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_715 ();
 DECAPx6_ASAP7_75t_R FILLER_0_18_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_740 ();
 FILLER_ASAP7_75t_R FILLER_0_18_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_749 ();
 DECAPx6_ASAP7_75t_R FILLER_0_18_761 ();
 DECAPx1_ASAP7_75t_R FILLER_0_18_775 ();
 FILLER_ASAP7_75t_R FILLER_0_18_790 ();
 FILLER_ASAP7_75t_R FILLER_0_18_798 ();
 DECAPx6_ASAP7_75t_R FILLER_0_18_821 ();
 DECAPx1_ASAP7_75t_R FILLER_0_18_835 ();
 FILLER_ASAP7_75t_R FILLER_0_18_849 ();
 FILLER_ASAP7_75t_R FILLER_0_18_861 ();
 FILLER_ASAP7_75t_R FILLER_0_18_873 ();
 FILLER_ASAP7_75t_R FILLER_0_18_885 ();
 FILLER_ASAP7_75t_R FILLER_0_18_897 ();
 DECAPx1_ASAP7_75t_R FILLER_0_18_904 ();
 FILLER_ASAP7_75t_R FILLER_0_18_913 ();
 FILLER_ASAP7_75t_R FILLER_0_18_921 ();
 DECAPx1_ASAP7_75t_R FILLER_0_18_933 ();
 FILLER_ASAP7_75t_R FILLER_0_18_947 ();
 DECAPx2_ASAP7_75t_R FILLER_0_18_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_960 ();
 DECAPx1_ASAP7_75t_R FILLER_0_18_967 ();
 DECAPx6_ASAP7_75t_R FILLER_0_18_977 ();
 DECAPx1_ASAP7_75t_R FILLER_0_18_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_995 ();
 FILLER_ASAP7_75t_R FILLER_0_18_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_1008 ();
 FILLER_ASAP7_75t_R FILLER_0_18_1015 ();
 DECAPx4_ASAP7_75t_R FILLER_0_18_1023 ();
 FILLER_ASAP7_75t_R FILLER_0_18_1039 ();
 FILLER_ASAP7_75t_R FILLER_0_18_1048 ();
 FILLER_ASAP7_75t_R FILLER_0_18_1053 ();
 FILLER_ASAP7_75t_R FILLER_0_18_1065 ();
 FILLER_ASAP7_75t_R FILLER_0_18_1077 ();
 FILLER_ASAP7_75t_R FILLER_0_18_1089 ();
 FILLER_ASAP7_75t_R FILLER_0_18_1101 ();
 DECAPx1_ASAP7_75t_R FILLER_0_18_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_1117 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_1138 ();
 FILLER_ASAP7_75t_R FILLER_0_18_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_1162 ();
 FILLER_ASAP7_75t_R FILLER_0_18_1169 ();
 DECAPx1_ASAP7_75t_R FILLER_0_18_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_1181 ();
 DECAPx1_ASAP7_75t_R FILLER_0_18_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_1192 ();
 FILLER_ASAP7_75t_R FILLER_0_18_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_1211 ();
 DECAPx6_ASAP7_75t_R FILLER_0_18_1218 ();
 FILLER_ASAP7_75t_R FILLER_0_18_1238 ();
 FILLER_ASAP7_75t_R FILLER_0_18_1246 ();
 DECAPx6_ASAP7_75t_R FILLER_0_18_1254 ();
 FILLER_ASAP7_75t_R FILLER_0_18_1268 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_1270 ();
 FILLER_ASAP7_75t_R FILLER_0_18_1279 ();
 FILLER_ASAP7_75t_R FILLER_0_18_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_1288 ();
 DECAPx6_ASAP7_75t_R FILLER_0_18_1295 ();
 FILLER_ASAP7_75t_R FILLER_0_18_1315 ();
 DECAPx1_ASAP7_75t_R FILLER_0_18_1323 ();
 DECAPx2_ASAP7_75t_R FILLER_0_18_1333 ();
 FILLER_ASAP7_75t_R FILLER_0_18_1339 ();
 FILLER_ASAP7_75t_R FILLER_0_18_1347 ();
 DECAPx4_ASAP7_75t_R FILLER_0_18_1355 ();
 FILLER_ASAP7_75t_R FILLER_0_18_1371 ();
 FILLER_ASAP7_75t_R FILLER_0_18_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_24 ();
 DECAPx6_ASAP7_75t_R FILLER_0_19_46 ();
 FILLER_ASAP7_75t_R FILLER_0_19_60 ();
 FILLER_ASAP7_75t_R FILLER_0_19_68 ();
 DECAPx1_ASAP7_75t_R FILLER_0_19_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_82 ();
 FILLER_ASAP7_75t_R FILLER_0_19_89 ();
 FILLER_ASAP7_75t_R FILLER_0_19_99 ();
 DECAPx1_ASAP7_75t_R FILLER_0_19_111 ();
 FILLER_ASAP7_75t_R FILLER_0_19_121 ();
 FILLER_ASAP7_75t_R FILLER_0_19_129 ();
 FILLER_ASAP7_75t_R FILLER_0_19_136 ();
 FILLER_ASAP7_75t_R FILLER_0_19_144 ();
 FILLER_ASAP7_75t_R FILLER_0_19_151 ();
 DECAPx1_ASAP7_75t_R FILLER_0_19_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_167 ();
 FILLER_ASAP7_75t_R FILLER_0_19_174 ();
 FILLER_ASAP7_75t_R FILLER_0_19_184 ();
 DECAPx6_ASAP7_75t_R FILLER_0_19_206 ();
 DECAPx1_ASAP7_75t_R FILLER_0_19_220 ();
 FILLER_ASAP7_75t_R FILLER_0_19_232 ();
 FILLER_ASAP7_75t_R FILLER_0_19_240 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_258 ();
 DECAPx1_ASAP7_75t_R FILLER_0_19_280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_294 ();
 DECAPx2_ASAP7_75t_R FILLER_0_19_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_322 ();
 FILLER_ASAP7_75t_R FILLER_0_19_329 ();
 DECAPx2_ASAP7_75t_R FILLER_0_19_337 ();
 FILLER_ASAP7_75t_R FILLER_0_19_343 ();
 DECAPx1_ASAP7_75t_R FILLER_0_19_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_357 ();
 DECAPx2_ASAP7_75t_R FILLER_0_19_364 ();
 FILLER_ASAP7_75t_R FILLER_0_19_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_372 ();
 DECAPx4_ASAP7_75t_R FILLER_0_19_379 ();
 FILLER_ASAP7_75t_R FILLER_0_19_389 ();
 FILLER_ASAP7_75t_R FILLER_0_19_399 ();
 DECAPx4_ASAP7_75t_R FILLER_0_19_411 ();
 FILLER_ASAP7_75t_R FILLER_0_19_427 ();
 FILLER_ASAP7_75t_R FILLER_0_19_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_437 ();
 FILLER_ASAP7_75t_R FILLER_0_19_444 ();
 FILLER_ASAP7_75t_R FILLER_0_19_452 ();
 FILLER_ASAP7_75t_R FILLER_0_19_462 ();
 FILLER_ASAP7_75t_R FILLER_0_19_470 ();
 DECAPx6_ASAP7_75t_R FILLER_0_19_478 ();
 DECAPx1_ASAP7_75t_R FILLER_0_19_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_496 ();
 FILLER_ASAP7_75t_R FILLER_0_19_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_505 ();
 FILLER_ASAP7_75t_R FILLER_0_19_526 ();
 DECAPx4_ASAP7_75t_R FILLER_0_19_531 ();
 FILLER_ASAP7_75t_R FILLER_0_19_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_549 ();
 FILLER_ASAP7_75t_R FILLER_0_19_556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_564 ();
 DECAPx2_ASAP7_75t_R FILLER_0_19_586 ();
 FILLER_ASAP7_75t_R FILLER_0_19_592 ();
 FILLER_ASAP7_75t_R FILLER_0_19_597 ();
 DECAPx2_ASAP7_75t_R FILLER_0_19_609 ();
 FILLER_ASAP7_75t_R FILLER_0_19_627 ();
 DECAPx2_ASAP7_75t_R FILLER_0_19_636 ();
 DECAPx1_ASAP7_75t_R FILLER_0_19_652 ();
 FILLER_ASAP7_75t_R FILLER_0_19_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_666 ();
 FILLER_ASAP7_75t_R FILLER_0_19_673 ();
 DECAPx6_ASAP7_75t_R FILLER_0_19_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_695 ();
 DECAPx1_ASAP7_75t_R FILLER_0_19_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_708 ();
 DECAPx2_ASAP7_75t_R FILLER_0_19_720 ();
 FILLER_ASAP7_75t_R FILLER_0_19_726 ();
 FILLER_ASAP7_75t_R FILLER_0_19_734 ();
 DECAPx6_ASAP7_75t_R FILLER_0_19_742 ();
 DECAPx1_ASAP7_75t_R FILLER_0_19_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_766 ();
 DECAPx1_ASAP7_75t_R FILLER_0_19_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_792 ();
 FILLER_ASAP7_75t_R FILLER_0_19_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_801 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_805 ();
 FILLER_ASAP7_75t_R FILLER_0_19_832 ();
 DECAPx1_ASAP7_75t_R FILLER_0_19_844 ();
 FILLER_ASAP7_75t_R FILLER_0_19_855 ();
 FILLER_ASAP7_75t_R FILLER_0_19_867 ();
 FILLER_ASAP7_75t_R FILLER_0_19_879 ();
 FILLER_ASAP7_75t_R FILLER_0_19_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_893 ();
 FILLER_ASAP7_75t_R FILLER_0_19_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_902 ();
 FILLER_ASAP7_75t_R FILLER_0_19_911 ();
 FILLER_ASAP7_75t_R FILLER_0_19_923 ();
 DECAPx1_ASAP7_75t_R FILLER_0_19_927 ();
 FILLER_ASAP7_75t_R FILLER_0_19_937 ();
 DECAPx1_ASAP7_75t_R FILLER_0_19_945 ();
 DECAPx4_ASAP7_75t_R FILLER_0_19_959 ();
 FILLER_ASAP7_75t_R FILLER_0_19_975 ();
 FILLER_ASAP7_75t_R FILLER_0_19_984 ();
 FILLER_ASAP7_75t_R FILLER_0_19_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_994 ();
 DECAPx4_ASAP7_75t_R FILLER_0_19_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_1011 ();
 FILLER_ASAP7_75t_R FILLER_0_19_1018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_1025 ();
 DECAPx6_ASAP7_75t_R FILLER_0_19_1047 ();
 FILLER_ASAP7_75t_R FILLER_0_19_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_1073 ();
 FILLER_ASAP7_75t_R FILLER_0_19_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_1086 ();
 FILLER_ASAP7_75t_R FILLER_0_19_1095 ();
 FILLER_ASAP7_75t_R FILLER_0_19_1115 ();
 FILLER_ASAP7_75t_R FILLER_0_19_1123 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_1130 ();
 DECAPx6_ASAP7_75t_R FILLER_0_19_1152 ();
 FILLER_ASAP7_75t_R FILLER_0_19_1171 ();
 FILLER_ASAP7_75t_R FILLER_0_19_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_1182 ();
 DECAPx4_ASAP7_75t_R FILLER_0_19_1193 ();
 FILLER_ASAP7_75t_R FILLER_0_19_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_1213 ();
 DECAPx1_ASAP7_75t_R FILLER_0_19_1235 ();
 FILLER_ASAP7_75t_R FILLER_0_19_1244 ();
 FILLER_ASAP7_75t_R FILLER_0_19_1252 ();
 FILLER_ASAP7_75t_R FILLER_0_19_1260 ();
 FILLER_ASAP7_75t_R FILLER_0_19_1268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_19_1276 ();
 DECAPx1_ASAP7_75t_R FILLER_0_19_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_1294 ();
 DECAPx6_ASAP7_75t_R FILLER_0_19_1305 ();
 FILLER_ASAP7_75t_R FILLER_0_19_1319 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_1321 ();
 FILLER_ASAP7_75t_R FILLER_0_19_1328 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_1335 ();
 FILLER_ASAP7_75t_R FILLER_0_19_1357 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_1359 ();
 FILLER_ASAP7_75t_R FILLER_0_19_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_19_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_20_24 ();
 FILLER_ASAP7_75t_R FILLER_0_20_44 ();
 FILLER_ASAP7_75t_R FILLER_0_20_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_54 ();
 DECAPx4_ASAP7_75t_R FILLER_0_20_61 ();
 FILLER_ASAP7_75t_R FILLER_0_20_77 ();
 FILLER_ASAP7_75t_R FILLER_0_20_86 ();
 DECAPx2_ASAP7_75t_R FILLER_0_20_94 ();
 FILLER_ASAP7_75t_R FILLER_0_20_100 ();
 FILLER_ASAP7_75t_R FILLER_0_20_108 ();
 FILLER_ASAP7_75t_R FILLER_0_20_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_122 ();
 DECAPx1_ASAP7_75t_R FILLER_0_20_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_133 ();
 FILLER_ASAP7_75t_R FILLER_0_20_140 ();
 DECAPx1_ASAP7_75t_R FILLER_0_20_148 ();
 DECAPx1_ASAP7_75t_R FILLER_0_20_160 ();
 FILLER_ASAP7_75t_R FILLER_0_20_170 ();
 FILLER_ASAP7_75t_R FILLER_0_20_178 ();
 FILLER_ASAP7_75t_R FILLER_0_20_186 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_194 ();
 DECAPx2_ASAP7_75t_R FILLER_0_20_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_222 ();
 FILLER_ASAP7_75t_R FILLER_0_20_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_233 ();
 FILLER_ASAP7_75t_R FILLER_0_20_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_242 ();
 FILLER_ASAP7_75t_R FILLER_0_20_250 ();
 FILLER_ASAP7_75t_R FILLER_0_20_272 ();
 DECAPx1_ASAP7_75t_R FILLER_0_20_277 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_287 ();
 DECAPx4_ASAP7_75t_R FILLER_0_20_309 ();
 DECAPx1_ASAP7_75t_R FILLER_0_20_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_335 ();
 FILLER_ASAP7_75t_R FILLER_0_20_344 ();
 DECAPx2_ASAP7_75t_R FILLER_0_20_352 ();
 DECAPx2_ASAP7_75t_R FILLER_0_20_365 ();
 DECAPx4_ASAP7_75t_R FILLER_0_20_377 ();
 FILLER_ASAP7_75t_R FILLER_0_20_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_389 ();
 DECAPx2_ASAP7_75t_R FILLER_0_20_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_404 ();
 FILLER_ASAP7_75t_R FILLER_0_20_415 ();
 FILLER_ASAP7_75t_R FILLER_0_20_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_429 ();
 FILLER_ASAP7_75t_R FILLER_0_20_436 ();
 DECAPx1_ASAP7_75t_R FILLER_0_20_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_449 ();
 FILLER_ASAP7_75t_R FILLER_0_20_460 ();
 DECAPx2_ASAP7_75t_R FILLER_0_20_464 ();
 FILLER_ASAP7_75t_R FILLER_0_20_470 ();
 FILLER_ASAP7_75t_R FILLER_0_20_478 ();
 DECAPx2_ASAP7_75t_R FILLER_0_20_486 ();
 FILLER_ASAP7_75t_R FILLER_0_20_492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_20_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_520 ();
 FILLER_ASAP7_75t_R FILLER_0_20_527 ();
 DECAPx2_ASAP7_75t_R FILLER_0_20_535 ();
 FILLER_ASAP7_75t_R FILLER_0_20_547 ();
 DECAPx4_ASAP7_75t_R FILLER_0_20_557 ();
 FILLER_ASAP7_75t_R FILLER_0_20_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_569 ();
 FILLER_ASAP7_75t_R FILLER_0_20_573 ();
 DECAPx4_ASAP7_75t_R FILLER_0_20_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_595 ();
 FILLER_ASAP7_75t_R FILLER_0_20_608 ();
 DECAPx1_ASAP7_75t_R FILLER_0_20_622 ();
 FILLER_ASAP7_75t_R FILLER_0_20_632 ();
 FILLER_ASAP7_75t_R FILLER_0_20_640 ();
 DECAPx2_ASAP7_75t_R FILLER_0_20_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_654 ();
 FILLER_ASAP7_75t_R FILLER_0_20_665 ();
 FILLER_ASAP7_75t_R FILLER_0_20_675 ();
 DECAPx1_ASAP7_75t_R FILLER_0_20_689 ();
 DECAPx6_ASAP7_75t_R FILLER_0_20_699 ();
 DECAPx1_ASAP7_75t_R FILLER_0_20_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_717 ();
 FILLER_ASAP7_75t_R FILLER_0_20_724 ();
 FILLER_ASAP7_75t_R FILLER_0_20_732 ();
 FILLER_ASAP7_75t_R FILLER_0_20_742 ();
 FILLER_ASAP7_75t_R FILLER_0_20_752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_20_766 ();
 FILLER_ASAP7_75t_R FILLER_0_20_772 ();
 FILLER_ASAP7_75t_R FILLER_0_20_786 ();
 FILLER_ASAP7_75t_R FILLER_0_20_800 ();
 DECAPx6_ASAP7_75t_R FILLER_0_20_823 ();
 FILLER_ASAP7_75t_R FILLER_0_20_837 ();
 FILLER_ASAP7_75t_R FILLER_0_20_849 ();
 DECAPx1_ASAP7_75t_R FILLER_0_20_861 ();
 FILLER_ASAP7_75t_R FILLER_0_20_875 ();
 FILLER_ASAP7_75t_R FILLER_0_20_887 ();
 DECAPx2_ASAP7_75t_R FILLER_0_20_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_901 ();
 DECAPx2_ASAP7_75t_R FILLER_0_20_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_928 ();
 FILLER_ASAP7_75t_R FILLER_0_20_940 ();
 DECAPx6_ASAP7_75t_R FILLER_0_20_947 ();
 DECAPx1_ASAP7_75t_R FILLER_0_20_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_965 ();
 DECAPx2_ASAP7_75t_R FILLER_0_20_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_975 ();
 FILLER_ASAP7_75t_R FILLER_0_20_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_984 ();
 DECAPx1_ASAP7_75t_R FILLER_0_20_1005 ();
 DECAPx2_ASAP7_75t_R FILLER_0_20_1019 ();
 DECAPx1_ASAP7_75t_R FILLER_0_20_1036 ();
 FILLER_ASAP7_75t_R FILLER_0_20_1044 ();
 FILLER_ASAP7_75t_R FILLER_0_20_1056 ();
 FILLER_ASAP7_75t_R FILLER_0_20_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_1066 ();
 FILLER_ASAP7_75t_R FILLER_0_20_1072 ();
 FILLER_ASAP7_75t_R FILLER_0_20_1080 ();
 FILLER_ASAP7_75t_R FILLER_0_20_1090 ();
 DECAPx2_ASAP7_75t_R FILLER_0_20_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_1104 ();
 FILLER_ASAP7_75t_R FILLER_0_20_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_1123 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_1145 ();
 DECAPx1_ASAP7_75t_R FILLER_0_20_1167 ();
 FILLER_ASAP7_75t_R FILLER_0_20_1177 ();
 FILLER_ASAP7_75t_R FILLER_0_20_1185 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_1187 ();
 FILLER_ASAP7_75t_R FILLER_0_20_1194 ();
 DECAPx2_ASAP7_75t_R FILLER_0_20_1202 ();
 FILLER_ASAP7_75t_R FILLER_0_20_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_1210 ();
 DECAPx4_ASAP7_75t_R FILLER_0_20_1217 ();
 FILLER_ASAP7_75t_R FILLER_0_20_1227 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_1229 ();
 DECAPx6_ASAP7_75t_R FILLER_0_20_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_1256 ();
 DECAPx4_ASAP7_75t_R FILLER_0_20_1278 ();
 FILLER_ASAP7_75t_R FILLER_0_20_1294 ();
 FILLER_ASAP7_75t_R FILLER_0_20_1302 ();
 DECAPx4_ASAP7_75t_R FILLER_0_20_1310 ();
 FILLER_ASAP7_75t_R FILLER_0_20_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_1327 ();
 DECAPx4_ASAP7_75t_R FILLER_0_20_1349 ();
 FILLER_ASAP7_75t_R FILLER_0_20_1359 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_1361 ();
 FILLER_ASAP7_75t_R FILLER_0_20_1368 ();
 DECAPx2_ASAP7_75t_R FILLER_0_20_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_21_24 ();
 FILLER_ASAP7_75t_R FILLER_0_21_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_40 ();
 FILLER_ASAP7_75t_R FILLER_0_21_47 ();
 FILLER_ASAP7_75t_R FILLER_0_21_55 ();
 DECAPx2_ASAP7_75t_R FILLER_0_21_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_69 ();
 FILLER_ASAP7_75t_R FILLER_0_21_76 ();
 DECAPx1_ASAP7_75t_R FILLER_0_21_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_89 ();
 FILLER_ASAP7_75t_R FILLER_0_21_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_100 ();
 FILLER_ASAP7_75t_R FILLER_0_21_108 ();
 FILLER_ASAP7_75t_R FILLER_0_21_113 ();
 FILLER_ASAP7_75t_R FILLER_0_21_125 ();
 FILLER_ASAP7_75t_R FILLER_0_21_133 ();
 DECAPx2_ASAP7_75t_R FILLER_0_21_140 ();
 FILLER_ASAP7_75t_R FILLER_0_21_146 ();
 FILLER_ASAP7_75t_R FILLER_0_21_154 ();
 DECAPx6_ASAP7_75t_R FILLER_0_21_166 ();
 FILLER_ASAP7_75t_R FILLER_0_21_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_182 ();
 DECAPx4_ASAP7_75t_R FILLER_0_21_189 ();
 FILLER_ASAP7_75t_R FILLER_0_21_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_201 ();
 FILLER_ASAP7_75t_R FILLER_0_21_208 ();
 FILLER_ASAP7_75t_R FILLER_0_21_216 ();
 DECAPx6_ASAP7_75t_R FILLER_0_21_223 ();
 DECAPx1_ASAP7_75t_R FILLER_0_21_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_241 ();
 DECAPx2_ASAP7_75t_R FILLER_0_21_248 ();
 FILLER_ASAP7_75t_R FILLER_0_21_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_266 ();
 FILLER_ASAP7_75t_R FILLER_0_21_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_287 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_309 ();
 FILLER_ASAP7_75t_R FILLER_0_21_331 ();
 FILLER_ASAP7_75t_R FILLER_0_21_339 ();
 FILLER_ASAP7_75t_R FILLER_0_21_346 ();
 FILLER_ASAP7_75t_R FILLER_0_21_354 ();
 DECAPx1_ASAP7_75t_R FILLER_0_21_362 ();
 DECAPx2_ASAP7_75t_R FILLER_0_21_369 ();
 DECAPx1_ASAP7_75t_R FILLER_0_21_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_385 ();
 FILLER_ASAP7_75t_R FILLER_0_21_392 ();
 FILLER_ASAP7_75t_R FILLER_0_21_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_404 ();
 DECAPx2_ASAP7_75t_R FILLER_0_21_415 ();
 DECAPx2_ASAP7_75t_R FILLER_0_21_431 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_443 ();
 DECAPx1_ASAP7_75t_R FILLER_0_21_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_469 ();
 FILLER_ASAP7_75t_R FILLER_0_21_476 ();
 FILLER_ASAP7_75t_R FILLER_0_21_486 ();
 FILLER_ASAP7_75t_R FILLER_0_21_494 ();
 DECAPx2_ASAP7_75t_R FILLER_0_21_508 ();
 FILLER_ASAP7_75t_R FILLER_0_21_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_516 ();
 FILLER_ASAP7_75t_R FILLER_0_21_523 ();
 DECAPx2_ASAP7_75t_R FILLER_0_21_532 ();
 DECAPx4_ASAP7_75t_R FILLER_0_21_558 ();
 DECAPx6_ASAP7_75t_R FILLER_0_21_578 ();
 FILLER_ASAP7_75t_R FILLER_0_21_592 ();
 FILLER_ASAP7_75t_R FILLER_0_21_615 ();
 DECAPx1_ASAP7_75t_R FILLER_0_21_629 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_644 ();
 DECAPx6_ASAP7_75t_R FILLER_0_21_672 ();
 FILLER_ASAP7_75t_R FILLER_0_21_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_688 ();
 FILLER_ASAP7_75t_R FILLER_0_21_695 ();
 DECAPx6_ASAP7_75t_R FILLER_0_21_703 ();
 DECAPx2_ASAP7_75t_R FILLER_0_21_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_723 ();
 DECAPx2_ASAP7_75t_R FILLER_0_21_727 ();
 FILLER_ASAP7_75t_R FILLER_0_21_733 ();
 FILLER_ASAP7_75t_R FILLER_0_21_743 ();
 DECAPx2_ASAP7_75t_R FILLER_0_21_748 ();
 FILLER_ASAP7_75t_R FILLER_0_21_754 ();
 FILLER_ASAP7_75t_R FILLER_0_21_778 ();
 DECAPx4_ASAP7_75t_R FILLER_0_21_792 ();
 FILLER_ASAP7_75t_R FILLER_0_21_802 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_807 ();
 DECAPx2_ASAP7_75t_R FILLER_0_21_829 ();
 FILLER_ASAP7_75t_R FILLER_0_21_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_837 ();
 FILLER_ASAP7_75t_R FILLER_0_21_842 ();
 DECAPx1_ASAP7_75t_R FILLER_0_21_849 ();
 FILLER_ASAP7_75t_R FILLER_0_21_858 ();
 FILLER_ASAP7_75t_R FILLER_0_21_870 ();
 FILLER_ASAP7_75t_R FILLER_0_21_882 ();
 FILLER_ASAP7_75t_R FILLER_0_21_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_894 ();
 FILLER_ASAP7_75t_R FILLER_0_21_902 ();
 FILLER_ASAP7_75t_R FILLER_0_21_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_913 ();
 DECAPx1_ASAP7_75t_R FILLER_0_21_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_924 ();
 DECAPx2_ASAP7_75t_R FILLER_0_21_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_933 ();
 DECAPx2_ASAP7_75t_R FILLER_0_21_940 ();
 FILLER_ASAP7_75t_R FILLER_0_21_946 ();
 DECAPx4_ASAP7_75t_R FILLER_0_21_955 ();
 FILLER_ASAP7_75t_R FILLER_0_21_972 ();
 DECAPx4_ASAP7_75t_R FILLER_0_21_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_990 ();
 FILLER_ASAP7_75t_R FILLER_0_21_997 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_1006 ();
 DECAPx6_ASAP7_75t_R FILLER_0_21_1013 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1027 ();
 DECAPx2_ASAP7_75t_R FILLER_0_21_1035 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1041 ();
 DECAPx2_ASAP7_75t_R FILLER_0_21_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_1059 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1067 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1075 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1083 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1088 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1096 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1110 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1118 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_1133 ();
 DECAPx6_ASAP7_75t_R FILLER_0_21_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_1169 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1176 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1184 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_1200 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1222 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_1224 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1228 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_1244 ();
 DECAPx2_ASAP7_75t_R FILLER_0_21_1266 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1272 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1290 ();
 DECAPx1_ASAP7_75t_R FILLER_0_21_1300 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1310 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1318 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1326 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1334 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1342 ();
 DECAPx4_ASAP7_75t_R FILLER_0_21_1350 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_21_1374 ();
 FILLER_ASAP7_75t_R FILLER_0_21_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_22_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_38 ();
 DECAPx4_ASAP7_75t_R FILLER_0_22_45 ();
 FILLER_ASAP7_75t_R FILLER_0_22_55 ();
 FILLER_ASAP7_75t_R FILLER_0_22_63 ();
 DECAPx6_ASAP7_75t_R FILLER_0_22_71 ();
 FILLER_ASAP7_75t_R FILLER_0_22_95 ();
 FILLER_ASAP7_75t_R FILLER_0_22_107 ();
 FILLER_ASAP7_75t_R FILLER_0_22_116 ();
 FILLER_ASAP7_75t_R FILLER_0_22_125 ();
 FILLER_ASAP7_75t_R FILLER_0_22_132 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_144 ();
 DECAPx4_ASAP7_75t_R FILLER_0_22_166 ();
 FILLER_ASAP7_75t_R FILLER_0_22_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_178 ();
 FILLER_ASAP7_75t_R FILLER_0_22_185 ();
 FILLER_ASAP7_75t_R FILLER_0_22_193 ();
 DECAPx2_ASAP7_75t_R FILLER_0_22_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_207 ();
 DECAPx4_ASAP7_75t_R FILLER_0_22_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_228 ();
 DECAPx2_ASAP7_75t_R FILLER_0_22_235 ();
 FILLER_ASAP7_75t_R FILLER_0_22_241 ();
 DECAPx4_ASAP7_75t_R FILLER_0_22_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_256 ();
 FILLER_ASAP7_75t_R FILLER_0_22_263 ();
 FILLER_ASAP7_75t_R FILLER_0_22_271 ();
 FILLER_ASAP7_75t_R FILLER_0_22_281 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_293 ();
 DECAPx6_ASAP7_75t_R FILLER_0_22_315 ();
 DECAPx2_ASAP7_75t_R FILLER_0_22_341 ();
 DECAPx2_ASAP7_75t_R FILLER_0_22_353 ();
 FILLER_ASAP7_75t_R FILLER_0_22_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_361 ();
 DECAPx6_ASAP7_75t_R FILLER_0_22_370 ();
 FILLER_ASAP7_75t_R FILLER_0_22_384 ();
 FILLER_ASAP7_75t_R FILLER_0_22_389 ();
 FILLER_ASAP7_75t_R FILLER_0_22_397 ();
 DECAPx2_ASAP7_75t_R FILLER_0_22_409 ();
 FILLER_ASAP7_75t_R FILLER_0_22_415 ();
 DECAPx2_ASAP7_75t_R FILLER_0_22_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_433 ();
 FILLER_ASAP7_75t_R FILLER_0_22_440 ();
 FILLER_ASAP7_75t_R FILLER_0_22_448 ();
 FILLER_ASAP7_75t_R FILLER_0_22_460 ();
 DECAPx1_ASAP7_75t_R FILLER_0_22_464 ();
 FILLER_ASAP7_75t_R FILLER_0_22_474 ();
 DECAPx2_ASAP7_75t_R FILLER_0_22_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_488 ();
 FILLER_ASAP7_75t_R FILLER_0_22_517 ();
 FILLER_ASAP7_75t_R FILLER_0_22_525 ();
 FILLER_ASAP7_75t_R FILLER_0_22_532 ();
 DECAPx2_ASAP7_75t_R FILLER_0_22_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_546 ();
 DECAPx1_ASAP7_75t_R FILLER_0_22_554 ();
 FILLER_ASAP7_75t_R FILLER_0_22_578 ();
 DECAPx4_ASAP7_75t_R FILLER_0_22_583 ();
 FILLER_ASAP7_75t_R FILLER_0_22_593 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_595 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_599 ();
 DECAPx6_ASAP7_75t_R FILLER_0_22_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_635 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_647 ();
 DECAPx4_ASAP7_75t_R FILLER_0_22_669 ();
 FILLER_ASAP7_75t_R FILLER_0_22_679 ();
 FILLER_ASAP7_75t_R FILLER_0_22_687 ();
 DECAPx1_ASAP7_75t_R FILLER_0_22_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_701 ();
 DECAPx6_ASAP7_75t_R FILLER_0_22_713 ();
 DECAPx2_ASAP7_75t_R FILLER_0_22_727 ();
 DECAPx6_ASAP7_75t_R FILLER_0_22_744 ();
 DECAPx2_ASAP7_75t_R FILLER_0_22_761 ();
 FILLER_ASAP7_75t_R FILLER_0_22_767 ();
 FILLER_ASAP7_75t_R FILLER_0_22_787 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_811 ();
 DECAPx6_ASAP7_75t_R FILLER_0_22_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_847 ();
 FILLER_ASAP7_75t_R FILLER_0_22_858 ();
 FILLER_ASAP7_75t_R FILLER_0_22_870 ();
 FILLER_ASAP7_75t_R FILLER_0_22_882 ();
 FILLER_ASAP7_75t_R FILLER_0_22_892 ();
 DECAPx1_ASAP7_75t_R FILLER_0_22_900 ();
 FILLER_ASAP7_75t_R FILLER_0_22_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_911 ();
 DECAPx6_ASAP7_75t_R FILLER_0_22_918 ();
 FILLER_ASAP7_75t_R FILLER_0_22_942 ();
 FILLER_ASAP7_75t_R FILLER_0_22_951 ();
 FILLER_ASAP7_75t_R FILLER_0_22_959 ();
 FILLER_ASAP7_75t_R FILLER_0_22_967 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_972 ();
 DECAPx1_ASAP7_75t_R FILLER_0_22_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_998 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_1041 ();
 FILLER_ASAP7_75t_R FILLER_0_22_1062 ();
 FILLER_ASAP7_75t_R FILLER_0_22_1072 ();
 FILLER_ASAP7_75t_R FILLER_0_22_1084 ();
 FILLER_ASAP7_75t_R FILLER_0_22_1096 ();
 DECAPx1_ASAP7_75t_R FILLER_0_22_1108 ();
 FILLER_ASAP7_75t_R FILLER_0_22_1119 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_1126 ();
 DECAPx4_ASAP7_75t_R FILLER_0_22_1148 ();
 DECAPx1_ASAP7_75t_R FILLER_0_22_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_1170 ();
 DECAPx2_ASAP7_75t_R FILLER_0_22_1176 ();
 DECAPx2_ASAP7_75t_R FILLER_0_22_1188 ();
 FILLER_ASAP7_75t_R FILLER_0_22_1194 ();
 DECAPx4_ASAP7_75t_R FILLER_0_22_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_1212 ();
 FILLER_ASAP7_75t_R FILLER_0_22_1220 ();
 FILLER_ASAP7_75t_R FILLER_0_22_1230 ();
 DECAPx1_ASAP7_75t_R FILLER_0_22_1238 ();
 DECAPx2_ASAP7_75t_R FILLER_0_22_1252 ();
 FILLER_ASAP7_75t_R FILLER_0_22_1258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_1266 ();
 FILLER_ASAP7_75t_R FILLER_0_22_1294 ();
 FILLER_ASAP7_75t_R FILLER_0_22_1302 ();
 DECAPx2_ASAP7_75t_R FILLER_0_22_1310 ();
 DECAPx1_ASAP7_75t_R FILLER_0_22_1326 ();
 FILLER_ASAP7_75t_R FILLER_0_22_1336 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_1338 ();
 FILLER_ASAP7_75t_R FILLER_0_22_1345 ();
 DECAPx2_ASAP7_75t_R FILLER_0_22_1355 ();
 FILLER_ASAP7_75t_R FILLER_0_22_1361 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_1363 ();
 DECAPx4_ASAP7_75t_R FILLER_0_22_1370 ();
 FILLER_ASAP7_75t_R FILLER_0_22_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_46 ();
 DECAPx1_ASAP7_75t_R FILLER_0_23_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_72 ();
 DECAPx1_ASAP7_75t_R FILLER_0_23_111 ();
 FILLER_ASAP7_75t_R FILLER_0_23_133 ();
 FILLER_ASAP7_75t_R FILLER_0_23_145 ();
 DECAPx2_ASAP7_75t_R FILLER_0_23_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_159 ();
 DECAPx1_ASAP7_75t_R FILLER_0_23_188 ();
 FILLER_ASAP7_75t_R FILLER_0_23_198 ();
 FILLER_ASAP7_75t_R FILLER_0_23_205 ();
 FILLER_ASAP7_75t_R FILLER_0_23_218 ();
 DECAPx1_ASAP7_75t_R FILLER_0_23_226 ();
 DECAPx1_ASAP7_75t_R FILLER_0_23_238 ();
 DECAPx2_ASAP7_75t_R FILLER_0_23_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_254 ();
 DECAPx6_ASAP7_75t_R FILLER_0_23_261 ();
 FILLER_ASAP7_75t_R FILLER_0_23_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_277 ();
 FILLER_ASAP7_75t_R FILLER_0_23_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_295 ();
 FILLER_ASAP7_75t_R FILLER_0_23_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_319 ();
 DECAPx2_ASAP7_75t_R FILLER_0_23_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_346 ();
 FILLER_ASAP7_75t_R FILLER_0_23_353 ();
 FILLER_ASAP7_75t_R FILLER_0_23_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_363 ();
 DECAPx4_ASAP7_75t_R FILLER_0_23_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_382 ();
 DECAPx2_ASAP7_75t_R FILLER_0_23_393 ();
 FILLER_ASAP7_75t_R FILLER_0_23_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_401 ();
 DECAPx1_ASAP7_75t_R FILLER_0_23_406 ();
 DECAPx2_ASAP7_75t_R FILLER_0_23_415 ();
 FILLER_ASAP7_75t_R FILLER_0_23_421 ();
 DECAPx4_ASAP7_75t_R FILLER_0_23_428 ();
 DECAPx2_ASAP7_75t_R FILLER_0_23_450 ();
 FILLER_ASAP7_75t_R FILLER_0_23_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_458 ();
 DECAPx4_ASAP7_75t_R FILLER_0_23_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_474 ();
 DECAPx1_ASAP7_75t_R FILLER_0_23_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_482 ();
 DECAPx2_ASAP7_75t_R FILLER_0_23_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_494 ();
 FILLER_ASAP7_75t_R FILLER_0_23_500 ();
 DECAPx4_ASAP7_75t_R FILLER_0_23_507 ();
 FILLER_ASAP7_75t_R FILLER_0_23_517 ();
 FILLER_ASAP7_75t_R FILLER_0_23_525 ();
 DECAPx1_ASAP7_75t_R FILLER_0_23_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_537 ();
 FILLER_ASAP7_75t_R FILLER_0_23_544 ();
 DECAPx6_ASAP7_75t_R FILLER_0_23_552 ();
 DECAPx1_ASAP7_75t_R FILLER_0_23_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_576 ();
 FILLER_ASAP7_75t_R FILLER_0_23_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_585 ();
 FILLER_ASAP7_75t_R FILLER_0_23_589 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_594 ();
 DECAPx4_ASAP7_75t_R FILLER_0_23_616 ();
 DECAPx2_ASAP7_75t_R FILLER_0_23_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_638 ();
 FILLER_ASAP7_75t_R FILLER_0_23_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_653 ();
 FILLER_ASAP7_75t_R FILLER_0_23_660 ();
 FILLER_ASAP7_75t_R FILLER_0_23_668 ();
 DECAPx2_ASAP7_75t_R FILLER_0_23_676 ();
 FILLER_ASAP7_75t_R FILLER_0_23_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_684 ();
 DECAPx1_ASAP7_75t_R FILLER_0_23_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_712 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_734 ();
 FILLER_ASAP7_75t_R FILLER_0_23_756 ();
 FILLER_ASAP7_75t_R FILLER_0_23_779 ();
 FILLER_ASAP7_75t_R FILLER_0_23_793 ();
 DECAPx4_ASAP7_75t_R FILLER_0_23_798 ();
 FILLER_ASAP7_75t_R FILLER_0_23_808 ();
 FILLER_ASAP7_75t_R FILLER_0_23_828 ();
 FILLER_ASAP7_75t_R FILLER_0_23_841 ();
 DECAPx1_ASAP7_75t_R FILLER_0_23_846 ();
 DECAPx6_ASAP7_75t_R FILLER_0_23_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_868 ();
 FILLER_ASAP7_75t_R FILLER_0_23_875 ();
 FILLER_ASAP7_75t_R FILLER_0_23_891 ();
 FILLER_ASAP7_75t_R FILLER_0_23_899 ();
 DECAPx2_ASAP7_75t_R FILLER_0_23_904 ();
 FILLER_ASAP7_75t_R FILLER_0_23_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_912 ();
 FILLER_ASAP7_75t_R FILLER_0_23_923 ();
 DECAPx6_ASAP7_75t_R FILLER_0_23_927 ();
 DECAPx1_ASAP7_75t_R FILLER_0_23_941 ();
 DECAPx6_ASAP7_75t_R FILLER_0_23_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_965 ();
 DECAPx1_ASAP7_75t_R FILLER_0_23_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_976 ();
 FILLER_ASAP7_75t_R FILLER_0_23_983 ();
 FILLER_ASAP7_75t_R FILLER_0_23_999 ();
 DECAPx4_ASAP7_75t_R FILLER_0_23_1011 ();
 DECAPx1_ASAP7_75t_R FILLER_0_23_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_1032 ();
 DECAPx2_ASAP7_75t_R FILLER_0_23_1039 ();
 FILLER_ASAP7_75t_R FILLER_0_23_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_1047 ();
 FILLER_ASAP7_75t_R FILLER_0_23_1053 ();
 FILLER_ASAP7_75t_R FILLER_0_23_1065 ();
 DECAPx4_ASAP7_75t_R FILLER_0_23_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_1082 ();
 DECAPx1_ASAP7_75t_R FILLER_0_23_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_1097 ();
 DECAPx1_ASAP7_75t_R FILLER_0_23_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_1117 ();
 DECAPx1_ASAP7_75t_R FILLER_0_23_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_1143 ();
 DECAPx1_ASAP7_75t_R FILLER_0_23_1150 ();
 FILLER_ASAP7_75t_R FILLER_0_23_1161 ();
 DECAPx4_ASAP7_75t_R FILLER_0_23_1169 ();
 FILLER_ASAP7_75t_R FILLER_0_23_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_1181 ();
 DECAPx2_ASAP7_75t_R FILLER_0_23_1188 ();
 FILLER_ASAP7_75t_R FILLER_0_23_1194 ();
 DECAPx1_ASAP7_75t_R FILLER_0_23_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_1206 ();
 FILLER_ASAP7_75t_R FILLER_0_23_1213 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_1221 ();
 DECAPx4_ASAP7_75t_R FILLER_0_23_1243 ();
 FILLER_ASAP7_75t_R FILLER_0_23_1259 ();
 DECAPx4_ASAP7_75t_R FILLER_0_23_1267 ();
 FILLER_ASAP7_75t_R FILLER_0_23_1277 ();
 FILLER_ASAP7_75t_R FILLER_0_23_1289 ();
 FILLER_ASAP7_75t_R FILLER_0_23_1297 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_1299 ();
 DECAPx2_ASAP7_75t_R FILLER_0_23_1306 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_1312 ();
 DECAPx1_ASAP7_75t_R FILLER_0_23_1319 ();
 DECAPx1_ASAP7_75t_R FILLER_0_23_1328 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_1332 ();
 DECAPx1_ASAP7_75t_R FILLER_0_23_1339 ();
 DECAPx6_ASAP7_75t_R FILLER_0_23_1349 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_1363 ();
 DECAPx2_ASAP7_75t_R FILLER_0_23_1374 ();
 FILLER_ASAP7_75t_R FILLER_0_23_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_24_24 ();
 FILLER_ASAP7_75t_R FILLER_0_24_38 ();
 DECAPx4_ASAP7_75t_R FILLER_0_24_46 ();
 FILLER_ASAP7_75t_R FILLER_0_24_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_58 ();
 DECAPx1_ASAP7_75t_R FILLER_0_24_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_69 ();
 FILLER_ASAP7_75t_R FILLER_0_24_76 ();
 FILLER_ASAP7_75t_R FILLER_0_24_84 ();
 FILLER_ASAP7_75t_R FILLER_0_24_96 ();
 FILLER_ASAP7_75t_R FILLER_0_24_108 ();
 FILLER_ASAP7_75t_R FILLER_0_24_120 ();
 FILLER_ASAP7_75t_R FILLER_0_24_128 ();
 FILLER_ASAP7_75t_R FILLER_0_24_140 ();
 FILLER_ASAP7_75t_R FILLER_0_24_148 ();
 DECAPx2_ASAP7_75t_R FILLER_0_24_157 ();
 FILLER_ASAP7_75t_R FILLER_0_24_163 ();
 FILLER_ASAP7_75t_R FILLER_0_24_172 ();
 FILLER_ASAP7_75t_R FILLER_0_24_180 ();
 DECAPx4_ASAP7_75t_R FILLER_0_24_188 ();
 FILLER_ASAP7_75t_R FILLER_0_24_204 ();
 FILLER_ASAP7_75t_R FILLER_0_24_212 ();
 FILLER_ASAP7_75t_R FILLER_0_24_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_222 ();
 FILLER_ASAP7_75t_R FILLER_0_24_229 ();
 DECAPx2_ASAP7_75t_R FILLER_0_24_237 ();
 FILLER_ASAP7_75t_R FILLER_0_24_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_245 ();
 FILLER_ASAP7_75t_R FILLER_0_24_252 ();
 DECAPx4_ASAP7_75t_R FILLER_0_24_260 ();
 FILLER_ASAP7_75t_R FILLER_0_24_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_278 ();
 FILLER_ASAP7_75t_R FILLER_0_24_289 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_301 ();
 DECAPx2_ASAP7_75t_R FILLER_0_24_323 ();
 FILLER_ASAP7_75t_R FILLER_0_24_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_341 ();
 DECAPx6_ASAP7_75t_R FILLER_0_24_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_377 ();
 DECAPx4_ASAP7_75t_R FILLER_0_24_398 ();
 FILLER_ASAP7_75t_R FILLER_0_24_416 ();
 FILLER_ASAP7_75t_R FILLER_0_24_428 ();
 FILLER_ASAP7_75t_R FILLER_0_24_436 ();
 FILLER_ASAP7_75t_R FILLER_0_24_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_451 ();
 DECAPx1_ASAP7_75t_R FILLER_0_24_458 ();
 DECAPx1_ASAP7_75t_R FILLER_0_24_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_468 ();
 FILLER_ASAP7_75t_R FILLER_0_24_476 ();
 FILLER_ASAP7_75t_R FILLER_0_24_485 ();
 FILLER_ASAP7_75t_R FILLER_0_24_490 ();
 DECAPx4_ASAP7_75t_R FILLER_0_24_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_512 ();
 FILLER_ASAP7_75t_R FILLER_0_24_519 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_529 ();
 DECAPx4_ASAP7_75t_R FILLER_0_24_551 ();
 FILLER_ASAP7_75t_R FILLER_0_24_561 ();
 DECAPx6_ASAP7_75t_R FILLER_0_24_569 ();
 DECAPx1_ASAP7_75t_R FILLER_0_24_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_587 ();
 FILLER_ASAP7_75t_R FILLER_0_24_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_593 ();
 FILLER_ASAP7_75t_R FILLER_0_24_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_607 ();
 DECAPx2_ASAP7_75t_R FILLER_0_24_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_622 ();
 FILLER_ASAP7_75t_R FILLER_0_24_629 ();
 FILLER_ASAP7_75t_R FILLER_0_24_637 ();
 DECAPx1_ASAP7_75t_R FILLER_0_24_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_655 ();
 DECAPx1_ASAP7_75t_R FILLER_0_24_664 ();
 FILLER_ASAP7_75t_R FILLER_0_24_676 ();
 DECAPx1_ASAP7_75t_R FILLER_0_24_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_699 ();
 FILLER_ASAP7_75t_R FILLER_0_24_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_723 ();
 DECAPx2_ASAP7_75t_R FILLER_0_24_729 ();
 FILLER_ASAP7_75t_R FILLER_0_24_735 ();
 FILLER_ASAP7_75t_R FILLER_0_24_743 ();
 DECAPx2_ASAP7_75t_R FILLER_0_24_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_757 ();
 FILLER_ASAP7_75t_R FILLER_0_24_761 ();
 FILLER_ASAP7_75t_R FILLER_0_24_775 ();
 FILLER_ASAP7_75t_R FILLER_0_24_782 ();
 DECAPx6_ASAP7_75t_R FILLER_0_24_790 ();
 DECAPx1_ASAP7_75t_R FILLER_0_24_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_820 ();
 FILLER_ASAP7_75t_R FILLER_0_24_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_826 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_835 ();
 DECAPx1_ASAP7_75t_R FILLER_0_24_857 ();
 DECAPx1_ASAP7_75t_R FILLER_0_24_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_873 ();
 FILLER_ASAP7_75t_R FILLER_0_24_880 ();
 FILLER_ASAP7_75t_R FILLER_0_24_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_895 ();
 DECAPx1_ASAP7_75t_R FILLER_0_24_902 ();
 FILLER_ASAP7_75t_R FILLER_0_24_914 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_922 ();
 DECAPx1_ASAP7_75t_R FILLER_0_24_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_948 ();
 FILLER_ASAP7_75t_R FILLER_0_24_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_965 ();
 FILLER_ASAP7_75t_R FILLER_0_24_972 ();
 DECAPx2_ASAP7_75t_R FILLER_0_24_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_24_993 ();
 FILLER_ASAP7_75t_R FILLER_0_24_999 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_1001 ();
 FILLER_ASAP7_75t_R FILLER_0_24_1008 ();
 DECAPx6_ASAP7_75t_R FILLER_0_24_1015 ();
 DECAPx4_ASAP7_75t_R FILLER_0_24_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_1050 ();
 DECAPx2_ASAP7_75t_R FILLER_0_24_1057 ();
 FILLER_ASAP7_75t_R FILLER_0_24_1073 ();
 FILLER_ASAP7_75t_R FILLER_0_24_1095 ();
 FILLER_ASAP7_75t_R FILLER_0_24_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_1105 ();
 DECAPx1_ASAP7_75t_R FILLER_0_24_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_1116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_24_1128 ();
 DECAPx1_ASAP7_75t_R FILLER_0_24_1142 ();
 DECAPx1_ASAP7_75t_R FILLER_0_24_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_1156 ();
 DECAPx2_ASAP7_75t_R FILLER_0_24_1169 ();
 FILLER_ASAP7_75t_R FILLER_0_24_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_1177 ();
 DECAPx4_ASAP7_75t_R FILLER_0_24_1185 ();
 FILLER_ASAP7_75t_R FILLER_0_24_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_1197 ();
 DECAPx2_ASAP7_75t_R FILLER_0_24_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_1210 ();
 DECAPx6_ASAP7_75t_R FILLER_0_24_1217 ();
 DECAPx2_ASAP7_75t_R FILLER_0_24_1237 ();
 FILLER_ASAP7_75t_R FILLER_0_24_1243 ();
 FILLER_ASAP7_75t_R FILLER_0_24_1251 ();
 DECAPx2_ASAP7_75t_R FILLER_0_24_1259 ();
 FILLER_ASAP7_75t_R FILLER_0_24_1271 ();
 DECAPx4_ASAP7_75t_R FILLER_0_24_1278 ();
 FILLER_ASAP7_75t_R FILLER_0_24_1295 ();
 FILLER_ASAP7_75t_R FILLER_0_24_1303 ();
 FILLER_ASAP7_75t_R FILLER_0_24_1310 ();
 FILLER_ASAP7_75t_R FILLER_0_24_1315 ();
 DECAPx6_ASAP7_75t_R FILLER_0_24_1328 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_1342 ();
 FILLER_ASAP7_75t_R FILLER_0_24_1351 ();
 DECAPx1_ASAP7_75t_R FILLER_0_24_1359 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_1363 ();
 DECAPx4_ASAP7_75t_R FILLER_0_24_1370 ();
 FILLER_ASAP7_75t_R FILLER_0_24_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_25_24 ();
 FILLER_ASAP7_75t_R FILLER_0_25_44 ();
 DECAPx1_ASAP7_75t_R FILLER_0_25_51 ();
 DECAPx1_ASAP7_75t_R FILLER_0_25_61 ();
 DECAPx1_ASAP7_75t_R FILLER_0_25_75 ();
 FILLER_ASAP7_75t_R FILLER_0_25_85 ();
 FILLER_ASAP7_75t_R FILLER_0_25_95 ();
 DECAPx1_ASAP7_75t_R FILLER_0_25_107 ();
 DECAPx1_ASAP7_75t_R FILLER_0_25_122 ();
 FILLER_ASAP7_75t_R FILLER_0_25_131 ();
 DECAPx2_ASAP7_75t_R FILLER_0_25_153 ();
 DECAPx4_ASAP7_75t_R FILLER_0_25_179 ();
 FILLER_ASAP7_75t_R FILLER_0_25_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_191 ();
 FILLER_ASAP7_75t_R FILLER_0_25_197 ();
 DECAPx2_ASAP7_75t_R FILLER_0_25_204 ();
 FILLER_ASAP7_75t_R FILLER_0_25_216 ();
 DECAPx2_ASAP7_75t_R FILLER_0_25_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_230 ();
 FILLER_ASAP7_75t_R FILLER_0_25_237 ();
 FILLER_ASAP7_75t_R FILLER_0_25_245 ();
 DECAPx4_ASAP7_75t_R FILLER_0_25_252 ();
 FILLER_ASAP7_75t_R FILLER_0_25_274 ();
 FILLER_ASAP7_75t_R FILLER_0_25_281 ();
 FILLER_ASAP7_75t_R FILLER_0_25_301 ();
 FILLER_ASAP7_75t_R FILLER_0_25_309 ();
 DECAPx4_ASAP7_75t_R FILLER_0_25_315 ();
 FILLER_ASAP7_75t_R FILLER_0_25_328 ();
 DECAPx1_ASAP7_75t_R FILLER_0_25_337 ();
 FILLER_ASAP7_75t_R FILLER_0_25_347 ();
 DECAPx1_ASAP7_75t_R FILLER_0_25_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_359 ();
 FILLER_ASAP7_75t_R FILLER_0_25_366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_25_374 ();
 FILLER_ASAP7_75t_R FILLER_0_25_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_382 ();
 FILLER_ASAP7_75t_R FILLER_0_25_391 ();
 DECAPx2_ASAP7_75t_R FILLER_0_25_399 ();
 FILLER_ASAP7_75t_R FILLER_0_25_405 ();
 DECAPx6_ASAP7_75t_R FILLER_0_25_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_429 ();
 DECAPx2_ASAP7_75t_R FILLER_0_25_436 ();
 FILLER_ASAP7_75t_R FILLER_0_25_442 ();
 FILLER_ASAP7_75t_R FILLER_0_25_449 ();
 DECAPx2_ASAP7_75t_R FILLER_0_25_456 ();
 FILLER_ASAP7_75t_R FILLER_0_25_462 ();
 DECAPx6_ASAP7_75t_R FILLER_0_25_470 ();
 DECAPx1_ASAP7_75t_R FILLER_0_25_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_488 ();
 FILLER_ASAP7_75t_R FILLER_0_25_495 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_505 ();
 DECAPx2_ASAP7_75t_R FILLER_0_25_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_533 ();
 FILLER_ASAP7_75t_R FILLER_0_25_540 ();
 FILLER_ASAP7_75t_R FILLER_0_25_548 ();
 FILLER_ASAP7_75t_R FILLER_0_25_556 ();
 DECAPx6_ASAP7_75t_R FILLER_0_25_569 ();
 FILLER_ASAP7_75t_R FILLER_0_25_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_585 ();
 FILLER_ASAP7_75t_R FILLER_0_25_594 ();
 DECAPx2_ASAP7_75t_R FILLER_0_25_602 ();
 FILLER_ASAP7_75t_R FILLER_0_25_620 ();
 DECAPx2_ASAP7_75t_R FILLER_0_25_634 ();
 DECAPx2_ASAP7_75t_R FILLER_0_25_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_657 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_686 ();
 DECAPx2_ASAP7_75t_R FILLER_0_25_708 ();
 FILLER_ASAP7_75t_R FILLER_0_25_714 ();
 FILLER_ASAP7_75t_R FILLER_0_25_719 ();
 DECAPx4_ASAP7_75t_R FILLER_0_25_727 ();
 FILLER_ASAP7_75t_R FILLER_0_25_745 ();
 FILLER_ASAP7_75t_R FILLER_0_25_753 ();
 DECAPx6_ASAP7_75t_R FILLER_0_25_766 ();
 DECAPx1_ASAP7_75t_R FILLER_0_25_780 ();
 FILLER_ASAP7_75t_R FILLER_0_25_789 ();
 FILLER_ASAP7_75t_R FILLER_0_25_802 ();
 DECAPx2_ASAP7_75t_R FILLER_0_25_815 ();
 FILLER_ASAP7_75t_R FILLER_0_25_821 ();
 FILLER_ASAP7_75t_R FILLER_0_25_828 ();
 DECAPx4_ASAP7_75t_R FILLER_0_25_836 ();
 DECAPx4_ASAP7_75t_R FILLER_0_25_866 ();
 FILLER_ASAP7_75t_R FILLER_0_25_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_878 ();
 DECAPx1_ASAP7_75t_R FILLER_0_25_885 ();
 DECAPx1_ASAP7_75t_R FILLER_0_25_892 ();
 FILLER_ASAP7_75t_R FILLER_0_25_903 ();
 FILLER_ASAP7_75t_R FILLER_0_25_911 ();
 FILLER_ASAP7_75t_R FILLER_0_25_923 ();
 DECAPx6_ASAP7_75t_R FILLER_0_25_927 ();
 DECAPx1_ASAP7_75t_R FILLER_0_25_941 ();
 DECAPx2_ASAP7_75t_R FILLER_0_25_955 ();
 FILLER_ASAP7_75t_R FILLER_0_25_967 ();
 DECAPx6_ASAP7_75t_R FILLER_0_25_975 ();
 FILLER_ASAP7_75t_R FILLER_0_25_989 ();
 DECAPx2_ASAP7_75t_R FILLER_0_25_997 ();
 FILLER_ASAP7_75t_R FILLER_0_25_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_1005 ();
 FILLER_ASAP7_75t_R FILLER_0_25_1012 ();
 DECAPx1_ASAP7_75t_R FILLER_0_25_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_1024 ();
 FILLER_ASAP7_75t_R FILLER_0_25_1031 ();
 DECAPx2_ASAP7_75t_R FILLER_0_25_1041 ();
 FILLER_ASAP7_75t_R FILLER_0_25_1053 ();
 DECAPx6_ASAP7_75t_R FILLER_0_25_1066 ();
 FILLER_ASAP7_75t_R FILLER_0_25_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_1082 ();
 DECAPx4_ASAP7_75t_R FILLER_0_25_1091 ();
 FILLER_ASAP7_75t_R FILLER_0_25_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_1103 ();
 FILLER_ASAP7_75t_R FILLER_0_25_1109 ();
 FILLER_ASAP7_75t_R FILLER_0_25_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_1119 ();
 FILLER_ASAP7_75t_R FILLER_0_25_1126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_1133 ();
 DECAPx1_ASAP7_75t_R FILLER_0_25_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_1164 ();
 FILLER_ASAP7_75t_R FILLER_0_25_1171 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_1180 ();
 FILLER_ASAP7_75t_R FILLER_0_25_1208 ();
 FILLER_ASAP7_75t_R FILLER_0_25_1216 ();
 DECAPx2_ASAP7_75t_R FILLER_0_25_1224 ();
 FILLER_ASAP7_75t_R FILLER_0_25_1230 ();
 DECAPx1_ASAP7_75t_R FILLER_0_25_1243 ();
 DECAPx6_ASAP7_75t_R FILLER_0_25_1253 ();
 FILLER_ASAP7_75t_R FILLER_0_25_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_0_25_1275 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_1279 ();
 DECAPx2_ASAP7_75t_R FILLER_0_25_1287 ();
 FILLER_ASAP7_75t_R FILLER_0_25_1293 ();
 FILLER_ASAP7_75t_R FILLER_0_25_1301 ();
 FILLER_ASAP7_75t_R FILLER_0_25_1308 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_1310 ();
 FILLER_ASAP7_75t_R FILLER_0_25_1317 ();
 DECAPx4_ASAP7_75t_R FILLER_0_25_1325 ();
 FILLER_ASAP7_75t_R FILLER_0_25_1335 ();
 FILLER_ASAP7_75t_R FILLER_0_25_1357 ();
 DECAPx1_ASAP7_75t_R FILLER_0_25_1365 ();
 FILLER_ASAP7_75t_R FILLER_0_25_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_26_24 ();
 FILLER_ASAP7_75t_R FILLER_0_26_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_36 ();
 DECAPx1_ASAP7_75t_R FILLER_0_26_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_47 ();
 FILLER_ASAP7_75t_R FILLER_0_26_54 ();
 FILLER_ASAP7_75t_R FILLER_0_26_76 ();
 DECAPx1_ASAP7_75t_R FILLER_0_26_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_88 ();
 FILLER_ASAP7_75t_R FILLER_0_26_109 ();
 FILLER_ASAP7_75t_R FILLER_0_26_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_118 ();
 FILLER_ASAP7_75t_R FILLER_0_26_124 ();
 DECAPx1_ASAP7_75t_R FILLER_0_26_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_135 ();
 FILLER_ASAP7_75t_R FILLER_0_26_141 ();
 FILLER_ASAP7_75t_R FILLER_0_26_150 ();
 DECAPx1_ASAP7_75t_R FILLER_0_26_157 ();
 FILLER_ASAP7_75t_R FILLER_0_26_167 ();
 FILLER_ASAP7_75t_R FILLER_0_26_175 ();
 FILLER_ASAP7_75t_R FILLER_0_26_184 ();
 FILLER_ASAP7_75t_R FILLER_0_26_196 ();
 FILLER_ASAP7_75t_R FILLER_0_26_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_210 ();
 FILLER_ASAP7_75t_R FILLER_0_26_217 ();
 FILLER_ASAP7_75t_R FILLER_0_26_226 ();
 DECAPx1_ASAP7_75t_R FILLER_0_26_238 ();
 FILLER_ASAP7_75t_R FILLER_0_26_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_250 ();
 FILLER_ASAP7_75t_R FILLER_0_26_258 ();
 FILLER_ASAP7_75t_R FILLER_0_26_270 ();
 FILLER_ASAP7_75t_R FILLER_0_26_282 ();
 FILLER_ASAP7_75t_R FILLER_0_26_290 ();
 FILLER_ASAP7_75t_R FILLER_0_26_302 ();
 FILLER_ASAP7_75t_R FILLER_0_26_310 ();
 FILLER_ASAP7_75t_R FILLER_0_26_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_319 ();
 FILLER_ASAP7_75t_R FILLER_0_26_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_334 ();
 FILLER_ASAP7_75t_R FILLER_0_26_341 ();
 FILLER_ASAP7_75t_R FILLER_0_26_351 ();
 FILLER_ASAP7_75t_R FILLER_0_26_359 ();
 FILLER_ASAP7_75t_R FILLER_0_26_369 ();
 DECAPx2_ASAP7_75t_R FILLER_0_26_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_383 ();
 FILLER_ASAP7_75t_R FILLER_0_26_392 ();
 FILLER_ASAP7_75t_R FILLER_0_26_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_402 ();
 DECAPx4_ASAP7_75t_R FILLER_0_26_415 ();
 FILLER_ASAP7_75t_R FILLER_0_26_425 ();
 FILLER_ASAP7_75t_R FILLER_0_26_437 ();
 FILLER_ASAP7_75t_R FILLER_0_26_449 ();
 DECAPx1_ASAP7_75t_R FILLER_0_26_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_461 ();
 DECAPx1_ASAP7_75t_R FILLER_0_26_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_468 ();
 DECAPx6_ASAP7_75t_R FILLER_0_26_475 ();
 FILLER_ASAP7_75t_R FILLER_0_26_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_497 ();
 DECAPx6_ASAP7_75t_R FILLER_0_26_504 ();
 DECAPx2_ASAP7_75t_R FILLER_0_26_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_26_532 ();
 FILLER_ASAP7_75t_R FILLER_0_26_544 ();
 DECAPx6_ASAP7_75t_R FILLER_0_26_552 ();
 FILLER_ASAP7_75t_R FILLER_0_26_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_568 ();
 DECAPx2_ASAP7_75t_R FILLER_0_26_572 ();
 FILLER_ASAP7_75t_R FILLER_0_26_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_580 ();
 DECAPx6_ASAP7_75t_R FILLER_0_26_602 ();
 DECAPx2_ASAP7_75t_R FILLER_0_26_616 ();
 FILLER_ASAP7_75t_R FILLER_0_26_628 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_638 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_666 ();
 DECAPx6_ASAP7_75t_R FILLER_0_26_688 ();
 FILLER_ASAP7_75t_R FILLER_0_26_713 ();
 FILLER_ASAP7_75t_R FILLER_0_26_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_723 ();
 FILLER_ASAP7_75t_R FILLER_0_26_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_732 ();
 FILLER_ASAP7_75t_R FILLER_0_26_741 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_751 ();
 DECAPx6_ASAP7_75t_R FILLER_0_26_773 ();
 DECAPx2_ASAP7_75t_R FILLER_0_26_787 ();
 FILLER_ASAP7_75t_R FILLER_0_26_799 ();
 DECAPx6_ASAP7_75t_R FILLER_0_26_807 ();
 DECAPx1_ASAP7_75t_R FILLER_0_26_821 ();
 FILLER_ASAP7_75t_R FILLER_0_26_828 ();
 FILLER_ASAP7_75t_R FILLER_0_26_851 ();
 FILLER_ASAP7_75t_R FILLER_0_26_858 ();
 DECAPx2_ASAP7_75t_R FILLER_0_26_865 ();
 FILLER_ASAP7_75t_R FILLER_0_26_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_873 ();
 FILLER_ASAP7_75t_R FILLER_0_26_880 ();
 FILLER_ASAP7_75t_R FILLER_0_26_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_891 ();
 DECAPx1_ASAP7_75t_R FILLER_0_26_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_904 ();
 DECAPx1_ASAP7_75t_R FILLER_0_26_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_915 ();
 DECAPx1_ASAP7_75t_R FILLER_0_26_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_926 ();
 DECAPx1_ASAP7_75t_R FILLER_0_26_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_937 ();
 DECAPx6_ASAP7_75t_R FILLER_0_26_946 ();
 FILLER_ASAP7_75t_R FILLER_0_26_966 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_974 ();
 DECAPx2_ASAP7_75t_R FILLER_0_26_996 ();
 DECAPx2_ASAP7_75t_R FILLER_0_26_1012 ();
 FILLER_ASAP7_75t_R FILLER_0_26_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_1020 ();
 FILLER_ASAP7_75t_R FILLER_0_26_1028 ();
 FILLER_ASAP7_75t_R FILLER_0_26_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_1037 ();
 DECAPx1_ASAP7_75t_R FILLER_0_26_1046 ();
 DECAPx2_ASAP7_75t_R FILLER_0_26_1060 ();
 FILLER_ASAP7_75t_R FILLER_0_26_1066 ();
 FILLER_ASAP7_75t_R FILLER_0_26_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_1075 ();
 DECAPx6_ASAP7_75t_R FILLER_0_26_1082 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_1096 ();
 DECAPx1_ASAP7_75t_R FILLER_0_26_1104 ();
 FILLER_ASAP7_75t_R FILLER_0_26_1118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_1126 ();
 DECAPx4_ASAP7_75t_R FILLER_0_26_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_1158 ();
 FILLER_ASAP7_75t_R FILLER_0_26_1165 ();
 DECAPx2_ASAP7_75t_R FILLER_0_26_1173 ();
 FILLER_ASAP7_75t_R FILLER_0_26_1179 ();
 FILLER_ASAP7_75t_R FILLER_0_26_1192 ();
 DECAPx1_ASAP7_75t_R FILLER_0_26_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_1214 ();
 DECAPx6_ASAP7_75t_R FILLER_0_26_1247 ();
 DECAPx1_ASAP7_75t_R FILLER_0_26_1261 ();
 FILLER_ASAP7_75t_R FILLER_0_26_1271 ();
 DECAPx6_ASAP7_75t_R FILLER_0_26_1279 ();
 FILLER_ASAP7_75t_R FILLER_0_26_1293 ();
 DECAPx4_ASAP7_75t_R FILLER_0_26_1301 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_1311 ();
 DECAPx2_ASAP7_75t_R FILLER_0_26_1320 ();
 FILLER_ASAP7_75t_R FILLER_0_26_1326 ();
 DECAPx1_ASAP7_75t_R FILLER_0_26_1336 ();
 FILLER_ASAP7_75t_R FILLER_0_26_1343 ();
 FILLER_ASAP7_75t_R FILLER_0_26_1350 ();
 FILLER_ASAP7_75t_R FILLER_0_26_1358 ();
 FILLER_ASAP7_75t_R FILLER_0_26_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_27_24 ();
 DECAPx2_ASAP7_75t_R FILLER_0_27_38 ();
 FILLER_ASAP7_75t_R FILLER_0_27_49 ();
 FILLER_ASAP7_75t_R FILLER_0_27_59 ();
 DECAPx2_ASAP7_75t_R FILLER_0_27_66 ();
 DECAPx1_ASAP7_75t_R FILLER_0_27_92 ();
 FILLER_ASAP7_75t_R FILLER_0_27_102 ();
 FILLER_ASAP7_75t_R FILLER_0_27_112 ();
 FILLER_ASAP7_75t_R FILLER_0_27_122 ();
 FILLER_ASAP7_75t_R FILLER_0_27_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_132 ();
 DECAPx2_ASAP7_75t_R FILLER_0_27_143 ();
 DECAPx2_ASAP7_75t_R FILLER_0_27_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_162 ();
 DECAPx1_ASAP7_75t_R FILLER_0_27_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_173 ();
 DECAPx2_ASAP7_75t_R FILLER_0_27_182 ();
 FILLER_ASAP7_75t_R FILLER_0_27_193 ();
 FILLER_ASAP7_75t_R FILLER_0_27_205 ();
 FILLER_ASAP7_75t_R FILLER_0_27_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_216 ();
 FILLER_ASAP7_75t_R FILLER_0_27_223 ();
 FILLER_ASAP7_75t_R FILLER_0_27_231 ();
 FILLER_ASAP7_75t_R FILLER_0_27_243 ();
 FILLER_ASAP7_75t_R FILLER_0_27_250 ();
 FILLER_ASAP7_75t_R FILLER_0_27_262 ();
 FILLER_ASAP7_75t_R FILLER_0_27_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_276 ();
 FILLER_ASAP7_75t_R FILLER_0_27_295 ();
 FILLER_ASAP7_75t_R FILLER_0_27_307 ();
 FILLER_ASAP7_75t_R FILLER_0_27_317 ();
 FILLER_ASAP7_75t_R FILLER_0_27_325 ();
 DECAPx2_ASAP7_75t_R FILLER_0_27_335 ();
 FILLER_ASAP7_75t_R FILLER_0_27_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_343 ();
 DECAPx2_ASAP7_75t_R FILLER_0_27_350 ();
 FILLER_ASAP7_75t_R FILLER_0_27_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_358 ();
 FILLER_ASAP7_75t_R FILLER_0_27_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_367 ();
 DECAPx6_ASAP7_75t_R FILLER_0_27_378 ();
 DECAPx2_ASAP7_75t_R FILLER_0_27_392 ();
 DECAPx2_ASAP7_75t_R FILLER_0_27_418 ();
 FILLER_ASAP7_75t_R FILLER_0_27_424 ();
 FILLER_ASAP7_75t_R FILLER_0_27_438 ();
 DECAPx2_ASAP7_75t_R FILLER_0_27_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_453 ();
 DECAPx6_ASAP7_75t_R FILLER_0_27_464 ();
 FILLER_ASAP7_75t_R FILLER_0_27_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_480 ();
 FILLER_ASAP7_75t_R FILLER_0_27_496 ();
 DECAPx4_ASAP7_75t_R FILLER_0_27_509 ();
 FILLER_ASAP7_75t_R FILLER_0_27_525 ();
 DECAPx1_ASAP7_75t_R FILLER_0_27_535 ();
 DECAPx4_ASAP7_75t_R FILLER_0_27_543 ();
 FILLER_ASAP7_75t_R FILLER_0_27_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_558 ();
 FILLER_ASAP7_75t_R FILLER_0_27_565 ();
 DECAPx6_ASAP7_75t_R FILLER_0_27_578 ();
 DECAPx1_ASAP7_75t_R FILLER_0_27_592 ();
 FILLER_ASAP7_75t_R FILLER_0_27_599 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_611 ();
 FILLER_ASAP7_75t_R FILLER_0_27_633 ();
 DECAPx2_ASAP7_75t_R FILLER_0_27_641 ();
 FILLER_ASAP7_75t_R FILLER_0_27_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_649 ();
 FILLER_ASAP7_75t_R FILLER_0_27_661 ();
 DECAPx4_ASAP7_75t_R FILLER_0_27_666 ();
 FILLER_ASAP7_75t_R FILLER_0_27_676 ();
 FILLER_ASAP7_75t_R FILLER_0_27_690 ();
 DECAPx4_ASAP7_75t_R FILLER_0_27_698 ();
 FILLER_ASAP7_75t_R FILLER_0_27_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_722 ();
 DECAPx6_ASAP7_75t_R FILLER_0_27_726 ();
 DECAPx1_ASAP7_75t_R FILLER_0_27_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_748 ();
 FILLER_ASAP7_75t_R FILLER_0_27_770 ();
 DECAPx2_ASAP7_75t_R FILLER_0_27_782 ();
 FILLER_ASAP7_75t_R FILLER_0_27_788 ();
 FILLER_ASAP7_75t_R FILLER_0_27_798 ();
 FILLER_ASAP7_75t_R FILLER_0_27_808 ();
 DECAPx4_ASAP7_75t_R FILLER_0_27_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_831 ();
 DECAPx2_ASAP7_75t_R FILLER_0_27_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_841 ();
 DECAPx4_ASAP7_75t_R FILLER_0_27_854 ();
 FILLER_ASAP7_75t_R FILLER_0_27_870 ();
 FILLER_ASAP7_75t_R FILLER_0_27_877 ();
 FILLER_ASAP7_75t_R FILLER_0_27_884 ();
 FILLER_ASAP7_75t_R FILLER_0_27_891 ();
 FILLER_ASAP7_75t_R FILLER_0_27_899 ();
 FILLER_ASAP7_75t_R FILLER_0_27_904 ();
 FILLER_ASAP7_75t_R FILLER_0_27_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_914 ();
 DECAPx1_ASAP7_75t_R FILLER_0_27_921 ();
 FILLER_ASAP7_75t_R FILLER_0_27_927 ();
 DECAPx2_ASAP7_75t_R FILLER_0_27_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_941 ();
 FILLER_ASAP7_75t_R FILLER_0_27_953 ();
 FILLER_ASAP7_75t_R FILLER_0_27_961 ();
 DECAPx2_ASAP7_75t_R FILLER_0_27_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_975 ();
 DECAPx2_ASAP7_75t_R FILLER_0_27_987 ();
 FILLER_ASAP7_75t_R FILLER_0_27_999 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_1001 ();
 DECAPx1_ASAP7_75t_R FILLER_0_27_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_1012 ();
 FILLER_ASAP7_75t_R FILLER_0_27_1019 ();
 DECAPx2_ASAP7_75t_R FILLER_0_27_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_1033 ();
 DECAPx1_ASAP7_75t_R FILLER_0_27_1044 ();
 FILLER_ASAP7_75t_R FILLER_0_27_1054 ();
 DECAPx4_ASAP7_75t_R FILLER_0_27_1062 ();
 FILLER_ASAP7_75t_R FILLER_0_27_1072 ();
 FILLER_ASAP7_75t_R FILLER_0_27_1084 ();
 FILLER_ASAP7_75t_R FILLER_0_27_1091 ();
 FILLER_ASAP7_75t_R FILLER_0_27_1099 ();
 FILLER_ASAP7_75t_R FILLER_0_27_1107 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_1114 ();
 DECAPx6_ASAP7_75t_R FILLER_0_27_1136 ();
 DECAPx1_ASAP7_75t_R FILLER_0_27_1150 ();
 FILLER_ASAP7_75t_R FILLER_0_27_1162 ();
 FILLER_ASAP7_75t_R FILLER_0_27_1170 ();
 DECAPx2_ASAP7_75t_R FILLER_0_27_1175 ();
 DECAPx1_ASAP7_75t_R FILLER_0_27_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_1197 ();
 FILLER_ASAP7_75t_R FILLER_0_27_1219 ();
 DECAPx1_ASAP7_75t_R FILLER_0_27_1227 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_1231 ();
 FILLER_ASAP7_75t_R FILLER_0_27_1242 ();
 DECAPx6_ASAP7_75t_R FILLER_0_27_1249 ();
 FILLER_ASAP7_75t_R FILLER_0_27_1263 ();
 FILLER_ASAP7_75t_R FILLER_0_27_1271 ();
 DECAPx4_ASAP7_75t_R FILLER_0_27_1279 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_1289 ();
 FILLER_ASAP7_75t_R FILLER_0_27_1296 ();
 DECAPx4_ASAP7_75t_R FILLER_0_27_1304 ();
 FILLER_ASAP7_75t_R FILLER_0_27_1324 ();
 FILLER_ASAP7_75t_R FILLER_0_27_1332 ();
 DECAPx4_ASAP7_75t_R FILLER_0_27_1340 ();
 FILLER_ASAP7_75t_R FILLER_0_27_1358 ();
 FILLER_ASAP7_75t_R FILLER_0_27_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_24 ();
 DECAPx6_ASAP7_75t_R FILLER_0_28_57 ();
 FILLER_ASAP7_75t_R FILLER_0_28_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_73 ();
 DECAPx4_ASAP7_75t_R FILLER_0_28_80 ();
 FILLER_ASAP7_75t_R FILLER_0_28_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_92 ();
 FILLER_ASAP7_75t_R FILLER_0_28_99 ();
 DECAPx1_ASAP7_75t_R FILLER_0_28_112 ();
 FILLER_ASAP7_75t_R FILLER_0_28_126 ();
 FILLER_ASAP7_75t_R FILLER_0_28_138 ();
 DECAPx1_ASAP7_75t_R FILLER_0_28_150 ();
 FILLER_ASAP7_75t_R FILLER_0_28_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_166 ();
 FILLER_ASAP7_75t_R FILLER_0_28_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_189 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_195 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_211 ();
 FILLER_ASAP7_75t_R FILLER_0_28_217 ();
 FILLER_ASAP7_75t_R FILLER_0_28_226 ();
 FILLER_ASAP7_75t_R FILLER_0_28_236 ();
 FILLER_ASAP7_75t_R FILLER_0_28_248 ();
 FILLER_ASAP7_75t_R FILLER_0_28_260 ();
 FILLER_ASAP7_75t_R FILLER_0_28_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_274 ();
 FILLER_ASAP7_75t_R FILLER_0_28_290 ();
 FILLER_ASAP7_75t_R FILLER_0_28_297 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_317 ();
 FILLER_ASAP7_75t_R FILLER_0_28_329 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_345 ();
 FILLER_ASAP7_75t_R FILLER_0_28_352 ();
 DECAPx4_ASAP7_75t_R FILLER_0_28_360 ();
 FILLER_ASAP7_75t_R FILLER_0_28_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_372 ();
 DECAPx6_ASAP7_75t_R FILLER_0_28_376 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_390 ();
 FILLER_ASAP7_75t_R FILLER_0_28_402 ();
 DECAPx6_ASAP7_75t_R FILLER_0_28_410 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_430 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_448 ();
 FILLER_ASAP7_75t_R FILLER_0_28_460 ();
 DECAPx1_ASAP7_75t_R FILLER_0_28_464 ();
 DECAPx1_ASAP7_75t_R FILLER_0_28_474 ();
 DECAPx1_ASAP7_75t_R FILLER_0_28_485 ();
 FILLER_ASAP7_75t_R FILLER_0_28_501 ();
 DECAPx1_ASAP7_75t_R FILLER_0_28_509 ();
 DECAPx1_ASAP7_75t_R FILLER_0_28_523 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_533 ();
 FILLER_ASAP7_75t_R FILLER_0_28_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_541 ();
 FILLER_ASAP7_75t_R FILLER_0_28_548 ();
 DECAPx6_ASAP7_75t_R FILLER_0_28_556 ();
 DECAPx1_ASAP7_75t_R FILLER_0_28_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_574 ();
 DECAPx6_ASAP7_75t_R FILLER_0_28_581 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_595 ();
 FILLER_ASAP7_75t_R FILLER_0_28_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_609 ();
 FILLER_ASAP7_75t_R FILLER_0_28_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_618 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_630 ();
 FILLER_ASAP7_75t_R FILLER_0_28_636 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_656 ();
 FILLER_ASAP7_75t_R FILLER_0_28_663 ();
 FILLER_ASAP7_75t_R FILLER_0_28_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_675 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_693 ();
 DECAPx1_ASAP7_75t_R FILLER_0_28_702 ();
 DECAPx6_ASAP7_75t_R FILLER_0_28_718 ();
 FILLER_ASAP7_75t_R FILLER_0_28_732 ();
 DECAPx4_ASAP7_75t_R FILLER_0_28_742 ();
 FILLER_ASAP7_75t_R FILLER_0_28_764 ();
 FILLER_ASAP7_75t_R FILLER_0_28_786 ();
 FILLER_ASAP7_75t_R FILLER_0_28_798 ();
 FILLER_ASAP7_75t_R FILLER_0_28_808 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_821 ();
 FILLER_ASAP7_75t_R FILLER_0_28_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_829 ();
 DECAPx6_ASAP7_75t_R FILLER_0_28_835 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_855 ();
 FILLER_ASAP7_75t_R FILLER_0_28_874 ();
 FILLER_ASAP7_75t_R FILLER_0_28_882 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_887 ();
 FILLER_ASAP7_75t_R FILLER_0_28_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_902 ();
 FILLER_ASAP7_75t_R FILLER_0_28_909 ();
 DECAPx1_ASAP7_75t_R FILLER_0_28_918 ();
 FILLER_ASAP7_75t_R FILLER_0_28_928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_936 ();
 DECAPx6_ASAP7_75t_R FILLER_0_28_958 ();
 DECAPx1_ASAP7_75t_R FILLER_0_28_972 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_982 ();
 FILLER_ASAP7_75t_R FILLER_0_28_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_996 ();
 FILLER_ASAP7_75t_R FILLER_0_28_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_1009 ();
 DECAPx6_ASAP7_75t_R FILLER_0_28_1014 ();
 FILLER_ASAP7_75t_R FILLER_0_28_1028 ();
 FILLER_ASAP7_75t_R FILLER_0_28_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_1038 ();
 FILLER_ASAP7_75t_R FILLER_0_28_1044 ();
 FILLER_ASAP7_75t_R FILLER_0_28_1053 ();
 FILLER_ASAP7_75t_R FILLER_0_28_1061 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_1069 ();
 FILLER_ASAP7_75t_R FILLER_0_28_1075 ();
 FILLER_ASAP7_75t_R FILLER_0_28_1084 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_1098 ();
 FILLER_ASAP7_75t_R FILLER_0_28_1105 ();
 FILLER_ASAP7_75t_R FILLER_0_28_1113 ();
 DECAPx6_ASAP7_75t_R FILLER_0_28_1121 ();
 DECAPx1_ASAP7_75t_R FILLER_0_28_1135 ();
 FILLER_ASAP7_75t_R FILLER_0_28_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_1151 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_1170 ();
 FILLER_ASAP7_75t_R FILLER_0_28_1176 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_1178 ();
 DECAPx1_ASAP7_75t_R FILLER_0_28_1185 ();
 DECAPx4_ASAP7_75t_R FILLER_0_28_1195 ();
 FILLER_ASAP7_75t_R FILLER_0_28_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_1207 ();
 FILLER_ASAP7_75t_R FILLER_0_28_1220 ();
 FILLER_ASAP7_75t_R FILLER_0_28_1228 ();
 DECAPx4_ASAP7_75t_R FILLER_0_28_1236 ();
 FILLER_ASAP7_75t_R FILLER_0_28_1249 ();
 FILLER_ASAP7_75t_R FILLER_0_28_1257 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_1264 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_1270 ();
 FILLER_ASAP7_75t_R FILLER_0_28_1283 ();
 FILLER_ASAP7_75t_R FILLER_0_28_1290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_1298 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_1304 ();
 FILLER_ASAP7_75t_R FILLER_0_28_1317 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_1325 ();
 FILLER_ASAP7_75t_R FILLER_0_28_1331 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_1333 ();
 DECAPx4_ASAP7_75t_R FILLER_0_28_1342 ();
 FILLER_ASAP7_75t_R FILLER_0_28_1352 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_1354 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_1361 ();
 DECAPx1_ASAP7_75t_R FILLER_0_28_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_24 ();
 DECAPx6_ASAP7_75t_R FILLER_0_29_46 ();
 DECAPx1_ASAP7_75t_R FILLER_0_29_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_64 ();
 FILLER_ASAP7_75t_R FILLER_0_29_70 ();
 DECAPx1_ASAP7_75t_R FILLER_0_29_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_81 ();
 FILLER_ASAP7_75t_R FILLER_0_29_87 ();
 FILLER_ASAP7_75t_R FILLER_0_29_99 ();
 FILLER_ASAP7_75t_R FILLER_0_29_109 ();
 DECAPx2_ASAP7_75t_R FILLER_0_29_122 ();
 DECAPx1_ASAP7_75t_R FILLER_0_29_139 ();
 FILLER_ASAP7_75t_R FILLER_0_29_148 ();
 FILLER_ASAP7_75t_R FILLER_0_29_170 ();
 FILLER_ASAP7_75t_R FILLER_0_29_182 ();
 FILLER_ASAP7_75t_R FILLER_0_29_192 ();
 FILLER_ASAP7_75t_R FILLER_0_29_204 ();
 DECAPx2_ASAP7_75t_R FILLER_0_29_213 ();
 FILLER_ASAP7_75t_R FILLER_0_29_219 ();
 FILLER_ASAP7_75t_R FILLER_0_29_229 ();
 DECAPx1_ASAP7_75t_R FILLER_0_29_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_241 ();
 DECAPx1_ASAP7_75t_R FILLER_0_29_252 ();
 FILLER_ASAP7_75t_R FILLER_0_29_294 ();
 DECAPx2_ASAP7_75t_R FILLER_0_29_306 ();
 FILLER_ASAP7_75t_R FILLER_0_29_312 ();
 DECAPx2_ASAP7_75t_R FILLER_0_29_326 ();
 DECAPx2_ASAP7_75t_R FILLER_0_29_342 ();
 FILLER_ASAP7_75t_R FILLER_0_29_354 ();
 DECAPx2_ASAP7_75t_R FILLER_0_29_363 ();
 FILLER_ASAP7_75t_R FILLER_0_29_375 ();
 DECAPx4_ASAP7_75t_R FILLER_0_29_384 ();
 FILLER_ASAP7_75t_R FILLER_0_29_394 ();
 DECAPx2_ASAP7_75t_R FILLER_0_29_402 ();
 FILLER_ASAP7_75t_R FILLER_0_29_418 ();
 FILLER_ASAP7_75t_R FILLER_0_29_430 ();
 DECAPx1_ASAP7_75t_R FILLER_0_29_444 ();
 DECAPx4_ASAP7_75t_R FILLER_0_29_458 ();
 FILLER_ASAP7_75t_R FILLER_0_29_468 ();
 DECAPx2_ASAP7_75t_R FILLER_0_29_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_482 ();
 FILLER_ASAP7_75t_R FILLER_0_29_487 ();
 DECAPx1_ASAP7_75t_R FILLER_0_29_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_498 ();
 DECAPx2_ASAP7_75t_R FILLER_0_29_515 ();
 FILLER_ASAP7_75t_R FILLER_0_29_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_523 ();
 DECAPx4_ASAP7_75t_R FILLER_0_29_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_544 ();
 FILLER_ASAP7_75t_R FILLER_0_29_551 ();
 DECAPx1_ASAP7_75t_R FILLER_0_29_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_576 ();
 DECAPx1_ASAP7_75t_R FILLER_0_29_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_602 ();
 FILLER_ASAP7_75t_R FILLER_0_29_611 ();
 DECAPx1_ASAP7_75t_R FILLER_0_29_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_627 ();
 DECAPx2_ASAP7_75t_R FILLER_0_29_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_655 ();
 FILLER_ASAP7_75t_R FILLER_0_29_664 ();
 DECAPx1_ASAP7_75t_R FILLER_0_29_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_680 ();
 FILLER_ASAP7_75t_R FILLER_0_29_687 ();
 DECAPx1_ASAP7_75t_R FILLER_0_29_695 ();
 DECAPx1_ASAP7_75t_R FILLER_0_29_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_706 ();
 DECAPx2_ASAP7_75t_R FILLER_0_29_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_725 ();
 FILLER_ASAP7_75t_R FILLER_0_29_732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_762 ();
 DECAPx6_ASAP7_75t_R FILLER_0_29_773 ();
 FILLER_ASAP7_75t_R FILLER_0_29_787 ();
 FILLER_ASAP7_75t_R FILLER_0_29_800 ();
 FILLER_ASAP7_75t_R FILLER_0_29_805 ();
 DECAPx2_ASAP7_75t_R FILLER_0_29_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_825 ();
 DECAPx1_ASAP7_75t_R FILLER_0_29_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_842 ();
 DECAPx4_ASAP7_75t_R FILLER_0_29_851 ();
 FILLER_ASAP7_75t_R FILLER_0_29_871 ();
 FILLER_ASAP7_75t_R FILLER_0_29_883 ();
 FILLER_ASAP7_75t_R FILLER_0_29_892 ();
 FILLER_ASAP7_75t_R FILLER_0_29_899 ();
 FILLER_ASAP7_75t_R FILLER_0_29_907 ();
 DECAPx1_ASAP7_75t_R FILLER_0_29_914 ();
 FILLER_ASAP7_75t_R FILLER_0_29_923 ();
 FILLER_ASAP7_75t_R FILLER_0_29_927 ();
 FILLER_ASAP7_75t_R FILLER_0_29_939 ();
 FILLER_ASAP7_75t_R FILLER_0_29_951 ();
 FILLER_ASAP7_75t_R FILLER_0_29_963 ();
 FILLER_ASAP7_75t_R FILLER_0_29_975 ();
 FILLER_ASAP7_75t_R FILLER_0_29_987 ();
 FILLER_ASAP7_75t_R FILLER_0_29_995 ();
 FILLER_ASAP7_75t_R FILLER_0_29_1003 ();
 DECAPx4_ASAP7_75t_R FILLER_0_29_1011 ();
 FILLER_ASAP7_75t_R FILLER_0_29_1021 ();
 FILLER_ASAP7_75t_R FILLER_0_29_1031 ();
 DECAPx2_ASAP7_75t_R FILLER_0_29_1039 ();
 FILLER_ASAP7_75t_R FILLER_0_29_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_1047 ();
 FILLER_ASAP7_75t_R FILLER_0_29_1058 ();
 FILLER_ASAP7_75t_R FILLER_0_29_1066 ();
 DECAPx2_ASAP7_75t_R FILLER_0_29_1074 ();
 FILLER_ASAP7_75t_R FILLER_0_29_1080 ();
 DECAPx1_ASAP7_75t_R FILLER_0_29_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_1095 ();
 DECAPx2_ASAP7_75t_R FILLER_0_29_1104 ();
 FILLER_ASAP7_75t_R FILLER_0_29_1116 ();
 DECAPx2_ASAP7_75t_R FILLER_0_29_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_1135 ();
 FILLER_ASAP7_75t_R FILLER_0_29_1156 ();
 DECAPx1_ASAP7_75t_R FILLER_0_29_1165 ();
 DECAPx4_ASAP7_75t_R FILLER_0_29_1175 ();
 FILLER_ASAP7_75t_R FILLER_0_29_1185 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_1187 ();
 DECAPx6_ASAP7_75t_R FILLER_0_29_1194 ();
 DECAPx1_ASAP7_75t_R FILLER_0_29_1208 ();
 FILLER_ASAP7_75t_R FILLER_0_29_1218 ();
 DECAPx2_ASAP7_75t_R FILLER_0_29_1226 ();
 FILLER_ASAP7_75t_R FILLER_0_29_1238 ();
 DECAPx2_ASAP7_75t_R FILLER_0_29_1245 ();
 FILLER_ASAP7_75t_R FILLER_0_29_1251 ();
 FILLER_ASAP7_75t_R FILLER_0_29_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_1269 ();
 FILLER_ASAP7_75t_R FILLER_0_29_1291 ();
 FILLER_ASAP7_75t_R FILLER_0_29_1303 ();
 DECAPx4_ASAP7_75t_R FILLER_0_29_1311 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_1321 ();
 DECAPx1_ASAP7_75t_R FILLER_0_29_1330 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_1334 ();
 FILLER_ASAP7_75t_R FILLER_0_29_1341 ();
 FILLER_ASAP7_75t_R FILLER_0_29_1354 ();
 DECAPx6_ASAP7_75t_R FILLER_0_29_1362 ();
 DECAPx2_ASAP7_75t_R FILLER_0_29_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_24 ();
 FILLER_ASAP7_75t_R FILLER_0_30_52 ();
 DECAPx1_ASAP7_75t_R FILLER_0_30_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_64 ();
 FILLER_ASAP7_75t_R FILLER_0_30_75 ();
 DECAPx1_ASAP7_75t_R FILLER_0_30_83 ();
 FILLER_ASAP7_75t_R FILLER_0_30_92 ();
 FILLER_ASAP7_75t_R FILLER_0_30_104 ();
 FILLER_ASAP7_75t_R FILLER_0_30_116 ();
 FILLER_ASAP7_75t_R FILLER_0_30_128 ();
 FILLER_ASAP7_75t_R FILLER_0_30_140 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_148 ();
 FILLER_ASAP7_75t_R FILLER_0_30_154 ();
 FILLER_ASAP7_75t_R FILLER_0_30_161 ();
 DECAPx1_ASAP7_75t_R FILLER_0_30_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_177 ();
 FILLER_ASAP7_75t_R FILLER_0_30_183 ();
 FILLER_ASAP7_75t_R FILLER_0_30_195 ();
 FILLER_ASAP7_75t_R FILLER_0_30_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_209 ();
 FILLER_ASAP7_75t_R FILLER_0_30_220 ();
 FILLER_ASAP7_75t_R FILLER_0_30_232 ();
 FILLER_ASAP7_75t_R FILLER_0_30_244 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_262 ();
 FILLER_ASAP7_75t_R FILLER_0_30_273 ();
 FILLER_ASAP7_75t_R FILLER_0_30_293 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_303 ();
 FILLER_ASAP7_75t_R FILLER_0_30_331 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_338 ();
 FILLER_ASAP7_75t_R FILLER_0_30_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_356 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_370 ();
 DECAPx1_ASAP7_75t_R FILLER_0_30_383 ();
 DECAPx1_ASAP7_75t_R FILLER_0_30_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_398 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_419 ();
 FILLER_ASAP7_75t_R FILLER_0_30_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_432 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_443 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_454 ();
 FILLER_ASAP7_75t_R FILLER_0_30_460 ();
 FILLER_ASAP7_75t_R FILLER_0_30_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_466 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_477 ();
 FILLER_ASAP7_75t_R FILLER_0_30_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_485 ();
 DECAPx6_ASAP7_75t_R FILLER_0_30_491 ();
 FILLER_ASAP7_75t_R FILLER_0_30_505 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_523 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_531 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_553 ();
 FILLER_ASAP7_75t_R FILLER_0_30_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_561 ();
 FILLER_ASAP7_75t_R FILLER_0_30_582 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_594 ();
 DECAPx4_ASAP7_75t_R FILLER_0_30_616 ();
 FILLER_ASAP7_75t_R FILLER_0_30_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_628 ();
 DECAPx1_ASAP7_75t_R FILLER_0_30_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_641 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_645 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_667 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_689 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_711 ();
 FILLER_ASAP7_75t_R FILLER_0_30_729 ();
 FILLER_ASAP7_75t_R FILLER_0_30_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_736 ();
 FILLER_ASAP7_75t_R FILLER_0_30_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_742 ();
 DECAPx4_ASAP7_75t_R FILLER_0_30_749 ();
 FILLER_ASAP7_75t_R FILLER_0_30_759 ();
 FILLER_ASAP7_75t_R FILLER_0_30_769 ();
 FILLER_ASAP7_75t_R FILLER_0_30_781 ();
 DECAPx6_ASAP7_75t_R FILLER_0_30_790 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_810 ();
 FILLER_ASAP7_75t_R FILLER_0_30_817 ();
 FILLER_ASAP7_75t_R FILLER_0_30_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_827 ();
 DECAPx1_ASAP7_75t_R FILLER_0_30_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_844 ();
 DECAPx1_ASAP7_75t_R FILLER_0_30_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_861 ();
 FILLER_ASAP7_75t_R FILLER_0_30_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_886 ();
 FILLER_ASAP7_75t_R FILLER_0_30_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_895 ();
 FILLER_ASAP7_75t_R FILLER_0_30_901 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_909 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_923 ();
 FILLER_ASAP7_75t_R FILLER_0_30_939 ();
 FILLER_ASAP7_75t_R FILLER_0_30_951 ();
 FILLER_ASAP7_75t_R FILLER_0_30_973 ();
 FILLER_ASAP7_75t_R FILLER_0_30_981 ();
 DECAPx1_ASAP7_75t_R FILLER_0_30_989 ();
 DECAPx4_ASAP7_75t_R FILLER_0_30_1003 ();
 FILLER_ASAP7_75t_R FILLER_0_30_1013 ();
 FILLER_ASAP7_75t_R FILLER_0_30_1021 ();
 DECAPx1_ASAP7_75t_R FILLER_0_30_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_1031 ();
 FILLER_ASAP7_75t_R FILLER_0_30_1043 ();
 FILLER_ASAP7_75t_R FILLER_0_30_1051 ();
 FILLER_ASAP7_75t_R FILLER_0_30_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_1067 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_1095 ();
 FILLER_ASAP7_75t_R FILLER_0_30_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_1110 ();
 FILLER_ASAP7_75t_R FILLER_0_30_1117 ();
 DECAPx4_ASAP7_75t_R FILLER_0_30_1130 ();
 FILLER_ASAP7_75t_R FILLER_0_30_1150 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_1161 ();
 FILLER_ASAP7_75t_R FILLER_0_30_1165 ();
 DECAPx1_ASAP7_75t_R FILLER_0_30_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_1182 ();
 FILLER_ASAP7_75t_R FILLER_0_30_1189 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_1198 ();
 DECAPx1_ASAP7_75t_R FILLER_0_30_1209 ();
 FILLER_ASAP7_75t_R FILLER_0_30_1224 ();
 FILLER_ASAP7_75t_R FILLER_0_30_1232 ();
 DECAPx4_ASAP7_75t_R FILLER_0_30_1240 ();
 FILLER_ASAP7_75t_R FILLER_0_30_1250 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_1252 ();
 FILLER_ASAP7_75t_R FILLER_0_30_1260 ();
 FILLER_ASAP7_75t_R FILLER_0_30_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_1295 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_1301 ();
 DECAPx4_ASAP7_75t_R FILLER_0_30_1308 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_1318 ();
 FILLER_ASAP7_75t_R FILLER_0_30_1325 ();
 FILLER_ASAP7_75t_R FILLER_0_30_1335 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_1343 ();
 FILLER_ASAP7_75t_R FILLER_0_30_1349 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_1351 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_1358 ();
 FILLER_ASAP7_75t_R FILLER_0_30_1370 ();
 DECAPx1_ASAP7_75t_R FILLER_0_30_1378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_46 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_53 ();
 DECAPx1_ASAP7_75t_R FILLER_0_31_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_69 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_78 ();
 FILLER_ASAP7_75t_R FILLER_0_31_84 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_92 ();
 FILLER_ASAP7_75t_R FILLER_0_31_98 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_112 ();
 DECAPx1_ASAP7_75t_R FILLER_0_31_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_123 ();
 FILLER_ASAP7_75t_R FILLER_0_31_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_136 ();
 FILLER_ASAP7_75t_R FILLER_0_31_147 ();
 FILLER_ASAP7_75t_R FILLER_0_31_155 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_173 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_186 ();
 FILLER_ASAP7_75t_R FILLER_0_31_192 ();
 FILLER_ASAP7_75t_R FILLER_0_31_200 ();
 FILLER_ASAP7_75t_R FILLER_0_31_208 ();
 FILLER_ASAP7_75t_R FILLER_0_31_220 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_238 ();
 FILLER_ASAP7_75t_R FILLER_0_31_249 ();
 FILLER_ASAP7_75t_R FILLER_0_31_261 ();
 FILLER_ASAP7_75t_R FILLER_0_31_273 ();
 FILLER_ASAP7_75t_R FILLER_0_31_293 ();
 FILLER_ASAP7_75t_R FILLER_0_31_303 ();
 FILLER_ASAP7_75t_R FILLER_0_31_311 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_319 ();
 FILLER_ASAP7_75t_R FILLER_0_31_333 ();
 DECAPx1_ASAP7_75t_R FILLER_0_31_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_349 ();
 DECAPx1_ASAP7_75t_R FILLER_0_31_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_360 ();
 FILLER_ASAP7_75t_R FILLER_0_31_367 ();
 DECAPx1_ASAP7_75t_R FILLER_0_31_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_379 ();
 FILLER_ASAP7_75t_R FILLER_0_31_392 ();
 DECAPx6_ASAP7_75t_R FILLER_0_31_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_418 ();
 FILLER_ASAP7_75t_R FILLER_0_31_429 ();
 DECAPx1_ASAP7_75t_R FILLER_0_31_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_440 ();
 DECAPx1_ASAP7_75t_R FILLER_0_31_447 ();
 FILLER_ASAP7_75t_R FILLER_0_31_456 ();
 FILLER_ASAP7_75t_R FILLER_0_31_463 ();
 DECAPx6_ASAP7_75t_R FILLER_0_31_469 ();
 FILLER_ASAP7_75t_R FILLER_0_31_483 ();
 FILLER_ASAP7_75t_R FILLER_0_31_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_495 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_502 ();
 DECAPx1_ASAP7_75t_R FILLER_0_31_514 ();
 FILLER_ASAP7_75t_R FILLER_0_31_525 ();
 DECAPx4_ASAP7_75t_R FILLER_0_31_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_545 ();
 FILLER_ASAP7_75t_R FILLER_0_31_552 ();
 FILLER_ASAP7_75t_R FILLER_0_31_561 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_566 ();
 FILLER_ASAP7_75t_R FILLER_0_31_572 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_584 ();
 FILLER_ASAP7_75t_R FILLER_0_31_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_600 ();
 FILLER_ASAP7_75t_R FILLER_0_31_622 ();
 FILLER_ASAP7_75t_R FILLER_0_31_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_632 ();
 FILLER_ASAP7_75t_R FILLER_0_31_641 ();
 FILLER_ASAP7_75t_R FILLER_0_31_654 ();
 FILLER_ASAP7_75t_R FILLER_0_31_668 ();
 DECAPx4_ASAP7_75t_R FILLER_0_31_678 ();
 FILLER_ASAP7_75t_R FILLER_0_31_694 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_708 ();
 DECAPx6_ASAP7_75t_R FILLER_0_31_720 ();
 FILLER_ASAP7_75t_R FILLER_0_31_734 ();
 FILLER_ASAP7_75t_R FILLER_0_31_746 ();
 FILLER_ASAP7_75t_R FILLER_0_31_759 ();
 FILLER_ASAP7_75t_R FILLER_0_31_767 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_811 ();
 DECAPx1_ASAP7_75t_R FILLER_0_31_820 ();
 DECAPx1_ASAP7_75t_R FILLER_0_31_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_836 ();
 DECAPx6_ASAP7_75t_R FILLER_0_31_843 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_863 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_867 ();
 FILLER_ASAP7_75t_R FILLER_0_31_893 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_901 ();
 FILLER_ASAP7_75t_R FILLER_0_31_915 ();
 FILLER_ASAP7_75t_R FILLER_0_31_923 ();
 FILLER_ASAP7_75t_R FILLER_0_31_927 ();
 FILLER_ASAP7_75t_R FILLER_0_31_939 ();
 FILLER_ASAP7_75t_R FILLER_0_31_951 ();
 FILLER_ASAP7_75t_R FILLER_0_31_963 ();
 FILLER_ASAP7_75t_R FILLER_0_31_971 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_978 ();
 FILLER_ASAP7_75t_R FILLER_0_31_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_986 ();
 DECAPx1_ASAP7_75t_R FILLER_0_31_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_1001 ();
 FILLER_ASAP7_75t_R FILLER_0_31_1012 ();
 FILLER_ASAP7_75t_R FILLER_0_31_1024 ();
 FILLER_ASAP7_75t_R FILLER_0_31_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_1034 ();
 DECAPx6_ASAP7_75t_R FILLER_0_31_1041 ();
 FILLER_ASAP7_75t_R FILLER_0_31_1055 ();
 DECAPx6_ASAP7_75t_R FILLER_0_31_1063 ();
 FILLER_ASAP7_75t_R FILLER_0_31_1077 ();
 FILLER_ASAP7_75t_R FILLER_0_31_1084 ();
 FILLER_ASAP7_75t_R FILLER_0_31_1092 ();
 FILLER_ASAP7_75t_R FILLER_0_31_1104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_1111 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_1139 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_1158 ();
 FILLER_ASAP7_75t_R FILLER_0_31_1165 ();
 FILLER_ASAP7_75t_R FILLER_0_31_1173 ();
 DECAPx1_ASAP7_75t_R FILLER_0_31_1180 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_1193 ();
 FILLER_ASAP7_75t_R FILLER_0_31_1205 ();
 FILLER_ASAP7_75t_R FILLER_0_31_1213 ();
 FILLER_ASAP7_75t_R FILLER_0_31_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_1223 ();
 DECAPx1_ASAP7_75t_R FILLER_0_31_1229 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_1233 ();
 DECAPx1_ASAP7_75t_R FILLER_0_31_1240 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_1255 ();
 FILLER_ASAP7_75t_R FILLER_0_31_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_1275 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_1297 ();
 FILLER_ASAP7_75t_R FILLER_0_31_1313 ();
 FILLER_ASAP7_75t_R FILLER_0_31_1321 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_1329 ();
 DECAPx6_ASAP7_75t_R FILLER_0_31_1338 ();
 DECAPx2_ASAP7_75t_R FILLER_0_31_1352 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_1358 ();
 FILLER_ASAP7_75t_R FILLER_0_31_1365 ();
 DECAPx1_ASAP7_75t_R FILLER_0_31_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_32_24 ();
 DECAPx1_ASAP7_75t_R FILLER_0_32_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_42 ();
 FILLER_ASAP7_75t_R FILLER_0_32_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_32_55 ();
 FILLER_ASAP7_75t_R FILLER_0_32_65 ();
 DECAPx2_ASAP7_75t_R FILLER_0_32_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_79 ();
 FILLER_ASAP7_75t_R FILLER_0_32_86 ();
 DECAPx2_ASAP7_75t_R FILLER_0_32_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_100 ();
 FILLER_ASAP7_75t_R FILLER_0_32_106 ();
 DECAPx2_ASAP7_75t_R FILLER_0_32_118 ();
 FILLER_ASAP7_75t_R FILLER_0_32_130 ();
 DECAPx2_ASAP7_75t_R FILLER_0_32_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_148 ();
 FILLER_ASAP7_75t_R FILLER_0_32_154 ();
 FILLER_ASAP7_75t_R FILLER_0_32_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_168 ();
 DECAPx2_ASAP7_75t_R FILLER_0_32_179 ();
 FILLER_ASAP7_75t_R FILLER_0_32_191 ();
 FILLER_ASAP7_75t_R FILLER_0_32_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_205 ();
 FILLER_ASAP7_75t_R FILLER_0_32_216 ();
 DECAPx2_ASAP7_75t_R FILLER_0_32_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_234 ();
 FILLER_ASAP7_75t_R FILLER_0_32_245 ();
 DECAPx1_ASAP7_75t_R FILLER_0_32_257 ();
 FILLER_ASAP7_75t_R FILLER_0_32_271 ();
 DECAPx1_ASAP7_75t_R FILLER_0_32_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_287 ();
 FILLER_ASAP7_75t_R FILLER_0_32_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_300 ();
 FILLER_ASAP7_75t_R FILLER_0_32_311 ();
 FILLER_ASAP7_75t_R FILLER_0_32_318 ();
 DECAPx1_ASAP7_75t_R FILLER_0_32_325 ();
 FILLER_ASAP7_75t_R FILLER_0_32_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_351 ();
 FILLER_ASAP7_75t_R FILLER_0_32_359 ();
 FILLER_ASAP7_75t_R FILLER_0_32_367 ();
 FILLER_ASAP7_75t_R FILLER_0_32_375 ();
 FILLER_ASAP7_75t_R FILLER_0_32_384 ();
 FILLER_ASAP7_75t_R FILLER_0_32_391 ();
 DECAPx2_ASAP7_75t_R FILLER_0_32_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_405 ();
 DECAPx1_ASAP7_75t_R FILLER_0_32_416 ();
 DECAPx2_ASAP7_75t_R FILLER_0_32_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_436 ();
 FILLER_ASAP7_75t_R FILLER_0_32_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_32_454 ();
 FILLER_ASAP7_75t_R FILLER_0_32_460 ();
 FILLER_ASAP7_75t_R FILLER_0_32_464 ();
 DECAPx1_ASAP7_75t_R FILLER_0_32_473 ();
 FILLER_ASAP7_75t_R FILLER_0_32_482 ();
 FILLER_ASAP7_75t_R FILLER_0_32_494 ();
 DECAPx2_ASAP7_75t_R FILLER_0_32_502 ();
 DECAPx4_ASAP7_75t_R FILLER_0_32_514 ();
 FILLER_ASAP7_75t_R FILLER_0_32_530 ();
 FILLER_ASAP7_75t_R FILLER_0_32_538 ();
 FILLER_ASAP7_75t_R FILLER_0_32_546 ();
 DECAPx1_ASAP7_75t_R FILLER_0_32_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_563 ();
 DECAPx6_ASAP7_75t_R FILLER_0_32_574 ();
 DECAPx2_ASAP7_75t_R FILLER_0_32_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_594 ();
 FILLER_ASAP7_75t_R FILLER_0_32_598 ();
 FILLER_ASAP7_75t_R FILLER_0_32_606 ();
 DECAPx4_ASAP7_75t_R FILLER_0_32_612 ();
 FILLER_ASAP7_75t_R FILLER_0_32_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_624 ();
 FILLER_ASAP7_75t_R FILLER_0_32_631 ();
 DECAPx1_ASAP7_75t_R FILLER_0_32_636 ();
 FILLER_ASAP7_75t_R FILLER_0_32_648 ();
 DECAPx1_ASAP7_75t_R FILLER_0_32_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_660 ();
 FILLER_ASAP7_75t_R FILLER_0_32_673 ();
 DECAPx4_ASAP7_75t_R FILLER_0_32_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_691 ();
 FILLER_ASAP7_75t_R FILLER_0_32_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_702 ();
 DECAPx6_ASAP7_75t_R FILLER_0_32_711 ();
 DECAPx2_ASAP7_75t_R FILLER_0_32_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_731 ();
 FILLER_ASAP7_75t_R FILLER_0_32_737 ();
 DECAPx6_ASAP7_75t_R FILLER_0_32_747 ();
 DECAPx2_ASAP7_75t_R FILLER_0_32_761 ();
 FILLER_ASAP7_75t_R FILLER_0_32_772 ();
 FILLER_ASAP7_75t_R FILLER_0_32_784 ();
 FILLER_ASAP7_75t_R FILLER_0_32_797 ();
 FILLER_ASAP7_75t_R FILLER_0_32_810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_822 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_844 ();
 DECAPx4_ASAP7_75t_R FILLER_0_32_866 ();
 FILLER_ASAP7_75t_R FILLER_0_32_876 ();
 DECAPx4_ASAP7_75t_R FILLER_0_32_886 ();
 DECAPx1_ASAP7_75t_R FILLER_0_32_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_906 ();
 FILLER_ASAP7_75t_R FILLER_0_32_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_915 ();
 FILLER_ASAP7_75t_R FILLER_0_32_926 ();
 FILLER_ASAP7_75t_R FILLER_0_32_934 ();
 DECAPx1_ASAP7_75t_R FILLER_0_32_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_946 ();
 DECAPx2_ASAP7_75t_R FILLER_0_32_952 ();
 FILLER_ASAP7_75t_R FILLER_0_32_972 ();
 FILLER_ASAP7_75t_R FILLER_0_32_984 ();
 DECAPx1_ASAP7_75t_R FILLER_0_32_992 ();
 FILLER_ASAP7_75t_R FILLER_0_32_1002 ();
 DECAPx2_ASAP7_75t_R FILLER_0_32_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_1015 ();
 FILLER_ASAP7_75t_R FILLER_0_32_1022 ();
 DECAPx6_ASAP7_75t_R FILLER_0_32_1030 ();
 DECAPx1_ASAP7_75t_R FILLER_0_32_1044 ();
 DECAPx1_ASAP7_75t_R FILLER_0_32_1056 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_1060 ();
 FILLER_ASAP7_75t_R FILLER_0_32_1067 ();
 FILLER_ASAP7_75t_R FILLER_0_32_1079 ();
 DECAPx6_ASAP7_75t_R FILLER_0_32_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_1101 ();
 FILLER_ASAP7_75t_R FILLER_0_32_1108 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_1117 ();
 DECAPx4_ASAP7_75t_R FILLER_0_32_1139 ();
 FILLER_ASAP7_75t_R FILLER_0_32_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_1151 ();
 FILLER_ASAP7_75t_R FILLER_0_32_1158 ();
 FILLER_ASAP7_75t_R FILLER_0_32_1163 ();
 FILLER_ASAP7_75t_R FILLER_0_32_1176 ();
 FILLER_ASAP7_75t_R FILLER_0_32_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_32_1194 ();
 FILLER_ASAP7_75t_R FILLER_0_32_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_1204 ();
 DECAPx6_ASAP7_75t_R FILLER_0_32_1215 ();
 DECAPx1_ASAP7_75t_R FILLER_0_32_1229 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_1245 ();
 DECAPx4_ASAP7_75t_R FILLER_0_32_1267 ();
 FILLER_ASAP7_75t_R FILLER_0_32_1277 ();
 FILLER_ASAP7_75t_R FILLER_0_32_1289 ();
 DECAPx2_ASAP7_75t_R FILLER_0_32_1296 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_1302 ();
 FILLER_ASAP7_75t_R FILLER_0_32_1316 ();
 DECAPx2_ASAP7_75t_R FILLER_0_32_1324 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32_1330 ();
 FILLER_ASAP7_75t_R FILLER_0_32_1337 ();
 DECAPx1_ASAP7_75t_R FILLER_0_32_1345 ();
 DECAPx4_ASAP7_75t_R FILLER_0_32_1352 ();
 DECAPx6_ASAP7_75t_R FILLER_0_32_1368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_33_24 ();
 FILLER_ASAP7_75t_R FILLER_0_33_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_36 ();
 FILLER_ASAP7_75t_R FILLER_0_33_43 ();
 DECAPx2_ASAP7_75t_R FILLER_0_33_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_57 ();
 DECAPx2_ASAP7_75t_R FILLER_0_33_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_70 ();
 DECAPx2_ASAP7_75t_R FILLER_0_33_78 ();
 FILLER_ASAP7_75t_R FILLER_0_33_90 ();
 DECAPx1_ASAP7_75t_R FILLER_0_33_98 ();
 FILLER_ASAP7_75t_R FILLER_0_33_107 ();
 FILLER_ASAP7_75t_R FILLER_0_33_119 ();
 DECAPx2_ASAP7_75t_R FILLER_0_33_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_137 ();
 DECAPx1_ASAP7_75t_R FILLER_0_33_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_148 ();
 FILLER_ASAP7_75t_R FILLER_0_33_159 ();
 FILLER_ASAP7_75t_R FILLER_0_33_171 ();
 FILLER_ASAP7_75t_R FILLER_0_33_183 ();
 FILLER_ASAP7_75t_R FILLER_0_33_211 ();
 FILLER_ASAP7_75t_R FILLER_0_33_223 ();
 FILLER_ASAP7_75t_R FILLER_0_33_233 ();
 DECAPx2_ASAP7_75t_R FILLER_0_33_245 ();
 DECAPx2_ASAP7_75t_R FILLER_0_33_257 ();
 FILLER_ASAP7_75t_R FILLER_0_33_273 ();
 FILLER_ASAP7_75t_R FILLER_0_33_285 ();
 FILLER_ASAP7_75t_R FILLER_0_33_297 ();
 DECAPx2_ASAP7_75t_R FILLER_0_33_309 ();
 FILLER_ASAP7_75t_R FILLER_0_33_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_322 ();
 FILLER_ASAP7_75t_R FILLER_0_33_329 ();
 FILLER_ASAP7_75t_R FILLER_0_33_337 ();
 FILLER_ASAP7_75t_R FILLER_0_33_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_349 ();
 FILLER_ASAP7_75t_R FILLER_0_33_356 ();
 FILLER_ASAP7_75t_R FILLER_0_33_364 ();
 FILLER_ASAP7_75t_R FILLER_0_33_372 ();
 FILLER_ASAP7_75t_R FILLER_0_33_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_381 ();
 FILLER_ASAP7_75t_R FILLER_0_33_388 ();
 DECAPx1_ASAP7_75t_R FILLER_0_33_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_400 ();
 FILLER_ASAP7_75t_R FILLER_0_33_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_413 ();
 FILLER_ASAP7_75t_R FILLER_0_33_424 ();
 DECAPx2_ASAP7_75t_R FILLER_0_33_432 ();
 FILLER_ASAP7_75t_R FILLER_0_33_444 ();
 FILLER_ASAP7_75t_R FILLER_0_33_456 ();
 FILLER_ASAP7_75t_R FILLER_0_33_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_465 ();
 FILLER_ASAP7_75t_R FILLER_0_33_474 ();
 DECAPx1_ASAP7_75t_R FILLER_0_33_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_487 ();
 FILLER_ASAP7_75t_R FILLER_0_33_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_496 ();
 FILLER_ASAP7_75t_R FILLER_0_33_503 ();
 DECAPx6_ASAP7_75t_R FILLER_0_33_511 ();
 FILLER_ASAP7_75t_R FILLER_0_33_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_527 ();
 DECAPx2_ASAP7_75t_R FILLER_0_33_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_540 ();
 FILLER_ASAP7_75t_R FILLER_0_33_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_548 ();
 FILLER_ASAP7_75t_R FILLER_0_33_555 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_563 ();
 DECAPx2_ASAP7_75t_R FILLER_0_33_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_591 ();
 DECAPx6_ASAP7_75t_R FILLER_0_33_604 ();
 DECAPx1_ASAP7_75t_R FILLER_0_33_618 ();
 DECAPx6_ASAP7_75t_R FILLER_0_33_627 ();
 FILLER_ASAP7_75t_R FILLER_0_33_647 ();
 DECAPx2_ASAP7_75t_R FILLER_0_33_661 ();
 FILLER_ASAP7_75t_R FILLER_0_33_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_669 ();
 FILLER_ASAP7_75t_R FILLER_0_33_676 ();
 FILLER_ASAP7_75t_R FILLER_0_33_681 ();
 DECAPx1_ASAP7_75t_R FILLER_0_33_695 ();
 FILLER_ASAP7_75t_R FILLER_0_33_705 ();
 DECAPx6_ASAP7_75t_R FILLER_0_33_713 ();
 DECAPx2_ASAP7_75t_R FILLER_0_33_727 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_744 ();
 DECAPx2_ASAP7_75t_R FILLER_0_33_766 ();
 FILLER_ASAP7_75t_R FILLER_0_33_778 ();
 FILLER_ASAP7_75t_R FILLER_0_33_786 ();
 DECAPx2_ASAP7_75t_R FILLER_0_33_794 ();
 FILLER_ASAP7_75t_R FILLER_0_33_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_802 ();
 FILLER_ASAP7_75t_R FILLER_0_33_815 ();
 DECAPx6_ASAP7_75t_R FILLER_0_33_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_837 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_844 ();
 DECAPx2_ASAP7_75t_R FILLER_0_33_866 ();
 FILLER_ASAP7_75t_R FILLER_0_33_882 ();
 DECAPx4_ASAP7_75t_R FILLER_0_33_891 ();
 DECAPx4_ASAP7_75t_R FILLER_0_33_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_917 ();
 FILLER_ASAP7_75t_R FILLER_0_33_923 ();
 FILLER_ASAP7_75t_R FILLER_0_33_927 ();
 FILLER_ASAP7_75t_R FILLER_0_33_935 ();
 DECAPx1_ASAP7_75t_R FILLER_0_33_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_946 ();
 FILLER_ASAP7_75t_R FILLER_0_33_957 ();
 DECAPx6_ASAP7_75t_R FILLER_0_33_970 ();
 FILLER_ASAP7_75t_R FILLER_0_33_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_986 ();
 FILLER_ASAP7_75t_R FILLER_0_33_1001 ();
 DECAPx1_ASAP7_75t_R FILLER_0_33_1013 ();
 DECAPx1_ASAP7_75t_R FILLER_0_33_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_1031 ();
 DECAPx4_ASAP7_75t_R FILLER_0_33_1039 ();
 FILLER_ASAP7_75t_R FILLER_0_33_1049 ();
 FILLER_ASAP7_75t_R FILLER_0_33_1056 ();
 FILLER_ASAP7_75t_R FILLER_0_33_1068 ();
 DECAPx1_ASAP7_75t_R FILLER_0_33_1082 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_1086 ();
 FILLER_ASAP7_75t_R FILLER_0_33_1090 ();
 DECAPx1_ASAP7_75t_R FILLER_0_33_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_1104 ();
 DECAPx1_ASAP7_75t_R FILLER_0_33_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_1122 ();
 FILLER_ASAP7_75t_R FILLER_0_33_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_1146 ();
 DECAPx2_ASAP7_75t_R FILLER_0_33_1158 ();
 FILLER_ASAP7_75t_R FILLER_0_33_1164 ();
 FILLER_ASAP7_75t_R FILLER_0_33_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_1182 ();
 DECAPx6_ASAP7_75t_R FILLER_0_33_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_1218 ();
 DECAPx1_ASAP7_75t_R FILLER_0_33_1225 ();
 DECAPx4_ASAP7_75t_R FILLER_0_33_1235 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33_1245 ();
 DECAPx1_ASAP7_75t_R FILLER_0_33_1256 ();
 FILLER_ASAP7_75t_R FILLER_0_33_1270 ();
 FILLER_ASAP7_75t_R FILLER_0_33_1278 ();
 FILLER_ASAP7_75t_R FILLER_0_33_1286 ();
 FILLER_ASAP7_75t_R FILLER_0_33_1294 ();
 FILLER_ASAP7_75t_R FILLER_0_33_1302 ();
 DECAPx2_ASAP7_75t_R FILLER_0_33_1310 ();
 FILLER_ASAP7_75t_R FILLER_0_33_1316 ();
 FILLER_ASAP7_75t_R FILLER_0_33_1328 ();
 DECAPx2_ASAP7_75t_R FILLER_0_33_1338 ();
 FILLER_ASAP7_75t_R FILLER_0_33_1347 ();
 DECAPx1_ASAP7_75t_R FILLER_0_33_1355 ();
 DECAPx4_ASAP7_75t_R FILLER_0_33_1370 ();
 FILLER_ASAP7_75t_R FILLER_0_33_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_24 ();
 FILLER_ASAP7_75t_R FILLER_0_34_31 ();
 FILLER_ASAP7_75t_R FILLER_0_34_39 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_47 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_69 ();
 DECAPx2_ASAP7_75t_R FILLER_0_34_91 ();
 FILLER_ASAP7_75t_R FILLER_0_34_97 ();
 FILLER_ASAP7_75t_R FILLER_0_34_104 ();
 FILLER_ASAP7_75t_R FILLER_0_34_111 ();
 FILLER_ASAP7_75t_R FILLER_0_34_119 ();
 FILLER_ASAP7_75t_R FILLER_0_34_131 ();
 DECAPx2_ASAP7_75t_R FILLER_0_34_143 ();
 FILLER_ASAP7_75t_R FILLER_0_34_155 ();
 FILLER_ASAP7_75t_R FILLER_0_34_165 ();
 FILLER_ASAP7_75t_R FILLER_0_34_177 ();
 FILLER_ASAP7_75t_R FILLER_0_34_189 ();
 FILLER_ASAP7_75t_R FILLER_0_34_196 ();
 DECAPx1_ASAP7_75t_R FILLER_0_34_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_210 ();
 FILLER_ASAP7_75t_R FILLER_0_34_218 ();
 FILLER_ASAP7_75t_R FILLER_0_34_228 ();
 FILLER_ASAP7_75t_R FILLER_0_34_240 ();
 FILLER_ASAP7_75t_R FILLER_0_34_248 ();
 DECAPx2_ASAP7_75t_R FILLER_0_34_261 ();
 DECAPx2_ASAP7_75t_R FILLER_0_34_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_281 ();
 FILLER_ASAP7_75t_R FILLER_0_34_292 ();
 FILLER_ASAP7_75t_R FILLER_0_34_304 ();
 DECAPx1_ASAP7_75t_R FILLER_0_34_316 ();
 DECAPx2_ASAP7_75t_R FILLER_0_34_323 ();
 FILLER_ASAP7_75t_R FILLER_0_34_334 ();
 FILLER_ASAP7_75t_R FILLER_0_34_346 ();
 FILLER_ASAP7_75t_R FILLER_0_34_358 ();
 FILLER_ASAP7_75t_R FILLER_0_34_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_370 ();
 FILLER_ASAP7_75t_R FILLER_0_34_381 ();
 FILLER_ASAP7_75t_R FILLER_0_34_388 ();
 FILLER_ASAP7_75t_R FILLER_0_34_397 ();
 DECAPx1_ASAP7_75t_R FILLER_0_34_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_413 ();
 DECAPx1_ASAP7_75t_R FILLER_0_34_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_428 ();
 FILLER_ASAP7_75t_R FILLER_0_34_436 ();
 DECAPx2_ASAP7_75t_R FILLER_0_34_448 ();
 FILLER_ASAP7_75t_R FILLER_0_34_460 ();
 FILLER_ASAP7_75t_R FILLER_0_34_464 ();
 FILLER_ASAP7_75t_R FILLER_0_34_476 ();
 DECAPx1_ASAP7_75t_R FILLER_0_34_485 ();
 DECAPx2_ASAP7_75t_R FILLER_0_34_495 ();
 FILLER_ASAP7_75t_R FILLER_0_34_501 ();
 FILLER_ASAP7_75t_R FILLER_0_34_508 ();
 DECAPx2_ASAP7_75t_R FILLER_0_34_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_526 ();
 FILLER_ASAP7_75t_R FILLER_0_34_533 ();
 DECAPx4_ASAP7_75t_R FILLER_0_34_541 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_572 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_594 ();
 FILLER_ASAP7_75t_R FILLER_0_34_616 ();
 FILLER_ASAP7_75t_R FILLER_0_34_630 ();
 DECAPx6_ASAP7_75t_R FILLER_0_34_644 ();
 FILLER_ASAP7_75t_R FILLER_0_34_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_660 ();
 FILLER_ASAP7_75t_R FILLER_0_34_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_668 ();
 DECAPx4_ASAP7_75t_R FILLER_0_34_681 ();
 FILLER_ASAP7_75t_R FILLER_0_34_697 ();
 DECAPx6_ASAP7_75t_R FILLER_0_34_711 ();
 DECAPx2_ASAP7_75t_R FILLER_0_34_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_731 ();
 FILLER_ASAP7_75t_R FILLER_0_34_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_737 ();
 DECAPx1_ASAP7_75t_R FILLER_0_34_744 ();
 FILLER_ASAP7_75t_R FILLER_0_34_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_762 ();
 DECAPx1_ASAP7_75t_R FILLER_0_34_769 ();
 FILLER_ASAP7_75t_R FILLER_0_34_776 ();
 FILLER_ASAP7_75t_R FILLER_0_34_786 ();
 DECAPx4_ASAP7_75t_R FILLER_0_34_796 ();
 FILLER_ASAP7_75t_R FILLER_0_34_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_808 ();
 FILLER_ASAP7_75t_R FILLER_0_34_815 ();
 FILLER_ASAP7_75t_R FILLER_0_34_823 ();
 FILLER_ASAP7_75t_R FILLER_0_34_831 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_839 ();
 DECAPx6_ASAP7_75t_R FILLER_0_34_861 ();
 FILLER_ASAP7_75t_R FILLER_0_34_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_877 ();
 FILLER_ASAP7_75t_R FILLER_0_34_888 ();
 FILLER_ASAP7_75t_R FILLER_0_34_896 ();
 FILLER_ASAP7_75t_R FILLER_0_34_904 ();
 FILLER_ASAP7_75t_R FILLER_0_34_912 ();
 FILLER_ASAP7_75t_R FILLER_0_34_919 ();
 DECAPx2_ASAP7_75t_R FILLER_0_34_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_932 ();
 DECAPx1_ASAP7_75t_R FILLER_0_34_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_943 ();
 FILLER_ASAP7_75t_R FILLER_0_34_955 ();
 FILLER_ASAP7_75t_R FILLER_0_34_963 ();
 DECAPx4_ASAP7_75t_R FILLER_0_34_968 ();
 FILLER_ASAP7_75t_R FILLER_0_34_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_980 ();
 DECAPx2_ASAP7_75t_R FILLER_0_34_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_994 ();
 DECAPx6_ASAP7_75t_R FILLER_0_34_1001 ();
 DECAPx2_ASAP7_75t_R FILLER_0_34_1015 ();
 FILLER_ASAP7_75t_R FILLER_0_34_1027 ();
 DECAPx2_ASAP7_75t_R FILLER_0_34_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_1046 ();
 DECAPx2_ASAP7_75t_R FILLER_0_34_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_1060 ();
 DECAPx1_ASAP7_75t_R FILLER_0_34_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_1070 ();
 FILLER_ASAP7_75t_R FILLER_0_34_1083 ();
 FILLER_ASAP7_75t_R FILLER_0_34_1095 ();
 DECAPx1_ASAP7_75t_R FILLER_0_34_1107 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_1131 ();
 DECAPx2_ASAP7_75t_R FILLER_0_34_1159 ();
 FILLER_ASAP7_75t_R FILLER_0_34_1165 ();
 FILLER_ASAP7_75t_R FILLER_0_34_1173 ();
 DECAPx6_ASAP7_75t_R FILLER_0_34_1180 ();
 FILLER_ASAP7_75t_R FILLER_0_34_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_1196 ();
 DECAPx1_ASAP7_75t_R FILLER_0_34_1203 ();
 FILLER_ASAP7_75t_R FILLER_0_34_1217 ();
 FILLER_ASAP7_75t_R FILLER_0_34_1230 ();
 FILLER_ASAP7_75t_R FILLER_0_34_1235 ();
 FILLER_ASAP7_75t_R FILLER_0_34_1243 ();
 DECAPx4_ASAP7_75t_R FILLER_0_34_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_0_34_1275 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_1289 ();
 FILLER_ASAP7_75t_R FILLER_0_34_1296 ();
 DECAPx1_ASAP7_75t_R FILLER_0_34_1304 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_1308 ();
 DECAPx1_ASAP7_75t_R FILLER_0_34_1315 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_1319 ();
 DECAPx2_ASAP7_75t_R FILLER_0_34_1330 ();
 FILLER_ASAP7_75t_R FILLER_0_34_1336 ();
 DECAPx4_ASAP7_75t_R FILLER_0_34_1344 ();
 FILLER_ASAP7_75t_R FILLER_0_34_1354 ();
 FILLER_ASAP7_75t_R FILLER_0_34_1362 ();
 DECAPx6_ASAP7_75t_R FILLER_0_34_1367 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_35_24 ();
 FILLER_ASAP7_75t_R FILLER_0_35_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_36 ();
 FILLER_ASAP7_75t_R FILLER_0_35_42 ();
 DECAPx1_ASAP7_75t_R FILLER_0_35_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_58 ();
 DECAPx6_ASAP7_75t_R FILLER_0_35_65 ();
 DECAPx1_ASAP7_75t_R FILLER_0_35_79 ();
 DECAPx1_ASAP7_75t_R FILLER_0_35_89 ();
 DECAPx1_ASAP7_75t_R FILLER_0_35_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_103 ();
 DECAPx1_ASAP7_75t_R FILLER_0_35_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_114 ();
 DECAPx1_ASAP7_75t_R FILLER_0_35_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_125 ();
 FILLER_ASAP7_75t_R FILLER_0_35_132 ();
 FILLER_ASAP7_75t_R FILLER_0_35_139 ();
 FILLER_ASAP7_75t_R FILLER_0_35_149 ();
 FILLER_ASAP7_75t_R FILLER_0_35_154 ();
 FILLER_ASAP7_75t_R FILLER_0_35_168 ();
 FILLER_ASAP7_75t_R FILLER_0_35_180 ();
 DECAPx1_ASAP7_75t_R FILLER_0_35_192 ();
 DECAPx2_ASAP7_75t_R FILLER_0_35_206 ();
 FILLER_ASAP7_75t_R FILLER_0_35_212 ();
 FILLER_ASAP7_75t_R FILLER_0_35_221 ();
 FILLER_ASAP7_75t_R FILLER_0_35_230 ();
 FILLER_ASAP7_75t_R FILLER_0_35_237 ();
 FILLER_ASAP7_75t_R FILLER_0_35_245 ();
 FILLER_ASAP7_75t_R FILLER_0_35_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_259 ();
 DECAPx1_ASAP7_75t_R FILLER_0_35_266 ();
 FILLER_ASAP7_75t_R FILLER_0_35_277 ();
 FILLER_ASAP7_75t_R FILLER_0_35_289 ();
 FILLER_ASAP7_75t_R FILLER_0_35_295 ();
 DECAPx4_ASAP7_75t_R FILLER_0_35_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_317 ();
 FILLER_ASAP7_75t_R FILLER_0_35_323 ();
 FILLER_ASAP7_75t_R FILLER_0_35_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_337 ();
 FILLER_ASAP7_75t_R FILLER_0_35_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_350 ();
 FILLER_ASAP7_75t_R FILLER_0_35_361 ();
 DECAPx1_ASAP7_75t_R FILLER_0_35_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_373 ();
 FILLER_ASAP7_75t_R FILLER_0_35_384 ();
 DECAPx2_ASAP7_75t_R FILLER_0_35_394 ();
 FILLER_ASAP7_75t_R FILLER_0_35_400 ();
 FILLER_ASAP7_75t_R FILLER_0_35_412 ();
 DECAPx2_ASAP7_75t_R FILLER_0_35_422 ();
 DECAPx1_ASAP7_75t_R FILLER_0_35_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_438 ();
 FILLER_ASAP7_75t_R FILLER_0_35_445 ();
 FILLER_ASAP7_75t_R FILLER_0_35_457 ();
 FILLER_ASAP7_75t_R FILLER_0_35_469 ();
 FILLER_ASAP7_75t_R FILLER_0_35_481 ();
 DECAPx1_ASAP7_75t_R FILLER_0_35_489 ();
 DECAPx2_ASAP7_75t_R FILLER_0_35_499 ();
 DECAPx2_ASAP7_75t_R FILLER_0_35_513 ();
 DECAPx2_ASAP7_75t_R FILLER_0_35_525 ();
 DECAPx1_ASAP7_75t_R FILLER_0_35_542 ();
 FILLER_ASAP7_75t_R FILLER_0_35_552 ();
 FILLER_ASAP7_75t_R FILLER_0_35_560 ();
 FILLER_ASAP7_75t_R FILLER_0_35_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_570 ();
 FILLER_ASAP7_75t_R FILLER_0_35_581 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_589 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_611 ();
 DECAPx2_ASAP7_75t_R FILLER_0_35_644 ();
 DECAPx6_ASAP7_75t_R FILLER_0_35_671 ();
 DECAPx1_ASAP7_75t_R FILLER_0_35_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_689 ();
 DECAPx6_ASAP7_75t_R FILLER_0_35_694 ();
 DECAPx1_ASAP7_75t_R FILLER_0_35_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_712 ();
 FILLER_ASAP7_75t_R FILLER_0_35_719 ();
 FILLER_ASAP7_75t_R FILLER_0_35_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_727 ();
 FILLER_ASAP7_75t_R FILLER_0_35_734 ();
 DECAPx4_ASAP7_75t_R FILLER_0_35_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_752 ();
 DECAPx1_ASAP7_75t_R FILLER_0_35_765 ();
 FILLER_ASAP7_75t_R FILLER_0_35_777 ();
 DECAPx2_ASAP7_75t_R FILLER_0_35_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_788 ();
 DECAPx4_ASAP7_75t_R FILLER_0_35_797 ();
 FILLER_ASAP7_75t_R FILLER_0_35_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_809 ();
 DECAPx1_ASAP7_75t_R FILLER_0_35_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_826 ();
 FILLER_ASAP7_75t_R FILLER_0_35_835 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_845 ();
 DECAPx1_ASAP7_75t_R FILLER_0_35_867 ();
 FILLER_ASAP7_75t_R FILLER_0_35_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_879 ();
 FILLER_ASAP7_75t_R FILLER_0_35_890 ();
 FILLER_ASAP7_75t_R FILLER_0_35_898 ();
 DECAPx2_ASAP7_75t_R FILLER_0_35_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_912 ();
 DECAPx2_ASAP7_75t_R FILLER_0_35_919 ();
 DECAPx2_ASAP7_75t_R FILLER_0_35_927 ();
 DECAPx6_ASAP7_75t_R FILLER_0_35_939 ();
 FILLER_ASAP7_75t_R FILLER_0_35_953 ();
 FILLER_ASAP7_75t_R FILLER_0_35_961 ();
 FILLER_ASAP7_75t_R FILLER_0_35_973 ();
 FILLER_ASAP7_75t_R FILLER_0_35_987 ();
 FILLER_ASAP7_75t_R FILLER_0_35_996 ();
 DECAPx6_ASAP7_75t_R FILLER_0_35_1004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_1023 ();
 FILLER_ASAP7_75t_R FILLER_0_35_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_1047 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_1054 ();
 DECAPx1_ASAP7_75t_R FILLER_0_35_1076 ();
 DECAPx2_ASAP7_75t_R FILLER_0_35_1088 ();
 FILLER_ASAP7_75t_R FILLER_0_35_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_1096 ();
 DECAPx2_ASAP7_75t_R FILLER_0_35_1102 ();
 FILLER_ASAP7_75t_R FILLER_0_35_1111 ();
 DECAPx4_ASAP7_75t_R FILLER_0_35_1123 ();
 FILLER_ASAP7_75t_R FILLER_0_35_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_1135 ();
 FILLER_ASAP7_75t_R FILLER_0_35_1142 ();
 FILLER_ASAP7_75t_R FILLER_0_35_1147 ();
 DECAPx6_ASAP7_75t_R FILLER_0_35_1152 ();
 FILLER_ASAP7_75t_R FILLER_0_35_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_1177 ();
 FILLER_ASAP7_75t_R FILLER_0_35_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_1201 ();
 FILLER_ASAP7_75t_R FILLER_0_35_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_1209 ();
 DECAPx2_ASAP7_75t_R FILLER_0_35_1217 ();
 FILLER_ASAP7_75t_R FILLER_0_35_1229 ();
 DECAPx1_ASAP7_75t_R FILLER_0_35_1237 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_1241 ();
 DECAPx2_ASAP7_75t_R FILLER_0_35_1254 ();
 FILLER_ASAP7_75t_R FILLER_0_35_1260 ();
 DECAPx4_ASAP7_75t_R FILLER_0_35_1274 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_1284 ();
 FILLER_ASAP7_75t_R FILLER_0_35_1291 ();
 DECAPx2_ASAP7_75t_R FILLER_0_35_1299 ();
 DECAPx6_ASAP7_75t_R FILLER_0_35_1325 ();
 DECAPx1_ASAP7_75t_R FILLER_0_35_1339 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_1343 ();
 FILLER_ASAP7_75t_R FILLER_0_35_1347 ();
 DECAPx2_ASAP7_75t_R FILLER_0_35_1355 ();
 FILLER_ASAP7_75t_R FILLER_0_35_1361 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_1363 ();
 DECAPx4_ASAP7_75t_R FILLER_0_35_1370 ();
 FILLER_ASAP7_75t_R FILLER_0_35_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_36_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_28 ();
 FILLER_ASAP7_75t_R FILLER_0_36_35 ();
 FILLER_ASAP7_75t_R FILLER_0_36_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_45 ();
 DECAPx1_ASAP7_75t_R FILLER_0_36_52 ();
 DECAPx1_ASAP7_75t_R FILLER_0_36_67 ();
 FILLER_ASAP7_75t_R FILLER_0_36_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_87 ();
 FILLER_ASAP7_75t_R FILLER_0_36_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_96 ();
 DECAPx1_ASAP7_75t_R FILLER_0_36_100 ();
 DECAPx1_ASAP7_75t_R FILLER_0_36_112 ();
 FILLER_ASAP7_75t_R FILLER_0_36_123 ();
 FILLER_ASAP7_75t_R FILLER_0_36_145 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_152 ();
 FILLER_ASAP7_75t_R FILLER_0_36_170 ();
 FILLER_ASAP7_75t_R FILLER_0_36_177 ();
 FILLER_ASAP7_75t_R FILLER_0_36_184 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_198 ();
 DECAPx1_ASAP7_75t_R FILLER_0_36_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_209 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_217 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_230 ();
 FILLER_ASAP7_75t_R FILLER_0_36_242 ();
 FILLER_ASAP7_75t_R FILLER_0_36_250 ();
 DECAPx1_ASAP7_75t_R FILLER_0_36_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_262 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_275 ();
 DECAPx1_ASAP7_75t_R FILLER_0_36_282 ();
 FILLER_ASAP7_75t_R FILLER_0_36_296 ();
 FILLER_ASAP7_75t_R FILLER_0_36_303 ();
 DECAPx6_ASAP7_75t_R FILLER_0_36_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_323 ();
 FILLER_ASAP7_75t_R FILLER_0_36_329 ();
 FILLER_ASAP7_75t_R FILLER_0_36_337 ();
 FILLER_ASAP7_75t_R FILLER_0_36_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_351 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_362 ();
 FILLER_ASAP7_75t_R FILLER_0_36_378 ();
 DECAPx1_ASAP7_75t_R FILLER_0_36_390 ();
 FILLER_ASAP7_75t_R FILLER_0_36_404 ();
 FILLER_ASAP7_75t_R FILLER_0_36_416 ();
 FILLER_ASAP7_75t_R FILLER_0_36_426 ();
 FILLER_ASAP7_75t_R FILLER_0_36_434 ();
 FILLER_ASAP7_75t_R FILLER_0_36_446 ();
 FILLER_ASAP7_75t_R FILLER_0_36_454 ();
 FILLER_ASAP7_75t_R FILLER_0_36_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_461 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_470 ();
 FILLER_ASAP7_75t_R FILLER_0_36_481 ();
 FILLER_ASAP7_75t_R FILLER_0_36_488 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_496 ();
 FILLER_ASAP7_75t_R FILLER_0_36_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_504 ();
 DECAPx1_ASAP7_75t_R FILLER_0_36_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_515 ();
 FILLER_ASAP7_75t_R FILLER_0_36_522 ();
 FILLER_ASAP7_75t_R FILLER_0_36_530 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_539 ();
 FILLER_ASAP7_75t_R FILLER_0_36_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_547 ();
 FILLER_ASAP7_75t_R FILLER_0_36_554 ();
 FILLER_ASAP7_75t_R FILLER_0_36_562 ();
 FILLER_ASAP7_75t_R FILLER_0_36_570 ();
 FILLER_ASAP7_75t_R FILLER_0_36_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_577 ();
 FILLER_ASAP7_75t_R FILLER_0_36_581 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_591 ();
 FILLER_ASAP7_75t_R FILLER_0_36_597 ();
 DECAPx1_ASAP7_75t_R FILLER_0_36_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_615 ();
 DECAPx4_ASAP7_75t_R FILLER_0_36_627 ();
 FILLER_ASAP7_75t_R FILLER_0_36_642 ();
 FILLER_ASAP7_75t_R FILLER_0_36_655 ();
 DECAPx4_ASAP7_75t_R FILLER_0_36_660 ();
 DECAPx6_ASAP7_75t_R FILLER_0_36_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_696 ();
 FILLER_ASAP7_75t_R FILLER_0_36_705 ();
 FILLER_ASAP7_75t_R FILLER_0_36_718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_730 ();
 FILLER_ASAP7_75t_R FILLER_0_36_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_754 ();
 DECAPx1_ASAP7_75t_R FILLER_0_36_761 ();
 DECAPx1_ASAP7_75t_R FILLER_0_36_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_775 ();
 DECAPx1_ASAP7_75t_R FILLER_0_36_784 ();
 DECAPx6_ASAP7_75t_R FILLER_0_36_791 ();
 FILLER_ASAP7_75t_R FILLER_0_36_805 ();
 FILLER_ASAP7_75t_R FILLER_0_36_819 ();
 FILLER_ASAP7_75t_R FILLER_0_36_827 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_837 ();
 FILLER_ASAP7_75t_R FILLER_0_36_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_845 ();
 FILLER_ASAP7_75t_R FILLER_0_36_867 ();
 FILLER_ASAP7_75t_R FILLER_0_36_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_877 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_889 ();
 FILLER_ASAP7_75t_R FILLER_0_36_895 ();
 FILLER_ASAP7_75t_R FILLER_0_36_903 ();
 FILLER_ASAP7_75t_R FILLER_0_36_911 ();
 FILLER_ASAP7_75t_R FILLER_0_36_919 ();
 FILLER_ASAP7_75t_R FILLER_0_36_931 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_940 ();
 FILLER_ASAP7_75t_R FILLER_0_36_956 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_972 ();
 FILLER_ASAP7_75t_R FILLER_0_36_984 ();
 DECAPx4_ASAP7_75t_R FILLER_0_36_993 ();
 FILLER_ASAP7_75t_R FILLER_0_36_1003 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_1015 ();
 DECAPx6_ASAP7_75t_R FILLER_0_36_1028 ();
 FILLER_ASAP7_75t_R FILLER_0_36_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_1044 ();
 FILLER_ASAP7_75t_R FILLER_0_36_1051 ();
 FILLER_ASAP7_75t_R FILLER_0_36_1059 ();
 FILLER_ASAP7_75t_R FILLER_0_36_1067 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_1075 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_1093 ();
 FILLER_ASAP7_75t_R FILLER_0_36_1100 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_1108 ();
 DECAPx6_ASAP7_75t_R FILLER_0_36_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_1144 ();
 FILLER_ASAP7_75t_R FILLER_0_36_1151 ();
 DECAPx4_ASAP7_75t_R FILLER_0_36_1163 ();
 FILLER_ASAP7_75t_R FILLER_0_36_1173 ();
 FILLER_ASAP7_75t_R FILLER_0_36_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_1183 ();
 DECAPx1_ASAP7_75t_R FILLER_0_36_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_1194 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_1207 ();
 DECAPx1_ASAP7_75t_R FILLER_0_36_1219 ();
 DECAPx6_ASAP7_75t_R FILLER_0_36_1229 ();
 DECAPx1_ASAP7_75t_R FILLER_0_36_1243 ();
 DECAPx1_ASAP7_75t_R FILLER_0_36_1253 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_1257 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_1264 ();
 DECAPx4_ASAP7_75t_R FILLER_0_36_1286 ();
 FILLER_ASAP7_75t_R FILLER_0_36_1302 ();
 FILLER_ASAP7_75t_R FILLER_0_36_1309 ();
 DECAPx1_ASAP7_75t_R FILLER_0_36_1317 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_1321 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_1333 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_1339 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_1346 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_1352 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_1356 ();
 FILLER_ASAP7_75t_R FILLER_0_36_1368 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_37_24 ();
 FILLER_ASAP7_75t_R FILLER_0_37_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_32 ();
 DECAPx1_ASAP7_75t_R FILLER_0_37_44 ();
 FILLER_ASAP7_75t_R FILLER_0_37_54 ();
 FILLER_ASAP7_75t_R FILLER_0_37_62 ();
 FILLER_ASAP7_75t_R FILLER_0_37_70 ();
 FILLER_ASAP7_75t_R FILLER_0_37_82 ();
 DECAPx1_ASAP7_75t_R FILLER_0_37_90 ();
 DECAPx1_ASAP7_75t_R FILLER_0_37_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_104 ();
 FILLER_ASAP7_75t_R FILLER_0_37_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_113 ();
 DECAPx1_ASAP7_75t_R FILLER_0_37_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_124 ();
 FILLER_ASAP7_75t_R FILLER_0_37_131 ();
 FILLER_ASAP7_75t_R FILLER_0_37_139 ();
 DECAPx2_ASAP7_75t_R FILLER_0_37_148 ();
 FILLER_ASAP7_75t_R FILLER_0_37_159 ();
 FILLER_ASAP7_75t_R FILLER_0_37_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_173 ();
 FILLER_ASAP7_75t_R FILLER_0_37_179 ();
 FILLER_ASAP7_75t_R FILLER_0_37_191 ();
 FILLER_ASAP7_75t_R FILLER_0_37_199 ();
 DECAPx1_ASAP7_75t_R FILLER_0_37_207 ();
 DECAPx2_ASAP7_75t_R FILLER_0_37_219 ();
 FILLER_ASAP7_75t_R FILLER_0_37_225 ();
 FILLER_ASAP7_75t_R FILLER_0_37_233 ();
 FILLER_ASAP7_75t_R FILLER_0_37_241 ();
 FILLER_ASAP7_75t_R FILLER_0_37_248 ();
 DECAPx4_ASAP7_75t_R FILLER_0_37_253 ();
 FILLER_ASAP7_75t_R FILLER_0_37_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_265 ();
 FILLER_ASAP7_75t_R FILLER_0_37_286 ();
 FILLER_ASAP7_75t_R FILLER_0_37_298 ();
 DECAPx6_ASAP7_75t_R FILLER_0_37_306 ();
 FILLER_ASAP7_75t_R FILLER_0_37_320 ();
 FILLER_ASAP7_75t_R FILLER_0_37_327 ();
 FILLER_ASAP7_75t_R FILLER_0_37_334 ();
 FILLER_ASAP7_75t_R FILLER_0_37_342 ();
 FILLER_ASAP7_75t_R FILLER_0_37_354 ();
 FILLER_ASAP7_75t_R FILLER_0_37_366 ();
 FILLER_ASAP7_75t_R FILLER_0_37_378 ();
 FILLER_ASAP7_75t_R FILLER_0_37_390 ();
 FILLER_ASAP7_75t_R FILLER_0_37_400 ();
 FILLER_ASAP7_75t_R FILLER_0_37_420 ();
 FILLER_ASAP7_75t_R FILLER_0_37_428 ();
 FILLER_ASAP7_75t_R FILLER_0_37_434 ();
 FILLER_ASAP7_75t_R FILLER_0_37_443 ();
 FILLER_ASAP7_75t_R FILLER_0_37_449 ();
 DECAPx4_ASAP7_75t_R FILLER_0_37_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_467 ();
 FILLER_ASAP7_75t_R FILLER_0_37_473 ();
 FILLER_ASAP7_75t_R FILLER_0_37_486 ();
 DECAPx4_ASAP7_75t_R FILLER_0_37_495 ();
 DECAPx6_ASAP7_75t_R FILLER_0_37_513 ();
 DECAPx1_ASAP7_75t_R FILLER_0_37_527 ();
 FILLER_ASAP7_75t_R FILLER_0_37_538 ();
 DECAPx6_ASAP7_75t_R FILLER_0_37_547 ();
 DECAPx2_ASAP7_75t_R FILLER_0_37_561 ();
 DECAPx2_ASAP7_75t_R FILLER_0_37_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_579 ();
 FILLER_ASAP7_75t_R FILLER_0_37_583 ();
 DECAPx1_ASAP7_75t_R FILLER_0_37_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_600 ();
 FILLER_ASAP7_75t_R FILLER_0_37_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_606 ();
 FILLER_ASAP7_75t_R FILLER_0_37_615 ();
 FILLER_ASAP7_75t_R FILLER_0_37_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_622 ();
 DECAPx6_ASAP7_75t_R FILLER_0_37_626 ();
 FILLER_ASAP7_75t_R FILLER_0_37_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_649 ();
 FILLER_ASAP7_75t_R FILLER_0_37_671 ();
 DECAPx1_ASAP7_75t_R FILLER_0_37_679 ();
 DECAPx1_ASAP7_75t_R FILLER_0_37_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_695 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_706 ();
 DECAPx2_ASAP7_75t_R FILLER_0_37_728 ();
 FILLER_ASAP7_75t_R FILLER_0_37_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_736 ();
 DECAPx1_ASAP7_75t_R FILLER_0_37_741 ();
 DECAPx6_ASAP7_75t_R FILLER_0_37_755 ();
 DECAPx2_ASAP7_75t_R FILLER_0_37_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_775 ();
 DECAPx2_ASAP7_75t_R FILLER_0_37_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_793 ();
 FILLER_ASAP7_75t_R FILLER_0_37_806 ();
 FILLER_ASAP7_75t_R FILLER_0_37_814 ();
 DECAPx2_ASAP7_75t_R FILLER_0_37_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_830 ();
 DECAPx1_ASAP7_75t_R FILLER_0_37_839 ();
 FILLER_ASAP7_75t_R FILLER_0_37_846 ();
 DECAPx6_ASAP7_75t_R FILLER_0_37_856 ();
 FILLER_ASAP7_75t_R FILLER_0_37_870 ();
 FILLER_ASAP7_75t_R FILLER_0_37_884 ();
 DECAPx2_ASAP7_75t_R FILLER_0_37_892 ();
 FILLER_ASAP7_75t_R FILLER_0_37_898 ();
 DECAPx2_ASAP7_75t_R FILLER_0_37_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_916 ();
 FILLER_ASAP7_75t_R FILLER_0_37_923 ();
 DECAPx1_ASAP7_75t_R FILLER_0_37_927 ();
 FILLER_ASAP7_75t_R FILLER_0_37_942 ();
 DECAPx2_ASAP7_75t_R FILLER_0_37_950 ();
 FILLER_ASAP7_75t_R FILLER_0_37_966 ();
 FILLER_ASAP7_75t_R FILLER_0_37_976 ();
 FILLER_ASAP7_75t_R FILLER_0_37_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_985 ();
 FILLER_ASAP7_75t_R FILLER_0_37_992 ();
 DECAPx1_ASAP7_75t_R FILLER_0_37_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_1004 ();
 FILLER_ASAP7_75t_R FILLER_0_37_1015 ();
 FILLER_ASAP7_75t_R FILLER_0_37_1027 ();
 DECAPx2_ASAP7_75t_R FILLER_0_37_1039 ();
 FILLER_ASAP7_75t_R FILLER_0_37_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_1047 ();
 FILLER_ASAP7_75t_R FILLER_0_37_1054 ();
 DECAPx4_ASAP7_75t_R FILLER_0_37_1063 ();
 FILLER_ASAP7_75t_R FILLER_0_37_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_1075 ();
 FILLER_ASAP7_75t_R FILLER_0_37_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_0_37_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_1102 ();
 DECAPx2_ASAP7_75t_R FILLER_0_37_1124 ();
 FILLER_ASAP7_75t_R FILLER_0_37_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_1132 ();
 DECAPx2_ASAP7_75t_R FILLER_0_37_1139 ();
 FILLER_ASAP7_75t_R FILLER_0_37_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_1147 ();
 FILLER_ASAP7_75t_R FILLER_0_37_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_1170 ();
 FILLER_ASAP7_75t_R FILLER_0_37_1177 ();
 DECAPx4_ASAP7_75t_R FILLER_0_37_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_37_1203 ();
 FILLER_ASAP7_75t_R FILLER_0_37_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_1223 ();
 DECAPx1_ASAP7_75t_R FILLER_0_37_1245 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_1249 ();
 FILLER_ASAP7_75t_R FILLER_0_37_1253 ();
 FILLER_ASAP7_75t_R FILLER_0_37_1262 ();
 DECAPx4_ASAP7_75t_R FILLER_0_37_1275 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_1285 ();
 FILLER_ASAP7_75t_R FILLER_0_37_1296 ();
 DECAPx1_ASAP7_75t_R FILLER_0_37_1304 ();
 DECAPx2_ASAP7_75t_R FILLER_0_37_1313 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_1319 ();
 FILLER_ASAP7_75t_R FILLER_0_37_1326 ();
 FILLER_ASAP7_75t_R FILLER_0_37_1333 ();
 FILLER_ASAP7_75t_R FILLER_0_37_1339 ();
 FILLER_ASAP7_75t_R FILLER_0_37_1347 ();
 DECAPx2_ASAP7_75t_R FILLER_0_37_1355 ();
 FILLER_ASAP7_75t_R FILLER_0_37_1361 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_1363 ();
 FILLER_ASAP7_75t_R FILLER_0_37_1370 ();
 DECAPx1_ASAP7_75t_R FILLER_0_37_1378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_38_24 ();
 FILLER_ASAP7_75t_R FILLER_0_38_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_32 ();
 FILLER_ASAP7_75t_R FILLER_0_38_39 ();
 DECAPx4_ASAP7_75t_R FILLER_0_38_47 ();
 DECAPx1_ASAP7_75t_R FILLER_0_38_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_67 ();
 FILLER_ASAP7_75t_R FILLER_0_38_73 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_81 ();
 DECAPx6_ASAP7_75t_R FILLER_0_38_103 ();
 DECAPx2_ASAP7_75t_R FILLER_0_38_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_123 ();
 FILLER_ASAP7_75t_R FILLER_0_38_129 ();
 FILLER_ASAP7_75t_R FILLER_0_38_136 ();
 DECAPx2_ASAP7_75t_R FILLER_0_38_148 ();
 FILLER_ASAP7_75t_R FILLER_0_38_154 ();
 FILLER_ASAP7_75t_R FILLER_0_38_164 ();
 DECAPx2_ASAP7_75t_R FILLER_0_38_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_182 ();
 FILLER_ASAP7_75t_R FILLER_0_38_193 ();
 FILLER_ASAP7_75t_R FILLER_0_38_206 ();
 DECAPx1_ASAP7_75t_R FILLER_0_38_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_217 ();
 FILLER_ASAP7_75t_R FILLER_0_38_224 ();
 DECAPx2_ASAP7_75t_R FILLER_0_38_232 ();
 FILLER_ASAP7_75t_R FILLER_0_38_244 ();
 DECAPx2_ASAP7_75t_R FILLER_0_38_254 ();
 FILLER_ASAP7_75t_R FILLER_0_38_260 ();
 FILLER_ASAP7_75t_R FILLER_0_38_268 ();
 FILLER_ASAP7_75t_R FILLER_0_38_278 ();
 FILLER_ASAP7_75t_R FILLER_0_38_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_288 ();
 FILLER_ASAP7_75t_R FILLER_0_38_299 ();
 FILLER_ASAP7_75t_R FILLER_0_38_309 ();
 DECAPx2_ASAP7_75t_R FILLER_0_38_316 ();
 FILLER_ASAP7_75t_R FILLER_0_38_322 ();
 FILLER_ASAP7_75t_R FILLER_0_38_329 ();
 FILLER_ASAP7_75t_R FILLER_0_38_361 ();
 FILLER_ASAP7_75t_R FILLER_0_38_371 ();
 FILLER_ASAP7_75t_R FILLER_0_38_383 ();
 FILLER_ASAP7_75t_R FILLER_0_38_395 ();
 DECAPx1_ASAP7_75t_R FILLER_0_38_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_411 ();
 FILLER_ASAP7_75t_R FILLER_0_38_418 ();
 FILLER_ASAP7_75t_R FILLER_0_38_426 ();
 FILLER_ASAP7_75t_R FILLER_0_38_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_438 ();
 DECAPx2_ASAP7_75t_R FILLER_0_38_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_451 ();
 FILLER_ASAP7_75t_R FILLER_0_38_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_461 ();
 DECAPx2_ASAP7_75t_R FILLER_0_38_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_470 ();
 FILLER_ASAP7_75t_R FILLER_0_38_481 ();
 FILLER_ASAP7_75t_R FILLER_0_38_489 ();
 DECAPx2_ASAP7_75t_R FILLER_0_38_497 ();
 DECAPx1_ASAP7_75t_R FILLER_0_38_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_527 ();
 DECAPx1_ASAP7_75t_R FILLER_0_38_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_552 ();
 DECAPx1_ASAP7_75t_R FILLER_0_38_559 ();
 DECAPx6_ASAP7_75t_R FILLER_0_38_573 ();
 FILLER_ASAP7_75t_R FILLER_0_38_595 ();
 FILLER_ASAP7_75t_R FILLER_0_38_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_607 ();
 FILLER_ASAP7_75t_R FILLER_0_38_619 ();
 FILLER_ASAP7_75t_R FILLER_0_38_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_629 ();
 DECAPx1_ASAP7_75t_R FILLER_0_38_642 ();
 DECAPx1_ASAP7_75t_R FILLER_0_38_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_656 ();
 DECAPx2_ASAP7_75t_R FILLER_0_38_668 ();
 FILLER_ASAP7_75t_R FILLER_0_38_681 ();
 DECAPx1_ASAP7_75t_R FILLER_0_38_695 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_699 ();
 FILLER_ASAP7_75t_R FILLER_0_38_711 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_719 ();
 FILLER_ASAP7_75t_R FILLER_0_38_752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_758 ();
 FILLER_ASAP7_75t_R FILLER_0_38_780 ();
 FILLER_ASAP7_75t_R FILLER_0_38_785 ();
 DECAPx6_ASAP7_75t_R FILLER_0_38_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_809 ();
 DECAPx6_ASAP7_75t_R FILLER_0_38_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_834 ();
 FILLER_ASAP7_75t_R FILLER_0_38_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_847 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_851 ();
 FILLER_ASAP7_75t_R FILLER_0_38_879 ();
 FILLER_ASAP7_75t_R FILLER_0_38_887 ();
 DECAPx1_ASAP7_75t_R FILLER_0_38_895 ();
 FILLER_ASAP7_75t_R FILLER_0_38_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_907 ();
 FILLER_ASAP7_75t_R FILLER_0_38_914 ();
 DECAPx4_ASAP7_75t_R FILLER_0_38_923 ();
 FILLER_ASAP7_75t_R FILLER_0_38_933 ();
 DECAPx2_ASAP7_75t_R FILLER_0_38_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_947 ();
 FILLER_ASAP7_75t_R FILLER_0_38_954 ();
 FILLER_ASAP7_75t_R FILLER_0_38_959 ();
 FILLER_ASAP7_75t_R FILLER_0_38_971 ();
 DECAPx1_ASAP7_75t_R FILLER_0_38_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_983 ();
 DECAPx2_ASAP7_75t_R FILLER_0_38_990 ();
 FILLER_ASAP7_75t_R FILLER_0_38_1007 ();
 FILLER_ASAP7_75t_R FILLER_0_38_1014 ();
 DECAPx2_ASAP7_75t_R FILLER_0_38_1022 ();
 DECAPx1_ASAP7_75t_R FILLER_0_38_1034 ();
 FILLER_ASAP7_75t_R FILLER_0_38_1044 ();
 FILLER_ASAP7_75t_R FILLER_0_38_1056 ();
 FILLER_ASAP7_75t_R FILLER_0_38_1064 ();
 FILLER_ASAP7_75t_R FILLER_0_38_1072 ();
 FILLER_ASAP7_75t_R FILLER_0_38_1084 ();
 FILLER_ASAP7_75t_R FILLER_0_38_1092 ();
 FILLER_ASAP7_75t_R FILLER_0_38_1100 ();
 DECAPx6_ASAP7_75t_R FILLER_0_38_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_1122 ();
 FILLER_ASAP7_75t_R FILLER_0_38_1133 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_1141 ();
 DECAPx2_ASAP7_75t_R FILLER_0_38_1163 ();
 FILLER_ASAP7_75t_R FILLER_0_38_1169 ();
 FILLER_ASAP7_75t_R FILLER_0_38_1178 ();
 FILLER_ASAP7_75t_R FILLER_0_38_1186 ();
 DECAPx6_ASAP7_75t_R FILLER_0_38_1194 ();
 FILLER_ASAP7_75t_R FILLER_0_38_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_1210 ();
 FILLER_ASAP7_75t_R FILLER_0_38_1217 ();
 FILLER_ASAP7_75t_R FILLER_0_38_1222 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_1224 ();
 FILLER_ASAP7_75t_R FILLER_0_38_1231 ();
 DECAPx1_ASAP7_75t_R FILLER_0_38_1244 ();
 DECAPx2_ASAP7_75t_R FILLER_0_38_1256 ();
 DECAPx6_ASAP7_75t_R FILLER_0_38_1273 ();
 FILLER_ASAP7_75t_R FILLER_0_38_1287 ();
 FILLER_ASAP7_75t_R FILLER_0_38_1309 ();
 FILLER_ASAP7_75t_R FILLER_0_38_1317 ();
 FILLER_ASAP7_75t_R FILLER_0_38_1325 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_1327 ();
 DECAPx1_ASAP7_75t_R FILLER_0_38_1334 ();
 DECAPx2_ASAP7_75t_R FILLER_0_38_1348 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_1354 ();
 FILLER_ASAP7_75t_R FILLER_0_38_1361 ();
 FILLER_ASAP7_75t_R FILLER_0_38_1369 ();
 DECAPx1_ASAP7_75t_R FILLER_0_38_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_24 ();
 DECAPx1_ASAP7_75t_R FILLER_0_39_52 ();
 DECAPx1_ASAP7_75t_R FILLER_0_39_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_66 ();
 FILLER_ASAP7_75t_R FILLER_0_39_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_72 ();
 DECAPx1_ASAP7_75t_R FILLER_0_39_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_83 ();
 DECAPx2_ASAP7_75t_R FILLER_0_39_94 ();
 FILLER_ASAP7_75t_R FILLER_0_39_100 ();
 FILLER_ASAP7_75t_R FILLER_0_39_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_116 ();
 DECAPx4_ASAP7_75t_R FILLER_0_39_124 ();
 DECAPx6_ASAP7_75t_R FILLER_0_39_141 ();
 FILLER_ASAP7_75t_R FILLER_0_39_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_157 ();
 FILLER_ASAP7_75t_R FILLER_0_39_168 ();
 FILLER_ASAP7_75t_R FILLER_0_39_180 ();
 FILLER_ASAP7_75t_R FILLER_0_39_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_190 ();
 DECAPx1_ASAP7_75t_R FILLER_0_39_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_203 ();
 FILLER_ASAP7_75t_R FILLER_0_39_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_212 ();
 FILLER_ASAP7_75t_R FILLER_0_39_219 ();
 DECAPx1_ASAP7_75t_R FILLER_0_39_227 ();
 FILLER_ASAP7_75t_R FILLER_0_39_241 ();
 DECAPx4_ASAP7_75t_R FILLER_0_39_249 ();
 FILLER_ASAP7_75t_R FILLER_0_39_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_269 ();
 FILLER_ASAP7_75t_R FILLER_0_39_276 ();
 DECAPx2_ASAP7_75t_R FILLER_0_39_286 ();
 FILLER_ASAP7_75t_R FILLER_0_39_292 ();
 FILLER_ASAP7_75t_R FILLER_0_39_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_306 ();
 FILLER_ASAP7_75t_R FILLER_0_39_345 ();
 FILLER_ASAP7_75t_R FILLER_0_39_355 ();
 FILLER_ASAP7_75t_R FILLER_0_39_367 ();
 FILLER_ASAP7_75t_R FILLER_0_39_378 ();
 FILLER_ASAP7_75t_R FILLER_0_39_390 ();
 FILLER_ASAP7_75t_R FILLER_0_39_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_401 ();
 FILLER_ASAP7_75t_R FILLER_0_39_412 ();
 DECAPx2_ASAP7_75t_R FILLER_0_39_420 ();
 FILLER_ASAP7_75t_R FILLER_0_39_432 ();
 DECAPx4_ASAP7_75t_R FILLER_0_39_439 ();
 FILLER_ASAP7_75t_R FILLER_0_39_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_451 ();
 DECAPx2_ASAP7_75t_R FILLER_0_39_458 ();
 FILLER_ASAP7_75t_R FILLER_0_39_464 ();
 DECAPx2_ASAP7_75t_R FILLER_0_39_472 ();
 FILLER_ASAP7_75t_R FILLER_0_39_484 ();
 DECAPx4_ASAP7_75t_R FILLER_0_39_492 ();
 FILLER_ASAP7_75t_R FILLER_0_39_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_504 ();
 DECAPx6_ASAP7_75t_R FILLER_0_39_515 ();
 FILLER_ASAP7_75t_R FILLER_0_39_529 ();
 DECAPx6_ASAP7_75t_R FILLER_0_39_537 ();
 FILLER_ASAP7_75t_R FILLER_0_39_551 ();
 DECAPx4_ASAP7_75t_R FILLER_0_39_559 ();
 DECAPx2_ASAP7_75t_R FILLER_0_39_579 ();
 FILLER_ASAP7_75t_R FILLER_0_39_585 ();
 DECAPx6_ASAP7_75t_R FILLER_0_39_593 ();
 DECAPx1_ASAP7_75t_R FILLER_0_39_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_611 ();
 FILLER_ASAP7_75t_R FILLER_0_39_615 ();
 FILLER_ASAP7_75t_R FILLER_0_39_628 ();
 DECAPx6_ASAP7_75t_R FILLER_0_39_641 ();
 DECAPx1_ASAP7_75t_R FILLER_0_39_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_659 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_668 ();
 DECAPx6_ASAP7_75t_R FILLER_0_39_690 ();
 DECAPx2_ASAP7_75t_R FILLER_0_39_704 ();
 FILLER_ASAP7_75t_R FILLER_0_39_731 ();
 DECAPx2_ASAP7_75t_R FILLER_0_39_744 ();
 FILLER_ASAP7_75t_R FILLER_0_39_760 ();
 DECAPx4_ASAP7_75t_R FILLER_0_39_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_775 ();
 DECAPx6_ASAP7_75t_R FILLER_0_39_796 ();
 FILLER_ASAP7_75t_R FILLER_0_39_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_812 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_821 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_855 ();
 FILLER_ASAP7_75t_R FILLER_0_39_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_879 ();
 DECAPx4_ASAP7_75t_R FILLER_0_39_886 ();
 FILLER_ASAP7_75t_R FILLER_0_39_902 ();
 DECAPx2_ASAP7_75t_R FILLER_0_39_909 ();
 FILLER_ASAP7_75t_R FILLER_0_39_915 ();
 FILLER_ASAP7_75t_R FILLER_0_39_923 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_927 ();
 FILLER_ASAP7_75t_R FILLER_0_39_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_951 ();
 DECAPx2_ASAP7_75t_R FILLER_0_39_958 ();
 FILLER_ASAP7_75t_R FILLER_0_39_964 ();
 FILLER_ASAP7_75t_R FILLER_0_39_972 ();
 FILLER_ASAP7_75t_R FILLER_0_39_980 ();
 DECAPx4_ASAP7_75t_R FILLER_0_39_988 ();
 FILLER_ASAP7_75t_R FILLER_0_39_998 ();
 DECAPx4_ASAP7_75t_R FILLER_0_39_1008 ();
 FILLER_ASAP7_75t_R FILLER_0_39_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_1020 ();
 FILLER_ASAP7_75t_R FILLER_0_39_1027 ();
 DECAPx2_ASAP7_75t_R FILLER_0_39_1035 ();
 FILLER_ASAP7_75t_R FILLER_0_39_1041 ();
 DECAPx2_ASAP7_75t_R FILLER_0_39_1049 ();
 FILLER_ASAP7_75t_R FILLER_0_39_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_0_39_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_1069 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_1076 ();
 FILLER_ASAP7_75t_R FILLER_0_39_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_1100 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_1107 ();
 DECAPx2_ASAP7_75t_R FILLER_0_39_1129 ();
 FILLER_ASAP7_75t_R FILLER_0_39_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_1137 ();
 DECAPx4_ASAP7_75t_R FILLER_0_39_1141 ();
 FILLER_ASAP7_75t_R FILLER_0_39_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_1153 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_1164 ();
 DECAPx6_ASAP7_75t_R FILLER_0_39_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_39_1200 ();
 FILLER_ASAP7_75t_R FILLER_0_39_1208 ();
 FILLER_ASAP7_75t_R FILLER_0_39_1216 ();
 FILLER_ASAP7_75t_R FILLER_0_39_1223 ();
 FILLER_ASAP7_75t_R FILLER_0_39_1233 ();
 FILLER_ASAP7_75t_R FILLER_0_39_1241 ();
 DECAPx1_ASAP7_75t_R FILLER_0_39_1254 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_1258 ();
 FILLER_ASAP7_75t_R FILLER_0_39_1266 ();
 DECAPx4_ASAP7_75t_R FILLER_0_39_1275 ();
 FILLER_ASAP7_75t_R FILLER_0_39_1285 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_1287 ();
 FILLER_ASAP7_75t_R FILLER_0_39_1298 ();
 FILLER_ASAP7_75t_R FILLER_0_39_1307 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_1309 ();
 FILLER_ASAP7_75t_R FILLER_0_39_1318 ();
 DECAPx1_ASAP7_75t_R FILLER_0_39_1326 ();
 DECAPx6_ASAP7_75t_R FILLER_0_39_1341 ();
 FILLER_ASAP7_75t_R FILLER_0_39_1355 ();
 FILLER_ASAP7_75t_R FILLER_0_39_1363 ();
 DECAPx4_ASAP7_75t_R FILLER_0_39_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_24 ();
 FILLER_ASAP7_75t_R FILLER_0_40_30 ();
 DECAPx6_ASAP7_75t_R FILLER_0_40_38 ();
 FILLER_ASAP7_75t_R FILLER_0_40_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_54 ();
 FILLER_ASAP7_75t_R FILLER_0_40_61 ();
 FILLER_ASAP7_75t_R FILLER_0_40_69 ();
 FILLER_ASAP7_75t_R FILLER_0_40_77 ();
 DECAPx6_ASAP7_75t_R FILLER_0_40_90 ();
 DECAPx1_ASAP7_75t_R FILLER_0_40_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_120 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_127 ();
 FILLER_ASAP7_75t_R FILLER_0_40_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_135 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_148 ();
 FILLER_ASAP7_75t_R FILLER_0_40_155 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_167 ();
 FILLER_ASAP7_75t_R FILLER_0_40_173 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_191 ();
 DECAPx1_ASAP7_75t_R FILLER_0_40_198 ();
 FILLER_ASAP7_75t_R FILLER_0_40_208 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_222 ();
 DECAPx1_ASAP7_75t_R FILLER_0_40_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_238 ();
 DECAPx1_ASAP7_75t_R FILLER_0_40_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_253 ();
 DECAPx1_ASAP7_75t_R FILLER_0_40_261 ();
 FILLER_ASAP7_75t_R FILLER_0_40_271 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_283 ();
 FILLER_ASAP7_75t_R FILLER_0_40_289 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_303 ();
 FILLER_ASAP7_75t_R FILLER_0_40_315 ();
 FILLER_ASAP7_75t_R FILLER_0_40_327 ();
 FILLER_ASAP7_75t_R FILLER_0_40_339 ();
 FILLER_ASAP7_75t_R FILLER_0_40_351 ();
 FILLER_ASAP7_75t_R FILLER_0_40_363 ();
 FILLER_ASAP7_75t_R FILLER_0_40_370 ();
 FILLER_ASAP7_75t_R FILLER_0_40_382 ();
 FILLER_ASAP7_75t_R FILLER_0_40_392 ();
 FILLER_ASAP7_75t_R FILLER_0_40_404 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_422 ();
 FILLER_ASAP7_75t_R FILLER_0_40_429 ();
 DECAPx4_ASAP7_75t_R FILLER_0_40_437 ();
 FILLER_ASAP7_75t_R FILLER_0_40_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_449 ();
 FILLER_ASAP7_75t_R FILLER_0_40_460 ();
 FILLER_ASAP7_75t_R FILLER_0_40_464 ();
 FILLER_ASAP7_75t_R FILLER_0_40_472 ();
 FILLER_ASAP7_75t_R FILLER_0_40_485 ();
 DECAPx6_ASAP7_75t_R FILLER_0_40_497 ();
 DECAPx1_ASAP7_75t_R FILLER_0_40_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_515 ();
 DECAPx6_ASAP7_75t_R FILLER_0_40_526 ();
 FILLER_ASAP7_75t_R FILLER_0_40_560 ();
 DECAPx1_ASAP7_75t_R FILLER_0_40_582 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_596 ();
 DECAPx4_ASAP7_75t_R FILLER_0_40_629 ();
 FILLER_ASAP7_75t_R FILLER_0_40_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_641 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_645 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_651 ();
 DECAPx1_ASAP7_75t_R FILLER_0_40_660 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_670 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_694 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_703 ();
 FILLER_ASAP7_75t_R FILLER_0_40_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_711 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_721 ();
 DECAPx4_ASAP7_75t_R FILLER_0_40_734 ();
 FILLER_ASAP7_75t_R FILLER_0_40_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_746 ();
 FILLER_ASAP7_75t_R FILLER_0_40_755 ();
 DECAPx1_ASAP7_75t_R FILLER_0_40_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_767 ();
 DECAPx4_ASAP7_75t_R FILLER_0_40_772 ();
 DECAPx6_ASAP7_75t_R FILLER_0_40_792 ();
 FILLER_ASAP7_75t_R FILLER_0_40_806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_816 ();
 DECAPx6_ASAP7_75t_R FILLER_0_40_838 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_861 ();
 DECAPx4_ASAP7_75t_R FILLER_0_40_883 ();
 FILLER_ASAP7_75t_R FILLER_0_40_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_895 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_902 ();
 DECAPx1_ASAP7_75t_R FILLER_0_40_924 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_928 ();
 FILLER_ASAP7_75t_R FILLER_0_40_935 ();
 DECAPx4_ASAP7_75t_R FILLER_0_40_943 ();
 DECAPx6_ASAP7_75t_R FILLER_0_40_963 ();
 FILLER_ASAP7_75t_R FILLER_0_40_977 ();
 DECAPx6_ASAP7_75t_R FILLER_0_40_985 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_999 ();
 FILLER_ASAP7_75t_R FILLER_0_40_1015 ();
 DECAPx4_ASAP7_75t_R FILLER_0_40_1025 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_1040 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_1062 ();
 FILLER_ASAP7_75t_R FILLER_0_40_1074 ();
 FILLER_ASAP7_75t_R FILLER_0_40_1082 ();
 DECAPx4_ASAP7_75t_R FILLER_0_40_1090 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_1100 ();
 FILLER_ASAP7_75t_R FILLER_0_40_1107 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_1115 ();
 FILLER_ASAP7_75t_R FILLER_0_40_1121 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_1126 ();
 DECAPx1_ASAP7_75t_R FILLER_0_40_1138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_1148 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_1160 ();
 DECAPx1_ASAP7_75t_R FILLER_0_40_1176 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_1180 ();
 FILLER_ASAP7_75t_R FILLER_0_40_1187 ();
 FILLER_ASAP7_75t_R FILLER_0_40_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_1197 ();
 FILLER_ASAP7_75t_R FILLER_0_40_1204 ();
 FILLER_ASAP7_75t_R FILLER_0_40_1214 ();
 FILLER_ASAP7_75t_R FILLER_0_40_1222 ();
 FILLER_ASAP7_75t_R FILLER_0_40_1230 ();
 FILLER_ASAP7_75t_R FILLER_0_40_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_1240 ();
 DECAPx4_ASAP7_75t_R FILLER_0_40_1247 ();
 FILLER_ASAP7_75t_R FILLER_0_40_1257 ();
 DECAPx4_ASAP7_75t_R FILLER_0_40_1266 ();
 FILLER_ASAP7_75t_R FILLER_0_40_1276 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_1278 ();
 FILLER_ASAP7_75t_R FILLER_0_40_1284 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_1294 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_1300 ();
 FILLER_ASAP7_75t_R FILLER_0_40_1307 ();
 FILLER_ASAP7_75t_R FILLER_0_40_1321 ();
 FILLER_ASAP7_75t_R FILLER_0_40_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_1337 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_1359 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_41_24 ();
 DECAPx1_ASAP7_75t_R FILLER_0_41_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_42 ();
 FILLER_ASAP7_75t_R FILLER_0_41_49 ();
 FILLER_ASAP7_75t_R FILLER_0_41_57 ();
 DECAPx4_ASAP7_75t_R FILLER_0_41_65 ();
 FILLER_ASAP7_75t_R FILLER_0_41_75 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_105 ();
 DECAPx1_ASAP7_75t_R FILLER_0_41_113 ();
 FILLER_ASAP7_75t_R FILLER_0_41_129 ();
 FILLER_ASAP7_75t_R FILLER_0_41_137 ();
 FILLER_ASAP7_75t_R FILLER_0_41_145 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_154 ();
 FILLER_ASAP7_75t_R FILLER_0_41_170 ();
 FILLER_ASAP7_75t_R FILLER_0_41_182 ();
 FILLER_ASAP7_75t_R FILLER_0_41_192 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_201 ();
 FILLER_ASAP7_75t_R FILLER_0_41_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_217 ();
 FILLER_ASAP7_75t_R FILLER_0_41_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_226 ();
 FILLER_ASAP7_75t_R FILLER_0_41_233 ();
 DECAPx1_ASAP7_75t_R FILLER_0_41_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_245 ();
 DECAPx1_ASAP7_75t_R FILLER_0_41_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_260 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_273 ();
 FILLER_ASAP7_75t_R FILLER_0_41_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_286 ();
 FILLER_ASAP7_75t_R FILLER_0_41_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_299 ();
 FILLER_ASAP7_75t_R FILLER_0_41_303 ();
 FILLER_ASAP7_75t_R FILLER_0_41_313 ();
 FILLER_ASAP7_75t_R FILLER_0_41_325 ();
 FILLER_ASAP7_75t_R FILLER_0_41_337 ();
 FILLER_ASAP7_75t_R FILLER_0_41_349 ();
 FILLER_ASAP7_75t_R FILLER_0_41_361 ();
 FILLER_ASAP7_75t_R FILLER_0_41_373 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_391 ();
 FILLER_ASAP7_75t_R FILLER_0_41_402 ();
 DECAPx1_ASAP7_75t_R FILLER_0_41_414 ();
 FILLER_ASAP7_75t_R FILLER_0_41_424 ();
 FILLER_ASAP7_75t_R FILLER_0_41_432 ();
 FILLER_ASAP7_75t_R FILLER_0_41_440 ();
 FILLER_ASAP7_75t_R FILLER_0_41_448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_466 ();
 DECAPx4_ASAP7_75t_R FILLER_0_41_470 ();
 FILLER_ASAP7_75t_R FILLER_0_41_480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_487 ();
 DECAPx4_ASAP7_75t_R FILLER_0_41_509 ();
 FILLER_ASAP7_75t_R FILLER_0_41_519 ();
 FILLER_ASAP7_75t_R FILLER_0_41_527 ();
 FILLER_ASAP7_75t_R FILLER_0_41_535 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_543 ();
 DECAPx6_ASAP7_75t_R FILLER_0_41_565 ();
 FILLER_ASAP7_75t_R FILLER_0_41_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_581 ();
 FILLER_ASAP7_75t_R FILLER_0_41_593 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_607 ();
 DECAPx4_ASAP7_75t_R FILLER_0_41_629 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_647 ();
 FILLER_ASAP7_75t_R FILLER_0_41_664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_671 ();
 DECAPx1_ASAP7_75t_R FILLER_0_41_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_705 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_718 ();
 DECAPx1_ASAP7_75t_R FILLER_0_41_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_744 ();
 FILLER_ASAP7_75t_R FILLER_0_41_753 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_763 ();
 DECAPx6_ASAP7_75t_R FILLER_0_41_781 ();
 FILLER_ASAP7_75t_R FILLER_0_41_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_797 ();
 FILLER_ASAP7_75t_R FILLER_0_41_808 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_818 ();
 FILLER_ASAP7_75t_R FILLER_0_41_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_826 ();
 DECAPx1_ASAP7_75t_R FILLER_0_41_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_841 ();
 FILLER_ASAP7_75t_R FILLER_0_41_845 ();
 FILLER_ASAP7_75t_R FILLER_0_41_857 ();
 DECAPx1_ASAP7_75t_R FILLER_0_41_879 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_889 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_907 ();
 FILLER_ASAP7_75t_R FILLER_0_41_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_916 ();
 FILLER_ASAP7_75t_R FILLER_0_41_923 ();
 FILLER_ASAP7_75t_R FILLER_0_41_927 ();
 FILLER_ASAP7_75t_R FILLER_0_41_934 ();
 FILLER_ASAP7_75t_R FILLER_0_41_946 ();
 FILLER_ASAP7_75t_R FILLER_0_41_954 ();
 FILLER_ASAP7_75t_R FILLER_0_41_962 ();
 DECAPx6_ASAP7_75t_R FILLER_0_41_974 ();
 DECAPx1_ASAP7_75t_R FILLER_0_41_988 ();
 FILLER_ASAP7_75t_R FILLER_0_41_1000 ();
 DECAPx1_ASAP7_75t_R FILLER_0_41_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_1017 ();
 FILLER_ASAP7_75t_R FILLER_0_41_1024 ();
 DECAPx1_ASAP7_75t_R FILLER_0_41_1029 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_1044 ();
 DECAPx4_ASAP7_75t_R FILLER_0_41_1053 ();
 FILLER_ASAP7_75t_R FILLER_0_41_1063 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_1071 ();
 DECAPx6_ASAP7_75t_R FILLER_0_41_1081 ();
 FILLER_ASAP7_75t_R FILLER_0_41_1101 ();
 DECAPx4_ASAP7_75t_R FILLER_0_41_1114 ();
 DECAPx1_ASAP7_75t_R FILLER_0_41_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_1134 ();
 DECAPx4_ASAP7_75t_R FILLER_0_41_1141 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_1157 ();
 FILLER_ASAP7_75t_R FILLER_0_41_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_1165 ();
 FILLER_ASAP7_75t_R FILLER_0_41_1172 ();
 FILLER_ASAP7_75t_R FILLER_0_41_1180 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_1188 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_1200 ();
 FILLER_ASAP7_75t_R FILLER_0_41_1206 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_1216 ();
 FILLER_ASAP7_75t_R FILLER_0_41_1222 ();
 FILLER_ASAP7_75t_R FILLER_0_41_1232 ();
 DECAPx1_ASAP7_75t_R FILLER_0_41_1240 ();
 DECAPx6_ASAP7_75t_R FILLER_0_41_1250 ();
 DECAPx1_ASAP7_75t_R FILLER_0_41_1264 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_1268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_41_1275 ();
 FILLER_ASAP7_75t_R FILLER_0_41_1289 ();
 FILLER_ASAP7_75t_R FILLER_0_41_1301 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_1313 ();
 DECAPx6_ASAP7_75t_R FILLER_0_41_1324 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_1348 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_1354 ();
 DECAPx6_ASAP7_75t_R FILLER_0_41_1361 ();
 DECAPx1_ASAP7_75t_R FILLER_0_41_1378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_42_24 ();
 FILLER_ASAP7_75t_R FILLER_0_42_38 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_68 ();
 DECAPx1_ASAP7_75t_R FILLER_0_42_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_94 ();
 FILLER_ASAP7_75t_R FILLER_0_42_107 ();
 DECAPx6_ASAP7_75t_R FILLER_0_42_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_130 ();
 FILLER_ASAP7_75t_R FILLER_0_42_137 ();
 DECAPx2_ASAP7_75t_R FILLER_0_42_145 ();
 DECAPx1_ASAP7_75t_R FILLER_0_42_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_161 ();
 FILLER_ASAP7_75t_R FILLER_0_42_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_169 ();
 FILLER_ASAP7_75t_R FILLER_0_42_180 ();
 FILLER_ASAP7_75t_R FILLER_0_42_188 ();
 FILLER_ASAP7_75t_R FILLER_0_42_196 ();
 FILLER_ASAP7_75t_R FILLER_0_42_206 ();
 FILLER_ASAP7_75t_R FILLER_0_42_213 ();
 FILLER_ASAP7_75t_R FILLER_0_42_220 ();
 FILLER_ASAP7_75t_R FILLER_0_42_229 ();
 DECAPx6_ASAP7_75t_R FILLER_0_42_237 ();
 FILLER_ASAP7_75t_R FILLER_0_42_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_253 ();
 FILLER_ASAP7_75t_R FILLER_0_42_274 ();
 FILLER_ASAP7_75t_R FILLER_0_42_282 ();
 DECAPx2_ASAP7_75t_R FILLER_0_42_294 ();
 FILLER_ASAP7_75t_R FILLER_0_42_310 ();
 FILLER_ASAP7_75t_R FILLER_0_42_322 ();
 FILLER_ASAP7_75t_R FILLER_0_42_334 ();
 FILLER_ASAP7_75t_R FILLER_0_42_346 ();
 DECAPx2_ASAP7_75t_R FILLER_0_42_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_364 ();
 FILLER_ASAP7_75t_R FILLER_0_42_375 ();
 DECAPx2_ASAP7_75t_R FILLER_0_42_395 ();
 FILLER_ASAP7_75t_R FILLER_0_42_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_413 ();
 FILLER_ASAP7_75t_R FILLER_0_42_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_426 ();
 FILLER_ASAP7_75t_R FILLER_0_42_433 ();
 FILLER_ASAP7_75t_R FILLER_0_42_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_42_454 ();
 FILLER_ASAP7_75t_R FILLER_0_42_460 ();
 FILLER_ASAP7_75t_R FILLER_0_42_464 ();
 FILLER_ASAP7_75t_R FILLER_0_42_472 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_480 ();
 DECAPx4_ASAP7_75t_R FILLER_0_42_502 ();
 DECAPx1_ASAP7_75t_R FILLER_0_42_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_536 ();
 FILLER_ASAP7_75t_R FILLER_0_42_543 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_551 ();
 DECAPx6_ASAP7_75t_R FILLER_0_42_573 ();
 FILLER_ASAP7_75t_R FILLER_0_42_587 ();
 DECAPx4_ASAP7_75t_R FILLER_0_42_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_602 ();
 DECAPx2_ASAP7_75t_R FILLER_0_42_609 ();
 DECAPx1_ASAP7_75t_R FILLER_0_42_621 ();
 DECAPx2_ASAP7_75t_R FILLER_0_42_629 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_640 ();
 FILLER_ASAP7_75t_R FILLER_0_42_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_664 ();
 FILLER_ASAP7_75t_R FILLER_0_42_675 ();
 DECAPx4_ASAP7_75t_R FILLER_0_42_682 ();
 FILLER_ASAP7_75t_R FILLER_0_42_692 ();
 FILLER_ASAP7_75t_R FILLER_0_42_702 ();
 DECAPx2_ASAP7_75t_R FILLER_0_42_707 ();
 FILLER_ASAP7_75t_R FILLER_0_42_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_715 ();
 DECAPx2_ASAP7_75t_R FILLER_0_42_721 ();
 FILLER_ASAP7_75t_R FILLER_0_42_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_729 ();
 FILLER_ASAP7_75t_R FILLER_0_42_736 ();
 FILLER_ASAP7_75t_R FILLER_0_42_744 ();
 FILLER_ASAP7_75t_R FILLER_0_42_754 ();
 DECAPx4_ASAP7_75t_R FILLER_0_42_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_781 ();
 DECAPx2_ASAP7_75t_R FILLER_0_42_803 ();
 FILLER_ASAP7_75t_R FILLER_0_42_815 ();
 FILLER_ASAP7_75t_R FILLER_0_42_823 ();
 FILLER_ASAP7_75t_R FILLER_0_42_833 ();
 FILLER_ASAP7_75t_R FILLER_0_42_845 ();
 DECAPx2_ASAP7_75t_R FILLER_0_42_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_861 ();
 DECAPx6_ASAP7_75t_R FILLER_0_42_873 ();
 FILLER_ASAP7_75t_R FILLER_0_42_893 ();
 FILLER_ASAP7_75t_R FILLER_0_42_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_903 ();
 DECAPx4_ASAP7_75t_R FILLER_0_42_911 ();
 FILLER_ASAP7_75t_R FILLER_0_42_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_923 ();
 FILLER_ASAP7_75t_R FILLER_0_42_930 ();
 DECAPx1_ASAP7_75t_R FILLER_0_42_938 ();
 DECAPx2_ASAP7_75t_R FILLER_0_42_953 ();
 DECAPx6_ASAP7_75t_R FILLER_0_42_965 ();
 FILLER_ASAP7_75t_R FILLER_0_42_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_981 ();
 FILLER_ASAP7_75t_R FILLER_0_42_988 ();
 DECAPx1_ASAP7_75t_R FILLER_0_42_996 ();
 DECAPx6_ASAP7_75t_R FILLER_0_42_1012 ();
 FILLER_ASAP7_75t_R FILLER_0_42_1026 ();
 DECAPx1_ASAP7_75t_R FILLER_0_42_1039 ();
 FILLER_ASAP7_75t_R FILLER_0_42_1054 ();
 FILLER_ASAP7_75t_R FILLER_0_42_1061 ();
 FILLER_ASAP7_75t_R FILLER_0_42_1069 ();
 DECAPx2_ASAP7_75t_R FILLER_0_42_1077 ();
 FILLER_ASAP7_75t_R FILLER_0_42_1083 ();
 DECAPx6_ASAP7_75t_R FILLER_0_42_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_1112 ();
 DECAPx2_ASAP7_75t_R FILLER_0_42_1144 ();
 FILLER_ASAP7_75t_R FILLER_0_42_1164 ();
 FILLER_ASAP7_75t_R FILLER_0_42_1176 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_1178 ();
 DECAPx4_ASAP7_75t_R FILLER_0_42_1192 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_1202 ();
 FILLER_ASAP7_75t_R FILLER_0_42_1213 ();
 FILLER_ASAP7_75t_R FILLER_0_42_1225 ();
 DECAPx2_ASAP7_75t_R FILLER_0_42_1235 ();
 FILLER_ASAP7_75t_R FILLER_0_42_1241 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_1243 ();
 DECAPx2_ASAP7_75t_R FILLER_0_42_1252 ();
 FILLER_ASAP7_75t_R FILLER_0_42_1258 ();
 FILLER_ASAP7_75t_R FILLER_0_42_1267 ();
 DECAPx1_ASAP7_75t_R FILLER_0_42_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_0_42_1289 ();
 FILLER_ASAP7_75t_R FILLER_0_42_1303 ();
 FILLER_ASAP7_75t_R FILLER_0_42_1310 ();
 DECAPx2_ASAP7_75t_R FILLER_0_42_1318 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_1324 ();
 DECAPx2_ASAP7_75t_R FILLER_0_42_1331 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_1337 ();
 FILLER_ASAP7_75t_R FILLER_0_42_1344 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_1346 ();
 FILLER_ASAP7_75t_R FILLER_0_42_1353 ();
 DECAPx1_ASAP7_75t_R FILLER_0_42_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_1367 ();
 FILLER_ASAP7_75t_R FILLER_0_42_1371 ();
 FILLER_ASAP7_75t_R FILLER_0_42_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_43_24 ();
 FILLER_ASAP7_75t_R FILLER_0_43_40 ();
 DECAPx1_ASAP7_75t_R FILLER_0_43_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_56 ();
 DECAPx1_ASAP7_75t_R FILLER_0_43_63 ();
 FILLER_ASAP7_75t_R FILLER_0_43_73 ();
 FILLER_ASAP7_75t_R FILLER_0_43_82 ();
 DECAPx2_ASAP7_75t_R FILLER_0_43_91 ();
 FILLER_ASAP7_75t_R FILLER_0_43_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_99 ();
 FILLER_ASAP7_75t_R FILLER_0_43_106 ();
 DECAPx2_ASAP7_75t_R FILLER_0_43_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_119 ();
 DECAPx4_ASAP7_75t_R FILLER_0_43_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_136 ();
 FILLER_ASAP7_75t_R FILLER_0_43_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_145 ();
 FILLER_ASAP7_75t_R FILLER_0_43_160 ();
 FILLER_ASAP7_75t_R FILLER_0_43_172 ();
 DECAPx4_ASAP7_75t_R FILLER_0_43_179 ();
 FILLER_ASAP7_75t_R FILLER_0_43_189 ();
 FILLER_ASAP7_75t_R FILLER_0_43_196 ();
 FILLER_ASAP7_75t_R FILLER_0_43_203 ();
 DECAPx6_ASAP7_75t_R FILLER_0_43_215 ();
 DECAPx2_ASAP7_75t_R FILLER_0_43_229 ();
 DECAPx6_ASAP7_75t_R FILLER_0_43_245 ();
 FILLER_ASAP7_75t_R FILLER_0_43_259 ();
 FILLER_ASAP7_75t_R FILLER_0_43_266 ();
 FILLER_ASAP7_75t_R FILLER_0_43_278 ();
 FILLER_ASAP7_75t_R FILLER_0_43_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_288 ();
 FILLER_ASAP7_75t_R FILLER_0_43_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_299 ();
 FILLER_ASAP7_75t_R FILLER_0_43_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_314 ();
 FILLER_ASAP7_75t_R FILLER_0_43_321 ();
 FILLER_ASAP7_75t_R FILLER_0_43_351 ();
 DECAPx2_ASAP7_75t_R FILLER_0_43_371 ();
 DECAPx1_ASAP7_75t_R FILLER_0_43_387 ();
 FILLER_ASAP7_75t_R FILLER_0_43_401 ();
 FILLER_ASAP7_75t_R FILLER_0_43_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_411 ();
 FILLER_ASAP7_75t_R FILLER_0_43_420 ();
 FILLER_ASAP7_75t_R FILLER_0_43_428 ();
 DECAPx6_ASAP7_75t_R FILLER_0_43_435 ();
 DECAPx1_ASAP7_75t_R FILLER_0_43_449 ();
 DECAPx6_ASAP7_75t_R FILLER_0_43_460 ();
 FILLER_ASAP7_75t_R FILLER_0_43_480 ();
 FILLER_ASAP7_75t_R FILLER_0_43_496 ();
 DECAPx2_ASAP7_75t_R FILLER_0_43_504 ();
 FILLER_ASAP7_75t_R FILLER_0_43_510 ();
 FILLER_ASAP7_75t_R FILLER_0_43_519 ();
 FILLER_ASAP7_75t_R FILLER_0_43_528 ();
 FILLER_ASAP7_75t_R FILLER_0_43_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_538 ();
 FILLER_ASAP7_75t_R FILLER_0_43_545 ();
 DECAPx2_ASAP7_75t_R FILLER_0_43_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_559 ();
 DECAPx6_ASAP7_75t_R FILLER_0_43_566 ();
 DECAPx1_ASAP7_75t_R FILLER_0_43_580 ();
 DECAPx2_ASAP7_75t_R FILLER_0_43_604 ();
 FILLER_ASAP7_75t_R FILLER_0_43_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_612 ();
 DECAPx1_ASAP7_75t_R FILLER_0_43_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_625 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_636 ();
 DECAPx1_ASAP7_75t_R FILLER_0_43_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_662 ();
 DECAPx2_ASAP7_75t_R FILLER_0_43_669 ();
 FILLER_ASAP7_75t_R FILLER_0_43_675 ();
 FILLER_ASAP7_75t_R FILLER_0_43_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_689 ();
 DECAPx6_ASAP7_75t_R FILLER_0_43_696 ();
 DECAPx1_ASAP7_75t_R FILLER_0_43_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_714 ();
 DECAPx4_ASAP7_75t_R FILLER_0_43_721 ();
 FILLER_ASAP7_75t_R FILLER_0_43_739 ();
 DECAPx1_ASAP7_75t_R FILLER_0_43_749 ();
 DECAPx4_ASAP7_75t_R FILLER_0_43_761 ();
 FILLER_ASAP7_75t_R FILLER_0_43_771 ();
 DECAPx1_ASAP7_75t_R FILLER_0_43_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_783 ();
 FILLER_ASAP7_75t_R FILLER_0_43_792 ();
 DECAPx2_ASAP7_75t_R FILLER_0_43_797 ();
 DECAPx4_ASAP7_75t_R FILLER_0_43_815 ();
 FILLER_ASAP7_75t_R FILLER_0_43_825 ();
 FILLER_ASAP7_75t_R FILLER_0_43_830 ();
 DECAPx1_ASAP7_75t_R FILLER_0_43_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_844 ();
 FILLER_ASAP7_75t_R FILLER_0_43_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_855 ();
 DECAPx1_ASAP7_75t_R FILLER_0_43_864 ();
 DECAPx6_ASAP7_75t_R FILLER_0_43_874 ();
 FILLER_ASAP7_75t_R FILLER_0_43_888 ();
 DECAPx1_ASAP7_75t_R FILLER_0_43_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_900 ();
 FILLER_ASAP7_75t_R FILLER_0_43_907 ();
 DECAPx4_ASAP7_75t_R FILLER_0_43_915 ();
 FILLER_ASAP7_75t_R FILLER_0_43_927 ();
 FILLER_ASAP7_75t_R FILLER_0_43_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_941 ();
 FILLER_ASAP7_75t_R FILLER_0_43_953 ();
 FILLER_ASAP7_75t_R FILLER_0_43_960 ();
 FILLER_ASAP7_75t_R FILLER_0_43_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_975 ();
 DECAPx1_ASAP7_75t_R FILLER_0_43_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_983 ();
 DECAPx4_ASAP7_75t_R FILLER_0_43_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_1002 ();
 FILLER_ASAP7_75t_R FILLER_0_43_1010 ();
 FILLER_ASAP7_75t_R FILLER_0_43_1018 ();
 FILLER_ASAP7_75t_R FILLER_0_43_1026 ();
 DECAPx2_ASAP7_75t_R FILLER_0_43_1038 ();
 FILLER_ASAP7_75t_R FILLER_0_43_1054 ();
 FILLER_ASAP7_75t_R FILLER_0_43_1066 ();
 DECAPx4_ASAP7_75t_R FILLER_0_43_1074 ();
 FILLER_ASAP7_75t_R FILLER_0_43_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_1086 ();
 DECAPx1_ASAP7_75t_R FILLER_0_43_1098 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_1108 ();
 DECAPx4_ASAP7_75t_R FILLER_0_43_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_1140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_1151 ();
 DECAPx6_ASAP7_75t_R FILLER_0_43_1173 ();
 DECAPx2_ASAP7_75t_R FILLER_0_43_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_1193 ();
 FILLER_ASAP7_75t_R FILLER_0_43_1200 ();
 FILLER_ASAP7_75t_R FILLER_0_43_1212 ();
 DECAPx1_ASAP7_75t_R FILLER_0_43_1232 ();
 DECAPx1_ASAP7_75t_R FILLER_0_43_1246 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_1250 ();
 FILLER_ASAP7_75t_R FILLER_0_43_1258 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_1260 ();
 FILLER_ASAP7_75t_R FILLER_0_43_1271 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_1273 ();
 FILLER_ASAP7_75t_R FILLER_0_43_1284 ();
 FILLER_ASAP7_75t_R FILLER_0_43_1296 ();
 FILLER_ASAP7_75t_R FILLER_0_43_1304 ();
 FILLER_ASAP7_75t_R FILLER_0_43_1312 ();
 FILLER_ASAP7_75t_R FILLER_0_43_1320 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_1322 ();
 DECAPx6_ASAP7_75t_R FILLER_0_43_1329 ();
 DECAPx2_ASAP7_75t_R FILLER_0_43_1343 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_1349 ();
 DECAPx6_ASAP7_75t_R FILLER_0_43_1356 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_1370 ();
 DECAPx1_ASAP7_75t_R FILLER_0_43_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_2 ();
 FILLER_ASAP7_75t_R FILLER_0_44_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_26 ();
 FILLER_ASAP7_75t_R FILLER_0_44_30 ();
 FILLER_ASAP7_75t_R FILLER_0_44_38 ();
 DECAPx2_ASAP7_75t_R FILLER_0_44_46 ();
 FILLER_ASAP7_75t_R FILLER_0_44_58 ();
 FILLER_ASAP7_75t_R FILLER_0_44_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_68 ();
 DECAPx2_ASAP7_75t_R FILLER_0_44_75 ();
 FILLER_ASAP7_75t_R FILLER_0_44_87 ();
 DECAPx2_ASAP7_75t_R FILLER_0_44_95 ();
 DECAPx2_ASAP7_75t_R FILLER_0_44_107 ();
 FILLER_ASAP7_75t_R FILLER_0_44_123 ();
 DECAPx1_ASAP7_75t_R FILLER_0_44_131 ();
 FILLER_ASAP7_75t_R FILLER_0_44_145 ();
 FILLER_ASAP7_75t_R FILLER_0_44_152 ();
 DECAPx1_ASAP7_75t_R FILLER_0_44_159 ();
 DECAPx1_ASAP7_75t_R FILLER_0_44_173 ();
 DECAPx6_ASAP7_75t_R FILLER_0_44_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_201 ();
 FILLER_ASAP7_75t_R FILLER_0_44_207 ();
 FILLER_ASAP7_75t_R FILLER_0_44_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_217 ();
 FILLER_ASAP7_75t_R FILLER_0_44_224 ();
 FILLER_ASAP7_75t_R FILLER_0_44_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_248 ();
 DECAPx4_ASAP7_75t_R FILLER_0_44_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_265 ();
 FILLER_ASAP7_75t_R FILLER_0_44_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_288 ();
 FILLER_ASAP7_75t_R FILLER_0_44_295 ();
 DECAPx1_ASAP7_75t_R FILLER_0_44_303 ();
 DECAPx1_ASAP7_75t_R FILLER_0_44_329 ();
 FILLER_ASAP7_75t_R FILLER_0_44_351 ();
 FILLER_ASAP7_75t_R FILLER_0_44_371 ();
 FILLER_ASAP7_75t_R FILLER_0_44_387 ();
 FILLER_ASAP7_75t_R FILLER_0_44_393 ();
 DECAPx1_ASAP7_75t_R FILLER_0_44_401 ();
 FILLER_ASAP7_75t_R FILLER_0_44_416 ();
 FILLER_ASAP7_75t_R FILLER_0_44_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_425 ();
 FILLER_ASAP7_75t_R FILLER_0_44_432 ();
 FILLER_ASAP7_75t_R FILLER_0_44_439 ();
 FILLER_ASAP7_75t_R FILLER_0_44_444 ();
 FILLER_ASAP7_75t_R FILLER_0_44_452 ();
 FILLER_ASAP7_75t_R FILLER_0_44_460 ();
 FILLER_ASAP7_75t_R FILLER_0_44_464 ();
 FILLER_ASAP7_75t_R FILLER_0_44_477 ();
 DECAPx2_ASAP7_75t_R FILLER_0_44_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_491 ();
 FILLER_ASAP7_75t_R FILLER_0_44_498 ();
 FILLER_ASAP7_75t_R FILLER_0_44_506 ();
 DECAPx1_ASAP7_75t_R FILLER_0_44_511 ();
 DECAPx2_ASAP7_75t_R FILLER_0_44_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_527 ();
 DECAPx4_ASAP7_75t_R FILLER_0_44_534 ();
 FILLER_ASAP7_75t_R FILLER_0_44_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_546 ();
 FILLER_ASAP7_75t_R FILLER_0_44_554 ();
 DECAPx6_ASAP7_75t_R FILLER_0_44_567 ();
 DECAPx2_ASAP7_75t_R FILLER_0_44_581 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_595 ();
 DECAPx2_ASAP7_75t_R FILLER_0_44_617 ();
 FILLER_ASAP7_75t_R FILLER_0_44_623 ();
 FILLER_ASAP7_75t_R FILLER_0_44_633 ();
 FILLER_ASAP7_75t_R FILLER_0_44_639 ();
 DECAPx2_ASAP7_75t_R FILLER_0_44_645 ();
 FILLER_ASAP7_75t_R FILLER_0_44_651 ();
 FILLER_ASAP7_75t_R FILLER_0_44_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_663 ();
 FILLER_ASAP7_75t_R FILLER_0_44_672 ();
 DECAPx4_ASAP7_75t_R FILLER_0_44_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_690 ();
 DECAPx2_ASAP7_75t_R FILLER_0_44_697 ();
 FILLER_ASAP7_75t_R FILLER_0_44_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_705 ();
 DECAPx4_ASAP7_75t_R FILLER_0_44_718 ();
 FILLER_ASAP7_75t_R FILLER_0_44_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_44_740 ();
 FILLER_ASAP7_75t_R FILLER_0_44_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_748 ();
 FILLER_ASAP7_75t_R FILLER_0_44_757 ();
 DECAPx4_ASAP7_75t_R FILLER_0_44_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_775 ();
 FILLER_ASAP7_75t_R FILLER_0_44_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_786 ();
 FILLER_ASAP7_75t_R FILLER_0_44_793 ();
 FILLER_ASAP7_75t_R FILLER_0_44_803 ();
 DECAPx6_ASAP7_75t_R FILLER_0_44_808 ();
 FILLER_ASAP7_75t_R FILLER_0_44_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_824 ();
 DECAPx1_ASAP7_75t_R FILLER_0_44_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_852 ();
 FILLER_ASAP7_75t_R FILLER_0_44_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_876 ();
 DECAPx6_ASAP7_75t_R FILLER_0_44_887 ();
 FILLER_ASAP7_75t_R FILLER_0_44_901 ();
 DECAPx6_ASAP7_75t_R FILLER_0_44_909 ();
 FILLER_ASAP7_75t_R FILLER_0_44_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_925 ();
 DECAPx1_ASAP7_75t_R FILLER_0_44_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_933 ();
 FILLER_ASAP7_75t_R FILLER_0_44_944 ();
 FILLER_ASAP7_75t_R FILLER_0_44_951 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_963 ();
 DECAPx4_ASAP7_75t_R FILLER_0_44_985 ();
 FILLER_ASAP7_75t_R FILLER_0_44_995 ();
 FILLER_ASAP7_75t_R FILLER_0_44_1002 ();
 DECAPx6_ASAP7_75t_R FILLER_0_44_1015 ();
 FILLER_ASAP7_75t_R FILLER_0_44_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_1031 ();
 FILLER_ASAP7_75t_R FILLER_0_44_1038 ();
 FILLER_ASAP7_75t_R FILLER_0_44_1050 ();
 FILLER_ASAP7_75t_R FILLER_0_44_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_1059 ();
 FILLER_ASAP7_75t_R FILLER_0_44_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_1069 ();
 FILLER_ASAP7_75t_R FILLER_0_44_1086 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_1094 ();
 DECAPx6_ASAP7_75t_R FILLER_0_44_1116 ();
 FILLER_ASAP7_75t_R FILLER_0_44_1133 ();
 DECAPx1_ASAP7_75t_R FILLER_0_44_1155 ();
 FILLER_ASAP7_75t_R FILLER_0_44_1165 ();
 FILLER_ASAP7_75t_R FILLER_0_44_1173 ();
 FILLER_ASAP7_75t_R FILLER_0_44_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_1180 ();
 DECAPx1_ASAP7_75t_R FILLER_0_44_1191 ();
 DECAPx2_ASAP7_75t_R FILLER_0_44_1201 ();
 DECAPx2_ASAP7_75t_R FILLER_0_44_1217 ();
 DECAPx1_ASAP7_75t_R FILLER_0_44_1233 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_1237 ();
 FILLER_ASAP7_75t_R FILLER_0_44_1244 ();
 FILLER_ASAP7_75t_R FILLER_0_44_1254 ();
 FILLER_ASAP7_75t_R FILLER_0_44_1261 ();
 DECAPx4_ASAP7_75t_R FILLER_0_44_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_1279 ();
 FILLER_ASAP7_75t_R FILLER_0_44_1290 ();
 FILLER_ASAP7_75t_R FILLER_0_44_1302 ();
 DECAPx1_ASAP7_75t_R FILLER_0_44_1310 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_1314 ();
 DECAPx1_ASAP7_75t_R FILLER_0_44_1320 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_1324 ();
 FILLER_ASAP7_75t_R FILLER_0_44_1333 ();
 FILLER_ASAP7_75t_R FILLER_0_44_1341 ();
 FILLER_ASAP7_75t_R FILLER_0_44_1349 ();
 DECAPx4_ASAP7_75t_R FILLER_0_44_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_44_1367 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_1369 ();
 FILLER_ASAP7_75t_R FILLER_0_44_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_45_24 ();
 DECAPx2_ASAP7_75t_R FILLER_0_45_38 ();
 DECAPx4_ASAP7_75t_R FILLER_0_45_50 ();
 DECAPx6_ASAP7_75t_R FILLER_0_45_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_79 ();
 FILLER_ASAP7_75t_R FILLER_0_45_86 ();
 FILLER_ASAP7_75t_R FILLER_0_45_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_95 ();
 DECAPx6_ASAP7_75t_R FILLER_0_45_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_116 ();
 FILLER_ASAP7_75t_R FILLER_0_45_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_125 ();
 DECAPx2_ASAP7_75t_R FILLER_0_45_131 ();
 FILLER_ASAP7_75t_R FILLER_0_45_147 ();
 FILLER_ASAP7_75t_R FILLER_0_45_154 ();
 FILLER_ASAP7_75t_R FILLER_0_45_162 ();
 DECAPx4_ASAP7_75t_R FILLER_0_45_174 ();
 FILLER_ASAP7_75t_R FILLER_0_45_184 ();
 FILLER_ASAP7_75t_R FILLER_0_45_192 ();
 FILLER_ASAP7_75t_R FILLER_0_45_200 ();
 FILLER_ASAP7_75t_R FILLER_0_45_213 ();
 FILLER_ASAP7_75t_R FILLER_0_45_225 ();
 DECAPx1_ASAP7_75t_R FILLER_0_45_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_251 ();
 DECAPx1_ASAP7_75t_R FILLER_0_45_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_262 ();
 FILLER_ASAP7_75t_R FILLER_0_45_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_271 ();
 DECAPx4_ASAP7_75t_R FILLER_0_45_276 ();
 FILLER_ASAP7_75t_R FILLER_0_45_286 ();
 FILLER_ASAP7_75t_R FILLER_0_45_296 ();
 FILLER_ASAP7_75t_R FILLER_0_45_301 ();
 DECAPx1_ASAP7_75t_R FILLER_0_45_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_313 ();
 FILLER_ASAP7_75t_R FILLER_0_45_319 ();
 FILLER_ASAP7_75t_R FILLER_0_45_326 ();
 FILLER_ASAP7_75t_R FILLER_0_45_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_340 ();
 FILLER_ASAP7_75t_R FILLER_0_45_351 ();
 FILLER_ASAP7_75t_R FILLER_0_45_363 ();
 FILLER_ASAP7_75t_R FILLER_0_45_377 ();
 DECAPx1_ASAP7_75t_R FILLER_0_45_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_393 ();
 FILLER_ASAP7_75t_R FILLER_0_45_404 ();
 DECAPx1_ASAP7_75t_R FILLER_0_45_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_418 ();
 DECAPx2_ASAP7_75t_R FILLER_0_45_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_432 ();
 FILLER_ASAP7_75t_R FILLER_0_45_439 ();
 DECAPx2_ASAP7_75t_R FILLER_0_45_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_450 ();
 DECAPx6_ASAP7_75t_R FILLER_0_45_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_470 ();
 FILLER_ASAP7_75t_R FILLER_0_45_477 ();
 FILLER_ASAP7_75t_R FILLER_0_45_485 ();
 DECAPx1_ASAP7_75t_R FILLER_0_45_493 ();
 DECAPx1_ASAP7_75t_R FILLER_0_45_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_507 ();
 FILLER_ASAP7_75t_R FILLER_0_45_514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_45_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_526 ();
 FILLER_ASAP7_75t_R FILLER_0_45_533 ();
 DECAPx2_ASAP7_75t_R FILLER_0_45_540 ();
 DECAPx6_ASAP7_75t_R FILLER_0_45_552 ();
 FILLER_ASAP7_75t_R FILLER_0_45_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_568 ();
 FILLER_ASAP7_75t_R FILLER_0_45_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_583 ();
 DECAPx1_ASAP7_75t_R FILLER_0_45_592 ();
 DECAPx1_ASAP7_75t_R FILLER_0_45_607 ();
 DECAPx1_ASAP7_75t_R FILLER_0_45_619 ();
 FILLER_ASAP7_75t_R FILLER_0_45_631 ();
 FILLER_ASAP7_75t_R FILLER_0_45_641 ();
 FILLER_ASAP7_75t_R FILLER_0_45_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_653 ();
 FILLER_ASAP7_75t_R FILLER_0_45_662 ();
 FILLER_ASAP7_75t_R FILLER_0_45_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_669 ();
 FILLER_ASAP7_75t_R FILLER_0_45_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_680 ();
 FILLER_ASAP7_75t_R FILLER_0_45_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_686 ();
 FILLER_ASAP7_75t_R FILLER_0_45_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_695 ();
 DECAPx1_ASAP7_75t_R FILLER_0_45_702 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_718 ();
 FILLER_ASAP7_75t_R FILLER_0_45_740 ();
 DECAPx1_ASAP7_75t_R FILLER_0_45_748 ();
 DECAPx2_ASAP7_75t_R FILLER_0_45_758 ();
 FILLER_ASAP7_75t_R FILLER_0_45_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_766 ();
 FILLER_ASAP7_75t_R FILLER_0_45_778 ();
 DECAPx1_ASAP7_75t_R FILLER_0_45_786 ();
 FILLER_ASAP7_75t_R FILLER_0_45_796 ();
 DECAPx4_ASAP7_75t_R FILLER_0_45_803 ();
 FILLER_ASAP7_75t_R FILLER_0_45_813 ();
 DECAPx4_ASAP7_75t_R FILLER_0_45_818 ();
 FILLER_ASAP7_75t_R FILLER_0_45_828 ();
 FILLER_ASAP7_75t_R FILLER_0_45_835 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_842 ();
 DECAPx6_ASAP7_75t_R FILLER_0_45_864 ();
 DECAPx2_ASAP7_75t_R FILLER_0_45_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_891 ();
 DECAPx4_ASAP7_75t_R FILLER_0_45_913 ();
 FILLER_ASAP7_75t_R FILLER_0_45_923 ();
 DECAPx2_ASAP7_75t_R FILLER_0_45_927 ();
 FILLER_ASAP7_75t_R FILLER_0_45_933 ();
 DECAPx2_ASAP7_75t_R FILLER_0_45_941 ();
 FILLER_ASAP7_75t_R FILLER_0_45_957 ();
 DECAPx6_ASAP7_75t_R FILLER_0_45_969 ();
 DECAPx2_ASAP7_75t_R FILLER_0_45_983 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_999 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_1021 ();
 DECAPx6_ASAP7_75t_R FILLER_0_45_1028 ();
 DECAPx1_ASAP7_75t_R FILLER_0_45_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_1046 ();
 FILLER_ASAP7_75t_R FILLER_0_45_1053 ();
 FILLER_ASAP7_75t_R FILLER_0_45_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_1063 ();
 DECAPx2_ASAP7_75t_R FILLER_0_45_1069 ();
 FILLER_ASAP7_75t_R FILLER_0_45_1081 ();
 FILLER_ASAP7_75t_R FILLER_0_45_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_0_45_1097 ();
 DECAPx4_ASAP7_75t_R FILLER_0_45_1111 ();
 FILLER_ASAP7_75t_R FILLER_0_45_1121 ();
 FILLER_ASAP7_75t_R FILLER_0_45_1133 ();
 FILLER_ASAP7_75t_R FILLER_0_45_1141 ();
 FILLER_ASAP7_75t_R FILLER_0_45_1149 ();
 DECAPx2_ASAP7_75t_R FILLER_0_45_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_1162 ();
 FILLER_ASAP7_75t_R FILLER_0_45_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_1171 ();
 DECAPx1_ASAP7_75t_R FILLER_0_45_1179 ();
 FILLER_ASAP7_75t_R FILLER_0_45_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_1195 ();
 DECAPx1_ASAP7_75t_R FILLER_0_45_1203 ();
 FILLER_ASAP7_75t_R FILLER_0_45_1217 ();
 FILLER_ASAP7_75t_R FILLER_0_45_1227 ();
 DECAPx4_ASAP7_75t_R FILLER_0_45_1235 ();
 FILLER_ASAP7_75t_R FILLER_0_45_1251 ();
 FILLER_ASAP7_75t_R FILLER_0_45_1259 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_1261 ();
 DECAPx2_ASAP7_75t_R FILLER_0_45_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_1275 ();
 FILLER_ASAP7_75t_R FILLER_0_45_1281 ();
 FILLER_ASAP7_75t_R FILLER_0_45_1289 ();
 FILLER_ASAP7_75t_R FILLER_0_45_1301 ();
 DECAPx6_ASAP7_75t_R FILLER_0_45_1308 ();
 DECAPx2_ASAP7_75t_R FILLER_0_45_1322 ();
 FILLER_ASAP7_75t_R FILLER_0_45_1334 ();
 DECAPx1_ASAP7_75t_R FILLER_0_45_1342 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_1346 ();
 DECAPx4_ASAP7_75t_R FILLER_0_45_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_45_1367 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_1369 ();
 FILLER_ASAP7_75t_R FILLER_0_45_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_46_24 ();
 FILLER_ASAP7_75t_R FILLER_0_46_46 ();
 FILLER_ASAP7_75t_R FILLER_0_46_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_61 ();
 DECAPx4_ASAP7_75t_R FILLER_0_46_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_93 ();
 DECAPx6_ASAP7_75t_R FILLER_0_46_100 ();
 FILLER_ASAP7_75t_R FILLER_0_46_130 ();
 FILLER_ASAP7_75t_R FILLER_0_46_138 ();
 DECAPx1_ASAP7_75t_R FILLER_0_46_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_155 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_163 ();
 DECAPx2_ASAP7_75t_R FILLER_0_46_192 ();
 FILLER_ASAP7_75t_R FILLER_0_46_204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_234 ();
 DECAPx4_ASAP7_75t_R FILLER_0_46_241 ();
 FILLER_ASAP7_75t_R FILLER_0_46_257 ();
 FILLER_ASAP7_75t_R FILLER_0_46_265 ();
 DECAPx1_ASAP7_75t_R FILLER_0_46_279 ();
 DECAPx4_ASAP7_75t_R FILLER_0_46_289 ();
 FILLER_ASAP7_75t_R FILLER_0_46_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_301 ();
 DECAPx2_ASAP7_75t_R FILLER_0_46_322 ();
 FILLER_ASAP7_75t_R FILLER_0_46_338 ();
 FILLER_ASAP7_75t_R FILLER_0_46_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_352 ();
 FILLER_ASAP7_75t_R FILLER_0_46_356 ();
 FILLER_ASAP7_75t_R FILLER_0_46_369 ();
 DECAPx2_ASAP7_75t_R FILLER_0_46_377 ();
 FILLER_ASAP7_75t_R FILLER_0_46_383 ();
 DECAPx1_ASAP7_75t_R FILLER_0_46_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_399 ();
 FILLER_ASAP7_75t_R FILLER_0_46_406 ();
 DECAPx1_ASAP7_75t_R FILLER_0_46_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_422 ();
 FILLER_ASAP7_75t_R FILLER_0_46_429 ();
 FILLER_ASAP7_75t_R FILLER_0_46_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_439 ();
 DECAPx1_ASAP7_75t_R FILLER_0_46_446 ();
 DECAPx1_ASAP7_75t_R FILLER_0_46_458 ();
 DECAPx1_ASAP7_75t_R FILLER_0_46_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_468 ();
 FILLER_ASAP7_75t_R FILLER_0_46_475 ();
 DECAPx4_ASAP7_75t_R FILLER_0_46_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_494 ();
 FILLER_ASAP7_75t_R FILLER_0_46_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_501 ();
 FILLER_ASAP7_75t_R FILLER_0_46_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_516 ();
 DECAPx1_ASAP7_75t_R FILLER_0_46_524 ();
 FILLER_ASAP7_75t_R FILLER_0_46_534 ();
 DECAPx2_ASAP7_75t_R FILLER_0_46_542 ();
 FILLER_ASAP7_75t_R FILLER_0_46_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_550 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_557 ();
 FILLER_ASAP7_75t_R FILLER_0_46_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_581 ();
 FILLER_ASAP7_75t_R FILLER_0_46_602 ();
 FILLER_ASAP7_75t_R FILLER_0_46_612 ();
 FILLER_ASAP7_75t_R FILLER_0_46_622 ();
 DECAPx1_ASAP7_75t_R FILLER_0_46_627 ();
 FILLER_ASAP7_75t_R FILLER_0_46_641 ();
 DECAPx2_ASAP7_75t_R FILLER_0_46_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_657 ();
 FILLER_ASAP7_75t_R FILLER_0_46_661 ();
 FILLER_ASAP7_75t_R FILLER_0_46_671 ();
 FILLER_ASAP7_75t_R FILLER_0_46_681 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_691 ();
 FILLER_ASAP7_75t_R FILLER_0_46_713 ();
 FILLER_ASAP7_75t_R FILLER_0_46_723 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_756 ();
 DECAPx2_ASAP7_75t_R FILLER_0_46_778 ();
 FILLER_ASAP7_75t_R FILLER_0_46_784 ();
 FILLER_ASAP7_75t_R FILLER_0_46_794 ();
 DECAPx4_ASAP7_75t_R FILLER_0_46_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_809 ();
 FILLER_ASAP7_75t_R FILLER_0_46_813 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_823 ();
 FILLER_ASAP7_75t_R FILLER_0_46_845 ();
 FILLER_ASAP7_75t_R FILLER_0_46_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_869 ();
 DECAPx6_ASAP7_75t_R FILLER_0_46_874 ();
 FILLER_ASAP7_75t_R FILLER_0_46_894 ();
 DECAPx2_ASAP7_75t_R FILLER_0_46_902 ();
 FILLER_ASAP7_75t_R FILLER_0_46_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_910 ();
 FILLER_ASAP7_75t_R FILLER_0_46_917 ();
 FILLER_ASAP7_75t_R FILLER_0_46_925 ();
 DECAPx2_ASAP7_75t_R FILLER_0_46_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_939 ();
 DECAPx6_ASAP7_75t_R FILLER_0_46_960 ();
 DECAPx1_ASAP7_75t_R FILLER_0_46_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_978 ();
 DECAPx1_ASAP7_75t_R FILLER_0_46_999 ();
 FILLER_ASAP7_75t_R FILLER_0_46_1009 ();
 FILLER_ASAP7_75t_R FILLER_0_46_1017 ();
 FILLER_ASAP7_75t_R FILLER_0_46_1025 ();
 DECAPx4_ASAP7_75t_R FILLER_0_46_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_1048 ();
 FILLER_ASAP7_75t_R FILLER_0_46_1059 ();
 FILLER_ASAP7_75t_R FILLER_0_46_1067 ();
 FILLER_ASAP7_75t_R FILLER_0_46_1075 ();
 FILLER_ASAP7_75t_R FILLER_0_46_1083 ();
 FILLER_ASAP7_75t_R FILLER_0_46_1091 ();
 DECAPx4_ASAP7_75t_R FILLER_0_46_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_1109 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_1120 ();
 FILLER_ASAP7_75t_R FILLER_0_46_1142 ();
 FILLER_ASAP7_75t_R FILLER_0_46_1164 ();
 FILLER_ASAP7_75t_R FILLER_0_46_1186 ();
 DECAPx4_ASAP7_75t_R FILLER_0_46_1194 ();
 FILLER_ASAP7_75t_R FILLER_0_46_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_1206 ();
 FILLER_ASAP7_75t_R FILLER_0_46_1217 ();
 FILLER_ASAP7_75t_R FILLER_0_46_1225 ();
 DECAPx6_ASAP7_75t_R FILLER_0_46_1230 ();
 FILLER_ASAP7_75t_R FILLER_0_46_1250 ();
 DECAPx2_ASAP7_75t_R FILLER_0_46_1257 ();
 FILLER_ASAP7_75t_R FILLER_0_46_1263 ();
 FILLER_ASAP7_75t_R FILLER_0_46_1271 ();
 DECAPx1_ASAP7_75t_R FILLER_0_46_1279 ();
 FILLER_ASAP7_75t_R FILLER_0_46_1293 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_1295 ();
 DECAPx1_ASAP7_75t_R FILLER_0_46_1306 ();
 FILLER_ASAP7_75t_R FILLER_0_46_1320 ();
 DECAPx2_ASAP7_75t_R FILLER_0_46_1327 ();
 DECAPx6_ASAP7_75t_R FILLER_0_46_1339 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_1353 ();
 DECAPx6_ASAP7_75t_R FILLER_0_46_1362 ();
 DECAPx2_ASAP7_75t_R FILLER_0_46_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_47_24 ();
 DECAPx2_ASAP7_75t_R FILLER_0_47_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_44 ();
 FILLER_ASAP7_75t_R FILLER_0_47_51 ();
 DECAPx2_ASAP7_75t_R FILLER_0_47_59 ();
 FILLER_ASAP7_75t_R FILLER_0_47_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_67 ();
 FILLER_ASAP7_75t_R FILLER_0_47_74 ();
 DECAPx2_ASAP7_75t_R FILLER_0_47_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_90 ();
 FILLER_ASAP7_75t_R FILLER_0_47_103 ();
 FILLER_ASAP7_75t_R FILLER_0_47_111 ();
 DECAPx1_ASAP7_75t_R FILLER_0_47_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_128 ();
 FILLER_ASAP7_75t_R FILLER_0_47_135 ();
 FILLER_ASAP7_75t_R FILLER_0_47_143 ();
 DECAPx1_ASAP7_75t_R FILLER_0_47_150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_160 ();
 DECAPx2_ASAP7_75t_R FILLER_0_47_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_188 ();
 FILLER_ASAP7_75t_R FILLER_0_47_195 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_207 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_229 ();
 DECAPx4_ASAP7_75t_R FILLER_0_47_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_261 ();
 FILLER_ASAP7_75t_R FILLER_0_47_268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_276 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_320 ();
 FILLER_ASAP7_75t_R FILLER_0_47_324 ();
 FILLER_ASAP7_75t_R FILLER_0_47_331 ();
 DECAPx2_ASAP7_75t_R FILLER_0_47_339 ();
 FILLER_ASAP7_75t_R FILLER_0_47_351 ();
 DECAPx1_ASAP7_75t_R FILLER_0_47_363 ();
 FILLER_ASAP7_75t_R FILLER_0_47_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_379 ();
 FILLER_ASAP7_75t_R FILLER_0_47_392 ();
 DECAPx1_ASAP7_75t_R FILLER_0_47_404 ();
 DECAPx1_ASAP7_75t_R FILLER_0_47_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_418 ();
 DECAPx1_ASAP7_75t_R FILLER_0_47_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_429 ();
 FILLER_ASAP7_75t_R FILLER_0_47_436 ();
 DECAPx4_ASAP7_75t_R FILLER_0_47_444 ();
 FILLER_ASAP7_75t_R FILLER_0_47_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_456 ();
 FILLER_ASAP7_75t_R FILLER_0_47_463 ();
 DECAPx2_ASAP7_75t_R FILLER_0_47_470 ();
 FILLER_ASAP7_75t_R FILLER_0_47_476 ();
 FILLER_ASAP7_75t_R FILLER_0_47_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_488 ();
 FILLER_ASAP7_75t_R FILLER_0_47_497 ();
 DECAPx2_ASAP7_75t_R FILLER_0_47_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_513 ();
 DECAPx1_ASAP7_75t_R FILLER_0_47_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_530 ();
 DECAPx4_ASAP7_75t_R FILLER_0_47_537 ();
 FILLER_ASAP7_75t_R FILLER_0_47_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_549 ();
 FILLER_ASAP7_75t_R FILLER_0_47_556 ();
 DECAPx6_ASAP7_75t_R FILLER_0_47_568 ();
 FILLER_ASAP7_75t_R FILLER_0_47_586 ();
 FILLER_ASAP7_75t_R FILLER_0_47_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_593 ();
 FILLER_ASAP7_75t_R FILLER_0_47_600 ();
 FILLER_ASAP7_75t_R FILLER_0_47_610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_620 ();
 DECAPx4_ASAP7_75t_R FILLER_0_47_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_664 ();
 DECAPx2_ASAP7_75t_R FILLER_0_47_686 ();
 FILLER_ASAP7_75t_R FILLER_0_47_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_700 ();
 FILLER_ASAP7_75t_R FILLER_0_47_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_715 ();
 FILLER_ASAP7_75t_R FILLER_0_47_720 ();
 FILLER_ASAP7_75t_R FILLER_0_47_733 ();
 DECAPx4_ASAP7_75t_R FILLER_0_47_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_751 ();
 DECAPx1_ASAP7_75t_R FILLER_0_47_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_777 ();
 FILLER_ASAP7_75t_R FILLER_0_47_790 ();
 FILLER_ASAP7_75t_R FILLER_0_47_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_802 ();
 FILLER_ASAP7_75t_R FILLER_0_47_806 ();
 FILLER_ASAP7_75t_R FILLER_0_47_819 ();
 DECAPx2_ASAP7_75t_R FILLER_0_47_827 ();
 DECAPx6_ASAP7_75t_R FILLER_0_47_845 ();
 DECAPx1_ASAP7_75t_R FILLER_0_47_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_863 ();
 FILLER_ASAP7_75t_R FILLER_0_47_874 ();
 FILLER_ASAP7_75t_R FILLER_0_47_882 ();
 DECAPx1_ASAP7_75t_R FILLER_0_47_887 ();
 FILLER_ASAP7_75t_R FILLER_0_47_897 ();
 DECAPx2_ASAP7_75t_R FILLER_0_47_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_911 ();
 DECAPx2_ASAP7_75t_R FILLER_0_47_919 ();
 DECAPx2_ASAP7_75t_R FILLER_0_47_927 ();
 FILLER_ASAP7_75t_R FILLER_0_47_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_955 ();
 DECAPx2_ASAP7_75t_R FILLER_0_47_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_968 ();
 FILLER_ASAP7_75t_R FILLER_0_47_977 ();
 FILLER_ASAP7_75t_R FILLER_0_47_999 ();
 DECAPx4_ASAP7_75t_R FILLER_0_47_1007 ();
 FILLER_ASAP7_75t_R FILLER_0_47_1017 ();
 FILLER_ASAP7_75t_R FILLER_0_47_1025 ();
 FILLER_ASAP7_75t_R FILLER_0_47_1033 ();
 FILLER_ASAP7_75t_R FILLER_0_47_1041 ();
 DECAPx2_ASAP7_75t_R FILLER_0_47_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_1055 ();
 FILLER_ASAP7_75t_R FILLER_0_47_1064 ();
 FILLER_ASAP7_75t_R FILLER_0_47_1074 ();
 DECAPx1_ASAP7_75t_R FILLER_0_47_1082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_1118 ();
 FILLER_ASAP7_75t_R FILLER_0_47_1152 ();
 DECAPx6_ASAP7_75t_R FILLER_0_47_1160 ();
 FILLER_ASAP7_75t_R FILLER_0_47_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_1176 ();
 DECAPx4_ASAP7_75t_R FILLER_0_47_1184 ();
 DECAPx4_ASAP7_75t_R FILLER_0_47_1200 ();
 FILLER_ASAP7_75t_R FILLER_0_47_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_1212 ();
 FILLER_ASAP7_75t_R FILLER_0_47_1219 ();
 FILLER_ASAP7_75t_R FILLER_0_47_1227 ();
 DECAPx4_ASAP7_75t_R FILLER_0_47_1234 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_1244 ();
 FILLER_ASAP7_75t_R FILLER_0_47_1251 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_1253 ();
 DECAPx2_ASAP7_75t_R FILLER_0_47_1261 ();
 FILLER_ASAP7_75t_R FILLER_0_47_1272 ();
 DECAPx1_ASAP7_75t_R FILLER_0_47_1284 ();
 FILLER_ASAP7_75t_R FILLER_0_47_1296 ();
 DECAPx1_ASAP7_75t_R FILLER_0_47_1303 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_1307 ();
 FILLER_ASAP7_75t_R FILLER_0_47_1313 ();
 FILLER_ASAP7_75t_R FILLER_0_47_1325 ();
 DECAPx1_ASAP7_75t_R FILLER_0_47_1330 ();
 DECAPx4_ASAP7_75t_R FILLER_0_47_1340 ();
 FILLER_ASAP7_75t_R FILLER_0_47_1350 ();
 DECAPx6_ASAP7_75t_R FILLER_0_47_1362 ();
 DECAPx2_ASAP7_75t_R FILLER_0_47_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_48_24 ();
 DECAPx2_ASAP7_75t_R FILLER_0_48_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_44 ();
 FILLER_ASAP7_75t_R FILLER_0_48_53 ();
 FILLER_ASAP7_75t_R FILLER_0_48_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_60 ();
 FILLER_ASAP7_75t_R FILLER_0_48_67 ();
 DECAPx1_ASAP7_75t_R FILLER_0_48_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_85 ();
 FILLER_ASAP7_75t_R FILLER_0_48_92 ();
 FILLER_ASAP7_75t_R FILLER_0_48_100 ();
 FILLER_ASAP7_75t_R FILLER_0_48_108 ();
 FILLER_ASAP7_75t_R FILLER_0_48_116 ();
 DECAPx2_ASAP7_75t_R FILLER_0_48_124 ();
 FILLER_ASAP7_75t_R FILLER_0_48_130 ();
 DECAPx2_ASAP7_75t_R FILLER_0_48_138 ();
 FILLER_ASAP7_75t_R FILLER_0_48_144 ();
 DECAPx2_ASAP7_75t_R FILLER_0_48_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_157 ();
 FILLER_ASAP7_75t_R FILLER_0_48_164 ();
 DECAPx4_ASAP7_75t_R FILLER_0_48_172 ();
 FILLER_ASAP7_75t_R FILLER_0_48_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_184 ();
 FILLER_ASAP7_75t_R FILLER_0_48_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_193 ();
 FILLER_ASAP7_75t_R FILLER_0_48_210 ();
 DECAPx1_ASAP7_75t_R FILLER_0_48_218 ();
 FILLER_ASAP7_75t_R FILLER_0_48_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_230 ();
 DECAPx2_ASAP7_75t_R FILLER_0_48_237 ();
 FILLER_ASAP7_75t_R FILLER_0_48_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_245 ();
 FILLER_ASAP7_75t_R FILLER_0_48_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_254 ();
 FILLER_ASAP7_75t_R FILLER_0_48_260 ();
 FILLER_ASAP7_75t_R FILLER_0_48_268 ();
 FILLER_ASAP7_75t_R FILLER_0_48_278 ();
 FILLER_ASAP7_75t_R FILLER_0_48_291 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_299 ();
 DECAPx6_ASAP7_75t_R FILLER_0_48_321 ();
 FILLER_ASAP7_75t_R FILLER_0_48_335 ();
 FILLER_ASAP7_75t_R FILLER_0_48_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_344 ();
 FILLER_ASAP7_75t_R FILLER_0_48_350 ();
 DECAPx1_ASAP7_75t_R FILLER_0_48_358 ();
 FILLER_ASAP7_75t_R FILLER_0_48_368 ();
 DECAPx1_ASAP7_75t_R FILLER_0_48_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_384 ();
 DECAPx1_ASAP7_75t_R FILLER_0_48_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_399 ();
 DECAPx1_ASAP7_75t_R FILLER_0_48_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_414 ();
 DECAPx6_ASAP7_75t_R FILLER_0_48_426 ();
 DECAPx2_ASAP7_75t_R FILLER_0_48_440 ();
 FILLER_ASAP7_75t_R FILLER_0_48_452 ();
 FILLER_ASAP7_75t_R FILLER_0_48_460 ();
 DECAPx6_ASAP7_75t_R FILLER_0_48_464 ();
 DECAPx2_ASAP7_75t_R FILLER_0_48_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_484 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_491 ();
 DECAPx2_ASAP7_75t_R FILLER_0_48_513 ();
 FILLER_ASAP7_75t_R FILLER_0_48_519 ();
 DECAPx1_ASAP7_75t_R FILLER_0_48_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_531 ();
 DECAPx2_ASAP7_75t_R FILLER_0_48_540 ();
 FILLER_ASAP7_75t_R FILLER_0_48_546 ();
 FILLER_ASAP7_75t_R FILLER_0_48_554 ();
 DECAPx4_ASAP7_75t_R FILLER_0_48_562 ();
 FILLER_ASAP7_75t_R FILLER_0_48_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_574 ();
 FILLER_ASAP7_75t_R FILLER_0_48_578 ();
 FILLER_ASAP7_75t_R FILLER_0_48_588 ();
 DECAPx6_ASAP7_75t_R FILLER_0_48_593 ();
 FILLER_ASAP7_75t_R FILLER_0_48_607 ();
 DECAPx4_ASAP7_75t_R FILLER_0_48_617 ();
 FILLER_ASAP7_75t_R FILLER_0_48_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_629 ();
 DECAPx6_ASAP7_75t_R FILLER_0_48_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_656 ();
 FILLER_ASAP7_75t_R FILLER_0_48_669 ();
 FILLER_ASAP7_75t_R FILLER_0_48_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_681 ();
 DECAPx1_ASAP7_75t_R FILLER_0_48_692 ();
 FILLER_ASAP7_75t_R FILLER_0_48_699 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_713 ();
 DECAPx6_ASAP7_75t_R FILLER_0_48_735 ();
 DECAPx1_ASAP7_75t_R FILLER_0_48_749 ();
 FILLER_ASAP7_75t_R FILLER_0_48_756 ();
 DECAPx1_ASAP7_75t_R FILLER_0_48_768 ();
 FILLER_ASAP7_75t_R FILLER_0_48_782 ();
 FILLER_ASAP7_75t_R FILLER_0_48_787 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_819 ();
 FILLER_ASAP7_75t_R FILLER_0_48_826 ();
 FILLER_ASAP7_75t_R FILLER_0_48_850 ();
 FILLER_ASAP7_75t_R FILLER_0_48_862 ();
 FILLER_ASAP7_75t_R FILLER_0_48_874 ();
 FILLER_ASAP7_75t_R FILLER_0_48_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_887 ();
 FILLER_ASAP7_75t_R FILLER_0_48_909 ();
 DECAPx4_ASAP7_75t_R FILLER_0_48_914 ();
 FILLER_ASAP7_75t_R FILLER_0_48_924 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_926 ();
 FILLER_ASAP7_75t_R FILLER_0_48_935 ();
 FILLER_ASAP7_75t_R FILLER_0_48_943 ();
 FILLER_ASAP7_75t_R FILLER_0_48_951 ();
 FILLER_ASAP7_75t_R FILLER_0_48_961 ();
 DECAPx6_ASAP7_75t_R FILLER_0_48_969 ();
 FILLER_ASAP7_75t_R FILLER_0_48_993 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1003 ();
 DECAPx4_ASAP7_75t_R FILLER_0_48_1011 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_1023 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1029 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1041 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1049 ();
 DECAPx1_ASAP7_75t_R FILLER_0_48_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_1065 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1070 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1078 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1090 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_1132 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1154 ();
 DECAPx1_ASAP7_75t_R FILLER_0_48_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_1166 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1177 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1191 ();
 DECAPx2_ASAP7_75t_R FILLER_0_48_1200 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1214 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1221 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1228 ();
 DECAPx1_ASAP7_75t_R FILLER_0_48_1235 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_1248 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_1270 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1275 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1284 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_1286 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1293 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1301 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_1303 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1314 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1323 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1329 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1334 ();
 DECAPx1_ASAP7_75t_R FILLER_0_48_1344 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1368 ();
 FILLER_ASAP7_75t_R FILLER_0_48_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_49_24 ();
 DECAPx6_ASAP7_75t_R FILLER_0_49_44 ();
 DECAPx2_ASAP7_75t_R FILLER_0_49_58 ();
 FILLER_ASAP7_75t_R FILLER_0_49_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_73 ();
 FILLER_ASAP7_75t_R FILLER_0_49_81 ();
 FILLER_ASAP7_75t_R FILLER_0_49_89 ();
 FILLER_ASAP7_75t_R FILLER_0_49_99 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_128 ();
 DECAPx2_ASAP7_75t_R FILLER_0_49_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_141 ();
 FILLER_ASAP7_75t_R FILLER_0_49_148 ();
 FILLER_ASAP7_75t_R FILLER_0_49_162 ();
 FILLER_ASAP7_75t_R FILLER_0_49_167 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_175 ();
 DECAPx6_ASAP7_75t_R FILLER_0_49_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_211 ();
 FILLER_ASAP7_75t_R FILLER_0_49_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_220 ();
 FILLER_ASAP7_75t_R FILLER_0_49_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_229 ();
 FILLER_ASAP7_75t_R FILLER_0_49_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_238 ();
 FILLER_ASAP7_75t_R FILLER_0_49_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_247 ();
 DECAPx1_ASAP7_75t_R FILLER_0_49_254 ();
 FILLER_ASAP7_75t_R FILLER_0_49_264 ();
 DECAPx2_ASAP7_75t_R FILLER_0_49_272 ();
 FILLER_ASAP7_75t_R FILLER_0_49_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_280 ();
 DECAPx4_ASAP7_75t_R FILLER_0_49_284 ();
 DECAPx4_ASAP7_75t_R FILLER_0_49_300 ();
 FILLER_ASAP7_75t_R FILLER_0_49_310 ();
 DECAPx2_ASAP7_75t_R FILLER_0_49_334 ();
 DECAPx1_ASAP7_75t_R FILLER_0_49_361 ();
 FILLER_ASAP7_75t_R FILLER_0_49_370 ();
 FILLER_ASAP7_75t_R FILLER_0_49_382 ();
 DECAPx2_ASAP7_75t_R FILLER_0_49_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_400 ();
 FILLER_ASAP7_75t_R FILLER_0_49_411 ();
 DECAPx6_ASAP7_75t_R FILLER_0_49_419 ();
 DECAPx1_ASAP7_75t_R FILLER_0_49_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_437 ();
 FILLER_ASAP7_75t_R FILLER_0_49_446 ();
 DECAPx2_ASAP7_75t_R FILLER_0_49_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_460 ();
 DECAPx6_ASAP7_75t_R FILLER_0_49_467 ();
 DECAPx1_ASAP7_75t_R FILLER_0_49_481 ();
 FILLER_ASAP7_75t_R FILLER_0_49_491 ();
 FILLER_ASAP7_75t_R FILLER_0_49_505 ();
 FILLER_ASAP7_75t_R FILLER_0_49_513 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_521 ();
 DECAPx4_ASAP7_75t_R FILLER_0_49_543 ();
 DECAPx6_ASAP7_75t_R FILLER_0_49_560 ();
 FILLER_ASAP7_75t_R FILLER_0_49_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_632 ();
 DECAPx1_ASAP7_75t_R FILLER_0_49_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_658 ();
 FILLER_ASAP7_75t_R FILLER_0_49_663 ();
 FILLER_ASAP7_75t_R FILLER_0_49_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_670 ();
 FILLER_ASAP7_75t_R FILLER_0_49_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_681 ();
 DECAPx1_ASAP7_75t_R FILLER_0_49_690 ();
 FILLER_ASAP7_75t_R FILLER_0_49_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_702 ();
 FILLER_ASAP7_75t_R FILLER_0_49_709 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_717 ();
 DECAPx6_ASAP7_75t_R FILLER_0_49_739 ();
 DECAPx4_ASAP7_75t_R FILLER_0_49_773 ();
 FILLER_ASAP7_75t_R FILLER_0_49_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_785 ();
 FILLER_ASAP7_75t_R FILLER_0_49_797 ();
 DECAPx2_ASAP7_75t_R FILLER_0_49_802 ();
 FILLER_ASAP7_75t_R FILLER_0_49_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_810 ();
 FILLER_ASAP7_75t_R FILLER_0_49_832 ();
 DECAPx4_ASAP7_75t_R FILLER_0_49_837 ();
 FILLER_ASAP7_75t_R FILLER_0_49_847 ();
 FILLER_ASAP7_75t_R FILLER_0_49_867 ();
 DECAPx6_ASAP7_75t_R FILLER_0_49_872 ();
 DECAPx2_ASAP7_75t_R FILLER_0_49_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_892 ();
 DECAPx2_ASAP7_75t_R FILLER_0_49_896 ();
 FILLER_ASAP7_75t_R FILLER_0_49_902 ();
 DECAPx6_ASAP7_75t_R FILLER_0_49_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_924 ();
 DECAPx1_ASAP7_75t_R FILLER_0_49_927 ();
 FILLER_ASAP7_75t_R FILLER_0_49_953 ();
 DECAPx6_ASAP7_75t_R FILLER_0_49_960 ();
 DECAPx1_ASAP7_75t_R FILLER_0_49_974 ();
 DECAPx4_ASAP7_75t_R FILLER_0_49_984 ();
 FILLER_ASAP7_75t_R FILLER_0_49_1004 ();
 DECAPx6_ASAP7_75t_R FILLER_0_49_1013 ();
 FILLER_ASAP7_75t_R FILLER_0_49_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_1029 ();
 DECAPx1_ASAP7_75t_R FILLER_0_49_1036 ();
 DECAPx4_ASAP7_75t_R FILLER_0_49_1046 ();
 DECAPx2_ASAP7_75t_R FILLER_0_49_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_1072 ();
 DECAPx1_ASAP7_75t_R FILLER_0_49_1093 ();
 DECAPx1_ASAP7_75t_R FILLER_0_49_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_1111 ();
 DECAPx6_ASAP7_75t_R FILLER_0_49_1115 ();
 DECAPx2_ASAP7_75t_R FILLER_0_49_1129 ();
 DECAPx4_ASAP7_75t_R FILLER_0_49_1141 ();
 FILLER_ASAP7_75t_R FILLER_0_49_1151 ();
 DECAPx1_ASAP7_75t_R FILLER_0_49_1156 ();
 FILLER_ASAP7_75t_R FILLER_0_49_1168 ();
 DECAPx1_ASAP7_75t_R FILLER_0_49_1178 ();
 FILLER_ASAP7_75t_R FILLER_0_49_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_1191 ();
 FILLER_ASAP7_75t_R FILLER_0_49_1197 ();
 FILLER_ASAP7_75t_R FILLER_0_49_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_1221 ();
 FILLER_ASAP7_75t_R FILLER_0_49_1227 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_1229 ();
 FILLER_ASAP7_75t_R FILLER_0_49_1240 ();
 FILLER_ASAP7_75t_R FILLER_0_49_1248 ();
 DECAPx2_ASAP7_75t_R FILLER_0_49_1255 ();
 FILLER_ASAP7_75t_R FILLER_0_49_1268 ();
 FILLER_ASAP7_75t_R FILLER_0_49_1276 ();
 FILLER_ASAP7_75t_R FILLER_0_49_1284 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_1286 ();
 DECAPx1_ASAP7_75t_R FILLER_0_49_1292 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_1296 ();
 FILLER_ASAP7_75t_R FILLER_0_49_1307 ();
 FILLER_ASAP7_75t_R FILLER_0_49_1319 ();
 FILLER_ASAP7_75t_R FILLER_0_49_1328 ();
 FILLER_ASAP7_75t_R FILLER_0_49_1336 ();
 DECAPx2_ASAP7_75t_R FILLER_0_49_1349 ();
 FILLER_ASAP7_75t_R FILLER_0_49_1355 ();
 DECAPx2_ASAP7_75t_R FILLER_0_49_1365 ();
 FILLER_ASAP7_75t_R FILLER_0_49_1371 ();
 FILLER_ASAP7_75t_R FILLER_0_49_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_50_24 ();
 FILLER_ASAP7_75t_R FILLER_0_50_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_40 ();
 DECAPx2_ASAP7_75t_R FILLER_0_50_47 ();
 FILLER_ASAP7_75t_R FILLER_0_50_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_55 ();
 DECAPx1_ASAP7_75t_R FILLER_0_50_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_66 ();
 DECAPx1_ASAP7_75t_R FILLER_0_50_73 ();
 DECAPx6_ASAP7_75t_R FILLER_0_50_81 ();
 DECAPx1_ASAP7_75t_R FILLER_0_50_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_99 ();
 DECAPx4_ASAP7_75t_R FILLER_0_50_112 ();
 FILLER_ASAP7_75t_R FILLER_0_50_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_124 ();
 FILLER_ASAP7_75t_R FILLER_0_50_135 ();
 FILLER_ASAP7_75t_R FILLER_0_50_140 ();
 FILLER_ASAP7_75t_R FILLER_0_50_148 ();
 FILLER_ASAP7_75t_R FILLER_0_50_162 ();
 FILLER_ASAP7_75t_R FILLER_0_50_171 ();
 DECAPx4_ASAP7_75t_R FILLER_0_50_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_187 ();
 DECAPx4_ASAP7_75t_R FILLER_0_50_194 ();
 FILLER_ASAP7_75t_R FILLER_0_50_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_206 ();
 DECAPx4_ASAP7_75t_R FILLER_0_50_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_229 ();
 DECAPx4_ASAP7_75t_R FILLER_0_50_240 ();
 FILLER_ASAP7_75t_R FILLER_0_50_250 ();
 DECAPx1_ASAP7_75t_R FILLER_0_50_258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_290 ();
 FILLER_ASAP7_75t_R FILLER_0_50_312 ();
 DECAPx6_ASAP7_75t_R FILLER_0_50_317 ();
 FILLER_ASAP7_75t_R FILLER_0_50_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_333 ();
 FILLER_ASAP7_75t_R FILLER_0_50_346 ();
 DECAPx4_ASAP7_75t_R FILLER_0_50_351 ();
 FILLER_ASAP7_75t_R FILLER_0_50_365 ();
 DECAPx2_ASAP7_75t_R FILLER_0_50_377 ();
 FILLER_ASAP7_75t_R FILLER_0_50_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_385 ();
 DECAPx2_ASAP7_75t_R FILLER_0_50_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_398 ();
 DECAPx1_ASAP7_75t_R FILLER_0_50_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_423 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_452 ();
 FILLER_ASAP7_75t_R FILLER_0_50_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_461 ();
 DECAPx2_ASAP7_75t_R FILLER_0_50_464 ();
 FILLER_ASAP7_75t_R FILLER_0_50_470 ();
 FILLER_ASAP7_75t_R FILLER_0_50_478 ();
 FILLER_ASAP7_75t_R FILLER_0_50_486 ();
 DECAPx6_ASAP7_75t_R FILLER_0_50_494 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_536 ();
 DECAPx6_ASAP7_75t_R FILLER_0_50_558 ();
 FILLER_ASAP7_75t_R FILLER_0_50_578 ();
 DECAPx1_ASAP7_75t_R FILLER_0_50_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_592 ();
 FILLER_ASAP7_75t_R FILLER_0_50_604 ();
 FILLER_ASAP7_75t_R FILLER_0_50_609 ();
 DECAPx4_ASAP7_75t_R FILLER_0_50_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_629 ();
 FILLER_ASAP7_75t_R FILLER_0_50_642 ();
 DECAPx2_ASAP7_75t_R FILLER_0_50_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_661 ();
 DECAPx2_ASAP7_75t_R FILLER_0_50_670 ();
 FILLER_ASAP7_75t_R FILLER_0_50_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_678 ();
 FILLER_ASAP7_75t_R FILLER_0_50_685 ();
 DECAPx2_ASAP7_75t_R FILLER_0_50_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_699 ();
 DECAPx4_ASAP7_75t_R FILLER_0_50_708 ();
 FILLER_ASAP7_75t_R FILLER_0_50_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_720 ();
 DECAPx4_ASAP7_75t_R FILLER_0_50_732 ();
 DECAPx2_ASAP7_75t_R FILLER_0_50_748 ();
 FILLER_ASAP7_75t_R FILLER_0_50_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_756 ();
 DECAPx6_ASAP7_75t_R FILLER_0_50_767 ();
 FILLER_ASAP7_75t_R FILLER_0_50_781 ();
 DECAPx1_ASAP7_75t_R FILLER_0_50_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_791 ();
 DECAPx6_ASAP7_75t_R FILLER_0_50_798 ();
 FILLER_ASAP7_75t_R FILLER_0_50_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_814 ();
 DECAPx2_ASAP7_75t_R FILLER_0_50_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_829 ();
 DECAPx6_ASAP7_75t_R FILLER_0_50_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_847 ();
 DECAPx2_ASAP7_75t_R FILLER_0_50_868 ();
 FILLER_ASAP7_75t_R FILLER_0_50_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_876 ();
 FILLER_ASAP7_75t_R FILLER_0_50_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_885 ();
 FILLER_ASAP7_75t_R FILLER_0_50_892 ();
 DECAPx4_ASAP7_75t_R FILLER_0_50_897 ();
 DECAPx1_ASAP7_75t_R FILLER_0_50_913 ();
 DECAPx1_ASAP7_75t_R FILLER_0_50_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_924 ();
 DECAPx1_ASAP7_75t_R FILLER_0_50_931 ();
 FILLER_ASAP7_75t_R FILLER_0_50_945 ();
 DECAPx2_ASAP7_75t_R FILLER_0_50_953 ();
 FILLER_ASAP7_75t_R FILLER_0_50_967 ();
 DECAPx6_ASAP7_75t_R FILLER_0_50_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_995 ();
 FILLER_ASAP7_75t_R FILLER_0_50_1001 ();
 DECAPx2_ASAP7_75t_R FILLER_0_50_1009 ();
 FILLER_ASAP7_75t_R FILLER_0_50_1021 ();
 FILLER_ASAP7_75t_R FILLER_0_50_1028 ();
 FILLER_ASAP7_75t_R FILLER_0_50_1036 ();
 DECAPx2_ASAP7_75t_R FILLER_0_50_1049 ();
 FILLER_ASAP7_75t_R FILLER_0_50_1055 ();
 FILLER_ASAP7_75t_R FILLER_0_50_1071 ();
 DECAPx2_ASAP7_75t_R FILLER_0_50_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_1085 ();
 FILLER_ASAP7_75t_R FILLER_0_50_1092 ();
 DECAPx4_ASAP7_75t_R FILLER_0_50_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_1110 ();
 FILLER_ASAP7_75t_R FILLER_0_50_1121 ();
 FILLER_ASAP7_75t_R FILLER_0_50_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_1131 ();
 DECAPx2_ASAP7_75t_R FILLER_0_50_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_1144 ();
 FILLER_ASAP7_75t_R FILLER_0_50_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_1150 ();
 DECAPx1_ASAP7_75t_R FILLER_0_50_1157 ();
 DECAPx2_ASAP7_75t_R FILLER_0_50_1167 ();
 DECAPx2_ASAP7_75t_R FILLER_0_50_1179 ();
 DECAPx1_ASAP7_75t_R FILLER_0_50_1200 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_1204 ();
 FILLER_ASAP7_75t_R FILLER_0_50_1215 ();
 FILLER_ASAP7_75t_R FILLER_0_50_1227 ();
 FILLER_ASAP7_75t_R FILLER_0_50_1239 ();
 DECAPx2_ASAP7_75t_R FILLER_0_50_1249 ();
 FILLER_ASAP7_75t_R FILLER_0_50_1255 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_1257 ();
 FILLER_ASAP7_75t_R FILLER_0_50_1265 ();
 FILLER_ASAP7_75t_R FILLER_0_50_1273 ();
 FILLER_ASAP7_75t_R FILLER_0_50_1281 ();
 DECAPx1_ASAP7_75t_R FILLER_0_50_1293 ();
 FILLER_ASAP7_75t_R FILLER_0_50_1303 ();
 DECAPx1_ASAP7_75t_R FILLER_0_50_1311 ();
 FILLER_ASAP7_75t_R FILLER_0_50_1325 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_1327 ();
 FILLER_ASAP7_75t_R FILLER_0_50_1334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_1342 ();
 FILLER_ASAP7_75t_R FILLER_0_50_1364 ();
 DECAPx1_ASAP7_75t_R FILLER_0_50_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_51_24 ();
 FILLER_ASAP7_75t_R FILLER_0_51_34 ();
 FILLER_ASAP7_75t_R FILLER_0_51_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_44 ();
 DECAPx2_ASAP7_75t_R FILLER_0_51_51 ();
 DECAPx1_ASAP7_75t_R FILLER_0_51_63 ();
 DECAPx1_ASAP7_75t_R FILLER_0_51_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_78 ();
 FILLER_ASAP7_75t_R FILLER_0_51_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_93 ();
 DECAPx1_ASAP7_75t_R FILLER_0_51_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_104 ();
 DECAPx2_ASAP7_75t_R FILLER_0_51_117 ();
 FILLER_ASAP7_75t_R FILLER_0_51_123 ();
 DECAPx2_ASAP7_75t_R FILLER_0_51_131 ();
 FILLER_ASAP7_75t_R FILLER_0_51_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_149 ();
 FILLER_ASAP7_75t_R FILLER_0_51_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_162 ();
 FILLER_ASAP7_75t_R FILLER_0_51_169 ();
 DECAPx2_ASAP7_75t_R FILLER_0_51_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_182 ();
 DECAPx1_ASAP7_75t_R FILLER_0_51_189 ();
 FILLER_ASAP7_75t_R FILLER_0_51_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_198 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_205 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_227 ();
 FILLER_ASAP7_75t_R FILLER_0_51_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_254 ();
 FILLER_ASAP7_75t_R FILLER_0_51_267 ();
 FILLER_ASAP7_75t_R FILLER_0_51_283 ();
 FILLER_ASAP7_75t_R FILLER_0_51_295 ();
 DECAPx1_ASAP7_75t_R FILLER_0_51_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_307 ();
 DECAPx4_ASAP7_75t_R FILLER_0_51_329 ();
 FILLER_ASAP7_75t_R FILLER_0_51_339 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_51_366 ();
 DECAPx1_ASAP7_75t_R FILLER_0_51_380 ();
 FILLER_ASAP7_75t_R FILLER_0_51_388 ();
 FILLER_ASAP7_75t_R FILLER_0_51_396 ();
 FILLER_ASAP7_75t_R FILLER_0_51_418 ();
 FILLER_ASAP7_75t_R FILLER_0_51_427 ();
 DECAPx4_ASAP7_75t_R FILLER_0_51_435 ();
 FILLER_ASAP7_75t_R FILLER_0_51_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_447 ();
 FILLER_ASAP7_75t_R FILLER_0_51_454 ();
 FILLER_ASAP7_75t_R FILLER_0_51_462 ();
 DECAPx6_ASAP7_75t_R FILLER_0_51_470 ();
 DECAPx2_ASAP7_75t_R FILLER_0_51_484 ();
 DECAPx1_ASAP7_75t_R FILLER_0_51_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_500 ();
 DECAPx6_ASAP7_75t_R FILLER_0_51_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_525 ();
 FILLER_ASAP7_75t_R FILLER_0_51_546 ();
 DECAPx4_ASAP7_75t_R FILLER_0_51_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_566 ();
 DECAPx6_ASAP7_75t_R FILLER_0_51_589 ();
 FILLER_ASAP7_75t_R FILLER_0_51_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_605 ();
 FILLER_ASAP7_75t_R FILLER_0_51_614 ();
 FILLER_ASAP7_75t_R FILLER_0_51_622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_630 ();
 FILLER_ASAP7_75t_R FILLER_0_51_652 ();
 FILLER_ASAP7_75t_R FILLER_0_51_662 ();
 FILLER_ASAP7_75t_R FILLER_0_51_672 ();
 DECAPx2_ASAP7_75t_R FILLER_0_51_680 ();
 FILLER_ASAP7_75t_R FILLER_0_51_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_688 ();
 FILLER_ASAP7_75t_R FILLER_0_51_699 ();
 FILLER_ASAP7_75t_R FILLER_0_51_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_708 ();
 DECAPx6_ASAP7_75t_R FILLER_0_51_721 ();
 DECAPx2_ASAP7_75t_R FILLER_0_51_735 ();
 DECAPx4_ASAP7_75t_R FILLER_0_51_747 ();
 FILLER_ASAP7_75t_R FILLER_0_51_757 ();
 DECAPx2_ASAP7_75t_R FILLER_0_51_765 ();
 FILLER_ASAP7_75t_R FILLER_0_51_771 ();
 FILLER_ASAP7_75t_R FILLER_0_51_794 ();
 DECAPx2_ASAP7_75t_R FILLER_0_51_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_810 ();
 DECAPx1_ASAP7_75t_R FILLER_0_51_823 ();
 DECAPx6_ASAP7_75t_R FILLER_0_51_830 ();
 DECAPx2_ASAP7_75t_R FILLER_0_51_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_850 ();
 DECAPx1_ASAP7_75t_R FILLER_0_51_871 ();
 FILLER_ASAP7_75t_R FILLER_0_51_885 ();
 FILLER_ASAP7_75t_R FILLER_0_51_893 ();
 DECAPx1_ASAP7_75t_R FILLER_0_51_901 ();
 DECAPx1_ASAP7_75t_R FILLER_0_51_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_915 ();
 FILLER_ASAP7_75t_R FILLER_0_51_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_924 ();
 FILLER_ASAP7_75t_R FILLER_0_51_927 ();
 FILLER_ASAP7_75t_R FILLER_0_51_939 ();
 FILLER_ASAP7_75t_R FILLER_0_51_951 ();
 FILLER_ASAP7_75t_R FILLER_0_51_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_961 ();
 FILLER_ASAP7_75t_R FILLER_0_51_968 ();
 FILLER_ASAP7_75t_R FILLER_0_51_978 ();
 FILLER_ASAP7_75t_R FILLER_0_51_986 ();
 FILLER_ASAP7_75t_R FILLER_0_51_991 ();
 FILLER_ASAP7_75t_R FILLER_0_51_997 ();
 FILLER_ASAP7_75t_R FILLER_0_51_1004 ();
 FILLER_ASAP7_75t_R FILLER_0_51_1011 ();
 FILLER_ASAP7_75t_R FILLER_0_51_1019 ();
 DECAPx6_ASAP7_75t_R FILLER_0_51_1027 ();
 DECAPx1_ASAP7_75t_R FILLER_0_51_1041 ();
 DECAPx2_ASAP7_75t_R FILLER_0_51_1051 ();
 FILLER_ASAP7_75t_R FILLER_0_51_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_1059 ();
 DECAPx1_ASAP7_75t_R FILLER_0_51_1065 ();
 DECAPx2_ASAP7_75t_R FILLER_0_51_1085 ();
 FILLER_ASAP7_75t_R FILLER_0_51_1091 ();
 FILLER_ASAP7_75t_R FILLER_0_51_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_1106 ();
 DECAPx6_ASAP7_75t_R FILLER_0_51_1113 ();
 FILLER_ASAP7_75t_R FILLER_0_51_1130 ();
 FILLER_ASAP7_75t_R FILLER_0_51_1138 ();
 FILLER_ASAP7_75t_R FILLER_0_51_1152 ();
 DECAPx2_ASAP7_75t_R FILLER_0_51_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_1184 ();
 DECAPx2_ASAP7_75t_R FILLER_0_51_1190 ();
 FILLER_ASAP7_75t_R FILLER_0_51_1196 ();
 FILLER_ASAP7_75t_R FILLER_0_51_1203 ();
 FILLER_ASAP7_75t_R FILLER_0_51_1211 ();
 DECAPx1_ASAP7_75t_R FILLER_0_51_1218 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_1222 ();
 FILLER_ASAP7_75t_R FILLER_0_51_1233 ();
 FILLER_ASAP7_75t_R FILLER_0_51_1240 ();
 FILLER_ASAP7_75t_R FILLER_0_51_1247 ();
 DECAPx2_ASAP7_75t_R FILLER_0_51_1254 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_1260 ();
 DECAPx1_ASAP7_75t_R FILLER_0_51_1267 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_1271 ();
 FILLER_ASAP7_75t_R FILLER_0_51_1283 ();
 FILLER_ASAP7_75t_R FILLER_0_51_1291 ();
 FILLER_ASAP7_75t_R FILLER_0_51_1298 ();
 FILLER_ASAP7_75t_R FILLER_0_51_1305 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_1311 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_1333 ();
 FILLER_ASAP7_75t_R FILLER_0_51_1340 ();
 DECAPx2_ASAP7_75t_R FILLER_0_51_1352 ();
 DECAPx2_ASAP7_75t_R FILLER_0_51_1374 ();
 FILLER_ASAP7_75t_R FILLER_0_51_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_52_24 ();
 FILLER_ASAP7_75t_R FILLER_0_52_38 ();
 FILLER_ASAP7_75t_R FILLER_0_52_46 ();
 FILLER_ASAP7_75t_R FILLER_0_52_54 ();
 FILLER_ASAP7_75t_R FILLER_0_52_61 ();
 DECAPx1_ASAP7_75t_R FILLER_0_52_83 ();
 DECAPx1_ASAP7_75t_R FILLER_0_52_93 ();
 FILLER_ASAP7_75t_R FILLER_0_52_109 ();
 DECAPx1_ASAP7_75t_R FILLER_0_52_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_118 ();
 FILLER_ASAP7_75t_R FILLER_0_52_125 ();
 DECAPx1_ASAP7_75t_R FILLER_0_52_133 ();
 DECAPx4_ASAP7_75t_R FILLER_0_52_143 ();
 FILLER_ASAP7_75t_R FILLER_0_52_153 ();
 FILLER_ASAP7_75t_R FILLER_0_52_160 ();
 DECAPx4_ASAP7_75t_R FILLER_0_52_168 ();
 FILLER_ASAP7_75t_R FILLER_0_52_178 ();
 DECAPx6_ASAP7_75t_R FILLER_0_52_192 ();
 FILLER_ASAP7_75t_R FILLER_0_52_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_208 ();
 FILLER_ASAP7_75t_R FILLER_0_52_217 ();
 FILLER_ASAP7_75t_R FILLER_0_52_225 ();
 DECAPx1_ASAP7_75t_R FILLER_0_52_238 ();
 DECAPx6_ASAP7_75t_R FILLER_0_52_248 ();
 FILLER_ASAP7_75t_R FILLER_0_52_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_264 ();
 DECAPx1_ASAP7_75t_R FILLER_0_52_271 ();
 FILLER_ASAP7_75t_R FILLER_0_52_281 ();
 FILLER_ASAP7_75t_R FILLER_0_52_289 ();
 DECAPx6_ASAP7_75t_R FILLER_0_52_294 ();
 FILLER_ASAP7_75t_R FILLER_0_52_308 ();
 DECAPx6_ASAP7_75t_R FILLER_0_52_313 ();
 FILLER_ASAP7_75t_R FILLER_0_52_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_329 ();
 FILLER_ASAP7_75t_R FILLER_0_52_336 ();
 DECAPx2_ASAP7_75t_R FILLER_0_52_341 ();
 FILLER_ASAP7_75t_R FILLER_0_52_353 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_358 ();
 DECAPx2_ASAP7_75t_R FILLER_0_52_380 ();
 FILLER_ASAP7_75t_R FILLER_0_52_386 ();
 FILLER_ASAP7_75t_R FILLER_0_52_395 ();
 FILLER_ASAP7_75t_R FILLER_0_52_417 ();
 DECAPx1_ASAP7_75t_R FILLER_0_52_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_428 ();
 FILLER_ASAP7_75t_R FILLER_0_52_439 ();
 DECAPx4_ASAP7_75t_R FILLER_0_52_444 ();
 FILLER_ASAP7_75t_R FILLER_0_52_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_456 ();
 FILLER_ASAP7_75t_R FILLER_0_52_460 ();
 FILLER_ASAP7_75t_R FILLER_0_52_464 ();
 DECAPx2_ASAP7_75t_R FILLER_0_52_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_478 ();
 DECAPx4_ASAP7_75t_R FILLER_0_52_485 ();
 FILLER_ASAP7_75t_R FILLER_0_52_515 ();
 DECAPx2_ASAP7_75t_R FILLER_0_52_537 ();
 FILLER_ASAP7_75t_R FILLER_0_52_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_545 ();
 FILLER_ASAP7_75t_R FILLER_0_52_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_569 ();
 FILLER_ASAP7_75t_R FILLER_0_52_576 ();
 DECAPx4_ASAP7_75t_R FILLER_0_52_600 ();
 FILLER_ASAP7_75t_R FILLER_0_52_610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_640 ();
 FILLER_ASAP7_75t_R FILLER_0_52_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_664 ();
 FILLER_ASAP7_75t_R FILLER_0_52_675 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_687 ();
 DECAPx2_ASAP7_75t_R FILLER_0_52_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_715 ();
 DECAPx2_ASAP7_75t_R FILLER_0_52_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_728 ();
 DECAPx1_ASAP7_75t_R FILLER_0_52_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_741 ();
 DECAPx4_ASAP7_75t_R FILLER_0_52_750 ();
 DECAPx1_ASAP7_75t_R FILLER_0_52_770 ();
 FILLER_ASAP7_75t_R FILLER_0_52_777 ();
 DECAPx1_ASAP7_75t_R FILLER_0_52_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_794 ();
 DECAPx6_ASAP7_75t_R FILLER_0_52_807 ();
 DECAPx1_ASAP7_75t_R FILLER_0_52_821 ();
 FILLER_ASAP7_75t_R FILLER_0_52_846 ();
 DECAPx6_ASAP7_75t_R FILLER_0_52_860 ();
 FILLER_ASAP7_75t_R FILLER_0_52_884 ();
 DECAPx2_ASAP7_75t_R FILLER_0_52_889 ();
 FILLER_ASAP7_75t_R FILLER_0_52_895 ();
 DECAPx2_ASAP7_75t_R FILLER_0_52_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_913 ();
 DECAPx2_ASAP7_75t_R FILLER_0_52_920 ();
 FILLER_ASAP7_75t_R FILLER_0_52_926 ();
 FILLER_ASAP7_75t_R FILLER_0_52_933 ();
 DECAPx2_ASAP7_75t_R FILLER_0_52_945 ();
 FILLER_ASAP7_75t_R FILLER_0_52_957 ();
 DECAPx1_ASAP7_75t_R FILLER_0_52_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_977 ();
 FILLER_ASAP7_75t_R FILLER_0_52_984 ();
 FILLER_ASAP7_75t_R FILLER_0_52_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_998 ();
 DECAPx6_ASAP7_75t_R FILLER_0_52_1005 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1019 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_1031 ();
 DECAPx6_ASAP7_75t_R FILLER_0_52_1038 ();
 DECAPx2_ASAP7_75t_R FILLER_0_52_1052 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1064 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1072 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1080 ();
 DECAPx2_ASAP7_75t_R FILLER_0_52_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_1093 ();
 DECAPx1_ASAP7_75t_R FILLER_0_52_1100 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_1110 ();
 DECAPx2_ASAP7_75t_R FILLER_0_52_1132 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1138 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1145 ();
 DECAPx2_ASAP7_75t_R FILLER_0_52_1157 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1163 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1171 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_1183 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1191 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1199 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1207 ();
 DECAPx2_ASAP7_75t_R FILLER_0_52_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_1221 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1232 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_1234 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1243 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1250 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1262 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1270 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1275 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1285 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1297 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1305 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1313 ();
 DECAPx6_ASAP7_75t_R FILLER_0_52_1321 ();
 DECAPx2_ASAP7_75t_R FILLER_0_52_1335 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_1341 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1362 ();
 FILLER_ASAP7_75t_R FILLER_0_52_1370 ();
 DECAPx1_ASAP7_75t_R FILLER_0_52_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_53_24 ();
 DECAPx1_ASAP7_75t_R FILLER_0_53_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_42 ();
 FILLER_ASAP7_75t_R FILLER_0_53_49 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_56 ();
 FILLER_ASAP7_75t_R FILLER_0_53_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_64 ();
 FILLER_ASAP7_75t_R FILLER_0_53_71 ();
 FILLER_ASAP7_75t_R FILLER_0_53_79 ();
 DECAPx6_ASAP7_75t_R FILLER_0_53_86 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_100 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_112 ();
 DECAPx4_ASAP7_75t_R FILLER_0_53_141 ();
 FILLER_ASAP7_75t_R FILLER_0_53_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_153 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_160 ();
 FILLER_ASAP7_75t_R FILLER_0_53_166 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_174 ();
 FILLER_ASAP7_75t_R FILLER_0_53_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_182 ();
 FILLER_ASAP7_75t_R FILLER_0_53_191 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_205 ();
 FILLER_ASAP7_75t_R FILLER_0_53_212 ();
 DECAPx1_ASAP7_75t_R FILLER_0_53_220 ();
 DECAPx6_ASAP7_75t_R FILLER_0_53_230 ();
 FILLER_ASAP7_75t_R FILLER_0_53_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_246 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_253 ();
 FILLER_ASAP7_75t_R FILLER_0_53_265 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_284 ();
 FILLER_ASAP7_75t_R FILLER_0_53_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_293 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_315 ();
 FILLER_ASAP7_75t_R FILLER_0_53_342 ();
 DECAPx1_ASAP7_75t_R FILLER_0_53_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_354 ();
 FILLER_ASAP7_75t_R FILLER_0_53_358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_366 ();
 DECAPx4_ASAP7_75t_R FILLER_0_53_388 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_431 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_459 ();
 FILLER_ASAP7_75t_R FILLER_0_53_463 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_475 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_484 ();
 DECAPx4_ASAP7_75t_R FILLER_0_53_506 ();
 DECAPx1_ASAP7_75t_R FILLER_0_53_519 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_523 ();
 DECAPx6_ASAP7_75t_R FILLER_0_53_530 ();
 DECAPx1_ASAP7_75t_R FILLER_0_53_544 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_562 ();
 FILLER_ASAP7_75t_R FILLER_0_53_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_570 ();
 FILLER_ASAP7_75t_R FILLER_0_53_579 ();
 DECAPx6_ASAP7_75t_R FILLER_0_53_587 ();
 FILLER_ASAP7_75t_R FILLER_0_53_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_603 ();
 DECAPx6_ASAP7_75t_R FILLER_0_53_625 ();
 DECAPx1_ASAP7_75t_R FILLER_0_53_639 ();
 DECAPx1_ASAP7_75t_R FILLER_0_53_646 ();
 FILLER_ASAP7_75t_R FILLER_0_53_656 ();
 FILLER_ASAP7_75t_R FILLER_0_53_664 ();
 DECAPx1_ASAP7_75t_R FILLER_0_53_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_675 ();
 DECAPx6_ASAP7_75t_R FILLER_0_53_688 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_702 ();
 DECAPx1_ASAP7_75t_R FILLER_0_53_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_723 ();
 FILLER_ASAP7_75t_R FILLER_0_53_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_730 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_737 ();
 FILLER_ASAP7_75t_R FILLER_0_53_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_745 ();
 DECAPx4_ASAP7_75t_R FILLER_0_53_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_762 ();
 DECAPx6_ASAP7_75t_R FILLER_0_53_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_787 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_799 ();
 FILLER_ASAP7_75t_R FILLER_0_53_805 ();
 FILLER_ASAP7_75t_R FILLER_0_53_815 ();
 DECAPx1_ASAP7_75t_R FILLER_0_53_825 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_835 ();
 DECAPx6_ASAP7_75t_R FILLER_0_53_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_861 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_868 ();
 DECAPx6_ASAP7_75t_R FILLER_0_53_890 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_911 ();
 FILLER_ASAP7_75t_R FILLER_0_53_923 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_933 ();
 FILLER_ASAP7_75t_R FILLER_0_53_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_941 ();
 FILLER_ASAP7_75t_R FILLER_0_53_952 ();
 FILLER_ASAP7_75t_R FILLER_0_53_961 ();
 FILLER_ASAP7_75t_R FILLER_0_53_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_970 ();
 FILLER_ASAP7_75t_R FILLER_0_53_977 ();
 DECAPx4_ASAP7_75t_R FILLER_0_53_985 ();
 FILLER_ASAP7_75t_R FILLER_0_53_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_997 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_1004 ();
 FILLER_ASAP7_75t_R FILLER_0_53_1010 ();
 FILLER_ASAP7_75t_R FILLER_0_53_1018 ();
 DECAPx6_ASAP7_75t_R FILLER_0_53_1026 ();
 DECAPx1_ASAP7_75t_R FILLER_0_53_1040 ();
 FILLER_ASAP7_75t_R FILLER_0_53_1050 ();
 FILLER_ASAP7_75t_R FILLER_0_53_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_1060 ();
 FILLER_ASAP7_75t_R FILLER_0_53_1067 ();
 DECAPx4_ASAP7_75t_R FILLER_0_53_1075 ();
 FILLER_ASAP7_75t_R FILLER_0_53_1091 ();
 FILLER_ASAP7_75t_R FILLER_0_53_1099 ();
 FILLER_ASAP7_75t_R FILLER_0_53_1107 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_1115 ();
 FILLER_ASAP7_75t_R FILLER_0_53_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_1123 ();
 DECAPx1_ASAP7_75t_R FILLER_0_53_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_1134 ();
 DECAPx1_ASAP7_75t_R FILLER_0_53_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_1145 ();
 DECAPx6_ASAP7_75t_R FILLER_0_53_1153 ();
 FILLER_ASAP7_75t_R FILLER_0_53_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_1180 ();
 FILLER_ASAP7_75t_R FILLER_0_53_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_1189 ();
 FILLER_ASAP7_75t_R FILLER_0_53_1197 ();
 FILLER_ASAP7_75t_R FILLER_0_53_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_1207 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_1225 ();
 FILLER_ASAP7_75t_R FILLER_0_53_1236 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_1238 ();
 FILLER_ASAP7_75t_R FILLER_0_53_1249 ();
 FILLER_ASAP7_75t_R FILLER_0_53_1261 ();
 FILLER_ASAP7_75t_R FILLER_0_53_1269 ();
 DECAPx1_ASAP7_75t_R FILLER_0_53_1291 ();
 DECAPx1_ASAP7_75t_R FILLER_0_53_1302 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_1306 ();
 FILLER_ASAP7_75t_R FILLER_0_53_1318 ();
 FILLER_ASAP7_75t_R FILLER_0_53_1326 ();
 FILLER_ASAP7_75t_R FILLER_0_53_1334 ();
 FILLER_ASAP7_75t_R FILLER_0_53_1342 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_1350 ();
 FILLER_ASAP7_75t_R FILLER_0_53_1356 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_1358 ();
 FILLER_ASAP7_75t_R FILLER_0_53_1365 ();
 FILLER_ASAP7_75t_R FILLER_0_53_1373 ();
 DECAPx1_ASAP7_75t_R FILLER_0_53_1378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_54_24 ();
 FILLER_ASAP7_75t_R FILLER_0_54_34 ();
 FILLER_ASAP7_75t_R FILLER_0_54_43 ();
 FILLER_ASAP7_75t_R FILLER_0_54_51 ();
 DECAPx1_ASAP7_75t_R FILLER_0_54_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_63 ();
 DECAPx2_ASAP7_75t_R FILLER_0_54_70 ();
 FILLER_ASAP7_75t_R FILLER_0_54_76 ();
 DECAPx2_ASAP7_75t_R FILLER_0_54_88 ();
 FILLER_ASAP7_75t_R FILLER_0_54_97 ();
 FILLER_ASAP7_75t_R FILLER_0_54_105 ();
 FILLER_ASAP7_75t_R FILLER_0_54_114 ();
 DECAPx6_ASAP7_75t_R FILLER_0_54_122 ();
 DECAPx2_ASAP7_75t_R FILLER_0_54_136 ();
 DECAPx2_ASAP7_75t_R FILLER_0_54_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_156 ();
 FILLER_ASAP7_75t_R FILLER_0_54_167 ();
 DECAPx2_ASAP7_75t_R FILLER_0_54_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_183 ();
 FILLER_ASAP7_75t_R FILLER_0_54_192 ();
 FILLER_ASAP7_75t_R FILLER_0_54_200 ();
 DECAPx1_ASAP7_75t_R FILLER_0_54_209 ();
 DECAPx2_ASAP7_75t_R FILLER_0_54_218 ();
 DECAPx1_ASAP7_75t_R FILLER_0_54_230 ();
 FILLER_ASAP7_75t_R FILLER_0_54_240 ();
 DECAPx2_ASAP7_75t_R FILLER_0_54_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_259 ();
 DECAPx6_ASAP7_75t_R FILLER_0_54_263 ();
 DECAPx1_ASAP7_75t_R FILLER_0_54_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_281 ();
 FILLER_ASAP7_75t_R FILLER_0_54_288 ();
 DECAPx1_ASAP7_75t_R FILLER_0_54_296 ();
 DECAPx2_ASAP7_75t_R FILLER_0_54_322 ();
 FILLER_ASAP7_75t_R FILLER_0_54_334 ();
 DECAPx2_ASAP7_75t_R FILLER_0_54_339 ();
 FILLER_ASAP7_75t_R FILLER_0_54_345 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_376 ();
 DECAPx6_ASAP7_75t_R FILLER_0_54_398 ();
 DECAPx2_ASAP7_75t_R FILLER_0_54_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_418 ();
 DECAPx4_ASAP7_75t_R FILLER_0_54_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_436 ();
 DECAPx1_ASAP7_75t_R FILLER_0_54_458 ();
 DECAPx4_ASAP7_75t_R FILLER_0_54_464 ();
 FILLER_ASAP7_75t_R FILLER_0_54_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_476 ();
 DECAPx6_ASAP7_75t_R FILLER_0_54_497 ();
 FILLER_ASAP7_75t_R FILLER_0_54_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_513 ();
 FILLER_ASAP7_75t_R FILLER_0_54_517 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_551 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_558 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_580 ();
 FILLER_ASAP7_75t_R FILLER_0_54_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_604 ();
 FILLER_ASAP7_75t_R FILLER_0_54_615 ();
 DECAPx2_ASAP7_75t_R FILLER_0_54_623 ();
 FILLER_ASAP7_75t_R FILLER_0_54_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_631 ();
 DECAPx1_ASAP7_75t_R FILLER_0_54_652 ();
 DECAPx1_ASAP7_75t_R FILLER_0_54_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_668 ();
 DECAPx2_ASAP7_75t_R FILLER_0_54_679 ();
 FILLER_ASAP7_75t_R FILLER_0_54_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_687 ();
 DECAPx2_ASAP7_75t_R FILLER_0_54_698 ();
 FILLER_ASAP7_75t_R FILLER_0_54_704 ();
 FILLER_ASAP7_75t_R FILLER_0_54_714 ();
 DECAPx1_ASAP7_75t_R FILLER_0_54_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_726 ();
 FILLER_ASAP7_75t_R FILLER_0_54_733 ();
 FILLER_ASAP7_75t_R FILLER_0_54_739 ();
 DECAPx4_ASAP7_75t_R FILLER_0_54_749 ();
 FILLER_ASAP7_75t_R FILLER_0_54_780 ();
 DECAPx2_ASAP7_75t_R FILLER_0_54_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_796 ();
 DECAPx2_ASAP7_75t_R FILLER_0_54_809 ();
 FILLER_ASAP7_75t_R FILLER_0_54_837 ();
 DECAPx6_ASAP7_75t_R FILLER_0_54_844 ();
 FILLER_ASAP7_75t_R FILLER_0_54_870 ();
 DECAPx4_ASAP7_75t_R FILLER_0_54_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_888 ();
 FILLER_ASAP7_75t_R FILLER_0_54_895 ();
 FILLER_ASAP7_75t_R FILLER_0_54_903 ();
 DECAPx2_ASAP7_75t_R FILLER_0_54_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_919 ();
 FILLER_ASAP7_75t_R FILLER_0_54_930 ();
 FILLER_ASAP7_75t_R FILLER_0_54_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_940 ();
 FILLER_ASAP7_75t_R FILLER_0_54_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_950 ();
 DECAPx1_ASAP7_75t_R FILLER_0_54_957 ();
 DECAPx4_ASAP7_75t_R FILLER_0_54_967 ();
 FILLER_ASAP7_75t_R FILLER_0_54_987 ();
 FILLER_ASAP7_75t_R FILLER_0_54_995 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_1005 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1014 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1024 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1032 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1040 ();
 DECAPx2_ASAP7_75t_R FILLER_0_54_1053 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_1096 ();
 DECAPx1_ASAP7_75t_R FILLER_0_54_1118 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1133 ();
 DECAPx2_ASAP7_75t_R FILLER_0_54_1138 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1150 ();
 DECAPx2_ASAP7_75t_R FILLER_0_54_1159 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_1165 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1177 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_1186 ();
 DECAPx2_ASAP7_75t_R FILLER_0_54_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_1199 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1206 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1214 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1222 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1234 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1241 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1250 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1262 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1274 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1286 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1294 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1302 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1310 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1318 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1326 ();
 DECAPx1_ASAP7_75t_R FILLER_0_54_1334 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_1338 ();
 DECAPx1_ASAP7_75t_R FILLER_0_54_1345 ();
 DECAPx1_ASAP7_75t_R FILLER_0_54_1359 ();
 DECAPx4_ASAP7_75t_R FILLER_0_54_1369 ();
 FILLER_ASAP7_75t_R FILLER_0_54_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_55_24 ();
 DECAPx2_ASAP7_75t_R FILLER_0_55_38 ();
 FILLER_ASAP7_75t_R FILLER_0_55_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_55_62 ();
 FILLER_ASAP7_75t_R FILLER_0_55_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_74 ();
 DECAPx2_ASAP7_75t_R FILLER_0_55_81 ();
 FILLER_ASAP7_75t_R FILLER_0_55_87 ();
 DECAPx1_ASAP7_75t_R FILLER_0_55_99 ();
 DECAPx1_ASAP7_75t_R FILLER_0_55_113 ();
 FILLER_ASAP7_75t_R FILLER_0_55_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_125 ();
 DECAPx1_ASAP7_75t_R FILLER_0_55_132 ();
 DECAPx4_ASAP7_75t_R FILLER_0_55_146 ();
 DECAPx4_ASAP7_75t_R FILLER_0_55_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_186 ();
 DECAPx1_ASAP7_75t_R FILLER_0_55_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_194 ();
 DECAPx2_ASAP7_75t_R FILLER_0_55_201 ();
 FILLER_ASAP7_75t_R FILLER_0_55_212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_217 ();
 DECAPx6_ASAP7_75t_R FILLER_0_55_239 ();
 DECAPx2_ASAP7_75t_R FILLER_0_55_253 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_265 ();
 DECAPx1_ASAP7_75t_R FILLER_0_55_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_301 ();
 DECAPx2_ASAP7_75t_R FILLER_0_55_305 ();
 FILLER_ASAP7_75t_R FILLER_0_55_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_313 ();
 FILLER_ASAP7_75t_R FILLER_0_55_319 ();
 DECAPx1_ASAP7_75t_R FILLER_0_55_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_335 ();
 FILLER_ASAP7_75t_R FILLER_0_55_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_344 ();
 FILLER_ASAP7_75t_R FILLER_0_55_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_354 ();
 FILLER_ASAP7_75t_R FILLER_0_55_358 ();
 DECAPx2_ASAP7_75t_R FILLER_0_55_366 ();
 FILLER_ASAP7_75t_R FILLER_0_55_378 ();
 DECAPx6_ASAP7_75t_R FILLER_0_55_383 ();
 FILLER_ASAP7_75t_R FILLER_0_55_403 ();
 DECAPx6_ASAP7_75t_R FILLER_0_55_411 ();
 DECAPx1_ASAP7_75t_R FILLER_0_55_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_429 ();
 FILLER_ASAP7_75t_R FILLER_0_55_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_438 ();
 FILLER_ASAP7_75t_R FILLER_0_55_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_447 ();
 FILLER_ASAP7_75t_R FILLER_0_55_451 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_456 ();
 DECAPx2_ASAP7_75t_R FILLER_0_55_478 ();
 FILLER_ASAP7_75t_R FILLER_0_55_484 ();
 DECAPx6_ASAP7_75t_R FILLER_0_55_492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_55_526 ();
 FILLER_ASAP7_75t_R FILLER_0_55_548 ();
 DECAPx2_ASAP7_75t_R FILLER_0_55_571 ();
 DECAPx4_ASAP7_75t_R FILLER_0_55_585 ();
 FILLER_ASAP7_75t_R FILLER_0_55_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_605 ();
 FILLER_ASAP7_75t_R FILLER_0_55_609 ();
 FILLER_ASAP7_75t_R FILLER_0_55_621 ();
 FILLER_ASAP7_75t_R FILLER_0_55_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_637 ();
 FILLER_ASAP7_75t_R FILLER_0_55_646 ();
 FILLER_ASAP7_75t_R FILLER_0_55_654 ();
 DECAPx1_ASAP7_75t_R FILLER_0_55_662 ();
 DECAPx1_ASAP7_75t_R FILLER_0_55_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_682 ();
 FILLER_ASAP7_75t_R FILLER_0_55_693 ();
 DECAPx1_ASAP7_75t_R FILLER_0_55_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_709 ();
 FILLER_ASAP7_75t_R FILLER_0_55_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_718 ();
 DECAPx1_ASAP7_75t_R FILLER_0_55_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_727 ();
 FILLER_ASAP7_75t_R FILLER_0_55_734 ();
 DECAPx6_ASAP7_75t_R FILLER_0_55_744 ();
 FILLER_ASAP7_75t_R FILLER_0_55_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_760 ();
 DECAPx4_ASAP7_75t_R FILLER_0_55_764 ();
 FILLER_ASAP7_75t_R FILLER_0_55_784 ();
 DECAPx4_ASAP7_75t_R FILLER_0_55_807 ();
 DECAPx6_ASAP7_75t_R FILLER_0_55_820 ();
 FILLER_ASAP7_75t_R FILLER_0_55_834 ();
 DECAPx6_ASAP7_75t_R FILLER_0_55_841 ();
 DECAPx2_ASAP7_75t_R FILLER_0_55_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_861 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_874 ();
 FILLER_ASAP7_75t_R FILLER_0_55_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_898 ();
 FILLER_ASAP7_75t_R FILLER_0_55_905 ();
 DECAPx1_ASAP7_75t_R FILLER_0_55_913 ();
 FILLER_ASAP7_75t_R FILLER_0_55_923 ();
 DECAPx1_ASAP7_75t_R FILLER_0_55_927 ();
 DECAPx4_ASAP7_75t_R FILLER_0_55_951 ();
 FILLER_ASAP7_75t_R FILLER_0_55_961 ();
 DECAPx2_ASAP7_75t_R FILLER_0_55_969 ();
 DECAPx1_ASAP7_75t_R FILLER_0_55_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_999 ();
 DECAPx4_ASAP7_75t_R FILLER_0_55_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_1016 ();
 DECAPx4_ASAP7_75t_R FILLER_0_55_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_1038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_1045 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_1067 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_1111 ();
 DECAPx1_ASAP7_75t_R FILLER_0_55_1133 ();
 FILLER_ASAP7_75t_R FILLER_0_55_1149 ();
 DECAPx2_ASAP7_75t_R FILLER_0_55_1156 ();
 FILLER_ASAP7_75t_R FILLER_0_55_1172 ();
 FILLER_ASAP7_75t_R FILLER_0_55_1179 ();
 DECAPx4_ASAP7_75t_R FILLER_0_55_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_1194 ();
 FILLER_ASAP7_75t_R FILLER_0_55_1200 ();
 DECAPx2_ASAP7_75t_R FILLER_0_55_1213 ();
 FILLER_ASAP7_75t_R FILLER_0_55_1219 ();
 FILLER_ASAP7_75t_R FILLER_0_55_1239 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_1241 ();
 FILLER_ASAP7_75t_R FILLER_0_55_1262 ();
 DECAPx2_ASAP7_75t_R FILLER_0_55_1274 ();
 FILLER_ASAP7_75t_R FILLER_0_55_1290 ();
 FILLER_ASAP7_75t_R FILLER_0_55_1299 ();
 FILLER_ASAP7_75t_R FILLER_0_55_1307 ();
 DECAPx1_ASAP7_75t_R FILLER_0_55_1315 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_1319 ();
 FILLER_ASAP7_75t_R FILLER_0_55_1327 ();
 FILLER_ASAP7_75t_R FILLER_0_55_1334 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_1336 ();
 FILLER_ASAP7_75t_R FILLER_0_55_1343 ();
 DECAPx4_ASAP7_75t_R FILLER_0_55_1351 ();
 FILLER_ASAP7_75t_R FILLER_0_55_1367 ();
 DECAPx2_ASAP7_75t_R FILLER_0_55_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_56_24 ();
 FILLER_ASAP7_75t_R FILLER_0_56_44 ();
 DECAPx2_ASAP7_75t_R FILLER_0_56_52 ();
 FILLER_ASAP7_75t_R FILLER_0_56_64 ();
 FILLER_ASAP7_75t_R FILLER_0_56_86 ();
 DECAPx2_ASAP7_75t_R FILLER_0_56_94 ();
 FILLER_ASAP7_75t_R FILLER_0_56_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_108 ();
 FILLER_ASAP7_75t_R FILLER_0_56_115 ();
 DECAPx2_ASAP7_75t_R FILLER_0_56_123 ();
 FILLER_ASAP7_75t_R FILLER_0_56_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_131 ();
 FILLER_ASAP7_75t_R FILLER_0_56_138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_56_148 ();
 FILLER_ASAP7_75t_R FILLER_0_56_154 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_184 ();
 FILLER_ASAP7_75t_R FILLER_0_56_196 ();
 DECAPx6_ASAP7_75t_R FILLER_0_56_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_218 ();
 FILLER_ASAP7_75t_R FILLER_0_56_228 ();
 FILLER_ASAP7_75t_R FILLER_0_56_235 ();
 FILLER_ASAP7_75t_R FILLER_0_56_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_251 ();
 FILLER_ASAP7_75t_R FILLER_0_56_258 ();
 FILLER_ASAP7_75t_R FILLER_0_56_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_274 ();
 DECAPx6_ASAP7_75t_R FILLER_0_56_296 ();
 FILLER_ASAP7_75t_R FILLER_0_56_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_312 ();
 FILLER_ASAP7_75t_R FILLER_0_56_320 ();
 FILLER_ASAP7_75t_R FILLER_0_56_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_330 ();
 DECAPx1_ASAP7_75t_R FILLER_0_56_337 ();
 DECAPx2_ASAP7_75t_R FILLER_0_56_347 ();
 DECAPx2_ASAP7_75t_R FILLER_0_56_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_367 ();
 FILLER_ASAP7_75t_R FILLER_0_56_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_376 ();
 DECAPx1_ASAP7_75t_R FILLER_0_56_384 ();
 DECAPx1_ASAP7_75t_R FILLER_0_56_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_416 ();
 FILLER_ASAP7_75t_R FILLER_0_56_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_425 ();
 FILLER_ASAP7_75t_R FILLER_0_56_434 ();
 FILLER_ASAP7_75t_R FILLER_0_56_460 ();
 FILLER_ASAP7_75t_R FILLER_0_56_464 ();
 DECAPx6_ASAP7_75t_R FILLER_0_56_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_486 ();
 FILLER_ASAP7_75t_R FILLER_0_56_493 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_500 ();
 DECAPx6_ASAP7_75t_R FILLER_0_56_522 ();
 DECAPx1_ASAP7_75t_R FILLER_0_56_536 ();
 DECAPx2_ASAP7_75t_R FILLER_0_56_546 ();
 DECAPx2_ASAP7_75t_R FILLER_0_56_555 ();
 FILLER_ASAP7_75t_R FILLER_0_56_573 ();
 DECAPx6_ASAP7_75t_R FILLER_0_56_581 ();
 DECAPx2_ASAP7_75t_R FILLER_0_56_595 ();
 FILLER_ASAP7_75t_R FILLER_0_56_609 ();
 DECAPx1_ASAP7_75t_R FILLER_0_56_619 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_629 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_651 ();
 DECAPx4_ASAP7_75t_R FILLER_0_56_673 ();
 FILLER_ASAP7_75t_R FILLER_0_56_683 ();
 FILLER_ASAP7_75t_R FILLER_0_56_691 ();
 DECAPx2_ASAP7_75t_R FILLER_0_56_697 ();
 FILLER_ASAP7_75t_R FILLER_0_56_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_705 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_718 ();
 DECAPx6_ASAP7_75t_R FILLER_0_56_740 ();
 DECAPx1_ASAP7_75t_R FILLER_0_56_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_758 ();
 DECAPx2_ASAP7_75t_R FILLER_0_56_769 ();
 FILLER_ASAP7_75t_R FILLER_0_56_781 ();
 FILLER_ASAP7_75t_R FILLER_0_56_786 ();
 DECAPx4_ASAP7_75t_R FILLER_0_56_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_801 ();
 FILLER_ASAP7_75t_R FILLER_0_56_814 ();
 DECAPx2_ASAP7_75t_R FILLER_0_56_824 ();
 FILLER_ASAP7_75t_R FILLER_0_56_842 ();
 FILLER_ASAP7_75t_R FILLER_0_56_865 ();
 FILLER_ASAP7_75t_R FILLER_0_56_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_877 ();
 FILLER_ASAP7_75t_R FILLER_0_56_890 ();
 DECAPx2_ASAP7_75t_R FILLER_0_56_900 ();
 FILLER_ASAP7_75t_R FILLER_0_56_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_908 ();
 DECAPx2_ASAP7_75t_R FILLER_0_56_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_921 ();
 FILLER_ASAP7_75t_R FILLER_0_56_928 ();
 FILLER_ASAP7_75t_R FILLER_0_56_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_942 ();
 FILLER_ASAP7_75t_R FILLER_0_56_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_951 ();
 FILLER_ASAP7_75t_R FILLER_0_56_958 ();
 FILLER_ASAP7_75t_R FILLER_0_56_971 ();
 FILLER_ASAP7_75t_R FILLER_0_56_976 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_1006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_1028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_1050 ();
 FILLER_ASAP7_75t_R FILLER_0_56_1075 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_1085 ();
 DECAPx6_ASAP7_75t_R FILLER_0_56_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_1121 ();
 FILLER_ASAP7_75t_R FILLER_0_56_1132 ();
 DECAPx1_ASAP7_75t_R FILLER_0_56_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_1144 ();
 DECAPx1_ASAP7_75t_R FILLER_0_56_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_1159 ();
 FILLER_ASAP7_75t_R FILLER_0_56_1172 ();
 DECAPx2_ASAP7_75t_R FILLER_0_56_1184 ();
 FILLER_ASAP7_75t_R FILLER_0_56_1190 ();
 DECAPx2_ASAP7_75t_R FILLER_0_56_1198 ();
 DECAPx1_ASAP7_75t_R FILLER_0_56_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_1214 ();
 FILLER_ASAP7_75t_R FILLER_0_56_1235 ();
 FILLER_ASAP7_75t_R FILLER_0_56_1247 ();
 DECAPx2_ASAP7_75t_R FILLER_0_56_1255 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_1261 ();
 FILLER_ASAP7_75t_R FILLER_0_56_1272 ();
 FILLER_ASAP7_75t_R FILLER_0_56_1279 ();
 FILLER_ASAP7_75t_R FILLER_0_56_1291 ();
 FILLER_ASAP7_75t_R FILLER_0_56_1303 ();
 FILLER_ASAP7_75t_R FILLER_0_56_1315 ();
 FILLER_ASAP7_75t_R FILLER_0_56_1323 ();
 FILLER_ASAP7_75t_R FILLER_0_56_1331 ();
 FILLER_ASAP7_75t_R FILLER_0_56_1339 ();
 DECAPx4_ASAP7_75t_R FILLER_0_56_1346 ();
 FILLER_ASAP7_75t_R FILLER_0_56_1356 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_1358 ();
 FILLER_ASAP7_75t_R FILLER_0_56_1365 ();
 DECAPx4_ASAP7_75t_R FILLER_0_56_1370 ();
 FILLER_ASAP7_75t_R FILLER_0_56_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_46 ();
 DECAPx6_ASAP7_75t_R FILLER_0_57_68 ();
 FILLER_ASAP7_75t_R FILLER_0_57_92 ();
 FILLER_ASAP7_75t_R FILLER_0_57_114 ();
 FILLER_ASAP7_75t_R FILLER_0_57_122 ();
 FILLER_ASAP7_75t_R FILLER_0_57_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_131 ();
 DECAPx2_ASAP7_75t_R FILLER_0_57_152 ();
 FILLER_ASAP7_75t_R FILLER_0_57_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_163 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_170 ();
 DECAPx1_ASAP7_75t_R FILLER_0_57_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_196 ();
 FILLER_ASAP7_75t_R FILLER_0_57_203 ();
 DECAPx1_ASAP7_75t_R FILLER_0_57_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_215 ();
 FILLER_ASAP7_75t_R FILLER_0_57_228 ();
 DECAPx1_ASAP7_75t_R FILLER_0_57_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_240 ();
 DECAPx4_ASAP7_75t_R FILLER_0_57_249 ();
 FILLER_ASAP7_75t_R FILLER_0_57_259 ();
 FILLER_ASAP7_75t_R FILLER_0_57_264 ();
 FILLER_ASAP7_75t_R FILLER_0_57_272 ();
 DECAPx2_ASAP7_75t_R FILLER_0_57_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_286 ();
 DECAPx2_ASAP7_75t_R FILLER_0_57_293 ();
 FILLER_ASAP7_75t_R FILLER_0_57_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_301 ();
 FILLER_ASAP7_75t_R FILLER_0_57_308 ();
 DECAPx1_ASAP7_75t_R FILLER_0_57_316 ();
 FILLER_ASAP7_75t_R FILLER_0_57_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_329 ();
 FILLER_ASAP7_75t_R FILLER_0_57_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_338 ();
 DECAPx2_ASAP7_75t_R FILLER_0_57_344 ();
 FILLER_ASAP7_75t_R FILLER_0_57_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_352 ();
 DECAPx2_ASAP7_75t_R FILLER_0_57_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_365 ();
 FILLER_ASAP7_75t_R FILLER_0_57_369 ();
 FILLER_ASAP7_75t_R FILLER_0_57_377 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_382 ();
 DECAPx1_ASAP7_75t_R FILLER_0_57_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_408 ();
 FILLER_ASAP7_75t_R FILLER_0_57_412 ();
 DECAPx1_ASAP7_75t_R FILLER_0_57_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_424 ();
 FILLER_ASAP7_75t_R FILLER_0_57_431 ();
 DECAPx6_ASAP7_75t_R FILLER_0_57_439 ();
 DECAPx1_ASAP7_75t_R FILLER_0_57_453 ();
 FILLER_ASAP7_75t_R FILLER_0_57_460 ();
 FILLER_ASAP7_75t_R FILLER_0_57_468 ();
 DECAPx4_ASAP7_75t_R FILLER_0_57_473 ();
 FILLER_ASAP7_75t_R FILLER_0_57_504 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_509 ();
 DECAPx2_ASAP7_75t_R FILLER_0_57_531 ();
 DECAPx6_ASAP7_75t_R FILLER_0_57_549 ();
 FILLER_ASAP7_75t_R FILLER_0_57_575 ();
 DECAPx4_ASAP7_75t_R FILLER_0_57_583 ();
 DECAPx2_ASAP7_75t_R FILLER_0_57_601 ();
 FILLER_ASAP7_75t_R FILLER_0_57_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_609 ();
 DECAPx6_ASAP7_75t_R FILLER_0_57_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_632 ();
 DECAPx6_ASAP7_75t_R FILLER_0_57_639 ();
 FILLER_ASAP7_75t_R FILLER_0_57_656 ();
 FILLER_ASAP7_75t_R FILLER_0_57_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_663 ();
 DECAPx2_ASAP7_75t_R FILLER_0_57_672 ();
 FILLER_ASAP7_75t_R FILLER_0_57_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_680 ();
 FILLER_ASAP7_75t_R FILLER_0_57_684 ();
 FILLER_ASAP7_75t_R FILLER_0_57_692 ();
 DECAPx2_ASAP7_75t_R FILLER_0_57_702 ();
 FILLER_ASAP7_75t_R FILLER_0_57_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_710 ();
 DECAPx1_ASAP7_75t_R FILLER_0_57_715 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_751 ();
 FILLER_ASAP7_75t_R FILLER_0_57_762 ();
 FILLER_ASAP7_75t_R FILLER_0_57_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_772 ();
 FILLER_ASAP7_75t_R FILLER_0_57_776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_784 ();
 DECAPx4_ASAP7_75t_R FILLER_0_57_806 ();
 FILLER_ASAP7_75t_R FILLER_0_57_816 ();
 DECAPx1_ASAP7_75t_R FILLER_0_57_828 ();
 DECAPx6_ASAP7_75t_R FILLER_0_57_844 ();
 FILLER_ASAP7_75t_R FILLER_0_57_869 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_883 ();
 DECAPx1_ASAP7_75t_R FILLER_0_57_905 ();
 DECAPx4_ASAP7_75t_R FILLER_0_57_915 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_927 ();
 DECAPx6_ASAP7_75t_R FILLER_0_57_949 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_969 ();
 DECAPx4_ASAP7_75t_R FILLER_0_57_991 ();
 FILLER_ASAP7_75t_R FILLER_0_57_1001 ();
 FILLER_ASAP7_75t_R FILLER_0_57_1006 ();
 DECAPx4_ASAP7_75t_R FILLER_0_57_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_1039 ();
 DECAPx6_ASAP7_75t_R FILLER_0_57_1043 ();
 FILLER_ASAP7_75t_R FILLER_0_57_1057 ();
 FILLER_ASAP7_75t_R FILLER_0_57_1062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_57_1069 ();
 DECAPx6_ASAP7_75t_R FILLER_0_57_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_1110 ();
 FILLER_ASAP7_75t_R FILLER_0_57_1131 ();
 FILLER_ASAP7_75t_R FILLER_0_57_1143 ();
 DECAPx1_ASAP7_75t_R FILLER_0_57_1155 ();
 FILLER_ASAP7_75t_R FILLER_0_57_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_1181 ();
 FILLER_ASAP7_75t_R FILLER_0_57_1192 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_1194 ();
 DECAPx2_ASAP7_75t_R FILLER_0_57_1201 ();
 DECAPx1_ASAP7_75t_R FILLER_0_57_1213 ();
 FILLER_ASAP7_75t_R FILLER_0_57_1225 ();
 FILLER_ASAP7_75t_R FILLER_0_57_1237 ();
 FILLER_ASAP7_75t_R FILLER_0_57_1249 ();
 FILLER_ASAP7_75t_R FILLER_0_57_1259 ();
 FILLER_ASAP7_75t_R FILLER_0_57_1267 ();
 FILLER_ASAP7_75t_R FILLER_0_57_1275 ();
 DECAPx2_ASAP7_75t_R FILLER_0_57_1283 ();
 FILLER_ASAP7_75t_R FILLER_0_57_1299 ();
 FILLER_ASAP7_75t_R FILLER_0_57_1311 ();
 FILLER_ASAP7_75t_R FILLER_0_57_1320 ();
 DECAPx2_ASAP7_75t_R FILLER_0_57_1328 ();
 FILLER_ASAP7_75t_R FILLER_0_57_1346 ();
 FILLER_ASAP7_75t_R FILLER_0_57_1354 ();
 FILLER_ASAP7_75t_R FILLER_0_57_1362 ();
 FILLER_ASAP7_75t_R FILLER_0_57_1370 ();
 DECAPx1_ASAP7_75t_R FILLER_0_57_1378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_58_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_58_24 ();
 FILLER_ASAP7_75t_R FILLER_0_58_38 ();
 DECAPx2_ASAP7_75t_R FILLER_0_58_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_52 ();
 DECAPx4_ASAP7_75t_R FILLER_0_58_59 ();
 FILLER_ASAP7_75t_R FILLER_0_58_69 ();
 DECAPx2_ASAP7_75t_R FILLER_0_58_77 ();
 FILLER_ASAP7_75t_R FILLER_0_58_89 ();
 FILLER_ASAP7_75t_R FILLER_0_58_96 ();
 DECAPx4_ASAP7_75t_R FILLER_0_58_104 ();
 FILLER_ASAP7_75t_R FILLER_0_58_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_116 ();
 DECAPx4_ASAP7_75t_R FILLER_0_58_123 ();
 FILLER_ASAP7_75t_R FILLER_0_58_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_135 ();
 FILLER_ASAP7_75t_R FILLER_0_58_142 ();
 DECAPx2_ASAP7_75t_R FILLER_0_58_150 ();
 FILLER_ASAP7_75t_R FILLER_0_58_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_158 ();
 FILLER_ASAP7_75t_R FILLER_0_58_165 ();
 DECAPx6_ASAP7_75t_R FILLER_0_58_178 ();
 FILLER_ASAP7_75t_R FILLER_0_58_192 ();
 FILLER_ASAP7_75t_R FILLER_0_58_197 ();
 DECAPx4_ASAP7_75t_R FILLER_0_58_205 ();
 FILLER_ASAP7_75t_R FILLER_0_58_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_217 ();
 FILLER_ASAP7_75t_R FILLER_0_58_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_228 ();
 DECAPx2_ASAP7_75t_R FILLER_0_58_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_242 ();
 DECAPx4_ASAP7_75t_R FILLER_0_58_251 ();
 FILLER_ASAP7_75t_R FILLER_0_58_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_263 ();
 DECAPx4_ASAP7_75t_R FILLER_0_58_270 ();
 FILLER_ASAP7_75t_R FILLER_0_58_280 ();
 FILLER_ASAP7_75t_R FILLER_0_58_288 ();
 DECAPx6_ASAP7_75t_R FILLER_0_58_297 ();
 DECAPx1_ASAP7_75t_R FILLER_0_58_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_315 ();
 FILLER_ASAP7_75t_R FILLER_0_58_322 ();
 FILLER_ASAP7_75t_R FILLER_0_58_330 ();
 DECAPx1_ASAP7_75t_R FILLER_0_58_338 ();
 FILLER_ASAP7_75t_R FILLER_0_58_350 ();
 DECAPx6_ASAP7_75t_R FILLER_0_58_358 ();
 DECAPx1_ASAP7_75t_R FILLER_0_58_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_382 ();
 FILLER_ASAP7_75t_R FILLER_0_58_390 ();
 FILLER_ASAP7_75t_R FILLER_0_58_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_400 ();
 DECAPx2_ASAP7_75t_R FILLER_0_58_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_410 ();
 DECAPx1_ASAP7_75t_R FILLER_0_58_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_421 ();
 FILLER_ASAP7_75t_R FILLER_0_58_442 ();
 FILLER_ASAP7_75t_R FILLER_0_58_450 ();
 FILLER_ASAP7_75t_R FILLER_0_58_460 ();
 DECAPx2_ASAP7_75t_R FILLER_0_58_464 ();
 FILLER_ASAP7_75t_R FILLER_0_58_470 ();
 FILLER_ASAP7_75t_R FILLER_0_58_475 ();
 FILLER_ASAP7_75t_R FILLER_0_58_498 ();
 FILLER_ASAP7_75t_R FILLER_0_58_506 ();
 FILLER_ASAP7_75t_R FILLER_0_58_514 ();
 FILLER_ASAP7_75t_R FILLER_0_58_522 ();
 FILLER_ASAP7_75t_R FILLER_0_58_530 ();
 FILLER_ASAP7_75t_R FILLER_0_58_536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_58_544 ();
 DECAPx2_ASAP7_75t_R FILLER_0_58_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_565 ();
 DECAPx6_ASAP7_75t_R FILLER_0_58_569 ();
 FILLER_ASAP7_75t_R FILLER_0_58_591 ();
 FILLER_ASAP7_75t_R FILLER_0_58_601 ();
 DECAPx6_ASAP7_75t_R FILLER_0_58_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_621 ();
 FILLER_ASAP7_75t_R FILLER_0_58_634 ();
 DECAPx4_ASAP7_75t_R FILLER_0_58_639 ();
 FILLER_ASAP7_75t_R FILLER_0_58_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_651 ();
 FILLER_ASAP7_75t_R FILLER_0_58_663 ();
 DECAPx4_ASAP7_75t_R FILLER_0_58_671 ();
 FILLER_ASAP7_75t_R FILLER_0_58_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_683 ();
 DECAPx6_ASAP7_75t_R FILLER_0_58_692 ();
 DECAPx1_ASAP7_75t_R FILLER_0_58_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_720 ();
 FILLER_ASAP7_75t_R FILLER_0_58_727 ();
 DECAPx6_ASAP7_75t_R FILLER_0_58_735 ();
 DECAPx2_ASAP7_75t_R FILLER_0_58_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_755 ();
 FILLER_ASAP7_75t_R FILLER_0_58_762 ();
 DECAPx2_ASAP7_75t_R FILLER_0_58_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_773 ();
 FILLER_ASAP7_75t_R FILLER_0_58_780 ();
 FILLER_ASAP7_75t_R FILLER_0_58_788 ();
 DECAPx4_ASAP7_75t_R FILLER_0_58_800 ();
 FILLER_ASAP7_75t_R FILLER_0_58_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_812 ();
 DECAPx4_ASAP7_75t_R FILLER_0_58_824 ();
 DECAPx6_ASAP7_75t_R FILLER_0_58_846 ();
 FILLER_ASAP7_75t_R FILLER_0_58_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_862 ();
 DECAPx4_ASAP7_75t_R FILLER_0_58_866 ();
 FILLER_ASAP7_75t_R FILLER_0_58_898 ();
 DECAPx2_ASAP7_75t_R FILLER_0_58_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_912 ();
 FILLER_ASAP7_75t_R FILLER_0_58_919 ();
 FILLER_ASAP7_75t_R FILLER_0_58_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_944 ();
 DECAPx10_ASAP7_75t_R FILLER_0_58_963 ();
 DECAPx1_ASAP7_75t_R FILLER_0_58_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_989 ();
 FILLER_ASAP7_75t_R FILLER_0_58_1000 ();
 FILLER_ASAP7_75t_R FILLER_0_58_1012 ();
 DECAPx6_ASAP7_75t_R FILLER_0_58_1017 ();
 DECAPx2_ASAP7_75t_R FILLER_0_58_1031 ();
 FILLER_ASAP7_75t_R FILLER_0_58_1058 ();
 FILLER_ASAP7_75t_R FILLER_0_58_1081 ();
 FILLER_ASAP7_75t_R FILLER_0_58_1105 ();
 FILLER_ASAP7_75t_R FILLER_0_58_1113 ();
 DECAPx1_ASAP7_75t_R FILLER_0_58_1118 ();
 FILLER_ASAP7_75t_R FILLER_0_58_1128 ();
 DECAPx2_ASAP7_75t_R FILLER_0_58_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_1141 ();
 FILLER_ASAP7_75t_R FILLER_0_58_1149 ();
 DECAPx1_ASAP7_75t_R FILLER_0_58_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_1165 ();
 FILLER_ASAP7_75t_R FILLER_0_58_1176 ();
 FILLER_ASAP7_75t_R FILLER_0_58_1186 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_1188 ();
 DECAPx2_ASAP7_75t_R FILLER_0_58_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_1201 ();
 DECAPx1_ASAP7_75t_R FILLER_0_58_1212 ();
 FILLER_ASAP7_75t_R FILLER_0_58_1226 ();
 FILLER_ASAP7_75t_R FILLER_0_58_1238 ();
 FILLER_ASAP7_75t_R FILLER_0_58_1250 ();
 FILLER_ASAP7_75t_R FILLER_0_58_1262 ();
 FILLER_ASAP7_75t_R FILLER_0_58_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_0_58_1287 ();
 FILLER_ASAP7_75t_R FILLER_0_58_1301 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_1303 ();
 FILLER_ASAP7_75t_R FILLER_0_58_1307 ();
 FILLER_ASAP7_75t_R FILLER_0_58_1319 ();
 DECAPx1_ASAP7_75t_R FILLER_0_58_1329 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_1333 ();
 FILLER_ASAP7_75t_R FILLER_0_58_1341 ();
 DECAPx2_ASAP7_75t_R FILLER_0_58_1349 ();
 FILLER_ASAP7_75t_R FILLER_0_58_1365 ();
 FILLER_ASAP7_75t_R FILLER_0_58_1372 ();
 FILLER_ASAP7_75t_R FILLER_0_58_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_59_24 ();
 FILLER_ASAP7_75t_R FILLER_0_59_34 ();
 FILLER_ASAP7_75t_R FILLER_0_59_42 ();
 DECAPx1_ASAP7_75t_R FILLER_0_59_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_54 ();
 DECAPx6_ASAP7_75t_R FILLER_0_59_61 ();
 FILLER_ASAP7_75t_R FILLER_0_59_75 ();
 FILLER_ASAP7_75t_R FILLER_0_59_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_89 ();
 FILLER_ASAP7_75t_R FILLER_0_59_96 ();
 FILLER_ASAP7_75t_R FILLER_0_59_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_110 ();
 FILLER_ASAP7_75t_R FILLER_0_59_117 ();
 DECAPx4_ASAP7_75t_R FILLER_0_59_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_136 ();
 FILLER_ASAP7_75t_R FILLER_0_59_143 ();
 FILLER_ASAP7_75t_R FILLER_0_59_153 ();
 DECAPx2_ASAP7_75t_R FILLER_0_59_165 ();
 DECAPx4_ASAP7_75t_R FILLER_0_59_177 ();
 FILLER_ASAP7_75t_R FILLER_0_59_187 ();
 FILLER_ASAP7_75t_R FILLER_0_59_200 ();
 DECAPx4_ASAP7_75t_R FILLER_0_59_208 ();
 FILLER_ASAP7_75t_R FILLER_0_59_218 ();
 DECAPx4_ASAP7_75t_R FILLER_0_59_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_240 ();
 DECAPx6_ASAP7_75t_R FILLER_0_59_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_263 ();
 FILLER_ASAP7_75t_R FILLER_0_59_267 ();
 DECAPx4_ASAP7_75t_R FILLER_0_59_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_285 ();
 DECAPx4_ASAP7_75t_R FILLER_0_59_292 ();
 DECAPx2_ASAP7_75t_R FILLER_0_59_308 ();
 DECAPx2_ASAP7_75t_R FILLER_0_59_320 ();
 DECAPx4_ASAP7_75t_R FILLER_0_59_333 ();
 FILLER_ASAP7_75t_R FILLER_0_59_349 ();
 FILLER_ASAP7_75t_R FILLER_0_59_357 ();
 DECAPx2_ASAP7_75t_R FILLER_0_59_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_371 ();
 DECAPx1_ASAP7_75t_R FILLER_0_59_379 ();
 DECAPx2_ASAP7_75t_R FILLER_0_59_407 ();
 DECAPx1_ASAP7_75t_R FILLER_0_59_420 ();
 DECAPx2_ASAP7_75t_R FILLER_0_59_430 ();
 FILLER_ASAP7_75t_R FILLER_0_59_442 ();
 DECAPx1_ASAP7_75t_R FILLER_0_59_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_456 ();
 FILLER_ASAP7_75t_R FILLER_0_59_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_491 ();
 FILLER_ASAP7_75t_R FILLER_0_59_495 ();
 FILLER_ASAP7_75t_R FILLER_0_59_507 ();
 DECAPx2_ASAP7_75t_R FILLER_0_59_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_523 ();
 DECAPx2_ASAP7_75t_R FILLER_0_59_530 ();
 FILLER_ASAP7_75t_R FILLER_0_59_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_582 ();
 FILLER_ASAP7_75t_R FILLER_0_59_591 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_601 ();
 DECAPx2_ASAP7_75t_R FILLER_0_59_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_629 ();
 DECAPx4_ASAP7_75t_R FILLER_0_59_651 ();
 DECAPx6_ASAP7_75t_R FILLER_0_59_667 ();
 FILLER_ASAP7_75t_R FILLER_0_59_681 ();
 DECAPx4_ASAP7_75t_R FILLER_0_59_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_700 ();
 DECAPx4_ASAP7_75t_R FILLER_0_59_707 ();
 FILLER_ASAP7_75t_R FILLER_0_59_717 ();
 FILLER_ASAP7_75t_R FILLER_0_59_722 ();
 DECAPx6_ASAP7_75t_R FILLER_0_59_735 ();
 FILLER_ASAP7_75t_R FILLER_0_59_749 ();
 FILLER_ASAP7_75t_R FILLER_0_59_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_773 ();
 FILLER_ASAP7_75t_R FILLER_0_59_780 ();
 DECAPx2_ASAP7_75t_R FILLER_0_59_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_794 ();
 DECAPx6_ASAP7_75t_R FILLER_0_59_798 ();
 FILLER_ASAP7_75t_R FILLER_0_59_812 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_821 ();
 DECAPx1_ASAP7_75t_R FILLER_0_59_843 ();
 FILLER_ASAP7_75t_R FILLER_0_59_853 ();
 FILLER_ASAP7_75t_R FILLER_0_59_861 ();
 DECAPx1_ASAP7_75t_R FILLER_0_59_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_877 ();
 DECAPx4_ASAP7_75t_R FILLER_0_59_881 ();
 FILLER_ASAP7_75t_R FILLER_0_59_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_893 ();
 FILLER_ASAP7_75t_R FILLER_0_59_899 ();
 FILLER_ASAP7_75t_R FILLER_0_59_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_924 ();
 FILLER_ASAP7_75t_R FILLER_0_59_927 ();
 DECAPx4_ASAP7_75t_R FILLER_0_59_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_942 ();
 DECAPx4_ASAP7_75t_R FILLER_0_59_971 ();
 FILLER_ASAP7_75t_R FILLER_0_59_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_983 ();
 FILLER_ASAP7_75t_R FILLER_0_59_990 ();
 DECAPx1_ASAP7_75t_R FILLER_0_59_998 ();
 DECAPx1_ASAP7_75t_R FILLER_0_59_1012 ();
 DECAPx2_ASAP7_75t_R FILLER_0_59_1020 ();
 DECAPx2_ASAP7_75t_R FILLER_0_59_1032 ();
 FILLER_ASAP7_75t_R FILLER_0_59_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_1050 ();
 FILLER_ASAP7_75t_R FILLER_0_59_1061 ();
 DECAPx1_ASAP7_75t_R FILLER_0_59_1068 ();
 DECAPx1_ASAP7_75t_R FILLER_0_59_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_0_59_1098 ();
 FILLER_ASAP7_75t_R FILLER_0_59_1114 ();
 FILLER_ASAP7_75t_R FILLER_0_59_1121 ();
 DECAPx1_ASAP7_75t_R FILLER_0_59_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_1137 ();
 DECAPx6_ASAP7_75t_R FILLER_0_59_1148 ();
 DECAPx1_ASAP7_75t_R FILLER_0_59_1162 ();
 DECAPx4_ASAP7_75t_R FILLER_0_59_1172 ();
 FILLER_ASAP7_75t_R FILLER_0_59_1182 ();
 FILLER_ASAP7_75t_R FILLER_0_59_1189 ();
 FILLER_ASAP7_75t_R FILLER_0_59_1197 ();
 DECAPx2_ASAP7_75t_R FILLER_0_59_1209 ();
 FILLER_ASAP7_75t_R FILLER_0_59_1215 ();
 FILLER_ASAP7_75t_R FILLER_0_59_1227 ();
 FILLER_ASAP7_75t_R FILLER_0_59_1247 ();
 FILLER_ASAP7_75t_R FILLER_0_59_1260 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_1262 ();
 FILLER_ASAP7_75t_R FILLER_0_59_1273 ();
 FILLER_ASAP7_75t_R FILLER_0_59_1283 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_1285 ();
 FILLER_ASAP7_75t_R FILLER_0_59_1294 ();
 FILLER_ASAP7_75t_R FILLER_0_59_1310 ();
 FILLER_ASAP7_75t_R FILLER_0_59_1322 ();
 FILLER_ASAP7_75t_R FILLER_0_59_1330 ();
 FILLER_ASAP7_75t_R FILLER_0_59_1338 ();
 DECAPx1_ASAP7_75t_R FILLER_0_59_1346 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_1350 ();
 FILLER_ASAP7_75t_R FILLER_0_59_1358 ();
 FILLER_ASAP7_75t_R FILLER_0_59_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_24 ();
 DECAPx4_ASAP7_75t_R FILLER_0_60_46 ();
 DECAPx2_ASAP7_75t_R FILLER_0_60_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_68 ();
 FILLER_ASAP7_75t_R FILLER_0_60_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_91 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_96 ();
 DECAPx6_ASAP7_75t_R FILLER_0_60_124 ();
 FILLER_ASAP7_75t_R FILLER_0_60_138 ();
 DECAPx4_ASAP7_75t_R FILLER_0_60_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_156 ();
 FILLER_ASAP7_75t_R FILLER_0_60_168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_180 ();
 DECAPx6_ASAP7_75t_R FILLER_0_60_202 ();
 DECAPx1_ASAP7_75t_R FILLER_0_60_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_220 ();
 DECAPx1_ASAP7_75t_R FILLER_0_60_227 ();
 DECAPx6_ASAP7_75t_R FILLER_0_60_237 ();
 DECAPx2_ASAP7_75t_R FILLER_0_60_251 ();
 FILLER_ASAP7_75t_R FILLER_0_60_263 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_271 ();
 DECAPx4_ASAP7_75t_R FILLER_0_60_293 ();
 FILLER_ASAP7_75t_R FILLER_0_60_303 ();
 DECAPx1_ASAP7_75t_R FILLER_0_60_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_315 ();
 DECAPx6_ASAP7_75t_R FILLER_0_60_322 ();
 DECAPx2_ASAP7_75t_R FILLER_0_60_336 ();
 DECAPx2_ASAP7_75t_R FILLER_0_60_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_355 ();
 DECAPx2_ASAP7_75t_R FILLER_0_60_362 ();
 FILLER_ASAP7_75t_R FILLER_0_60_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_370 ();
 DECAPx6_ASAP7_75t_R FILLER_0_60_378 ();
 FILLER_ASAP7_75t_R FILLER_0_60_392 ();
 DECAPx1_ASAP7_75t_R FILLER_0_60_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_411 ();
 DECAPx1_ASAP7_75t_R FILLER_0_60_433 ();
 FILLER_ASAP7_75t_R FILLER_0_60_440 ();
 DECAPx6_ASAP7_75t_R FILLER_0_60_448 ();
 FILLER_ASAP7_75t_R FILLER_0_60_464 ();
 FILLER_ASAP7_75t_R FILLER_0_60_472 ();
 DECAPx4_ASAP7_75t_R FILLER_0_60_484 ();
 FILLER_ASAP7_75t_R FILLER_0_60_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_496 ();
 FILLER_ASAP7_75t_R FILLER_0_60_505 ();
 FILLER_ASAP7_75t_R FILLER_0_60_513 ();
 FILLER_ASAP7_75t_R FILLER_0_60_523 ();
 DECAPx2_ASAP7_75t_R FILLER_0_60_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_535 ();
 FILLER_ASAP7_75t_R FILLER_0_60_543 ();
 DECAPx2_ASAP7_75t_R FILLER_0_60_548 ();
 FILLER_ASAP7_75t_R FILLER_0_60_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_563 ();
 FILLER_ASAP7_75t_R FILLER_0_60_585 ();
 FILLER_ASAP7_75t_R FILLER_0_60_595 ();
 DECAPx6_ASAP7_75t_R FILLER_0_60_603 ();
 DECAPx1_ASAP7_75t_R FILLER_0_60_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_621 ();
 DECAPx2_ASAP7_75t_R FILLER_0_60_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_631 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_635 ();
 DECAPx2_ASAP7_75t_R FILLER_0_60_657 ();
 FILLER_ASAP7_75t_R FILLER_0_60_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_698 ();
 DECAPx4_ASAP7_75t_R FILLER_0_60_720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_736 ();
 DECAPx6_ASAP7_75t_R FILLER_0_60_758 ();
 FILLER_ASAP7_75t_R FILLER_0_60_772 ();
 FILLER_ASAP7_75t_R FILLER_0_60_777 ();
 DECAPx4_ASAP7_75t_R FILLER_0_60_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_800 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_807 ();
 DECAPx2_ASAP7_75t_R FILLER_0_60_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_835 ();
 FILLER_ASAP7_75t_R FILLER_0_60_842 ();
 DECAPx2_ASAP7_75t_R FILLER_0_60_855 ();
 FILLER_ASAP7_75t_R FILLER_0_60_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_863 ();
 DECAPx6_ASAP7_75t_R FILLER_0_60_870 ();
 DECAPx2_ASAP7_75t_R FILLER_0_60_884 ();
 FILLER_ASAP7_75t_R FILLER_0_60_895 ();
 FILLER_ASAP7_75t_R FILLER_0_60_911 ();
 FILLER_ASAP7_75t_R FILLER_0_60_919 ();
 FILLER_ASAP7_75t_R FILLER_0_60_927 ();
 DECAPx1_ASAP7_75t_R FILLER_0_60_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_939 ();
 FILLER_ASAP7_75t_R FILLER_0_60_943 ();
 FILLER_ASAP7_75t_R FILLER_0_60_950 ();
 DECAPx6_ASAP7_75t_R FILLER_0_60_973 ();
 DECAPx2_ASAP7_75t_R FILLER_0_60_987 ();
 DECAPx1_ASAP7_75t_R FILLER_0_60_999 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_1003 ();
 DECAPx1_ASAP7_75t_R FILLER_0_60_1012 ();
 DECAPx1_ASAP7_75t_R FILLER_0_60_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_1030 ();
 FILLER_ASAP7_75t_R FILLER_0_60_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_1040 ();
 FILLER_ASAP7_75t_R FILLER_0_60_1046 ();
 DECAPx2_ASAP7_75t_R FILLER_0_60_1058 ();
 DECAPx1_ASAP7_75t_R FILLER_0_60_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_1078 ();
 FILLER_ASAP7_75t_R FILLER_0_60_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_1105 ();
 DECAPx6_ASAP7_75t_R FILLER_0_60_1117 ();
 DECAPx2_ASAP7_75t_R FILLER_0_60_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_1137 ();
 DECAPx4_ASAP7_75t_R FILLER_0_60_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_1158 ();
 DECAPx4_ASAP7_75t_R FILLER_0_60_1165 ();
 FILLER_ASAP7_75t_R FILLER_0_60_1183 ();
 FILLER_ASAP7_75t_R FILLER_0_60_1191 ();
 FILLER_ASAP7_75t_R FILLER_0_60_1198 ();
 DECAPx1_ASAP7_75t_R FILLER_0_60_1206 ();
 FILLER_ASAP7_75t_R FILLER_0_60_1220 ();
 FILLER_ASAP7_75t_R FILLER_0_60_1232 ();
 FILLER_ASAP7_75t_R FILLER_0_60_1244 ();
 DECAPx1_ASAP7_75t_R FILLER_0_60_1254 ();
 FILLER_ASAP7_75t_R FILLER_0_60_1268 ();
 DECAPx2_ASAP7_75t_R FILLER_0_60_1280 ();
 FILLER_ASAP7_75t_R FILLER_0_60_1294 ();
 FILLER_ASAP7_75t_R FILLER_0_60_1306 ();
 FILLER_ASAP7_75t_R FILLER_0_60_1314 ();
 FILLER_ASAP7_75t_R FILLER_0_60_1322 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_1324 ();
 FILLER_ASAP7_75t_R FILLER_0_60_1333 ();
 FILLER_ASAP7_75t_R FILLER_0_60_1346 ();
 DECAPx2_ASAP7_75t_R FILLER_0_60_1353 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_1359 ();
 FILLER_ASAP7_75t_R FILLER_0_60_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_24 ();
 DECAPx2_ASAP7_75t_R FILLER_0_61_46 ();
 FILLER_ASAP7_75t_R FILLER_0_61_52 ();
 DECAPx1_ASAP7_75t_R FILLER_0_61_65 ();
 DECAPx6_ASAP7_75t_R FILLER_0_61_79 ();
 FILLER_ASAP7_75t_R FILLER_0_61_113 ();
 FILLER_ASAP7_75t_R FILLER_0_61_126 ();
 DECAPx1_ASAP7_75t_R FILLER_0_61_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_138 ();
 DECAPx6_ASAP7_75t_R FILLER_0_61_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_156 ();
 FILLER_ASAP7_75t_R FILLER_0_61_163 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_169 ();
 FILLER_ASAP7_75t_R FILLER_0_61_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_193 ();
 DECAPx4_ASAP7_75t_R FILLER_0_61_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_207 ();
 DECAPx4_ASAP7_75t_R FILLER_0_61_214 ();
 FILLER_ASAP7_75t_R FILLER_0_61_224 ();
 FILLER_ASAP7_75t_R FILLER_0_61_232 ();
 FILLER_ASAP7_75t_R FILLER_0_61_237 ();
 FILLER_ASAP7_75t_R FILLER_0_61_245 ();
 DECAPx1_ASAP7_75t_R FILLER_0_61_253 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_260 ();
 FILLER_ASAP7_75t_R FILLER_0_61_288 ();
 FILLER_ASAP7_75t_R FILLER_0_61_298 ();
 DECAPx1_ASAP7_75t_R FILLER_0_61_306 ();
 FILLER_ASAP7_75t_R FILLER_0_61_317 ();
 FILLER_ASAP7_75t_R FILLER_0_61_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_324 ();
 DECAPx4_ASAP7_75t_R FILLER_0_61_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_341 ();
 DECAPx4_ASAP7_75t_R FILLER_0_61_348 ();
 DECAPx2_ASAP7_75t_R FILLER_0_61_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_372 ();
 FILLER_ASAP7_75t_R FILLER_0_61_376 ();
 DECAPx4_ASAP7_75t_R FILLER_0_61_381 ();
 FILLER_ASAP7_75t_R FILLER_0_61_391 ();
 FILLER_ASAP7_75t_R FILLER_0_61_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_401 ();
 FILLER_ASAP7_75t_R FILLER_0_61_408 ();
 DECAPx6_ASAP7_75t_R FILLER_0_61_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_432 ();
 FILLER_ASAP7_75t_R FILLER_0_61_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_441 ();
 DECAPx4_ASAP7_75t_R FILLER_0_61_445 ();
 FILLER_ASAP7_75t_R FILLER_0_61_455 ();
 FILLER_ASAP7_75t_R FILLER_0_61_463 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_471 ();
 DECAPx4_ASAP7_75t_R FILLER_0_61_493 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_511 ();
 DECAPx1_ASAP7_75t_R FILLER_0_61_533 ();
 DECAPx1_ASAP7_75t_R FILLER_0_61_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_551 ();
 FILLER_ASAP7_75t_R FILLER_0_61_555 ();
 FILLER_ASAP7_75t_R FILLER_0_61_563 ();
 FILLER_ASAP7_75t_R FILLER_0_61_571 ();
 DECAPx6_ASAP7_75t_R FILLER_0_61_583 ();
 FILLER_ASAP7_75t_R FILLER_0_61_607 ();
 DECAPx1_ASAP7_75t_R FILLER_0_61_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_619 ();
 DECAPx6_ASAP7_75t_R FILLER_0_61_628 ();
 DECAPx1_ASAP7_75t_R FILLER_0_61_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_646 ();
 DECAPx2_ASAP7_75t_R FILLER_0_61_659 ();
 FILLER_ASAP7_75t_R FILLER_0_61_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_670 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_679 ();
 DECAPx2_ASAP7_75t_R FILLER_0_61_701 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_713 ();
 DECAPx6_ASAP7_75t_R FILLER_0_61_735 ();
 DECAPx2_ASAP7_75t_R FILLER_0_61_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_755 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_766 ();
 DECAPx2_ASAP7_75t_R FILLER_0_61_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_794 ();
 FILLER_ASAP7_75t_R FILLER_0_61_800 ();
 FILLER_ASAP7_75t_R FILLER_0_61_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_815 ();
 FILLER_ASAP7_75t_R FILLER_0_61_822 ();
 DECAPx4_ASAP7_75t_R FILLER_0_61_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_837 ();
 DECAPx2_ASAP7_75t_R FILLER_0_61_844 ();
 FILLER_ASAP7_75t_R FILLER_0_61_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_856 ();
 DECAPx6_ASAP7_75t_R FILLER_0_61_878 ();
 FILLER_ASAP7_75t_R FILLER_0_61_892 ();
 FILLER_ASAP7_75t_R FILLER_0_61_897 ();
 DECAPx1_ASAP7_75t_R FILLER_0_61_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_924 ();
 DECAPx4_ASAP7_75t_R FILLER_0_61_927 ();
 FILLER_ASAP7_75t_R FILLER_0_61_937 ();
 FILLER_ASAP7_75t_R FILLER_0_61_977 ();
 FILLER_ASAP7_75t_R FILLER_0_61_991 ();
 FILLER_ASAP7_75t_R FILLER_0_61_999 ();
 DECAPx1_ASAP7_75t_R FILLER_0_61_1013 ();
 FILLER_ASAP7_75t_R FILLER_0_61_1022 ();
 FILLER_ASAP7_75t_R FILLER_0_61_1029 ();
 FILLER_ASAP7_75t_R FILLER_0_61_1036 ();
 FILLER_ASAP7_75t_R FILLER_0_61_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_1050 ();
 FILLER_ASAP7_75t_R FILLER_0_61_1061 ();
 FILLER_ASAP7_75t_R FILLER_0_61_1073 ();
 DECAPx1_ASAP7_75t_R FILLER_0_61_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_1091 ();
 FILLER_ASAP7_75t_R FILLER_0_61_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_1106 ();
 DECAPx1_ASAP7_75t_R FILLER_0_61_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_1119 ();
 DECAPx1_ASAP7_75t_R FILLER_0_61_1142 ();
 FILLER_ASAP7_75t_R FILLER_0_61_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_61_1197 ();
 FILLER_ASAP7_75t_R FILLER_0_61_1205 ();
 FILLER_ASAP7_75t_R FILLER_0_61_1213 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_1215 ();
 DECAPx2_ASAP7_75t_R FILLER_0_61_1226 ();
 FILLER_ASAP7_75t_R FILLER_0_61_1242 ();
 FILLER_ASAP7_75t_R FILLER_0_61_1254 ();
 FILLER_ASAP7_75t_R FILLER_0_61_1266 ();
 FILLER_ASAP7_75t_R FILLER_0_61_1278 ();
 FILLER_ASAP7_75t_R FILLER_0_61_1290 ();
 FILLER_ASAP7_75t_R FILLER_0_61_1298 ();
 DECAPx1_ASAP7_75t_R FILLER_0_61_1310 ();
 FILLER_ASAP7_75t_R FILLER_0_61_1324 ();
 FILLER_ASAP7_75t_R FILLER_0_61_1332 ();
 FILLER_ASAP7_75t_R FILLER_0_61_1340 ();
 DECAPx1_ASAP7_75t_R FILLER_0_61_1348 ();
 FILLER_ASAP7_75t_R FILLER_0_61_1358 ();
 FILLER_ASAP7_75t_R FILLER_0_61_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_61_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_62_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_9 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_53 ();
 FILLER_ASAP7_75t_R FILLER_0_62_59 ();
 DECAPx4_ASAP7_75t_R FILLER_0_62_81 ();
 FILLER_ASAP7_75t_R FILLER_0_62_91 ();
 DECAPx6_ASAP7_75t_R FILLER_0_62_96 ();
 FILLER_ASAP7_75t_R FILLER_0_62_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_112 ();
 DECAPx6_ASAP7_75t_R FILLER_0_62_116 ();
 FILLER_ASAP7_75t_R FILLER_0_62_130 ();
 DECAPx6_ASAP7_75t_R FILLER_0_62_138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_62_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_158 ();
 FILLER_ASAP7_75t_R FILLER_0_62_165 ();
 DECAPx2_ASAP7_75t_R FILLER_0_62_173 ();
 FILLER_ASAP7_75t_R FILLER_0_62_185 ();
 FILLER_ASAP7_75t_R FILLER_0_62_193 ();
 DECAPx4_ASAP7_75t_R FILLER_0_62_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_208 ();
 DECAPx6_ASAP7_75t_R FILLER_0_62_212 ();
 DECAPx2_ASAP7_75t_R FILLER_0_62_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_232 ();
 FILLER_ASAP7_75t_R FILLER_0_62_253 ();
 DECAPx4_ASAP7_75t_R FILLER_0_62_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_275 ();
 DECAPx2_ASAP7_75t_R FILLER_0_62_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_289 ();
 FILLER_ASAP7_75t_R FILLER_0_62_296 ();
 FILLER_ASAP7_75t_R FILLER_0_62_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_306 ();
 DECAPx6_ASAP7_75t_R FILLER_0_62_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_328 ();
 DECAPx2_ASAP7_75t_R FILLER_0_62_335 ();
 FILLER_ASAP7_75t_R FILLER_0_62_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_343 ();
 DECAPx2_ASAP7_75t_R FILLER_0_62_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_353 ();
 DECAPx4_ASAP7_75t_R FILLER_0_62_360 ();
 FILLER_ASAP7_75t_R FILLER_0_62_370 ();
 DECAPx4_ASAP7_75t_R FILLER_0_62_378 ();
 FILLER_ASAP7_75t_R FILLER_0_62_395 ();
 DECAPx2_ASAP7_75t_R FILLER_0_62_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_409 ();
 DECAPx1_ASAP7_75t_R FILLER_0_62_416 ();
 DECAPx1_ASAP7_75t_R FILLER_0_62_426 ();
 FILLER_ASAP7_75t_R FILLER_0_62_436 ();
 FILLER_ASAP7_75t_R FILLER_0_62_444 ();
 DECAPx2_ASAP7_75t_R FILLER_0_62_454 ();
 FILLER_ASAP7_75t_R FILLER_0_62_460 ();
 DECAPx6_ASAP7_75t_R FILLER_0_62_464 ();
 DECAPx1_ASAP7_75t_R FILLER_0_62_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_482 ();
 DECAPx4_ASAP7_75t_R FILLER_0_62_493 ();
 FILLER_ASAP7_75t_R FILLER_0_62_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_505 ();
 DECAPx2_ASAP7_75t_R FILLER_0_62_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_518 ();
 DECAPx4_ASAP7_75t_R FILLER_0_62_540 ();
 FILLER_ASAP7_75t_R FILLER_0_62_550 ();
 DECAPx2_ASAP7_75t_R FILLER_0_62_564 ();
 FILLER_ASAP7_75t_R FILLER_0_62_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_572 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_581 ();
 FILLER_ASAP7_75t_R FILLER_0_62_625 ();
 DECAPx4_ASAP7_75t_R FILLER_0_62_630 ();
 DECAPx1_ASAP7_75t_R FILLER_0_62_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_652 ();
 FILLER_ASAP7_75t_R FILLER_0_62_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_667 ();
 DECAPx1_ASAP7_75t_R FILLER_0_62_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_693 ();
 FILLER_ASAP7_75t_R FILLER_0_62_700 ();
 DECAPx2_ASAP7_75t_R FILLER_0_62_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_714 ();
 DECAPx2_ASAP7_75t_R FILLER_0_62_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_727 ();
 DECAPx1_ASAP7_75t_R FILLER_0_62_731 ();
 FILLER_ASAP7_75t_R FILLER_0_62_746 ();
 DECAPx2_ASAP7_75t_R FILLER_0_62_754 ();
 FILLER_ASAP7_75t_R FILLER_0_62_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_762 ();
 FILLER_ASAP7_75t_R FILLER_0_62_772 ();
 FILLER_ASAP7_75t_R FILLER_0_62_780 ();
 DECAPx1_ASAP7_75t_R FILLER_0_62_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_792 ();
 FILLER_ASAP7_75t_R FILLER_0_62_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_801 ();
 DECAPx6_ASAP7_75t_R FILLER_0_62_808 ();
 DECAPx1_ASAP7_75t_R FILLER_0_62_822 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_837 ();
 DECAPx1_ASAP7_75t_R FILLER_0_62_859 ();
 DECAPx2_ASAP7_75t_R FILLER_0_62_869 ();
 FILLER_ASAP7_75t_R FILLER_0_62_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_877 ();
 DECAPx2_ASAP7_75t_R FILLER_0_62_885 ();
 FILLER_ASAP7_75t_R FILLER_0_62_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_893 ();
 FILLER_ASAP7_75t_R FILLER_0_62_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_902 ();
 FILLER_ASAP7_75t_R FILLER_0_62_909 ();
 DECAPx6_ASAP7_75t_R FILLER_0_62_914 ();
 DECAPx2_ASAP7_75t_R FILLER_0_62_928 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_934 ();
 FILLER_ASAP7_75t_R FILLER_0_62_945 ();
 FILLER_ASAP7_75t_R FILLER_0_62_957 ();
 FILLER_ASAP7_75t_R FILLER_0_62_971 ();
 FILLER_ASAP7_75t_R FILLER_0_62_983 ();
 FILLER_ASAP7_75t_R FILLER_0_62_991 ();
 FILLER_ASAP7_75t_R FILLER_0_62_997 ();
 DECAPx1_ASAP7_75t_R FILLER_0_62_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_1013 ();
 DECAPx1_ASAP7_75t_R FILLER_0_62_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_1028 ();
 FILLER_ASAP7_75t_R FILLER_0_62_1037 ();
 FILLER_ASAP7_75t_R FILLER_0_62_1049 ();
 FILLER_ASAP7_75t_R FILLER_0_62_1061 ();
 FILLER_ASAP7_75t_R FILLER_0_62_1069 ();
 FILLER_ASAP7_75t_R FILLER_0_62_1077 ();
 FILLER_ASAP7_75t_R FILLER_0_62_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_1089 ();
 DECAPx2_ASAP7_75t_R FILLER_0_62_1100 ();
 DECAPx2_ASAP7_75t_R FILLER_0_62_1113 ();
 FILLER_ASAP7_75t_R FILLER_0_62_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_1121 ();
 DECAPx1_ASAP7_75t_R FILLER_0_62_1125 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_1129 ();
 DECAPx1_ASAP7_75t_R FILLER_0_62_1137 ();
 FILLER_ASAP7_75t_R FILLER_0_62_1155 ();
 FILLER_ASAP7_75t_R FILLER_0_62_1162 ();
 FILLER_ASAP7_75t_R FILLER_0_62_1182 ();
 FILLER_ASAP7_75t_R FILLER_0_62_1189 ();
 FILLER_ASAP7_75t_R FILLER_0_62_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_1201 ();
 FILLER_ASAP7_75t_R FILLER_0_62_1212 ();
 DECAPx1_ASAP7_75t_R FILLER_0_62_1224 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_1228 ();
 FILLER_ASAP7_75t_R FILLER_0_62_1239 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_1241 ();
 DECAPx1_ASAP7_75t_R FILLER_0_62_1252 ();
 FILLER_ASAP7_75t_R FILLER_0_62_1266 ();
 FILLER_ASAP7_75t_R FILLER_0_62_1278 ();
 DECAPx1_ASAP7_75t_R FILLER_0_62_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_1292 ();
 FILLER_ASAP7_75t_R FILLER_0_62_1303 ();
 FILLER_ASAP7_75t_R FILLER_0_62_1313 ();
 FILLER_ASAP7_75t_R FILLER_0_62_1320 ();
 FILLER_ASAP7_75t_R FILLER_0_62_1332 ();
 FILLER_ASAP7_75t_R FILLER_0_62_1340 ();
 DECAPx2_ASAP7_75t_R FILLER_0_62_1348 ();
 FILLER_ASAP7_75t_R FILLER_0_62_1360 ();
 FILLER_ASAP7_75t_R FILLER_0_62_1368 ();
 DECAPx2_ASAP7_75t_R FILLER_0_62_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_1381 ();
 DECAPx2_ASAP7_75t_R FILLER_0_63_2 ();
 FILLER_ASAP7_75t_R FILLER_0_63_13 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_20 ();
 DECAPx4_ASAP7_75t_R FILLER_0_63_42 ();
 FILLER_ASAP7_75t_R FILLER_0_63_52 ();
 FILLER_ASAP7_75t_R FILLER_0_63_57 ();
 DECAPx1_ASAP7_75t_R FILLER_0_63_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_69 ();
 FILLER_ASAP7_75t_R FILLER_0_63_76 ();
 DECAPx2_ASAP7_75t_R FILLER_0_63_81 ();
 FILLER_ASAP7_75t_R FILLER_0_63_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_89 ();
 FILLER_ASAP7_75t_R FILLER_0_63_96 ();
 DECAPx4_ASAP7_75t_R FILLER_0_63_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_111 ();
 DECAPx4_ASAP7_75t_R FILLER_0_63_118 ();
 FILLER_ASAP7_75t_R FILLER_0_63_131 ();
 DECAPx6_ASAP7_75t_R FILLER_0_63_139 ();
 FILLER_ASAP7_75t_R FILLER_0_63_153 ();
 FILLER_ASAP7_75t_R FILLER_0_63_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_167 ();
 FILLER_ASAP7_75t_R FILLER_0_63_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_180 ();
 FILLER_ASAP7_75t_R FILLER_0_63_191 ();
 FILLER_ASAP7_75t_R FILLER_0_63_199 ();
 FILLER_ASAP7_75t_R FILLER_0_63_207 ();
 FILLER_ASAP7_75t_R FILLER_0_63_215 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_220 ();
 FILLER_ASAP7_75t_R FILLER_0_63_242 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_249 ();
 DECAPx4_ASAP7_75t_R FILLER_0_63_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_281 ();
 FILLER_ASAP7_75t_R FILLER_0_63_288 ();
 DECAPx2_ASAP7_75t_R FILLER_0_63_295 ();
 FILLER_ASAP7_75t_R FILLER_0_63_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_303 ();
 DECAPx1_ASAP7_75t_R FILLER_0_63_310 ();
 DECAPx4_ASAP7_75t_R FILLER_0_63_320 ();
 FILLER_ASAP7_75t_R FILLER_0_63_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_332 ();
 FILLER_ASAP7_75t_R FILLER_0_63_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_342 ();
 DECAPx1_ASAP7_75t_R FILLER_0_63_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_353 ();
 DECAPx4_ASAP7_75t_R FILLER_0_63_362 ();
 FILLER_ASAP7_75t_R FILLER_0_63_372 ();
 DECAPx1_ASAP7_75t_R FILLER_0_63_377 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_387 ();
 FILLER_ASAP7_75t_R FILLER_0_63_417 ();
 DECAPx2_ASAP7_75t_R FILLER_0_63_427 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_440 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_468 ();
 DECAPx1_ASAP7_75t_R FILLER_0_63_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_494 ();
 DECAPx1_ASAP7_75t_R FILLER_0_63_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_520 ();
 DECAPx2_ASAP7_75t_R FILLER_0_63_527 ();
 FILLER_ASAP7_75t_R FILLER_0_63_554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_568 ();
 FILLER_ASAP7_75t_R FILLER_0_63_590 ();
 FILLER_ASAP7_75t_R FILLER_0_63_598 ();
 FILLER_ASAP7_75t_R FILLER_0_63_608 ();
 DECAPx4_ASAP7_75t_R FILLER_0_63_613 ();
 FILLER_ASAP7_75t_R FILLER_0_63_634 ();
 FILLER_ASAP7_75t_R FILLER_0_63_642 ();
 DECAPx1_ASAP7_75t_R FILLER_0_63_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_654 ();
 FILLER_ASAP7_75t_R FILLER_0_63_667 ();
 FILLER_ASAP7_75t_R FILLER_0_63_672 ();
 DECAPx2_ASAP7_75t_R FILLER_0_63_684 ();
 FILLER_ASAP7_75t_R FILLER_0_63_696 ();
 FILLER_ASAP7_75t_R FILLER_0_63_708 ();
 DECAPx1_ASAP7_75t_R FILLER_0_63_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_725 ();
 FILLER_ASAP7_75t_R FILLER_0_63_732 ();
 DECAPx2_ASAP7_75t_R FILLER_0_63_739 ();
 FILLER_ASAP7_75t_R FILLER_0_63_745 ();
 FILLER_ASAP7_75t_R FILLER_0_63_753 ();
 DECAPx1_ASAP7_75t_R FILLER_0_63_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_767 ();
 FILLER_ASAP7_75t_R FILLER_0_63_774 ();
 FILLER_ASAP7_75t_R FILLER_0_63_784 ();
 FILLER_ASAP7_75t_R FILLER_0_63_792 ();
 FILLER_ASAP7_75t_R FILLER_0_63_800 ();
 FILLER_ASAP7_75t_R FILLER_0_63_808 ();
 DECAPx2_ASAP7_75t_R FILLER_0_63_815 ();
 FILLER_ASAP7_75t_R FILLER_0_63_821 ();
 FILLER_ASAP7_75t_R FILLER_0_63_829 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_837 ();
 DECAPx1_ASAP7_75t_R FILLER_0_63_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_863 ();
 FILLER_ASAP7_75t_R FILLER_0_63_870 ();
 FILLER_ASAP7_75t_R FILLER_0_63_878 ();
 FILLER_ASAP7_75t_R FILLER_0_63_886 ();
 FILLER_ASAP7_75t_R FILLER_0_63_891 ();
 FILLER_ASAP7_75t_R FILLER_0_63_899 ();
 DECAPx6_ASAP7_75t_R FILLER_0_63_908 ();
 FILLER_ASAP7_75t_R FILLER_0_63_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_924 ();
 DECAPx2_ASAP7_75t_R FILLER_0_63_927 ();
 DECAPx1_ASAP7_75t_R FILLER_0_63_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_947 ();
 FILLER_ASAP7_75t_R FILLER_0_63_953 ();
 FILLER_ASAP7_75t_R FILLER_0_63_973 ();
 DECAPx1_ASAP7_75t_R FILLER_0_63_987 ();
 FILLER_ASAP7_75t_R FILLER_0_63_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_999 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1010 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1025 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1037 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1049 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1061 ();
 DECAPx1_ASAP7_75t_R FILLER_0_63_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_1087 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1096 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1104 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1112 ();
 DECAPx2_ASAP7_75t_R FILLER_0_63_1119 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_1147 ();
 DECAPx1_ASAP7_75t_R FILLER_0_63_1160 ();
 DECAPx1_ASAP7_75t_R FILLER_0_63_1170 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1180 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1188 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1196 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_1206 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1217 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1229 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1237 ();
 DECAPx1_ASAP7_75t_R FILLER_0_63_1245 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1255 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1267 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1279 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1291 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1303 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1315 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1325 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1333 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1341 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1349 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1364 ();
 FILLER_ASAP7_75t_R FILLER_0_63_1371 ();
 DECAPx1_ASAP7_75t_R FILLER_0_63_1378 ();
 FILLER_ASAP7_75t_R FILLER_0_64_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_4 ();
 DECAPx2_ASAP7_75t_R FILLER_0_64_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_46 ();
 DECAPx2_ASAP7_75t_R FILLER_0_64_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_74 ();
 FILLER_ASAP7_75t_R FILLER_0_64_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_87 ();
 DECAPx1_ASAP7_75t_R FILLER_0_64_94 ();
 FILLER_ASAP7_75t_R FILLER_0_64_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_106 ();
 DECAPx1_ASAP7_75t_R FILLER_0_64_127 ();
 FILLER_ASAP7_75t_R FILLER_0_64_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_139 ();
 FILLER_ASAP7_75t_R FILLER_0_64_150 ();
 DECAPx2_ASAP7_75t_R FILLER_0_64_172 ();
 FILLER_ASAP7_75t_R FILLER_0_64_181 ();
 DECAPx2_ASAP7_75t_R FILLER_0_64_186 ();
 FILLER_ASAP7_75t_R FILLER_0_64_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_194 ();
 FILLER_ASAP7_75t_R FILLER_0_64_205 ();
 DECAPx6_ASAP7_75t_R FILLER_0_64_210 ();
 DECAPx1_ASAP7_75t_R FILLER_0_64_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_239 ();
 DECAPx2_ASAP7_75t_R FILLER_0_64_261 ();
 FILLER_ASAP7_75t_R FILLER_0_64_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_269 ();
 FILLER_ASAP7_75t_R FILLER_0_64_276 ();
 FILLER_ASAP7_75t_R FILLER_0_64_284 ();
 DECAPx1_ASAP7_75t_R FILLER_0_64_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_297 ();
 FILLER_ASAP7_75t_R FILLER_0_64_304 ();
 DECAPx6_ASAP7_75t_R FILLER_0_64_312 ();
 DECAPx2_ASAP7_75t_R FILLER_0_64_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_332 ();
 FILLER_ASAP7_75t_R FILLER_0_64_339 ();
 DECAPx4_ASAP7_75t_R FILLER_0_64_347 ();
 FILLER_ASAP7_75t_R FILLER_0_64_357 ();
 FILLER_ASAP7_75t_R FILLER_0_64_366 ();
 FILLER_ASAP7_75t_R FILLER_0_64_390 ();
 FILLER_ASAP7_75t_R FILLER_0_64_398 ();
 FILLER_ASAP7_75t_R FILLER_0_64_408 ();
 FILLER_ASAP7_75t_R FILLER_0_64_416 ();
 DECAPx4_ASAP7_75t_R FILLER_0_64_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_431 ();
 DECAPx2_ASAP7_75t_R FILLER_0_64_438 ();
 FILLER_ASAP7_75t_R FILLER_0_64_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_452 ();
 FILLER_ASAP7_75t_R FILLER_0_64_460 ();
 FILLER_ASAP7_75t_R FILLER_0_64_464 ();
 FILLER_ASAP7_75t_R FILLER_0_64_472 ();
 DECAPx2_ASAP7_75t_R FILLER_0_64_481 ();
 DECAPx6_ASAP7_75t_R FILLER_0_64_493 ();
 FILLER_ASAP7_75t_R FILLER_0_64_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_509 ();
 FILLER_ASAP7_75t_R FILLER_0_64_522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_527 ();
 FILLER_ASAP7_75t_R FILLER_0_64_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_551 ();
 DECAPx1_ASAP7_75t_R FILLER_0_64_555 ();
 DECAPx2_ASAP7_75t_R FILLER_0_64_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_586 ();
 FILLER_ASAP7_75t_R FILLER_0_64_595 ();
 DECAPx6_ASAP7_75t_R FILLER_0_64_605 ();
 DECAPx1_ASAP7_75t_R FILLER_0_64_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_623 ();
 DECAPx2_ASAP7_75t_R FILLER_0_64_629 ();
 FILLER_ASAP7_75t_R FILLER_0_64_635 ();
 FILLER_ASAP7_75t_R FILLER_0_64_643 ();
 FILLER_ASAP7_75t_R FILLER_0_64_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_655 ();
 FILLER_ASAP7_75t_R FILLER_0_64_667 ();
 FILLER_ASAP7_75t_R FILLER_0_64_679 ();
 FILLER_ASAP7_75t_R FILLER_0_64_691 ();
 DECAPx2_ASAP7_75t_R FILLER_0_64_699 ();
 DECAPx2_ASAP7_75t_R FILLER_0_64_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_717 ();
 FILLER_ASAP7_75t_R FILLER_0_64_726 ();
 FILLER_ASAP7_75t_R FILLER_0_64_734 ();
 DECAPx1_ASAP7_75t_R FILLER_0_64_742 ();
 FILLER_ASAP7_75t_R FILLER_0_64_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_753 ();
 FILLER_ASAP7_75t_R FILLER_0_64_760 ();
 FILLER_ASAP7_75t_R FILLER_0_64_768 ();
 FILLER_ASAP7_75t_R FILLER_0_64_778 ();
 DECAPx6_ASAP7_75t_R FILLER_0_64_785 ();
 DECAPx2_ASAP7_75t_R FILLER_0_64_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_811 ();
 DECAPx6_ASAP7_75t_R FILLER_0_64_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_832 ();
 FILLER_ASAP7_75t_R FILLER_0_64_841 ();
 FILLER_ASAP7_75t_R FILLER_0_64_849 ();
 FILLER_ASAP7_75t_R FILLER_0_64_857 ();
 DECAPx6_ASAP7_75t_R FILLER_0_64_865 ();
 DECAPx1_ASAP7_75t_R FILLER_0_64_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_883 ();
 FILLER_ASAP7_75t_R FILLER_0_64_890 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_898 ();
 DECAPx6_ASAP7_75t_R FILLER_0_64_920 ();
 DECAPx2_ASAP7_75t_R FILLER_0_64_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_940 ();
 FILLER_ASAP7_75t_R FILLER_0_64_946 ();
 FILLER_ASAP7_75t_R FILLER_0_64_953 ();
 DECAPx4_ASAP7_75t_R FILLER_0_64_967 ();
 DECAPx1_ASAP7_75t_R FILLER_0_64_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_987 ();
 DECAPx1_ASAP7_75t_R FILLER_0_64_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_1002 ();
 FILLER_ASAP7_75t_R FILLER_0_64_1013 ();
 FILLER_ASAP7_75t_R FILLER_0_64_1020 ();
 FILLER_ASAP7_75t_R FILLER_0_64_1032 ();
 FILLER_ASAP7_75t_R FILLER_0_64_1044 ();
 FILLER_ASAP7_75t_R FILLER_0_64_1056 ();
 FILLER_ASAP7_75t_R FILLER_0_64_1068 ();
 FILLER_ASAP7_75t_R FILLER_0_64_1080 ();
 FILLER_ASAP7_75t_R FILLER_0_64_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_1090 ();
 DECAPx2_ASAP7_75t_R FILLER_0_64_1101 ();
 FILLER_ASAP7_75t_R FILLER_0_64_1107 ();
 FILLER_ASAP7_75t_R FILLER_0_64_1117 ();
 DECAPx1_ASAP7_75t_R FILLER_0_64_1124 ();
 DECAPx4_ASAP7_75t_R FILLER_0_64_1134 ();
 FILLER_ASAP7_75t_R FILLER_0_64_1144 ();
 DECAPx1_ASAP7_75t_R FILLER_0_64_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_1155 ();
 DECAPx1_ASAP7_75t_R FILLER_0_64_1159 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_1163 ();
 DECAPx6_ASAP7_75t_R FILLER_0_64_1169 ();
 DECAPx1_ASAP7_75t_R FILLER_0_64_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_1187 ();
 FILLER_ASAP7_75t_R FILLER_0_64_1193 ();
 FILLER_ASAP7_75t_R FILLER_0_64_1200 ();
 FILLER_ASAP7_75t_R FILLER_0_64_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_1209 ();
 FILLER_ASAP7_75t_R FILLER_0_64_1218 ();
 FILLER_ASAP7_75t_R FILLER_0_64_1225 ();
 FILLER_ASAP7_75t_R FILLER_0_64_1233 ();
 DECAPx2_ASAP7_75t_R FILLER_0_64_1241 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_1247 ();
 FILLER_ASAP7_75t_R FILLER_0_64_1270 ();
 FILLER_ASAP7_75t_R FILLER_0_64_1282 ();
 DECAPx1_ASAP7_75t_R FILLER_0_64_1291 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_1295 ();
 FILLER_ASAP7_75t_R FILLER_0_64_1306 ();
 FILLER_ASAP7_75t_R FILLER_0_64_1311 ();
 DECAPx1_ASAP7_75t_R FILLER_0_64_1325 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_1329 ();
 DECAPx2_ASAP7_75t_R FILLER_0_64_1338 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_1344 ();
 DECAPx2_ASAP7_75t_R FILLER_0_64_1351 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_1357 ();
 DECAPx1_ASAP7_75t_R FILLER_0_64_1364 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_1368 ();
 FILLER_ASAP7_75t_R FILLER_0_64_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_1381 ();
 DECAPx1_ASAP7_75t_R FILLER_0_65_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_27 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_49 ();
 FILLER_ASAP7_75t_R FILLER_0_65_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_73 ();
 DECAPx1_ASAP7_75t_R FILLER_0_65_84 ();
 DECAPx2_ASAP7_75t_R FILLER_0_65_91 ();
 DECAPx2_ASAP7_75t_R FILLER_0_65_107 ();
 DECAPx1_ASAP7_75t_R FILLER_0_65_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_123 ();
 FILLER_ASAP7_75t_R FILLER_0_65_130 ();
 DECAPx2_ASAP7_75t_R FILLER_0_65_142 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_154 ();
 DECAPx2_ASAP7_75t_R FILLER_0_65_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_182 ();
 DECAPx4_ASAP7_75t_R FILLER_0_65_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_199 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_210 ();
 DECAPx6_ASAP7_75t_R FILLER_0_65_232 ();
 DECAPx6_ASAP7_75t_R FILLER_0_65_252 ();
 DECAPx1_ASAP7_75t_R FILLER_0_65_266 ();
 FILLER_ASAP7_75t_R FILLER_0_65_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_293 ();
 FILLER_ASAP7_75t_R FILLER_0_65_300 ();
 FILLER_ASAP7_75t_R FILLER_0_65_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_312 ();
 FILLER_ASAP7_75t_R FILLER_0_65_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_321 ();
 FILLER_ASAP7_75t_R FILLER_0_65_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_330 ();
 DECAPx1_ASAP7_75t_R FILLER_0_65_337 ();
 FILLER_ASAP7_75t_R FILLER_0_65_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_351 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_358 ();
 DECAPx6_ASAP7_75t_R FILLER_0_65_380 ();
 DECAPx1_ASAP7_75t_R FILLER_0_65_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_404 ();
 FILLER_ASAP7_75t_R FILLER_0_65_408 ();
 FILLER_ASAP7_75t_R FILLER_0_65_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_420 ();
 FILLER_ASAP7_75t_R FILLER_0_65_427 ();
 DECAPx2_ASAP7_75t_R FILLER_0_65_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_443 ();
 FILLER_ASAP7_75t_R FILLER_0_65_452 ();
 FILLER_ASAP7_75t_R FILLER_0_65_460 ();
 FILLER_ASAP7_75t_R FILLER_0_65_468 ();
 DECAPx6_ASAP7_75t_R FILLER_0_65_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_491 ();
 DECAPx6_ASAP7_75t_R FILLER_0_65_495 ();
 DECAPx1_ASAP7_75t_R FILLER_0_65_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_513 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_539 ();
 DECAPx2_ASAP7_75t_R FILLER_0_65_546 ();
 FILLER_ASAP7_75t_R FILLER_0_65_552 ();
 FILLER_ASAP7_75t_R FILLER_0_65_566 ();
 FILLER_ASAP7_75t_R FILLER_0_65_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_573 ();
 FILLER_ASAP7_75t_R FILLER_0_65_580 ();
 FILLER_ASAP7_75t_R FILLER_0_65_592 ();
 DECAPx2_ASAP7_75t_R FILLER_0_65_600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_65_612 ();
 FILLER_ASAP7_75t_R FILLER_0_65_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_628 ();
 DECAPx6_ASAP7_75t_R FILLER_0_65_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_671 ();
 DECAPx2_ASAP7_75t_R FILLER_0_65_684 ();
 FILLER_ASAP7_75t_R FILLER_0_65_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_692 ();
 DECAPx2_ASAP7_75t_R FILLER_0_65_699 ();
 FILLER_ASAP7_75t_R FILLER_0_65_705 ();
 FILLER_ASAP7_75t_R FILLER_0_65_713 ();
 FILLER_ASAP7_75t_R FILLER_0_65_720 ();
 DECAPx4_ASAP7_75t_R FILLER_0_65_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_737 ();
 DECAPx2_ASAP7_75t_R FILLER_0_65_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_750 ();
 FILLER_ASAP7_75t_R FILLER_0_65_756 ();
 DECAPx1_ASAP7_75t_R FILLER_0_65_764 ();
 FILLER_ASAP7_75t_R FILLER_0_65_774 ();
 FILLER_ASAP7_75t_R FILLER_0_65_783 ();
 DECAPx1_ASAP7_75t_R FILLER_0_65_793 ();
 FILLER_ASAP7_75t_R FILLER_0_65_803 ();
 DECAPx1_ASAP7_75t_R FILLER_0_65_811 ();
 DECAPx1_ASAP7_75t_R FILLER_0_65_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_825 ();
 FILLER_ASAP7_75t_R FILLER_0_65_833 ();
 FILLER_ASAP7_75t_R FILLER_0_65_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_843 ();
 DECAPx4_ASAP7_75t_R FILLER_0_65_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_860 ();
 FILLER_ASAP7_75t_R FILLER_0_65_867 ();
 DECAPx4_ASAP7_75t_R FILLER_0_65_875 ();
 DECAPx4_ASAP7_75t_R FILLER_0_65_891 ();
 FILLER_ASAP7_75t_R FILLER_0_65_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_903 ();
 DECAPx6_ASAP7_75t_R FILLER_0_65_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_924 ();
 DECAPx2_ASAP7_75t_R FILLER_0_65_927 ();
 FILLER_ASAP7_75t_R FILLER_0_65_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_935 ();
 FILLER_ASAP7_75t_R FILLER_0_65_946 ();
 DECAPx1_ASAP7_75t_R FILLER_0_65_958 ();
 DECAPx6_ASAP7_75t_R FILLER_0_65_965 ();
 FILLER_ASAP7_75t_R FILLER_0_65_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_981 ();
 FILLER_ASAP7_75t_R FILLER_0_65_988 ();
 FILLER_ASAP7_75t_R FILLER_0_65_996 ();
 FILLER_ASAP7_75t_R FILLER_0_65_1008 ();
 DECAPx2_ASAP7_75t_R FILLER_0_65_1020 ();
 FILLER_ASAP7_75t_R FILLER_0_65_1026 ();
 DECAPx1_ASAP7_75t_R FILLER_0_65_1038 ();
 FILLER_ASAP7_75t_R FILLER_0_65_1052 ();
 FILLER_ASAP7_75t_R FILLER_0_65_1064 ();
 FILLER_ASAP7_75t_R FILLER_0_65_1076 ();
 DECAPx1_ASAP7_75t_R FILLER_0_65_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_1092 ();
 FILLER_ASAP7_75t_R FILLER_0_65_1103 ();
 FILLER_ASAP7_75t_R FILLER_0_65_1115 ();
 FILLER_ASAP7_75t_R FILLER_0_65_1123 ();
 FILLER_ASAP7_75t_R FILLER_0_65_1133 ();
 DECAPx2_ASAP7_75t_R FILLER_0_65_1138 ();
 FILLER_ASAP7_75t_R FILLER_0_65_1154 ();
 FILLER_ASAP7_75t_R FILLER_0_65_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_1164 ();
 FILLER_ASAP7_75t_R FILLER_0_65_1171 ();
 FILLER_ASAP7_75t_R FILLER_0_65_1181 ();
 DECAPx2_ASAP7_75t_R FILLER_0_65_1189 ();
 FILLER_ASAP7_75t_R FILLER_0_65_1195 ();
 FILLER_ASAP7_75t_R FILLER_0_65_1207 ();
 FILLER_ASAP7_75t_R FILLER_0_65_1213 ();
 FILLER_ASAP7_75t_R FILLER_0_65_1225 ();
 DECAPx1_ASAP7_75t_R FILLER_0_65_1237 ();
 DECAPx1_ASAP7_75t_R FILLER_0_65_1251 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_1255 ();
 DECAPx2_ASAP7_75t_R FILLER_0_65_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_1284 ();
 FILLER_ASAP7_75t_R FILLER_0_65_1297 ();
 FILLER_ASAP7_75t_R FILLER_0_65_1305 ();
 FILLER_ASAP7_75t_R FILLER_0_65_1313 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_1315 ();
 FILLER_ASAP7_75t_R FILLER_0_65_1322 ();
 FILLER_ASAP7_75t_R FILLER_0_65_1330 ();
 DECAPx2_ASAP7_75t_R FILLER_0_65_1352 ();
 FILLER_ASAP7_75t_R FILLER_0_65_1358 ();
 FILLER_ASAP7_75t_R FILLER_0_65_1380 ();
 DECAPx1_ASAP7_75t_R FILLER_0_66_2 ();
 FILLER_ASAP7_75t_R FILLER_0_66_9 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_38 ();
 DECAPx6_ASAP7_75t_R FILLER_0_66_60 ();
 DECAPx1_ASAP7_75t_R FILLER_0_66_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_78 ();
 DECAPx2_ASAP7_75t_R FILLER_0_66_82 ();
 DECAPx6_ASAP7_75t_R FILLER_0_66_98 ();
 DECAPx2_ASAP7_75t_R FILLER_0_66_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_118 ();
 DECAPx1_ASAP7_75t_R FILLER_0_66_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_133 ();
 FILLER_ASAP7_75t_R FILLER_0_66_139 ();
 FILLER_ASAP7_75t_R FILLER_0_66_151 ();
 FILLER_ASAP7_75t_R FILLER_0_66_159 ();
 DECAPx1_ASAP7_75t_R FILLER_0_66_167 ();
 DECAPx2_ASAP7_75t_R FILLER_0_66_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_183 ();
 FILLER_ASAP7_75t_R FILLER_0_66_194 ();
 FILLER_ASAP7_75t_R FILLER_0_66_217 ();
 FILLER_ASAP7_75t_R FILLER_0_66_225 ();
 FILLER_ASAP7_75t_R FILLER_0_66_237 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_260 ();
 DECAPx2_ASAP7_75t_R FILLER_0_66_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_288 ();
 DECAPx1_ASAP7_75t_R FILLER_0_66_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_296 ();
 FILLER_ASAP7_75t_R FILLER_0_66_303 ();
 FILLER_ASAP7_75t_R FILLER_0_66_311 ();
 DECAPx2_ASAP7_75t_R FILLER_0_66_320 ();
 FILLER_ASAP7_75t_R FILLER_0_66_326 ();
 DECAPx6_ASAP7_75t_R FILLER_0_66_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_349 ();
 FILLER_ASAP7_75t_R FILLER_0_66_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_360 ();
 FILLER_ASAP7_75t_R FILLER_0_66_369 ();
 DECAPx6_ASAP7_75t_R FILLER_0_66_377 ();
 DECAPx2_ASAP7_75t_R FILLER_0_66_391 ();
 FILLER_ASAP7_75t_R FILLER_0_66_421 ();
 DECAPx2_ASAP7_75t_R FILLER_0_66_426 ();
 FILLER_ASAP7_75t_R FILLER_0_66_432 ();
 DECAPx1_ASAP7_75t_R FILLER_0_66_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_444 ();
 FILLER_ASAP7_75t_R FILLER_0_66_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_453 ();
 FILLER_ASAP7_75t_R FILLER_0_66_460 ();
 DECAPx1_ASAP7_75t_R FILLER_0_66_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_475 ();
 DECAPx4_ASAP7_75t_R FILLER_0_66_497 ();
 FILLER_ASAP7_75t_R FILLER_0_66_519 ();
 DECAPx2_ASAP7_75t_R FILLER_0_66_527 ();
 FILLER_ASAP7_75t_R FILLER_0_66_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_535 ();
 DECAPx6_ASAP7_75t_R FILLER_0_66_557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_66_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_575 ();
 FILLER_ASAP7_75t_R FILLER_0_66_582 ();
 DECAPx4_ASAP7_75t_R FILLER_0_66_592 ();
 FILLER_ASAP7_75t_R FILLER_0_66_602 ();
 FILLER_ASAP7_75t_R FILLER_0_66_610 ();
 FILLER_ASAP7_75t_R FILLER_0_66_620 ();
 FILLER_ASAP7_75t_R FILLER_0_66_628 ();
 DECAPx6_ASAP7_75t_R FILLER_0_66_651 ();
 DECAPx2_ASAP7_75t_R FILLER_0_66_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_671 ();
 FILLER_ASAP7_75t_R FILLER_0_66_678 ();
 FILLER_ASAP7_75t_R FILLER_0_66_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_687 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_694 ();
 DECAPx1_ASAP7_75t_R FILLER_0_66_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_720 ();
 FILLER_ASAP7_75t_R FILLER_0_66_727 ();
 FILLER_ASAP7_75t_R FILLER_0_66_735 ();
 DECAPx4_ASAP7_75t_R FILLER_0_66_743 ();
 FILLER_ASAP7_75t_R FILLER_0_66_758 ();
 DECAPx4_ASAP7_75t_R FILLER_0_66_765 ();
 FILLER_ASAP7_75t_R FILLER_0_66_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_777 ();
 DECAPx6_ASAP7_75t_R FILLER_0_66_784 ();
 DECAPx4_ASAP7_75t_R FILLER_0_66_804 ();
 FILLER_ASAP7_75t_R FILLER_0_66_814 ();
 DECAPx2_ASAP7_75t_R FILLER_0_66_821 ();
 DECAPx2_ASAP7_75t_R FILLER_0_66_832 ();
 FILLER_ASAP7_75t_R FILLER_0_66_843 ();
 FILLER_ASAP7_75t_R FILLER_0_66_851 ();
 DECAPx4_ASAP7_75t_R FILLER_0_66_859 ();
 FILLER_ASAP7_75t_R FILLER_0_66_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_871 ();
 DECAPx4_ASAP7_75t_R FILLER_0_66_878 ();
 FILLER_ASAP7_75t_R FILLER_0_66_893 ();
 DECAPx2_ASAP7_75t_R FILLER_0_66_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_904 ();
 FILLER_ASAP7_75t_R FILLER_0_66_911 ();
 DECAPx6_ASAP7_75t_R FILLER_0_66_919 ();
 DECAPx1_ASAP7_75t_R FILLER_0_66_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_937 ();
 DECAPx1_ASAP7_75t_R FILLER_0_66_944 ();
 DECAPx2_ASAP7_75t_R FILLER_0_66_958 ();
 FILLER_ASAP7_75t_R FILLER_0_66_970 ();
 DECAPx2_ASAP7_75t_R FILLER_0_66_978 ();
 DECAPx2_ASAP7_75t_R FILLER_0_66_995 ();
 FILLER_ASAP7_75t_R FILLER_0_66_1011 ();
 DECAPx1_ASAP7_75t_R FILLER_0_66_1023 ();
 FILLER_ASAP7_75t_R FILLER_0_66_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_1039 ();
 FILLER_ASAP7_75t_R FILLER_0_66_1046 ();
 FILLER_ASAP7_75t_R FILLER_0_66_1066 ();
 FILLER_ASAP7_75t_R FILLER_0_66_1078 ();
 FILLER_ASAP7_75t_R FILLER_0_66_1088 ();
 DECAPx1_ASAP7_75t_R FILLER_0_66_1108 ();
 FILLER_ASAP7_75t_R FILLER_0_66_1119 ();
 DECAPx1_ASAP7_75t_R FILLER_0_66_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_1137 ();
 FILLER_ASAP7_75t_R FILLER_0_66_1150 ();
 DECAPx2_ASAP7_75t_R FILLER_0_66_1163 ();
 FILLER_ASAP7_75t_R FILLER_0_66_1169 ();
 FILLER_ASAP7_75t_R FILLER_0_66_1177 ();
 FILLER_ASAP7_75t_R FILLER_0_66_1185 ();
 DECAPx4_ASAP7_75t_R FILLER_0_66_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_1203 ();
 FILLER_ASAP7_75t_R FILLER_0_66_1214 ();
 DECAPx1_ASAP7_75t_R FILLER_0_66_1226 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_1230 ();
 FILLER_ASAP7_75t_R FILLER_0_66_1241 ();
 DECAPx2_ASAP7_75t_R FILLER_0_66_1253 ();
 FILLER_ASAP7_75t_R FILLER_0_66_1259 ();
 DECAPx1_ASAP7_75t_R FILLER_0_66_1267 ();
 FILLER_ASAP7_75t_R FILLER_0_66_1281 ();
 FILLER_ASAP7_75t_R FILLER_0_66_1289 ();
 FILLER_ASAP7_75t_R FILLER_0_66_1301 ();
 DECAPx1_ASAP7_75t_R FILLER_0_66_1308 ();
 FILLER_ASAP7_75t_R FILLER_0_66_1324 ();
 FILLER_ASAP7_75t_R FILLER_0_66_1334 ();
 FILLER_ASAP7_75t_R FILLER_0_66_1342 ();
 FILLER_ASAP7_75t_R FILLER_0_66_1350 ();
 FILLER_ASAP7_75t_R FILLER_0_66_1355 ();
 FILLER_ASAP7_75t_R FILLER_0_66_1362 ();
 DECAPx4_ASAP7_75t_R FILLER_0_66_1370 ();
 FILLER_ASAP7_75t_R FILLER_0_66_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_30 ();
 FILLER_ASAP7_75t_R FILLER_0_67_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_36 ();
 DECAPx6_ASAP7_75t_R FILLER_0_67_43 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_60 ();
 FILLER_ASAP7_75t_R FILLER_0_67_72 ();
 FILLER_ASAP7_75t_R FILLER_0_67_80 ();
 FILLER_ASAP7_75t_R FILLER_0_67_87 ();
 FILLER_ASAP7_75t_R FILLER_0_67_94 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_99 ();
 FILLER_ASAP7_75t_R FILLER_0_67_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_107 ();
 FILLER_ASAP7_75t_R FILLER_0_67_113 ();
 FILLER_ASAP7_75t_R FILLER_0_67_120 ();
 FILLER_ASAP7_75t_R FILLER_0_67_132 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_152 ();
 FILLER_ASAP7_75t_R FILLER_0_67_164 ();
 FILLER_ASAP7_75t_R FILLER_0_67_172 ();
 FILLER_ASAP7_75t_R FILLER_0_67_180 ();
 DECAPx4_ASAP7_75t_R FILLER_0_67_185 ();
 FILLER_ASAP7_75t_R FILLER_0_67_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_197 ();
 DECAPx4_ASAP7_75t_R FILLER_0_67_201 ();
 FILLER_ASAP7_75t_R FILLER_0_67_211 ();
 FILLER_ASAP7_75t_R FILLER_0_67_219 ();
 FILLER_ASAP7_75t_R FILLER_0_67_224 ();
 FILLER_ASAP7_75t_R FILLER_0_67_232 ();
 FILLER_ASAP7_75t_R FILLER_0_67_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_239 ();
 FILLER_ASAP7_75t_R FILLER_0_67_246 ();
 DECAPx6_ASAP7_75t_R FILLER_0_67_251 ();
 DECAPx1_ASAP7_75t_R FILLER_0_67_265 ();
 FILLER_ASAP7_75t_R FILLER_0_67_275 ();
 FILLER_ASAP7_75t_R FILLER_0_67_285 ();
 FILLER_ASAP7_75t_R FILLER_0_67_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_295 ();
 DECAPx4_ASAP7_75t_R FILLER_0_67_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_312 ();
 DECAPx4_ASAP7_75t_R FILLER_0_67_319 ();
 FILLER_ASAP7_75t_R FILLER_0_67_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_331 ();
 FILLER_ASAP7_75t_R FILLER_0_67_338 ();
 FILLER_ASAP7_75t_R FILLER_0_67_346 ();
 FILLER_ASAP7_75t_R FILLER_0_67_354 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_362 ();
 FILLER_ASAP7_75t_R FILLER_0_67_378 ();
 FILLER_ASAP7_75t_R FILLER_0_67_388 ();
 FILLER_ASAP7_75t_R FILLER_0_67_396 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_404 ();
 FILLER_ASAP7_75t_R FILLER_0_67_416 ();
 FILLER_ASAP7_75t_R FILLER_0_67_424 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_431 ();
 FILLER_ASAP7_75t_R FILLER_0_67_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_439 ();
 DECAPx1_ASAP7_75t_R FILLER_0_67_447 ();
 DECAPx1_ASAP7_75t_R FILLER_0_67_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_461 ();
 DECAPx1_ASAP7_75t_R FILLER_0_67_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_472 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_480 ();
 DECAPx1_ASAP7_75t_R FILLER_0_67_502 ();
 FILLER_ASAP7_75t_R FILLER_0_67_518 ();
 FILLER_ASAP7_75t_R FILLER_0_67_541 ();
 DECAPx4_ASAP7_75t_R FILLER_0_67_546 ();
 FILLER_ASAP7_75t_R FILLER_0_67_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_558 ();
 FILLER_ASAP7_75t_R FILLER_0_67_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_564 ();
 FILLER_ASAP7_75t_R FILLER_0_67_571 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_594 ();
 DECAPx6_ASAP7_75t_R FILLER_0_67_616 ();
 FILLER_ASAP7_75t_R FILLER_0_67_630 ();
 DECAPx1_ASAP7_75t_R FILLER_0_67_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_639 ();
 FILLER_ASAP7_75t_R FILLER_0_67_644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_654 ();
 DECAPx1_ASAP7_75t_R FILLER_0_67_676 ();
 FILLER_ASAP7_75t_R FILLER_0_67_686 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_694 ();
 FILLER_ASAP7_75t_R FILLER_0_67_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_702 ();
 DECAPx1_ASAP7_75t_R FILLER_0_67_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_713 ();
 FILLER_ASAP7_75t_R FILLER_0_67_720 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_728 ();
 FILLER_ASAP7_75t_R FILLER_0_67_740 ();
 FILLER_ASAP7_75t_R FILLER_0_67_748 ();
 FILLER_ASAP7_75t_R FILLER_0_67_756 ();
 FILLER_ASAP7_75t_R FILLER_0_67_762 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_770 ();
 FILLER_ASAP7_75t_R FILLER_0_67_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_778 ();
 FILLER_ASAP7_75t_R FILLER_0_67_786 ();
 FILLER_ASAP7_75t_R FILLER_0_67_794 ();
 DECAPx6_ASAP7_75t_R FILLER_0_67_802 ();
 DECAPx1_ASAP7_75t_R FILLER_0_67_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_820 ();
 FILLER_ASAP7_75t_R FILLER_0_67_827 ();
 DECAPx4_ASAP7_75t_R FILLER_0_67_836 ();
 DECAPx6_ASAP7_75t_R FILLER_0_67_853 ();
 FILLER_ASAP7_75t_R FILLER_0_67_867 ();
 FILLER_ASAP7_75t_R FILLER_0_67_876 ();
 DECAPx4_ASAP7_75t_R FILLER_0_67_883 ();
 FILLER_ASAP7_75t_R FILLER_0_67_893 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_901 ();
 FILLER_ASAP7_75t_R FILLER_0_67_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_909 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_916 ();
 FILLER_ASAP7_75t_R FILLER_0_67_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_924 ();
 DECAPx1_ASAP7_75t_R FILLER_0_67_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_931 ();
 FILLER_ASAP7_75t_R FILLER_0_67_942 ();
 FILLER_ASAP7_75t_R FILLER_0_67_949 ();
 FILLER_ASAP7_75t_R FILLER_0_67_958 ();
 FILLER_ASAP7_75t_R FILLER_0_67_966 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_968 ();
 FILLER_ASAP7_75t_R FILLER_0_67_975 ();
 FILLER_ASAP7_75t_R FILLER_0_67_983 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_994 ();
 FILLER_ASAP7_75t_R FILLER_0_67_1005 ();
 FILLER_ASAP7_75t_R FILLER_0_67_1017 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_1030 ();
 DECAPx1_ASAP7_75t_R FILLER_0_67_1055 ();
 FILLER_ASAP7_75t_R FILLER_0_67_1069 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_1091 ();
 FILLER_ASAP7_75t_R FILLER_0_67_1105 ();
 FILLER_ASAP7_75t_R FILLER_0_67_1113 ();
 DECAPx1_ASAP7_75t_R FILLER_0_67_1120 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_1132 ();
 FILLER_ASAP7_75t_R FILLER_0_67_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_1140 ();
 DECAPx1_ASAP7_75t_R FILLER_0_67_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_1151 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_1158 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_1180 ();
 DECAPx6_ASAP7_75t_R FILLER_0_67_1197 ();
 FILLER_ASAP7_75t_R FILLER_0_67_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_1213 ();
 FILLER_ASAP7_75t_R FILLER_0_67_1224 ();
 DECAPx1_ASAP7_75t_R FILLER_0_67_1231 ();
 FILLER_ASAP7_75t_R FILLER_0_67_1240 ();
 FILLER_ASAP7_75t_R FILLER_0_67_1252 ();
 FILLER_ASAP7_75t_R FILLER_0_67_1264 ();
 FILLER_ASAP7_75t_R FILLER_0_67_1276 ();
 DECAPx1_ASAP7_75t_R FILLER_0_67_1283 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_1287 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_1304 ();
 FILLER_ASAP7_75t_R FILLER_0_67_1310 ();
 FILLER_ASAP7_75t_R FILLER_0_67_1322 ();
 FILLER_ASAP7_75t_R FILLER_0_67_1329 ();
 FILLER_ASAP7_75t_R FILLER_0_67_1336 ();
 FILLER_ASAP7_75t_R FILLER_0_67_1343 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_1345 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_1356 ();
 FILLER_ASAP7_75t_R FILLER_0_67_1368 ();
 FILLER_ASAP7_75t_R FILLER_0_67_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_68_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_39 ();
 FILLER_ASAP7_75t_R FILLER_0_68_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_45 ();
 FILLER_ASAP7_75t_R FILLER_0_68_52 ();
 FILLER_ASAP7_75t_R FILLER_0_68_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_68 ();
 FILLER_ASAP7_75t_R FILLER_0_68_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_83 ();
 FILLER_ASAP7_75t_R FILLER_0_68_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_98 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_119 ();
 FILLER_ASAP7_75t_R FILLER_0_68_125 ();
 FILLER_ASAP7_75t_R FILLER_0_68_145 ();
 DECAPx1_ASAP7_75t_R FILLER_0_68_155 ();
 FILLER_ASAP7_75t_R FILLER_0_68_165 ();
 FILLER_ASAP7_75t_R FILLER_0_68_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_175 ();
 FILLER_ASAP7_75t_R FILLER_0_68_182 ();
 FILLER_ASAP7_75t_R FILLER_0_68_190 ();
 DECAPx6_ASAP7_75t_R FILLER_0_68_197 ();
 DECAPx1_ASAP7_75t_R FILLER_0_68_211 ();
 DECAPx1_ASAP7_75t_R FILLER_0_68_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_229 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_251 ();
 FILLER_ASAP7_75t_R FILLER_0_68_273 ();
 FILLER_ASAP7_75t_R FILLER_0_68_281 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_295 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_299 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_321 ();
 FILLER_ASAP7_75t_R FILLER_0_68_327 ();
 DECAPx6_ASAP7_75t_R FILLER_0_68_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_350 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_359 ();
 FILLER_ASAP7_75t_R FILLER_0_68_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_367 ();
 FILLER_ASAP7_75t_R FILLER_0_68_371 ();
 FILLER_ASAP7_75t_R FILLER_0_68_379 ();
 DECAPx6_ASAP7_75t_R FILLER_0_68_386 ();
 FILLER_ASAP7_75t_R FILLER_0_68_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_402 ();
 FILLER_ASAP7_75t_R FILLER_0_68_409 ();
 DECAPx1_ASAP7_75t_R FILLER_0_68_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_422 ();
 FILLER_ASAP7_75t_R FILLER_0_68_429 ();
 FILLER_ASAP7_75t_R FILLER_0_68_441 ();
 FILLER_ASAP7_75t_R FILLER_0_68_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_451 ();
 FILLER_ASAP7_75t_R FILLER_0_68_460 ();
 FILLER_ASAP7_75t_R FILLER_0_68_464 ();
 FILLER_ASAP7_75t_R FILLER_0_68_472 ();
 FILLER_ASAP7_75t_R FILLER_0_68_479 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_484 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_506 ();
 FILLER_ASAP7_75t_R FILLER_0_68_512 ();
 FILLER_ASAP7_75t_R FILLER_0_68_517 ();
 FILLER_ASAP7_75t_R FILLER_0_68_529 ();
 DECAPx4_ASAP7_75t_R FILLER_0_68_543 ();
 FILLER_ASAP7_75t_R FILLER_0_68_553 ();
 FILLER_ASAP7_75t_R FILLER_0_68_566 ();
 DECAPx1_ASAP7_75t_R FILLER_0_68_571 ();
 DECAPx6_ASAP7_75t_R FILLER_0_68_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_592 ();
 FILLER_ASAP7_75t_R FILLER_0_68_603 ();
 FILLER_ASAP7_75t_R FILLER_0_68_613 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_643 ();
 DECAPx6_ASAP7_75t_R FILLER_0_68_650 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_664 ();
 DECAPx1_ASAP7_75t_R FILLER_0_68_675 ();
 FILLER_ASAP7_75t_R FILLER_0_68_685 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_692 ();
 FILLER_ASAP7_75t_R FILLER_0_68_698 ();
 FILLER_ASAP7_75t_R FILLER_0_68_711 ();
 FILLER_ASAP7_75t_R FILLER_0_68_719 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_726 ();
 FILLER_ASAP7_75t_R FILLER_0_68_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_734 ();
 FILLER_ASAP7_75t_R FILLER_0_68_741 ();
 FILLER_ASAP7_75t_R FILLER_0_68_749 ();
 FILLER_ASAP7_75t_R FILLER_0_68_757 ();
 DECAPx4_ASAP7_75t_R FILLER_0_68_779 ();
 FILLER_ASAP7_75t_R FILLER_0_68_795 ();
 DECAPx6_ASAP7_75t_R FILLER_0_68_803 ();
 DECAPx1_ASAP7_75t_R FILLER_0_68_817 ();
 FILLER_ASAP7_75t_R FILLER_0_68_831 ();
 FILLER_ASAP7_75t_R FILLER_0_68_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_841 ();
 FILLER_ASAP7_75t_R FILLER_0_68_848 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_856 ();
 FILLER_ASAP7_75t_R FILLER_0_68_868 ();
 FILLER_ASAP7_75t_R FILLER_0_68_875 ();
 FILLER_ASAP7_75t_R FILLER_0_68_881 ();
 FILLER_ASAP7_75t_R FILLER_0_68_889 ();
 FILLER_ASAP7_75t_R FILLER_0_68_897 ();
 FILLER_ASAP7_75t_R FILLER_0_68_905 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_917 ();
 FILLER_ASAP7_75t_R FILLER_0_68_945 ();
 DECAPx1_ASAP7_75t_R FILLER_0_68_967 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_977 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_989 ();
 FILLER_ASAP7_75t_R FILLER_0_68_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_997 ();
 FILLER_ASAP7_75t_R FILLER_0_68_1004 ();
 FILLER_ASAP7_75t_R FILLER_0_68_1016 ();
 FILLER_ASAP7_75t_R FILLER_0_68_1023 ();
 FILLER_ASAP7_75t_R FILLER_0_68_1035 ();
 FILLER_ASAP7_75t_R FILLER_0_68_1047 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_1059 ();
 FILLER_ASAP7_75t_R FILLER_0_68_1083 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_1091 ();
 FILLER_ASAP7_75t_R FILLER_0_68_1097 ();
 FILLER_ASAP7_75t_R FILLER_0_68_1106 ();
 FILLER_ASAP7_75t_R FILLER_0_68_1118 ();
 DECAPx4_ASAP7_75t_R FILLER_0_68_1125 ();
 FILLER_ASAP7_75t_R FILLER_0_68_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_1137 ();
 DECAPx1_ASAP7_75t_R FILLER_0_68_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_1153 ();
 FILLER_ASAP7_75t_R FILLER_0_68_1157 ();
 DECAPx6_ASAP7_75t_R FILLER_0_68_1165 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_1192 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_1214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_1225 ();
 FILLER_ASAP7_75t_R FILLER_0_68_1231 ();
 FILLER_ASAP7_75t_R FILLER_0_68_1238 ();
 DECAPx1_ASAP7_75t_R FILLER_0_68_1250 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_1254 ();
 FILLER_ASAP7_75t_R FILLER_0_68_1265 ();
 FILLER_ASAP7_75t_R FILLER_0_68_1280 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_1287 ();
 FILLER_ASAP7_75t_R FILLER_0_68_1305 ();
 FILLER_ASAP7_75t_R FILLER_0_68_1313 ();
 FILLER_ASAP7_75t_R FILLER_0_68_1320 ();
 DECAPx1_ASAP7_75t_R FILLER_0_68_1327 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_1331 ();
 FILLER_ASAP7_75t_R FILLER_0_68_1338 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_1350 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_1376 ();
 DECAPx4_ASAP7_75t_R FILLER_0_69_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_12 ();
 FILLER_ASAP7_75t_R FILLER_0_69_23 ();
 DECAPx4_ASAP7_75t_R FILLER_0_69_45 ();
 FILLER_ASAP7_75t_R FILLER_0_69_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_57 ();
 DECAPx1_ASAP7_75t_R FILLER_0_69_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_100 ();
 FILLER_ASAP7_75t_R FILLER_0_69_111 ();
 FILLER_ASAP7_75t_R FILLER_0_69_151 ();
 DECAPx1_ASAP7_75t_R FILLER_0_69_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_165 ();
 FILLER_ASAP7_75t_R FILLER_0_69_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_174 ();
 FILLER_ASAP7_75t_R FILLER_0_69_185 ();
 FILLER_ASAP7_75t_R FILLER_0_69_193 ();
 DECAPx4_ASAP7_75t_R FILLER_0_69_201 ();
 FILLER_ASAP7_75t_R FILLER_0_69_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_213 ();
 FILLER_ASAP7_75t_R FILLER_0_69_220 ();
 DECAPx1_ASAP7_75t_R FILLER_0_69_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_232 ();
 FILLER_ASAP7_75t_R FILLER_0_69_239 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_247 ();
 FILLER_ASAP7_75t_R FILLER_0_69_269 ();
 FILLER_ASAP7_75t_R FILLER_0_69_274 ();
 DECAPx1_ASAP7_75t_R FILLER_0_69_284 ();
 FILLER_ASAP7_75t_R FILLER_0_69_291 ();
 FILLER_ASAP7_75t_R FILLER_0_69_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_301 ();
 DECAPx2_ASAP7_75t_R FILLER_0_69_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_314 ();
 FILLER_ASAP7_75t_R FILLER_0_69_321 ();
 DECAPx4_ASAP7_75t_R FILLER_0_69_333 ();
 FILLER_ASAP7_75t_R FILLER_0_69_348 ();
 FILLER_ASAP7_75t_R FILLER_0_69_356 ();
 DECAPx4_ASAP7_75t_R FILLER_0_69_361 ();
 FILLER_ASAP7_75t_R FILLER_0_69_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_373 ();
 DECAPx1_ASAP7_75t_R FILLER_0_69_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_384 ();
 FILLER_ASAP7_75t_R FILLER_0_69_395 ();
 DECAPx4_ASAP7_75t_R FILLER_0_69_402 ();
 FILLER_ASAP7_75t_R FILLER_0_69_418 ();
 FILLER_ASAP7_75t_R FILLER_0_69_428 ();
 DECAPx1_ASAP7_75t_R FILLER_0_69_436 ();
 DECAPx6_ASAP7_75t_R FILLER_0_69_446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_488 ();
 FILLER_ASAP7_75t_R FILLER_0_69_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_512 ();
 DECAPx6_ASAP7_75t_R FILLER_0_69_534 ();
 DECAPx1_ASAP7_75t_R FILLER_0_69_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_552 ();
 FILLER_ASAP7_75t_R FILLER_0_69_556 ();
 DECAPx6_ASAP7_75t_R FILLER_0_69_566 ();
 FILLER_ASAP7_75t_R FILLER_0_69_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_582 ();
 FILLER_ASAP7_75t_R FILLER_0_69_595 ();
 DECAPx2_ASAP7_75t_R FILLER_0_69_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_615 ();
 DECAPx2_ASAP7_75t_R FILLER_0_69_624 ();
 FILLER_ASAP7_75t_R FILLER_0_69_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_632 ();
 FILLER_ASAP7_75t_R FILLER_0_69_639 ();
 DECAPx1_ASAP7_75t_R FILLER_0_69_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_651 ();
 DECAPx1_ASAP7_75t_R FILLER_0_69_658 ();
 FILLER_ASAP7_75t_R FILLER_0_69_683 ();
 DECAPx2_ASAP7_75t_R FILLER_0_69_691 ();
 FILLER_ASAP7_75t_R FILLER_0_69_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_699 ();
 DECAPx4_ASAP7_75t_R FILLER_0_69_706 ();
 FILLER_ASAP7_75t_R FILLER_0_69_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_718 ();
 FILLER_ASAP7_75t_R FILLER_0_69_725 ();
 FILLER_ASAP7_75t_R FILLER_0_69_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_734 ();
 FILLER_ASAP7_75t_R FILLER_0_69_741 ();
 FILLER_ASAP7_75t_R FILLER_0_69_749 ();
 DECAPx1_ASAP7_75t_R FILLER_0_69_756 ();
 DECAPx4_ASAP7_75t_R FILLER_0_69_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_790 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_802 ();
 DECAPx6_ASAP7_75t_R FILLER_0_69_824 ();
 FILLER_ASAP7_75t_R FILLER_0_69_838 ();
 DECAPx2_ASAP7_75t_R FILLER_0_69_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_852 ();
 DECAPx1_ASAP7_75t_R FILLER_0_69_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_863 ();
 FILLER_ASAP7_75t_R FILLER_0_69_874 ();
 FILLER_ASAP7_75t_R FILLER_0_69_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_888 ();
 FILLER_ASAP7_75t_R FILLER_0_69_894 ();
 FILLER_ASAP7_75t_R FILLER_0_69_903 ();
 DECAPx6_ASAP7_75t_R FILLER_0_69_911 ();
 DECAPx4_ASAP7_75t_R FILLER_0_69_927 ();
 FILLER_ASAP7_75t_R FILLER_0_69_937 ();
 DECAPx4_ASAP7_75t_R FILLER_0_69_944 ();
 FILLER_ASAP7_75t_R FILLER_0_69_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_956 ();
 FILLER_ASAP7_75t_R FILLER_0_69_967 ();
 DECAPx1_ASAP7_75t_R FILLER_0_69_976 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_986 ();
 DECAPx1_ASAP7_75t_R FILLER_0_69_1008 ();
 FILLER_ASAP7_75t_R FILLER_0_69_1018 ();
 FILLER_ASAP7_75t_R FILLER_0_69_1028 ();
 FILLER_ASAP7_75t_R FILLER_0_69_1048 ();
 FILLER_ASAP7_75t_R FILLER_0_69_1060 ();
 FILLER_ASAP7_75t_R FILLER_0_69_1067 ();
 FILLER_ASAP7_75t_R FILLER_0_69_1083 ();
 DECAPx1_ASAP7_75t_R FILLER_0_69_1091 ();
 FILLER_ASAP7_75t_R FILLER_0_69_1103 ();
 FILLER_ASAP7_75t_R FILLER_0_69_1125 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_1127 ();
 DECAPx2_ASAP7_75t_R FILLER_0_69_1134 ();
 DECAPx2_ASAP7_75t_R FILLER_0_69_1146 ();
 DECAPx1_ASAP7_75t_R FILLER_0_69_1160 ();
 FILLER_ASAP7_75t_R FILLER_0_69_1170 ();
 DECAPx2_ASAP7_75t_R FILLER_0_69_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_1184 ();
 FILLER_ASAP7_75t_R FILLER_0_69_1188 ();
 DECAPx4_ASAP7_75t_R FILLER_0_69_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_1206 ();
 FILLER_ASAP7_75t_R FILLER_0_69_1237 ();
 DECAPx2_ASAP7_75t_R FILLER_0_69_1249 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_1255 ();
 FILLER_ASAP7_75t_R FILLER_0_69_1268 ();
 FILLER_ASAP7_75t_R FILLER_0_69_1275 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_1277 ();
 DECAPx2_ASAP7_75t_R FILLER_0_69_1284 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_1290 ();
 FILLER_ASAP7_75t_R FILLER_0_69_1303 ();
 DECAPx1_ASAP7_75t_R FILLER_0_69_1315 ();
 DECAPx1_ASAP7_75t_R FILLER_0_69_1329 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_1333 ();
 FILLER_ASAP7_75t_R FILLER_0_69_1340 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_1342 ();
 DECAPx1_ASAP7_75t_R FILLER_0_69_1346 ();
 FILLER_ASAP7_75t_R FILLER_0_69_1360 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_1362 ();
 DECAPx1_ASAP7_75t_R FILLER_0_69_1369 ();
 FILLER_ASAP7_75t_R FILLER_0_69_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_70_34 ();
 FILLER_ASAP7_75t_R FILLER_0_70_44 ();
 DECAPx2_ASAP7_75t_R FILLER_0_70_56 ();
 FILLER_ASAP7_75t_R FILLER_0_70_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_64 ();
 FILLER_ASAP7_75t_R FILLER_0_70_75 ();
 DECAPx1_ASAP7_75t_R FILLER_0_70_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_91 ();
 DECAPx1_ASAP7_75t_R FILLER_0_70_100 ();
 FILLER_ASAP7_75t_R FILLER_0_70_109 ();
 FILLER_ASAP7_75t_R FILLER_0_70_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_141 ();
 FILLER_ASAP7_75t_R FILLER_0_70_152 ();
 FILLER_ASAP7_75t_R FILLER_0_70_164 ();
 DECAPx2_ASAP7_75t_R FILLER_0_70_172 ();
 FILLER_ASAP7_75t_R FILLER_0_70_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_190 ();
 FILLER_ASAP7_75t_R FILLER_0_70_197 ();
 FILLER_ASAP7_75t_R FILLER_0_70_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_213 ();
 DECAPx1_ASAP7_75t_R FILLER_0_70_217 ();
 FILLER_ASAP7_75t_R FILLER_0_70_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_229 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_242 ();
 DECAPx1_ASAP7_75t_R FILLER_0_70_264 ();
 FILLER_ASAP7_75t_R FILLER_0_70_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_276 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_283 ();
 DECAPx2_ASAP7_75t_R FILLER_0_70_305 ();
 FILLER_ASAP7_75t_R FILLER_0_70_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_313 ();
 DECAPx2_ASAP7_75t_R FILLER_0_70_321 ();
 FILLER_ASAP7_75t_R FILLER_0_70_334 ();
 FILLER_ASAP7_75t_R FILLER_0_70_346 ();
 FILLER_ASAP7_75t_R FILLER_0_70_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_356 ();
 DECAPx4_ASAP7_75t_R FILLER_0_70_363 ();
 FILLER_ASAP7_75t_R FILLER_0_70_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_375 ();
 FILLER_ASAP7_75t_R FILLER_0_70_382 ();
 FILLER_ASAP7_75t_R FILLER_0_70_387 ();
 FILLER_ASAP7_75t_R FILLER_0_70_409 ();
 FILLER_ASAP7_75t_R FILLER_0_70_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_416 ();
 DECAPx1_ASAP7_75t_R FILLER_0_70_423 ();
 FILLER_ASAP7_75t_R FILLER_0_70_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_435 ();
 DECAPx6_ASAP7_75t_R FILLER_0_70_444 ();
 DECAPx1_ASAP7_75t_R FILLER_0_70_458 ();
 FILLER_ASAP7_75t_R FILLER_0_70_464 ();
 DECAPx1_ASAP7_75t_R FILLER_0_70_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_476 ();
 DECAPx6_ASAP7_75t_R FILLER_0_70_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_494 ();
 DECAPx6_ASAP7_75t_R FILLER_0_70_505 ();
 DECAPx1_ASAP7_75t_R FILLER_0_70_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_544 ();
 DECAPx1_ASAP7_75t_R FILLER_0_70_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_555 ();
 DECAPx6_ASAP7_75t_R FILLER_0_70_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_582 ();
 FILLER_ASAP7_75t_R FILLER_0_70_586 ();
 FILLER_ASAP7_75t_R FILLER_0_70_600 ();
 FILLER_ASAP7_75t_R FILLER_0_70_614 ();
 FILLER_ASAP7_75t_R FILLER_0_70_637 ();
 FILLER_ASAP7_75t_R FILLER_0_70_650 ();
 FILLER_ASAP7_75t_R FILLER_0_70_664 ();
 DECAPx4_ASAP7_75t_R FILLER_0_70_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_679 ();
 DECAPx4_ASAP7_75t_R FILLER_0_70_691 ();
 FILLER_ASAP7_75t_R FILLER_0_70_701 ();
 DECAPx1_ASAP7_75t_R FILLER_0_70_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_712 ();
 FILLER_ASAP7_75t_R FILLER_0_70_719 ();
 DECAPx2_ASAP7_75t_R FILLER_0_70_727 ();
 FILLER_ASAP7_75t_R FILLER_0_70_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_735 ();
 FILLER_ASAP7_75t_R FILLER_0_70_742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_750 ();
 DECAPx4_ASAP7_75t_R FILLER_0_70_772 ();
 FILLER_ASAP7_75t_R FILLER_0_70_789 ();
 FILLER_ASAP7_75t_R FILLER_0_70_799 ();
 DECAPx2_ASAP7_75t_R FILLER_0_70_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_813 ();
 FILLER_ASAP7_75t_R FILLER_0_70_825 ();
 DECAPx1_ASAP7_75t_R FILLER_0_70_833 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_840 ();
 DECAPx2_ASAP7_75t_R FILLER_0_70_862 ();
 FILLER_ASAP7_75t_R FILLER_0_70_868 ();
 DECAPx1_ASAP7_75t_R FILLER_0_70_890 ();
 DECAPx1_ASAP7_75t_R FILLER_0_70_900 ();
 FILLER_ASAP7_75t_R FILLER_0_70_910 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_918 ();
 DECAPx2_ASAP7_75t_R FILLER_0_70_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_946 ();
 FILLER_ASAP7_75t_R FILLER_0_70_957 ();
 FILLER_ASAP7_75t_R FILLER_0_70_965 ();
 FILLER_ASAP7_75t_R FILLER_0_70_973 ();
 DECAPx2_ASAP7_75t_R FILLER_0_70_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_987 ();
 FILLER_ASAP7_75t_R FILLER_0_70_999 ();
 FILLER_ASAP7_75t_R FILLER_0_70_1007 ();
 DECAPx2_ASAP7_75t_R FILLER_0_70_1020 ();
 FILLER_ASAP7_75t_R FILLER_0_70_1026 ();
 FILLER_ASAP7_75t_R FILLER_0_70_1038 ();
 DECAPx2_ASAP7_75t_R FILLER_0_70_1050 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_1056 ();
 DECAPx1_ASAP7_75t_R FILLER_0_70_1067 ();
 FILLER_ASAP7_75t_R FILLER_0_70_1091 ();
 DECAPx2_ASAP7_75t_R FILLER_0_70_1099 ();
 FILLER_ASAP7_75t_R FILLER_0_70_1125 ();
 DECAPx1_ASAP7_75t_R FILLER_0_70_1137 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_1141 ();
 DECAPx1_ASAP7_75t_R FILLER_0_70_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_1156 ();
 DECAPx2_ASAP7_75t_R FILLER_0_70_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_1169 ();
 DECAPx2_ASAP7_75t_R FILLER_0_70_1176 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_1182 ();
 DECAPx2_ASAP7_75t_R FILLER_0_70_1189 ();
 FILLER_ASAP7_75t_R FILLER_0_70_1205 ();
 DECAPx1_ASAP7_75t_R FILLER_0_70_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_1221 ();
 FILLER_ASAP7_75t_R FILLER_0_70_1232 ();
 FILLER_ASAP7_75t_R FILLER_0_70_1244 ();
 FILLER_ASAP7_75t_R FILLER_0_70_1254 ();
 DECAPx2_ASAP7_75t_R FILLER_0_70_1268 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_1274 ();
 DECAPx1_ASAP7_75t_R FILLER_0_70_1283 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_1287 ();
 FILLER_ASAP7_75t_R FILLER_0_70_1300 ();
 FILLER_ASAP7_75t_R FILLER_0_70_1322 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_1324 ();
 FILLER_ASAP7_75t_R FILLER_0_70_1331 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_1333 ();
 FILLER_ASAP7_75t_R FILLER_0_70_1337 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_1339 ();
 FILLER_ASAP7_75t_R FILLER_0_70_1350 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_1352 ();
 DECAPx2_ASAP7_75t_R FILLER_0_70_1359 ();
 FILLER_ASAP7_75t_R FILLER_0_70_1365 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_1367 ();
 DECAPx4_ASAP7_75t_R FILLER_0_70_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_71_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_30 ();
 FILLER_ASAP7_75t_R FILLER_0_71_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_41 ();
 FILLER_ASAP7_75t_R FILLER_0_71_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_64 ();
 FILLER_ASAP7_75t_R FILLER_0_71_75 ();
 FILLER_ASAP7_75t_R FILLER_0_71_97 ();
 FILLER_ASAP7_75t_R FILLER_0_71_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_121 ();
 FILLER_ASAP7_75t_R FILLER_0_71_132 ();
 FILLER_ASAP7_75t_R FILLER_0_71_152 ();
 FILLER_ASAP7_75t_R FILLER_0_71_164 ();
 FILLER_ASAP7_75t_R FILLER_0_71_174 ();
 FILLER_ASAP7_75t_R FILLER_0_71_181 ();
 DECAPx2_ASAP7_75t_R FILLER_0_71_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_203 ();
 DECAPx2_ASAP7_75t_R FILLER_0_71_210 ();
 FILLER_ASAP7_75t_R FILLER_0_71_216 ();
 DECAPx2_ASAP7_75t_R FILLER_0_71_224 ();
 FILLER_ASAP7_75t_R FILLER_0_71_240 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_270 ();
 FILLER_ASAP7_75t_R FILLER_0_71_274 ();
 DECAPx2_ASAP7_75t_R FILLER_0_71_284 ();
 FILLER_ASAP7_75t_R FILLER_0_71_290 ();
 FILLER_ASAP7_75t_R FILLER_0_71_299 ();
 DECAPx2_ASAP7_75t_R FILLER_0_71_305 ();
 FILLER_ASAP7_75t_R FILLER_0_71_311 ();
 FILLER_ASAP7_75t_R FILLER_0_71_319 ();
 FILLER_ASAP7_75t_R FILLER_0_71_331 ();
 DECAPx2_ASAP7_75t_R FILLER_0_71_339 ();
 FILLER_ASAP7_75t_R FILLER_0_71_355 ();
 DECAPx1_ASAP7_75t_R FILLER_0_71_365 ();
 FILLER_ASAP7_75t_R FILLER_0_71_375 ();
 FILLER_ASAP7_75t_R FILLER_0_71_387 ();
 DECAPx4_ASAP7_75t_R FILLER_0_71_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_405 ();
 DECAPx1_ASAP7_75t_R FILLER_0_71_413 ();
 FILLER_ASAP7_75t_R FILLER_0_71_424 ();
 DECAPx1_ASAP7_75t_R FILLER_0_71_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_436 ();
 DECAPx2_ASAP7_75t_R FILLER_0_71_445 ();
 FILLER_ASAP7_75t_R FILLER_0_71_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_453 ();
 FILLER_ASAP7_75t_R FILLER_0_71_461 ();
 FILLER_ASAP7_75t_R FILLER_0_71_469 ();
 FILLER_ASAP7_75t_R FILLER_0_71_479 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_484 ();
 DECAPx4_ASAP7_75t_R FILLER_0_71_506 ();
 FILLER_ASAP7_75t_R FILLER_0_71_516 ();
 FILLER_ASAP7_75t_R FILLER_0_71_521 ();
 FILLER_ASAP7_75t_R FILLER_0_71_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_531 ();
 FILLER_ASAP7_75t_R FILLER_0_71_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_537 ();
 DECAPx2_ASAP7_75t_R FILLER_0_71_541 ();
 FILLER_ASAP7_75t_R FILLER_0_71_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_549 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_556 ();
 FILLER_ASAP7_75t_R FILLER_0_71_578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_592 ();
 DECAPx1_ASAP7_75t_R FILLER_0_71_614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_621 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_643 ();
 DECAPx2_ASAP7_75t_R FILLER_0_71_665 ();
 FILLER_ASAP7_75t_R FILLER_0_71_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_673 ();
 FILLER_ASAP7_75t_R FILLER_0_71_680 ();
 DECAPx2_ASAP7_75t_R FILLER_0_71_692 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_703 ();
 DECAPx1_ASAP7_75t_R FILLER_0_71_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_729 ();
 FILLER_ASAP7_75t_R FILLER_0_71_733 ();
 FILLER_ASAP7_75t_R FILLER_0_71_745 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_753 ();
 DECAPx2_ASAP7_75t_R FILLER_0_71_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_781 ();
 FILLER_ASAP7_75t_R FILLER_0_71_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_791 ();
 FILLER_ASAP7_75t_R FILLER_0_71_812 ();
 DECAPx2_ASAP7_75t_R FILLER_0_71_820 ();
 FILLER_ASAP7_75t_R FILLER_0_71_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_828 ();
 FILLER_ASAP7_75t_R FILLER_0_71_835 ();
 DECAPx2_ASAP7_75t_R FILLER_0_71_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_854 ();
 DECAPx1_ASAP7_75t_R FILLER_0_71_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_870 ();
 FILLER_ASAP7_75t_R FILLER_0_71_879 ();
 FILLER_ASAP7_75t_R FILLER_0_71_891 ();
 FILLER_ASAP7_75t_R FILLER_0_71_899 ();
 DECAPx1_ASAP7_75t_R FILLER_0_71_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_911 ();
 DECAPx1_ASAP7_75t_R FILLER_0_71_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_924 ();
 DECAPx4_ASAP7_75t_R FILLER_0_71_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_937 ();
 FILLER_ASAP7_75t_R FILLER_0_71_943 ();
 FILLER_ASAP7_75t_R FILLER_0_71_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_952 ();
 FILLER_ASAP7_75t_R FILLER_0_71_959 ();
 DECAPx1_ASAP7_75t_R FILLER_0_71_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_971 ();
 FILLER_ASAP7_75t_R FILLER_0_71_982 ();
 FILLER_ASAP7_75t_R FILLER_0_71_989 ();
 DECAPx6_ASAP7_75t_R FILLER_0_71_997 ();
 DECAPx4_ASAP7_75t_R FILLER_0_71_1017 ();
 DECAPx1_ASAP7_75t_R FILLER_0_71_1037 ();
 FILLER_ASAP7_75t_R FILLER_0_71_1046 ();
 FILLER_ASAP7_75t_R FILLER_0_71_1054 ();
 FILLER_ASAP7_75t_R FILLER_0_71_1067 ();
 DECAPx2_ASAP7_75t_R FILLER_0_71_1079 ();
 FILLER_ASAP7_75t_R FILLER_0_71_1085 ();
 FILLER_ASAP7_75t_R FILLER_0_71_1093 ();
 DECAPx6_ASAP7_75t_R FILLER_0_71_1101 ();
 FILLER_ASAP7_75t_R FILLER_0_71_1115 ();
 FILLER_ASAP7_75t_R FILLER_0_71_1125 ();
 FILLER_ASAP7_75t_R FILLER_0_71_1133 ();
 FILLER_ASAP7_75t_R FILLER_0_71_1140 ();
 FILLER_ASAP7_75t_R FILLER_0_71_1145 ();
 FILLER_ASAP7_75t_R FILLER_0_71_1150 ();
 DECAPx6_ASAP7_75t_R FILLER_0_71_1158 ();
 FILLER_ASAP7_75t_R FILLER_0_71_1178 ();
 DECAPx6_ASAP7_75t_R FILLER_0_71_1186 ();
 DECAPx1_ASAP7_75t_R FILLER_0_71_1208 ();
 DECAPx4_ASAP7_75t_R FILLER_0_71_1217 ();
 FILLER_ASAP7_75t_R FILLER_0_71_1227 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_1229 ();
 FILLER_ASAP7_75t_R FILLER_0_71_1240 ();
 FILLER_ASAP7_75t_R FILLER_0_71_1247 ();
 DECAPx2_ASAP7_75t_R FILLER_0_71_1254 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_1260 ();
 DECAPx2_ASAP7_75t_R FILLER_0_71_1267 ();
 FILLER_ASAP7_75t_R FILLER_0_71_1279 ();
 FILLER_ASAP7_75t_R FILLER_0_71_1287 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_1289 ();
 FILLER_ASAP7_75t_R FILLER_0_71_1296 ();
 DECAPx1_ASAP7_75t_R FILLER_0_71_1308 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_1312 ();
 FILLER_ASAP7_75t_R FILLER_0_71_1316 ();
 FILLER_ASAP7_75t_R FILLER_0_71_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_1337 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_1359 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_72_24 ();
 FILLER_ASAP7_75t_R FILLER_0_72_34 ();
 FILLER_ASAP7_75t_R FILLER_0_72_42 ();
 FILLER_ASAP7_75t_R FILLER_0_72_50 ();
 FILLER_ASAP7_75t_R FILLER_0_72_55 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_69 ();
 FILLER_ASAP7_75t_R FILLER_0_72_75 ();
 FILLER_ASAP7_75t_R FILLER_0_72_85 ();
 FILLER_ASAP7_75t_R FILLER_0_72_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_96 ();
 FILLER_ASAP7_75t_R FILLER_0_72_105 ();
 FILLER_ASAP7_75t_R FILLER_0_72_117 ();
 FILLER_ASAP7_75t_R FILLER_0_72_129 ();
 FILLER_ASAP7_75t_R FILLER_0_72_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_143 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_164 ();
 FILLER_ASAP7_75t_R FILLER_0_72_180 ();
 DECAPx1_ASAP7_75t_R FILLER_0_72_192 ();
 FILLER_ASAP7_75t_R FILLER_0_72_202 ();
 FILLER_ASAP7_75t_R FILLER_0_72_211 ();
 FILLER_ASAP7_75t_R FILLER_0_72_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_218 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_229 ();
 DECAPx4_ASAP7_75t_R FILLER_0_72_251 ();
 FILLER_ASAP7_75t_R FILLER_0_72_261 ();
 FILLER_ASAP7_75t_R FILLER_0_72_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_289 ();
 DECAPx1_ASAP7_75t_R FILLER_0_72_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_302 ();
 FILLER_ASAP7_75t_R FILLER_0_72_309 ();
 DECAPx1_ASAP7_75t_R FILLER_0_72_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_321 ();
 FILLER_ASAP7_75t_R FILLER_0_72_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_330 ();
 DECAPx1_ASAP7_75t_R FILLER_0_72_337 ();
 FILLER_ASAP7_75t_R FILLER_0_72_346 ();
 FILLER_ASAP7_75t_R FILLER_0_72_353 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_365 ();
 FILLER_ASAP7_75t_R FILLER_0_72_383 ();
 DECAPx4_ASAP7_75t_R FILLER_0_72_390 ();
 FILLER_ASAP7_75t_R FILLER_0_72_400 ();
 DECAPx1_ASAP7_75t_R FILLER_0_72_408 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_422 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_434 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_446 ();
 FILLER_ASAP7_75t_R FILLER_0_72_460 ();
 FILLER_ASAP7_75t_R FILLER_0_72_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_466 ();
 FILLER_ASAP7_75t_R FILLER_0_72_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_476 ();
 DECAPx6_ASAP7_75t_R FILLER_0_72_483 ();
 DECAPx1_ASAP7_75t_R FILLER_0_72_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_501 ();
 FILLER_ASAP7_75t_R FILLER_0_72_508 ();
 DECAPx1_ASAP7_75t_R FILLER_0_72_516 ();
 DECAPx6_ASAP7_75t_R FILLER_0_72_526 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_540 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_586 ();
 DECAPx6_ASAP7_75t_R FILLER_0_72_608 ();
 FILLER_ASAP7_75t_R FILLER_0_72_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_624 ();
 DECAPx1_ASAP7_75t_R FILLER_0_72_637 ();
 FILLER_ASAP7_75t_R FILLER_0_72_649 ();
 FILLER_ASAP7_75t_R FILLER_0_72_663 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_677 ();
 FILLER_ASAP7_75t_R FILLER_0_72_689 ();
 FILLER_ASAP7_75t_R FILLER_0_72_697 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_705 ();
 FILLER_ASAP7_75t_R FILLER_0_72_711 ();
 DECAPx1_ASAP7_75t_R FILLER_0_72_719 ();
 DECAPx4_ASAP7_75t_R FILLER_0_72_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_739 ();
 DECAPx6_ASAP7_75t_R FILLER_0_72_746 ();
 FILLER_ASAP7_75t_R FILLER_0_72_766 ();
 FILLER_ASAP7_75t_R FILLER_0_72_774 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_779 ();
 FILLER_ASAP7_75t_R FILLER_0_72_785 ();
 FILLER_ASAP7_75t_R FILLER_0_72_793 ();
 DECAPx1_ASAP7_75t_R FILLER_0_72_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_806 ();
 FILLER_ASAP7_75t_R FILLER_0_72_814 ();
 FILLER_ASAP7_75t_R FILLER_0_72_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_824 ();
 FILLER_ASAP7_75t_R FILLER_0_72_831 ();
 FILLER_ASAP7_75t_R FILLER_0_72_843 ();
 FILLER_ASAP7_75t_R FILLER_0_72_851 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_865 ();
 FILLER_ASAP7_75t_R FILLER_0_72_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_879 ();
 FILLER_ASAP7_75t_R FILLER_0_72_890 ();
 DECAPx6_ASAP7_75t_R FILLER_0_72_898 ();
 FILLER_ASAP7_75t_R FILLER_0_72_912 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_920 ();
 DECAPx1_ASAP7_75t_R FILLER_0_72_942 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_953 ();
 DECAPx1_ASAP7_75t_R FILLER_0_72_965 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_969 ();
 DECAPx4_ASAP7_75t_R FILLER_0_72_976 ();
 FILLER_ASAP7_75t_R FILLER_0_72_986 ();
 DECAPx4_ASAP7_75t_R FILLER_0_72_991 ();
 FILLER_ASAP7_75t_R FILLER_0_72_1008 ();
 DECAPx6_ASAP7_75t_R FILLER_0_72_1015 ();
 FILLER_ASAP7_75t_R FILLER_0_72_1029 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_1037 ();
 FILLER_ASAP7_75t_R FILLER_0_72_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_1045 ();
 FILLER_ASAP7_75t_R FILLER_0_72_1051 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_1067 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_1074 ();
 FILLER_ASAP7_75t_R FILLER_0_72_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_1087 ();
 FILLER_ASAP7_75t_R FILLER_0_72_1101 ();
 FILLER_ASAP7_75t_R FILLER_0_72_1109 ();
 FILLER_ASAP7_75t_R FILLER_0_72_1117 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_1125 ();
 DECAPx1_ASAP7_75t_R FILLER_0_72_1137 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_1153 ();
 DECAPx6_ASAP7_75t_R FILLER_0_72_1160 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_1174 ();
 DECAPx1_ASAP7_75t_R FILLER_0_72_1186 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_1190 ();
 FILLER_ASAP7_75t_R FILLER_0_72_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_1202 ();
 DECAPx4_ASAP7_75t_R FILLER_0_72_1224 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_1245 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_1267 ();
 FILLER_ASAP7_75t_R FILLER_0_72_1273 ();
 FILLER_ASAP7_75t_R FILLER_0_72_1281 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_1332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_1354 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_2 ();
 FILLER_ASAP7_75t_R FILLER_0_73_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_26 ();
 FILLER_ASAP7_75t_R FILLER_0_73_30 ();
 FILLER_ASAP7_75t_R FILLER_0_73_38 ();
 FILLER_ASAP7_75t_R FILLER_0_73_46 ();
 DECAPx6_ASAP7_75t_R FILLER_0_73_54 ();
 FILLER_ASAP7_75t_R FILLER_0_73_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_70 ();
 FILLER_ASAP7_75t_R FILLER_0_73_77 ();
 FILLER_ASAP7_75t_R FILLER_0_73_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_101 ();
 FILLER_ASAP7_75t_R FILLER_0_73_110 ();
 FILLER_ASAP7_75t_R FILLER_0_73_122 ();
 FILLER_ASAP7_75t_R FILLER_0_73_134 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_146 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_162 ();
 FILLER_ASAP7_75t_R FILLER_0_73_173 ();
 FILLER_ASAP7_75t_R FILLER_0_73_185 ();
 FILLER_ASAP7_75t_R FILLER_0_73_201 ();
 FILLER_ASAP7_75t_R FILLER_0_73_211 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_219 ();
 DECAPx2_ASAP7_75t_R FILLER_0_73_229 ();
 FILLER_ASAP7_75t_R FILLER_0_73_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_237 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_241 ();
 FILLER_ASAP7_75t_R FILLER_0_73_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_271 ();
 FILLER_ASAP7_75t_R FILLER_0_73_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_280 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_284 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_302 ();
 FILLER_ASAP7_75t_R FILLER_0_73_309 ();
 FILLER_ASAP7_75t_R FILLER_0_73_321 ();
 FILLER_ASAP7_75t_R FILLER_0_73_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_331 ();
 FILLER_ASAP7_75t_R FILLER_0_73_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_342 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_346 ();
 DECAPx2_ASAP7_75t_R FILLER_0_73_360 ();
 FILLER_ASAP7_75t_R FILLER_0_73_366 ();
 FILLER_ASAP7_75t_R FILLER_0_73_374 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_385 ();
 FILLER_ASAP7_75t_R FILLER_0_73_390 ();
 FILLER_ASAP7_75t_R FILLER_0_73_398 ();
 DECAPx4_ASAP7_75t_R FILLER_0_73_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_416 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_423 ();
 FILLER_ASAP7_75t_R FILLER_0_73_445 ();
 FILLER_ASAP7_75t_R FILLER_0_73_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_455 ();
 FILLER_ASAP7_75t_R FILLER_0_73_462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_470 ();
 DECAPx2_ASAP7_75t_R FILLER_0_73_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_504 ();
 DECAPx2_ASAP7_75t_R FILLER_0_73_516 ();
 FILLER_ASAP7_75t_R FILLER_0_73_528 ();
 FILLER_ASAP7_75t_R FILLER_0_73_536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_544 ();
 FILLER_ASAP7_75t_R FILLER_0_73_554 ();
 FILLER_ASAP7_75t_R FILLER_0_73_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_565 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_576 ();
 DECAPx2_ASAP7_75t_R FILLER_0_73_583 ();
 FILLER_ASAP7_75t_R FILLER_0_73_595 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_603 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_625 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_645 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_661 ();
 FILLER_ASAP7_75t_R FILLER_0_73_673 ();
 FILLER_ASAP7_75t_R FILLER_0_73_678 ();
 DECAPx2_ASAP7_75t_R FILLER_0_73_686 ();
 FILLER_ASAP7_75t_R FILLER_0_73_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_694 ();
 FILLER_ASAP7_75t_R FILLER_0_73_701 ();
 FILLER_ASAP7_75t_R FILLER_0_73_709 ();
 FILLER_ASAP7_75t_R FILLER_0_73_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_719 ();
 FILLER_ASAP7_75t_R FILLER_0_73_726 ();
 DECAPx6_ASAP7_75t_R FILLER_0_73_734 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_748 ();
 FILLER_ASAP7_75t_R FILLER_0_73_762 ();
 DECAPx6_ASAP7_75t_R FILLER_0_73_770 ();
 FILLER_ASAP7_75t_R FILLER_0_73_784 ();
 FILLER_ASAP7_75t_R FILLER_0_73_796 ();
 DECAPx4_ASAP7_75t_R FILLER_0_73_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_816 ();
 DECAPx4_ASAP7_75t_R FILLER_0_73_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_833 ();
 DECAPx6_ASAP7_75t_R FILLER_0_73_844 ();
 FILLER_ASAP7_75t_R FILLER_0_73_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_860 ();
 FILLER_ASAP7_75t_R FILLER_0_73_867 ();
 DECAPx2_ASAP7_75t_R FILLER_0_73_875 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_908 ();
 DECAPx4_ASAP7_75t_R FILLER_0_73_915 ();
 DECAPx4_ASAP7_75t_R FILLER_0_73_927 ();
 FILLER_ASAP7_75t_R FILLER_0_73_937 ();
 FILLER_ASAP7_75t_R FILLER_0_73_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_953 ();
 FILLER_ASAP7_75t_R FILLER_0_73_959 ();
 DECAPx2_ASAP7_75t_R FILLER_0_73_967 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_980 ();
 DECAPx2_ASAP7_75t_R FILLER_0_73_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_994 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_1005 ();
 DECAPx2_ASAP7_75t_R FILLER_0_73_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_1018 ();
 DECAPx2_ASAP7_75t_R FILLER_0_73_1029 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_1049 ();
 FILLER_ASAP7_75t_R FILLER_0_73_1056 ();
 DECAPx2_ASAP7_75t_R FILLER_0_73_1066 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_1079 ();
 DECAPx6_ASAP7_75t_R FILLER_0_73_1088 ();
 FILLER_ASAP7_75t_R FILLER_0_73_1102 ();
 DECAPx4_ASAP7_75t_R FILLER_0_73_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_1120 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_1126 ();
 FILLER_ASAP7_75t_R FILLER_0_73_1140 ();
 DECAPx2_ASAP7_75t_R FILLER_0_73_1148 ();
 FILLER_ASAP7_75t_R FILLER_0_73_1154 ();
 FILLER_ASAP7_75t_R FILLER_0_73_1163 ();
 DECAPx2_ASAP7_75t_R FILLER_0_73_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_1181 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_1266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_1332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_1354 ();
 DECAPx2_ASAP7_75t_R FILLER_0_73_1376 ();
 DECAPx2_ASAP7_75t_R FILLER_0_74_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_8 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_15 ();
 DECAPx2_ASAP7_75t_R FILLER_0_74_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_74_49 ();
 FILLER_ASAP7_75t_R FILLER_0_74_67 ();
 FILLER_ASAP7_75t_R FILLER_0_74_74 ();
 FILLER_ASAP7_75t_R FILLER_0_74_81 ();
 DECAPx2_ASAP7_75t_R FILLER_0_74_93 ();
 FILLER_ASAP7_75t_R FILLER_0_74_99 ();
 DECAPx1_ASAP7_75t_R FILLER_0_74_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_115 ();
 DECAPx2_ASAP7_75t_R FILLER_0_74_126 ();
 FILLER_ASAP7_75t_R FILLER_0_74_142 ();
 FILLER_ASAP7_75t_R FILLER_0_74_154 ();
 FILLER_ASAP7_75t_R FILLER_0_74_164 ();
 DECAPx2_ASAP7_75t_R FILLER_0_74_172 ();
 FILLER_ASAP7_75t_R FILLER_0_74_188 ();
 DECAPx1_ASAP7_75t_R FILLER_0_74_198 ();
 FILLER_ASAP7_75t_R FILLER_0_74_208 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_260 ();
 DECAPx4_ASAP7_75t_R FILLER_0_74_282 ();
 DECAPx1_ASAP7_75t_R FILLER_0_74_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_301 ();
 DECAPx1_ASAP7_75t_R FILLER_0_74_312 ();
 FILLER_ASAP7_75t_R FILLER_0_74_319 ();
 DECAPx2_ASAP7_75t_R FILLER_0_74_331 ();
 DECAPx1_ASAP7_75t_R FILLER_0_74_345 ();
 FILLER_ASAP7_75t_R FILLER_0_74_359 ();
 FILLER_ASAP7_75t_R FILLER_0_74_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_375 ();
 DECAPx6_ASAP7_75t_R FILLER_0_74_397 ();
 DECAPx1_ASAP7_75t_R FILLER_0_74_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_415 ();
 DECAPx1_ASAP7_75t_R FILLER_0_74_426 ();
 DECAPx1_ASAP7_75t_R FILLER_0_74_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_74_446 ();
 FILLER_ASAP7_75t_R FILLER_0_74_460 ();
 DECAPx1_ASAP7_75t_R FILLER_0_74_464 ();
 DECAPx6_ASAP7_75t_R FILLER_0_74_476 ();
 DECAPx2_ASAP7_75t_R FILLER_0_74_490 ();
 FILLER_ASAP7_75t_R FILLER_0_74_502 ();
 FILLER_ASAP7_75t_R FILLER_0_74_510 ();
 FILLER_ASAP7_75t_R FILLER_0_74_518 ();
 FILLER_ASAP7_75t_R FILLER_0_74_526 ();
 FILLER_ASAP7_75t_R FILLER_0_74_534 ();
 DECAPx1_ASAP7_75t_R FILLER_0_74_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_546 ();
 DECAPx2_ASAP7_75t_R FILLER_0_74_557 ();
 FILLER_ASAP7_75t_R FILLER_0_74_563 ();
 DECAPx1_ASAP7_75t_R FILLER_0_74_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_589 ();
 FILLER_ASAP7_75t_R FILLER_0_74_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_599 ();
 FILLER_ASAP7_75t_R FILLER_0_74_606 ();
 FILLER_ASAP7_75t_R FILLER_0_74_614 ();
 FILLER_ASAP7_75t_R FILLER_0_74_622 ();
 FILLER_ASAP7_75t_R FILLER_0_74_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_633 ();
 DECAPx2_ASAP7_75t_R FILLER_0_74_655 ();
 FILLER_ASAP7_75t_R FILLER_0_74_664 ();
 FILLER_ASAP7_75t_R FILLER_0_74_674 ();
 DECAPx1_ASAP7_75t_R FILLER_0_74_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_686 ();
 DECAPx2_ASAP7_75t_R FILLER_0_74_693 ();
 FILLER_ASAP7_75t_R FILLER_0_74_699 ();
 DECAPx1_ASAP7_75t_R FILLER_0_74_709 ();
 DECAPx2_ASAP7_75t_R FILLER_0_74_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_725 ();
 FILLER_ASAP7_75t_R FILLER_0_74_732 ();
 FILLER_ASAP7_75t_R FILLER_0_74_740 ();
 FILLER_ASAP7_75t_R FILLER_0_74_748 ();
 FILLER_ASAP7_75t_R FILLER_0_74_756 ();
 FILLER_ASAP7_75t_R FILLER_0_74_764 ();
 DECAPx6_ASAP7_75t_R FILLER_0_74_769 ();
 DECAPx2_ASAP7_75t_R FILLER_0_74_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_789 ();
 DECAPx2_ASAP7_75t_R FILLER_0_74_796 ();
 DECAPx4_ASAP7_75t_R FILLER_0_74_808 ();
 FILLER_ASAP7_75t_R FILLER_0_74_824 ();
 FILLER_ASAP7_75t_R FILLER_0_74_829 ();
 FILLER_ASAP7_75t_R FILLER_0_74_838 ();
 DECAPx4_ASAP7_75t_R FILLER_0_74_850 ();
 FILLER_ASAP7_75t_R FILLER_0_74_868 ();
 DECAPx2_ASAP7_75t_R FILLER_0_74_876 ();
 DECAPx1_ASAP7_75t_R FILLER_0_74_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_896 ();
 FILLER_ASAP7_75t_R FILLER_0_74_903 ();
 FILLER_ASAP7_75t_R FILLER_0_74_911 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_919 ();
 DECAPx2_ASAP7_75t_R FILLER_0_74_941 ();
 DECAPx1_ASAP7_75t_R FILLER_0_74_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_959 ();
 DECAPx2_ASAP7_75t_R FILLER_0_74_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_976 ();
 FILLER_ASAP7_75t_R FILLER_0_74_983 ();
 DECAPx4_ASAP7_75t_R FILLER_0_74_991 ();
 FILLER_ASAP7_75t_R FILLER_0_74_1001 ();
 FILLER_ASAP7_75t_R FILLER_0_74_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_1015 ();
 DECAPx4_ASAP7_75t_R FILLER_0_74_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_1030 ();
 FILLER_ASAP7_75t_R FILLER_0_74_1035 ();
 DECAPx1_ASAP7_75t_R FILLER_0_74_1041 ();
 DECAPx6_ASAP7_75t_R FILLER_0_74_1050 ();
 FILLER_ASAP7_75t_R FILLER_0_74_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_1086 ();
 DECAPx1_ASAP7_75t_R FILLER_0_74_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_1098 ();
 FILLER_ASAP7_75t_R FILLER_0_74_1119 ();
 FILLER_ASAP7_75t_R FILLER_0_74_1127 ();
 DECAPx2_ASAP7_75t_R FILLER_0_74_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_1141 ();
 FILLER_ASAP7_75t_R FILLER_0_74_1148 ();
 DECAPx2_ASAP7_75t_R FILLER_0_74_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_1162 ();
 DECAPx6_ASAP7_75t_R FILLER_0_74_1169 ();
 DECAPx1_ASAP7_75t_R FILLER_0_74_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_1251 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_1273 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_1295 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_1317 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_1339 ();
 DECAPx6_ASAP7_75t_R FILLER_0_74_1361 ();
 DECAPx2_ASAP7_75t_R FILLER_0_74_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_75_2 ();
 FILLER_ASAP7_75t_R FILLER_0_75_25 ();
 FILLER_ASAP7_75t_R FILLER_0_75_33 ();
 DECAPx1_ASAP7_75t_R FILLER_0_75_41 ();
 DECAPx2_ASAP7_75t_R FILLER_0_75_51 ();
 DECAPx1_ASAP7_75t_R FILLER_0_75_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_71 ();
 FILLER_ASAP7_75t_R FILLER_0_75_77 ();
 FILLER_ASAP7_75t_R FILLER_0_75_84 ();
 DECAPx2_ASAP7_75t_R FILLER_0_75_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_98 ();
 FILLER_ASAP7_75t_R FILLER_0_75_104 ();
 FILLER_ASAP7_75t_R FILLER_0_75_111 ();
 FILLER_ASAP7_75t_R FILLER_0_75_118 ();
 FILLER_ASAP7_75t_R FILLER_0_75_130 ();
 FILLER_ASAP7_75t_R FILLER_0_75_135 ();
 FILLER_ASAP7_75t_R FILLER_0_75_155 ();
 FILLER_ASAP7_75t_R FILLER_0_75_162 ();
 FILLER_ASAP7_75t_R FILLER_0_75_174 ();
 FILLER_ASAP7_75t_R FILLER_0_75_182 ();
 DECAPx1_ASAP7_75t_R FILLER_0_75_194 ();
 FILLER_ASAP7_75t_R FILLER_0_75_204 ();
 FILLER_ASAP7_75t_R FILLER_0_75_212 ();
 FILLER_ASAP7_75t_R FILLER_0_75_220 ();
 FILLER_ASAP7_75t_R FILLER_0_75_228 ();
 FILLER_ASAP7_75t_R FILLER_0_75_236 ();
 FILLER_ASAP7_75t_R FILLER_0_75_241 ();
 DECAPx1_ASAP7_75t_R FILLER_0_75_249 ();
 DECAPx2_ASAP7_75t_R FILLER_0_75_259 ();
 FILLER_ASAP7_75t_R FILLER_0_75_273 ();
 FILLER_ASAP7_75t_R FILLER_0_75_278 ();
 FILLER_ASAP7_75t_R FILLER_0_75_285 ();
 FILLER_ASAP7_75t_R FILLER_0_75_297 ();
 FILLER_ASAP7_75t_R FILLER_0_75_305 ();
 DECAPx1_ASAP7_75t_R FILLER_0_75_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_321 ();
 FILLER_ASAP7_75t_R FILLER_0_75_328 ();
 DECAPx6_ASAP7_75t_R FILLER_0_75_336 ();
 DECAPx1_ASAP7_75t_R FILLER_0_75_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_354 ();
 DECAPx4_ASAP7_75t_R FILLER_0_75_363 ();
 FILLER_ASAP7_75t_R FILLER_0_75_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_385 ();
 FILLER_ASAP7_75t_R FILLER_0_75_392 ();
 DECAPx2_ASAP7_75t_R FILLER_0_75_402 ();
 FILLER_ASAP7_75t_R FILLER_0_75_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_410 ();
 FILLER_ASAP7_75t_R FILLER_0_75_417 ();
 FILLER_ASAP7_75t_R FILLER_0_75_425 ();
 FILLER_ASAP7_75t_R FILLER_0_75_435 ();
 DECAPx6_ASAP7_75t_R FILLER_0_75_442 ();
 FILLER_ASAP7_75t_R FILLER_0_75_456 ();
 FILLER_ASAP7_75t_R FILLER_0_75_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_466 ();
 FILLER_ASAP7_75t_R FILLER_0_75_470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_478 ();
 DECAPx6_ASAP7_75t_R FILLER_0_75_506 ();
 FILLER_ASAP7_75t_R FILLER_0_75_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_522 ();
 DECAPx1_ASAP7_75t_R FILLER_0_75_528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_75_538 ();
 FILLER_ASAP7_75t_R FILLER_0_75_544 ();
 DECAPx2_ASAP7_75t_R FILLER_0_75_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_562 ();
 FILLER_ASAP7_75t_R FILLER_0_75_569 ();
 FILLER_ASAP7_75t_R FILLER_0_75_577 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_579 ();
 FILLER_ASAP7_75t_R FILLER_0_75_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_588 ();
 DECAPx1_ASAP7_75t_R FILLER_0_75_595 ();
 DECAPx2_ASAP7_75t_R FILLER_0_75_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_608 ();
 FILLER_ASAP7_75t_R FILLER_0_75_615 ();
 DECAPx4_ASAP7_75t_R FILLER_0_75_624 ();
 FILLER_ASAP7_75t_R FILLER_0_75_634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_639 ();
 DECAPx4_ASAP7_75t_R FILLER_0_75_661 ();
 DECAPx6_ASAP7_75t_R FILLER_0_75_677 ();
 DECAPx2_ASAP7_75t_R FILLER_0_75_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_697 ();
 FILLER_ASAP7_75t_R FILLER_0_75_704 ();
 DECAPx2_ASAP7_75t_R FILLER_0_75_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_718 ();
 FILLER_ASAP7_75t_R FILLER_0_75_724 ();
 FILLER_ASAP7_75t_R FILLER_0_75_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_733 ();
 FILLER_ASAP7_75t_R FILLER_0_75_740 ();
 DECAPx2_ASAP7_75t_R FILLER_0_75_748 ();
 DECAPx4_ASAP7_75t_R FILLER_0_75_759 ();
 FILLER_ASAP7_75t_R FILLER_0_75_769 ();
 DECAPx1_ASAP7_75t_R FILLER_0_75_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_781 ();
 FILLER_ASAP7_75t_R FILLER_0_75_788 ();
 FILLER_ASAP7_75t_R FILLER_0_75_793 ();
 FILLER_ASAP7_75t_R FILLER_0_75_805 ();
 FILLER_ASAP7_75t_R FILLER_0_75_814 ();
 DECAPx2_ASAP7_75t_R FILLER_0_75_822 ();
 DECAPx1_ASAP7_75t_R FILLER_0_75_834 ();
 DECAPx2_ASAP7_75t_R FILLER_0_75_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_849 ();
 DECAPx1_ASAP7_75t_R FILLER_0_75_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_874 ();
 DECAPx2_ASAP7_75t_R FILLER_0_75_895 ();
 FILLER_ASAP7_75t_R FILLER_0_75_907 ();
 DECAPx1_ASAP7_75t_R FILLER_0_75_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_924 ();
 DECAPx6_ASAP7_75t_R FILLER_0_75_927 ();
 FILLER_ASAP7_75t_R FILLER_0_75_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_943 ();
 FILLER_ASAP7_75t_R FILLER_0_75_954 ();
 DECAPx1_ASAP7_75t_R FILLER_0_75_964 ();
 FILLER_ASAP7_75t_R FILLER_0_75_974 ();
 DECAPx1_ASAP7_75t_R FILLER_0_75_986 ();
 DECAPx6_ASAP7_75t_R FILLER_0_75_996 ();
 DECAPx2_ASAP7_75t_R FILLER_0_75_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_1016 ();
 DECAPx2_ASAP7_75t_R FILLER_0_75_1027 ();
 FILLER_ASAP7_75t_R FILLER_0_75_1033 ();
 FILLER_ASAP7_75t_R FILLER_0_75_1055 ();
 FILLER_ASAP7_75t_R FILLER_0_75_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_1065 ();
 FILLER_ASAP7_75t_R FILLER_0_75_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_1074 ();
 DECAPx1_ASAP7_75t_R FILLER_0_75_1081 ();
 FILLER_ASAP7_75t_R FILLER_0_75_1093 ();
 DECAPx1_ASAP7_75t_R FILLER_0_75_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_1106 ();
 DECAPx1_ASAP7_75t_R FILLER_0_75_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_1117 ();
 DECAPx1_ASAP7_75t_R FILLER_0_75_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_1128 ();
 DECAPx2_ASAP7_75t_R FILLER_0_75_1135 ();
 FILLER_ASAP7_75t_R FILLER_0_75_1141 ();
 FILLER_ASAP7_75t_R FILLER_0_75_1149 ();
 DECAPx4_ASAP7_75t_R FILLER_0_75_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_1167 ();
 DECAPx6_ASAP7_75t_R FILLER_0_75_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_1240 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_1262 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_1284 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_1306 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_1328 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_1350 ();
 DECAPx4_ASAP7_75t_R FILLER_0_75_1372 ();
 FILLER_ASAP7_75t_R FILLER_0_76_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_4 ();
 FILLER_ASAP7_75t_R FILLER_0_76_11 ();
 FILLER_ASAP7_75t_R FILLER_0_76_18 ();
 DECAPx2_ASAP7_75t_R FILLER_0_76_23 ();
 FILLER_ASAP7_75t_R FILLER_0_76_29 ();
 FILLER_ASAP7_75t_R FILLER_0_76_39 ();
 DECAPx1_ASAP7_75t_R FILLER_0_76_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_56 ();
 DECAPx4_ASAP7_75t_R FILLER_0_76_69 ();
 FILLER_ASAP7_75t_R FILLER_0_76_85 ();
 DECAPx1_ASAP7_75t_R FILLER_0_76_97 ();
 DECAPx2_ASAP7_75t_R FILLER_0_76_113 ();
 FILLER_ASAP7_75t_R FILLER_0_76_125 ();
 FILLER_ASAP7_75t_R FILLER_0_76_133 ();
 FILLER_ASAP7_75t_R FILLER_0_76_145 ();
 FILLER_ASAP7_75t_R FILLER_0_76_153 ();
 FILLER_ASAP7_75t_R FILLER_0_76_161 ();
 FILLER_ASAP7_75t_R FILLER_0_76_166 ();
 FILLER_ASAP7_75t_R FILLER_0_76_188 ();
 FILLER_ASAP7_75t_R FILLER_0_76_197 ();
 DECAPx4_ASAP7_75t_R FILLER_0_76_204 ();
 FILLER_ASAP7_75t_R FILLER_0_76_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_216 ();
 FILLER_ASAP7_75t_R FILLER_0_76_227 ();
 DECAPx2_ASAP7_75t_R FILLER_0_76_235 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_252 ();
 DECAPx2_ASAP7_75t_R FILLER_0_76_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_280 ();
 DECAPx1_ASAP7_75t_R FILLER_0_76_291 ();
 FILLER_ASAP7_75t_R FILLER_0_76_323 ();
 FILLER_ASAP7_75t_R FILLER_0_76_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_332 ();
 FILLER_ASAP7_75t_R FILLER_0_76_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_341 ();
 DECAPx2_ASAP7_75t_R FILLER_0_76_348 ();
 FILLER_ASAP7_75t_R FILLER_0_76_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_356 ();
 DECAPx4_ASAP7_75t_R FILLER_0_76_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_373 ();
 FILLER_ASAP7_75t_R FILLER_0_76_380 ();
 FILLER_ASAP7_75t_R FILLER_0_76_388 ();
 DECAPx4_ASAP7_75t_R FILLER_0_76_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_410 ();
 DECAPx1_ASAP7_75t_R FILLER_0_76_421 ();
 DECAPx2_ASAP7_75t_R FILLER_0_76_435 ();
 DECAPx6_ASAP7_75t_R FILLER_0_76_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_461 ();
 FILLER_ASAP7_75t_R FILLER_0_76_464 ();
 FILLER_ASAP7_75t_R FILLER_0_76_469 ();
 DECAPx6_ASAP7_75t_R FILLER_0_76_477 ();
 DECAPx1_ASAP7_75t_R FILLER_0_76_491 ();
 DECAPx4_ASAP7_75t_R FILLER_0_76_501 ();
 FILLER_ASAP7_75t_R FILLER_0_76_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_519 ();
 FILLER_ASAP7_75t_R FILLER_0_76_523 ();
 DECAPx4_ASAP7_75t_R FILLER_0_76_531 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_561 ();
 DECAPx6_ASAP7_75t_R FILLER_0_76_583 ();
 FILLER_ASAP7_75t_R FILLER_0_76_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_599 ();
 DECAPx2_ASAP7_75t_R FILLER_0_76_606 ();
 FILLER_ASAP7_75t_R FILLER_0_76_612 ();
 DECAPx2_ASAP7_75t_R FILLER_0_76_620 ();
 FILLER_ASAP7_75t_R FILLER_0_76_632 ();
 DECAPx2_ASAP7_75t_R FILLER_0_76_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_661 ();
 DECAPx1_ASAP7_75t_R FILLER_0_76_668 ();
 DECAPx2_ASAP7_75t_R FILLER_0_76_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_686 ();
 FILLER_ASAP7_75t_R FILLER_0_76_693 ();
 DECAPx2_ASAP7_75t_R FILLER_0_76_701 ();
 FILLER_ASAP7_75t_R FILLER_0_76_707 ();
 DECAPx1_ASAP7_75t_R FILLER_0_76_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_719 ();
 DECAPx6_ASAP7_75t_R FILLER_0_76_730 ();
 FILLER_ASAP7_75t_R FILLER_0_76_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_746 ();
 DECAPx6_ASAP7_75t_R FILLER_0_76_751 ();
 FILLER_ASAP7_75t_R FILLER_0_76_771 ();
 DECAPx4_ASAP7_75t_R FILLER_0_76_783 ();
 FILLER_ASAP7_75t_R FILLER_0_76_793 ();
 FILLER_ASAP7_75t_R FILLER_0_76_801 ();
 DECAPx2_ASAP7_75t_R FILLER_0_76_823 ();
 FILLER_ASAP7_75t_R FILLER_0_76_829 ();
 DECAPx4_ASAP7_75t_R FILLER_0_76_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_851 ();
 FILLER_ASAP7_75t_R FILLER_0_76_862 ();
 FILLER_ASAP7_75t_R FILLER_0_76_874 ();
 DECAPx1_ASAP7_75t_R FILLER_0_76_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_883 ();
 DECAPx2_ASAP7_75t_R FILLER_0_76_890 ();
 DECAPx4_ASAP7_75t_R FILLER_0_76_902 ();
 FILLER_ASAP7_75t_R FILLER_0_76_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_914 ();
 DECAPx6_ASAP7_75t_R FILLER_0_76_921 ();
 FILLER_ASAP7_75t_R FILLER_0_76_947 ();
 FILLER_ASAP7_75t_R FILLER_0_76_957 ();
 FILLER_ASAP7_75t_R FILLER_0_76_965 ();
 FILLER_ASAP7_75t_R FILLER_0_76_974 ();
 DECAPx4_ASAP7_75t_R FILLER_0_76_981 ();
 DECAPx2_ASAP7_75t_R FILLER_0_76_1002 ();
 FILLER_ASAP7_75t_R FILLER_0_76_1008 ();
 DECAPx2_ASAP7_75t_R FILLER_0_76_1016 ();
 DECAPx1_ASAP7_75t_R FILLER_0_76_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_1031 ();
 DECAPx2_ASAP7_75t_R FILLER_0_76_1037 ();
 FILLER_ASAP7_75t_R FILLER_0_76_1053 ();
 FILLER_ASAP7_75t_R FILLER_0_76_1060 ();
 FILLER_ASAP7_75t_R FILLER_0_76_1068 ();
 DECAPx1_ASAP7_75t_R FILLER_0_76_1080 ();
 FILLER_ASAP7_75t_R FILLER_0_76_1090 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_1092 ();
 DECAPx1_ASAP7_75t_R FILLER_0_76_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_1102 ();
 DECAPx1_ASAP7_75t_R FILLER_0_76_1123 ();
 FILLER_ASAP7_75t_R FILLER_0_76_1133 ();
 DECAPx4_ASAP7_75t_R FILLER_0_76_1141 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_1151 ();
 FILLER_ASAP7_75t_R FILLER_0_76_1158 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_1160 ();
 DECAPx6_ASAP7_75t_R FILLER_0_76_1169 ();
 FILLER_ASAP7_75t_R FILLER_0_76_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_1185 ();
 FILLER_ASAP7_75t_R FILLER_0_76_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_1244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_1266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_1332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_1354 ();
 DECAPx2_ASAP7_75t_R FILLER_0_76_1376 ();
 DECAPx2_ASAP7_75t_R FILLER_0_77_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_77_13 ();
 FILLER_ASAP7_75t_R FILLER_0_77_19 ();
 FILLER_ASAP7_75t_R FILLER_0_77_27 ();
 FILLER_ASAP7_75t_R FILLER_0_77_35 ();
 FILLER_ASAP7_75t_R FILLER_0_77_43 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_51 ();
 DECAPx2_ASAP7_75t_R FILLER_0_77_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_79 ();
 FILLER_ASAP7_75t_R FILLER_0_77_100 ();
 FILLER_ASAP7_75t_R FILLER_0_77_108 ();
 FILLER_ASAP7_75t_R FILLER_0_77_116 ();
 DECAPx2_ASAP7_75t_R FILLER_0_77_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_134 ();
 DECAPx1_ASAP7_75t_R FILLER_0_77_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_147 ();
 DECAPx1_ASAP7_75t_R FILLER_0_77_154 ();
 DECAPx1_ASAP7_75t_R FILLER_0_77_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_168 ();
 DECAPx2_ASAP7_75t_R FILLER_0_77_175 ();
 FILLER_ASAP7_75t_R FILLER_0_77_181 ();
 FILLER_ASAP7_75t_R FILLER_0_77_193 ();
 DECAPx2_ASAP7_75t_R FILLER_0_77_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_207 ();
 FILLER_ASAP7_75t_R FILLER_0_77_214 ();
 DECAPx1_ASAP7_75t_R FILLER_0_77_221 ();
 DECAPx2_ASAP7_75t_R FILLER_0_77_231 ();
 FILLER_ASAP7_75t_R FILLER_0_77_243 ();
 FILLER_ASAP7_75t_R FILLER_0_77_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_253 ();
 DECAPx6_ASAP7_75t_R FILLER_0_77_264 ();
 DECAPx1_ASAP7_75t_R FILLER_0_77_278 ();
 FILLER_ASAP7_75t_R FILLER_0_77_292 ();
 FILLER_ASAP7_75t_R FILLER_0_77_316 ();
 DECAPx1_ASAP7_75t_R FILLER_0_77_325 ();
 FILLER_ASAP7_75t_R FILLER_0_77_338 ();
 FILLER_ASAP7_75t_R FILLER_0_77_346 ();
 DECAPx2_ASAP7_75t_R FILLER_0_77_354 ();
 FILLER_ASAP7_75t_R FILLER_0_77_360 ();
 DECAPx4_ASAP7_75t_R FILLER_0_77_370 ();
 DECAPx2_ASAP7_75t_R FILLER_0_77_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_392 ();
 FILLER_ASAP7_75t_R FILLER_0_77_399 ();
 DECAPx6_ASAP7_75t_R FILLER_0_77_409 ();
 DECAPx1_ASAP7_75t_R FILLER_0_77_433 ();
 FILLER_ASAP7_75t_R FILLER_0_77_443 ();
 FILLER_ASAP7_75t_R FILLER_0_77_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_453 ();
 FILLER_ASAP7_75t_R FILLER_0_77_461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_470 ();
 DECAPx1_ASAP7_75t_R FILLER_0_77_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_496 ();
 FILLER_ASAP7_75t_R FILLER_0_77_504 ();
 DECAPx2_ASAP7_75t_R FILLER_0_77_512 ();
 FILLER_ASAP7_75t_R FILLER_0_77_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_520 ();
 DECAPx1_ASAP7_75t_R FILLER_0_77_527 ();
 FILLER_ASAP7_75t_R FILLER_0_77_537 ();
 DECAPx2_ASAP7_75t_R FILLER_0_77_545 ();
 FILLER_ASAP7_75t_R FILLER_0_77_551 ();
 DECAPx2_ASAP7_75t_R FILLER_0_77_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_565 ();
 DECAPx1_ASAP7_75t_R FILLER_0_77_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_576 ();
 DECAPx2_ASAP7_75t_R FILLER_0_77_583 ();
 DECAPx1_ASAP7_75t_R FILLER_0_77_595 ();
 FILLER_ASAP7_75t_R FILLER_0_77_607 ();
 DECAPx6_ASAP7_75t_R FILLER_0_77_619 ();
 FILLER_ASAP7_75t_R FILLER_0_77_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_635 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_639 ();
 DECAPx1_ASAP7_75t_R FILLER_0_77_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_665 ();
 DECAPx1_ASAP7_75t_R FILLER_0_77_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_676 ();
 FILLER_ASAP7_75t_R FILLER_0_77_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_685 ();
 FILLER_ASAP7_75t_R FILLER_0_77_692 ();
 DECAPx2_ASAP7_75t_R FILLER_0_77_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_705 ();
 DECAPx1_ASAP7_75t_R FILLER_0_77_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_716 ();
 FILLER_ASAP7_75t_R FILLER_0_77_728 ();
 FILLER_ASAP7_75t_R FILLER_0_77_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_738 ();
 FILLER_ASAP7_75t_R FILLER_0_77_745 ();
 DECAPx6_ASAP7_75t_R FILLER_0_77_758 ();
 DECAPx1_ASAP7_75t_R FILLER_0_77_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_781 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_789 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_811 ();
 FILLER_ASAP7_75t_R FILLER_0_77_833 ();
 FILLER_ASAP7_75t_R FILLER_0_77_841 ();
 FILLER_ASAP7_75t_R FILLER_0_77_849 ();
 FILLER_ASAP7_75t_R FILLER_0_77_871 ();
 DECAPx1_ASAP7_75t_R FILLER_0_77_879 ();
 FILLER_ASAP7_75t_R FILLER_0_77_893 ();
 DECAPx4_ASAP7_75t_R FILLER_0_77_901 ();
 FILLER_ASAP7_75t_R FILLER_0_77_911 ();
 DECAPx2_ASAP7_75t_R FILLER_0_77_919 ();
 DECAPx6_ASAP7_75t_R FILLER_0_77_927 ();
 DECAPx1_ASAP7_75t_R FILLER_0_77_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_945 ();
 DECAPx1_ASAP7_75t_R FILLER_0_77_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_955 ();
 FILLER_ASAP7_75t_R FILLER_0_77_966 ();
 DECAPx2_ASAP7_75t_R FILLER_0_77_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_980 ();
 FILLER_ASAP7_75t_R FILLER_0_77_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_995 ();
 DECAPx2_ASAP7_75t_R FILLER_0_77_999 ();
 FILLER_ASAP7_75t_R FILLER_0_77_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_1007 ();
 FILLER_ASAP7_75t_R FILLER_0_77_1018 ();
 FILLER_ASAP7_75t_R FILLER_0_77_1030 ();
 FILLER_ASAP7_75t_R FILLER_0_77_1042 ();
 FILLER_ASAP7_75t_R FILLER_0_77_1054 ();
 FILLER_ASAP7_75t_R FILLER_0_77_1066 ();
 DECAPx2_ASAP7_75t_R FILLER_0_77_1076 ();
 DECAPx4_ASAP7_75t_R FILLER_0_77_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_1098 ();
 FILLER_ASAP7_75t_R FILLER_0_77_1104 ();
 DECAPx2_ASAP7_75t_R FILLER_0_77_1112 ();
 FILLER_ASAP7_75t_R FILLER_0_77_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_1120 ();
 DECAPx1_ASAP7_75t_R FILLER_0_77_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_1131 ();
 DECAPx6_ASAP7_75t_R FILLER_0_77_1137 ();
 DECAPx2_ASAP7_75t_R FILLER_0_77_1159 ();
 FILLER_ASAP7_75t_R FILLER_0_77_1165 ();
 FILLER_ASAP7_75t_R FILLER_0_77_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_1240 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_1262 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_1284 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_1306 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_1328 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_1350 ();
 DECAPx4_ASAP7_75t_R FILLER_0_77_1372 ();
 FILLER_ASAP7_75t_R FILLER_0_78_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_78_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_19 ();
 FILLER_ASAP7_75t_R FILLER_0_78_30 ();
 FILLER_ASAP7_75t_R FILLER_0_78_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_37 ();
 FILLER_ASAP7_75t_R FILLER_0_78_48 ();
 DECAPx4_ASAP7_75t_R FILLER_0_78_56 ();
 FILLER_ASAP7_75t_R FILLER_0_78_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_68 ();
 FILLER_ASAP7_75t_R FILLER_0_78_77 ();
 DECAPx1_ASAP7_75t_R FILLER_0_78_85 ();
 DECAPx1_ASAP7_75t_R FILLER_0_78_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_103 ();
 DECAPx2_ASAP7_75t_R FILLER_0_78_112 ();
 FILLER_ASAP7_75t_R FILLER_0_78_128 ();
 FILLER_ASAP7_75t_R FILLER_0_78_140 ();
 FILLER_ASAP7_75t_R FILLER_0_78_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_150 ();
 FILLER_ASAP7_75t_R FILLER_0_78_157 ();
 FILLER_ASAP7_75t_R FILLER_0_78_165 ();
 FILLER_ASAP7_75t_R FILLER_0_78_177 ();
 FILLER_ASAP7_75t_R FILLER_0_78_199 ();
 FILLER_ASAP7_75t_R FILLER_0_78_207 ();
 FILLER_ASAP7_75t_R FILLER_0_78_215 ();
 FILLER_ASAP7_75t_R FILLER_0_78_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_225 ();
 DECAPx2_ASAP7_75t_R FILLER_0_78_236 ();
 FILLER_ASAP7_75t_R FILLER_0_78_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_244 ();
 FILLER_ASAP7_75t_R FILLER_0_78_251 ();
 FILLER_ASAP7_75t_R FILLER_0_78_256 ();
 DECAPx6_ASAP7_75t_R FILLER_0_78_264 ();
 DECAPx1_ASAP7_75t_R FILLER_0_78_278 ();
 FILLER_ASAP7_75t_R FILLER_0_78_292 ();
 DECAPx2_ASAP7_75t_R FILLER_0_78_304 ();
 FILLER_ASAP7_75t_R FILLER_0_78_310 ();
 FILLER_ASAP7_75t_R FILLER_0_78_318 ();
 FILLER_ASAP7_75t_R FILLER_0_78_328 ();
 DECAPx4_ASAP7_75t_R FILLER_0_78_340 ();
 DECAPx6_ASAP7_75t_R FILLER_0_78_356 ();
 FILLER_ASAP7_75t_R FILLER_0_78_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_372 ();
 DECAPx4_ASAP7_75t_R FILLER_0_78_383 ();
 FILLER_ASAP7_75t_R FILLER_0_78_397 ();
 DECAPx1_ASAP7_75t_R FILLER_0_78_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_413 ();
 DECAPx2_ASAP7_75t_R FILLER_0_78_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_427 ();
 DECAPx1_ASAP7_75t_R FILLER_0_78_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_442 ();
 FILLER_ASAP7_75t_R FILLER_0_78_449 ();
 FILLER_ASAP7_75t_R FILLER_0_78_454 ();
 FILLER_ASAP7_75t_R FILLER_0_78_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_461 ();
 DECAPx1_ASAP7_75t_R FILLER_0_78_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_474 ();
 DECAPx6_ASAP7_75t_R FILLER_0_78_502 ();
 DECAPx2_ASAP7_75t_R FILLER_0_78_516 ();
 DECAPx1_ASAP7_75t_R FILLER_0_78_530 ();
 FILLER_ASAP7_75t_R FILLER_0_78_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_78_549 ();
 FILLER_ASAP7_75t_R FILLER_0_78_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_561 ();
 FILLER_ASAP7_75t_R FILLER_0_78_570 ();
 FILLER_ASAP7_75t_R FILLER_0_78_578 ();
 DECAPx1_ASAP7_75t_R FILLER_0_78_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_587 ();
 DECAPx4_ASAP7_75t_R FILLER_0_78_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_610 ();
 FILLER_ASAP7_75t_R FILLER_0_78_617 ();
 FILLER_ASAP7_75t_R FILLER_0_78_625 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_633 ();
 DECAPx2_ASAP7_75t_R FILLER_0_78_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_661 ();
 FILLER_ASAP7_75t_R FILLER_0_78_668 ();
 DECAPx1_ASAP7_75t_R FILLER_0_78_676 ();
 FILLER_ASAP7_75t_R FILLER_0_78_686 ();
 DECAPx6_ASAP7_75t_R FILLER_0_78_694 ();
 FILLER_ASAP7_75t_R FILLER_0_78_714 ();
 FILLER_ASAP7_75t_R FILLER_0_78_721 ();
 DECAPx4_ASAP7_75t_R FILLER_0_78_730 ();
 FILLER_ASAP7_75t_R FILLER_0_78_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_742 ();
 DECAPx2_ASAP7_75t_R FILLER_0_78_749 ();
 FILLER_ASAP7_75t_R FILLER_0_78_755 ();
 DECAPx1_ASAP7_75t_R FILLER_0_78_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_767 ();
 DECAPx1_ASAP7_75t_R FILLER_0_78_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_782 ();
 DECAPx2_ASAP7_75t_R FILLER_0_78_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_799 ();
 DECAPx2_ASAP7_75t_R FILLER_0_78_820 ();
 FILLER_ASAP7_75t_R FILLER_0_78_826 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_835 ();
 DECAPx4_ASAP7_75t_R FILLER_0_78_857 ();
 FILLER_ASAP7_75t_R FILLER_0_78_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_869 ();
 DECAPx6_ASAP7_75t_R FILLER_0_78_882 ();
 FILLER_ASAP7_75t_R FILLER_0_78_896 ();
 FILLER_ASAP7_75t_R FILLER_0_78_904 ();
 FILLER_ASAP7_75t_R FILLER_0_78_912 ();
 FILLER_ASAP7_75t_R FILLER_0_78_920 ();
 DECAPx4_ASAP7_75t_R FILLER_0_78_928 ();
 FILLER_ASAP7_75t_R FILLER_0_78_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_940 ();
 FILLER_ASAP7_75t_R FILLER_0_78_951 ();
 DECAPx2_ASAP7_75t_R FILLER_0_78_959 ();
 FILLER_ASAP7_75t_R FILLER_0_78_973 ();
 DECAPx6_ASAP7_75t_R FILLER_0_78_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_994 ();
 DECAPx1_ASAP7_75t_R FILLER_0_78_1006 ();
 DECAPx2_ASAP7_75t_R FILLER_0_78_1020 ();
 FILLER_ASAP7_75t_R FILLER_0_78_1036 ();
 FILLER_ASAP7_75t_R FILLER_0_78_1048 ();
 DECAPx1_ASAP7_75t_R FILLER_0_78_1056 ();
 DECAPx1_ASAP7_75t_R FILLER_0_78_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_1074 ();
 FILLER_ASAP7_75t_R FILLER_0_78_1080 ();
 FILLER_ASAP7_75t_R FILLER_0_78_1087 ();
 FILLER_ASAP7_75t_R FILLER_0_78_1095 ();
 DECAPx2_ASAP7_75t_R FILLER_0_78_1103 ();
 FILLER_ASAP7_75t_R FILLER_0_78_1109 ();
 DECAPx1_ASAP7_75t_R FILLER_0_78_1121 ();
 FILLER_ASAP7_75t_R FILLER_0_78_1131 ();
 DECAPx1_ASAP7_75t_R FILLER_0_78_1138 ();
 FILLER_ASAP7_75t_R FILLER_0_78_1148 ();
 DECAPx2_ASAP7_75t_R FILLER_0_78_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_1162 ();
 DECAPx6_ASAP7_75t_R FILLER_0_78_1169 ();
 DECAPx1_ASAP7_75t_R FILLER_0_78_1183 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_1259 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_1281 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_1303 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_1325 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_1347 ();
 DECAPx4_ASAP7_75t_R FILLER_0_78_1369 ();
 FILLER_ASAP7_75t_R FILLER_0_78_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_79_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_9 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_26 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_33 ();
 FILLER_ASAP7_75t_R FILLER_0_79_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_41 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_53 ();
 DECAPx4_ASAP7_75t_R FILLER_0_79_71 ();
 DECAPx1_ASAP7_75t_R FILLER_0_79_87 ();
 FILLER_ASAP7_75t_R FILLER_0_79_97 ();
 FILLER_ASAP7_75t_R FILLER_0_79_106 ();
 FILLER_ASAP7_75t_R FILLER_0_79_118 ();
 FILLER_ASAP7_75t_R FILLER_0_79_130 ();
 FILLER_ASAP7_75t_R FILLER_0_79_142 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_158 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_171 ();
 FILLER_ASAP7_75t_R FILLER_0_79_177 ();
 DECAPx4_ASAP7_75t_R FILLER_0_79_187 ();
 FILLER_ASAP7_75t_R FILLER_0_79_209 ();
 DECAPx1_ASAP7_75t_R FILLER_0_79_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_221 ();
 FILLER_ASAP7_75t_R FILLER_0_79_230 ();
 FILLER_ASAP7_75t_R FILLER_0_79_238 ();
 FILLER_ASAP7_75t_R FILLER_0_79_246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_254 ();
 FILLER_ASAP7_75t_R FILLER_0_79_276 ();
 FILLER_ASAP7_75t_R FILLER_0_79_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_290 ();
 FILLER_ASAP7_75t_R FILLER_0_79_300 ();
 DECAPx4_ASAP7_75t_R FILLER_0_79_307 ();
 FILLER_ASAP7_75t_R FILLER_0_79_321 ();
 DECAPx1_ASAP7_75t_R FILLER_0_79_327 ();
 DECAPx1_ASAP7_75t_R FILLER_0_79_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_345 ();
 FILLER_ASAP7_75t_R FILLER_0_79_354 ();
 FILLER_ASAP7_75t_R FILLER_0_79_362 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_377 ();
 FILLER_ASAP7_75t_R FILLER_0_79_383 ();
 DECAPx1_ASAP7_75t_R FILLER_0_79_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_399 ();
 FILLER_ASAP7_75t_R FILLER_0_79_403 ();
 FILLER_ASAP7_75t_R FILLER_0_79_427 ();
 FILLER_ASAP7_75t_R FILLER_0_79_453 ();
 FILLER_ASAP7_75t_R FILLER_0_79_458 ();
 DECAPx6_ASAP7_75t_R FILLER_0_79_466 ();
 FILLER_ASAP7_75t_R FILLER_0_79_480 ();
 FILLER_ASAP7_75t_R FILLER_0_79_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_490 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_497 ();
 FILLER_ASAP7_75t_R FILLER_0_79_510 ();
 FILLER_ASAP7_75t_R FILLER_0_79_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_517 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_529 ();
 FILLER_ASAP7_75t_R FILLER_0_79_535 ();
 FILLER_ASAP7_75t_R FILLER_0_79_547 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_556 ();
 DECAPx4_ASAP7_75t_R FILLER_0_79_568 ();
 FILLER_ASAP7_75t_R FILLER_0_79_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_580 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_598 ();
 FILLER_ASAP7_75t_R FILLER_0_79_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_622 ();
 FILLER_ASAP7_75t_R FILLER_0_79_629 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_637 ();
 DECAPx6_ASAP7_75t_R FILLER_0_79_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_673 ();
 FILLER_ASAP7_75t_R FILLER_0_79_680 ();
 DECAPx6_ASAP7_75t_R FILLER_0_79_688 ();
 FILLER_ASAP7_75t_R FILLER_0_79_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_704 ();
 DECAPx1_ASAP7_75t_R FILLER_0_79_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_715 ();
 FILLER_ASAP7_75t_R FILLER_0_79_722 ();
 FILLER_ASAP7_75t_R FILLER_0_79_734 ();
 DECAPx1_ASAP7_75t_R FILLER_0_79_739 ();
 DECAPx4_ASAP7_75t_R FILLER_0_79_751 ();
 FILLER_ASAP7_75t_R FILLER_0_79_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_763 ();
 FILLER_ASAP7_75t_R FILLER_0_79_784 ();
 FILLER_ASAP7_75t_R FILLER_0_79_792 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_808 ();
 FILLER_ASAP7_75t_R FILLER_0_79_815 ();
 FILLER_ASAP7_75t_R FILLER_0_79_823 ();
 FILLER_ASAP7_75t_R FILLER_0_79_831 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_839 ();
 DECAPx1_ASAP7_75t_R FILLER_0_79_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_865 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_872 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_884 ();
 FILLER_ASAP7_75t_R FILLER_0_79_890 ();
 FILLER_ASAP7_75t_R FILLER_0_79_897 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_911 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_919 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_927 ();
 FILLER_ASAP7_75t_R FILLER_0_79_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_935 ();
 FILLER_ASAP7_75t_R FILLER_0_79_941 ();
 DECAPx1_ASAP7_75t_R FILLER_0_79_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_967 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_974 ();
 DECAPx6_ASAP7_75t_R FILLER_0_79_996 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_1016 ();
 FILLER_ASAP7_75t_R FILLER_0_79_1023 ();
 FILLER_ASAP7_75t_R FILLER_0_79_1030 ();
 FILLER_ASAP7_75t_R FILLER_0_79_1042 ();
 FILLER_ASAP7_75t_R FILLER_0_79_1056 ();
 FILLER_ASAP7_75t_R FILLER_0_79_1063 ();
 FILLER_ASAP7_75t_R FILLER_0_79_1073 ();
 DECAPx1_ASAP7_75t_R FILLER_0_79_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_1084 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_1091 ();
 FILLER_ASAP7_75t_R FILLER_0_79_1097 ();
 FILLER_ASAP7_75t_R FILLER_0_79_1105 ();
 FILLER_ASAP7_75t_R FILLER_0_79_1119 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_1127 ();
 FILLER_ASAP7_75t_R FILLER_0_79_1133 ();
 DECAPx6_ASAP7_75t_R FILLER_0_79_1155 ();
 FILLER_ASAP7_75t_R FILLER_0_79_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_1171 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_1219 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_1263 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_1285 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_1307 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_1351 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_79_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_1381 ();
 DECAPx6_ASAP7_75t_R FILLER_0_80_2 ();
 FILLER_ASAP7_75t_R FILLER_0_80_16 ();
 FILLER_ASAP7_75t_R FILLER_0_80_21 ();
 FILLER_ASAP7_75t_R FILLER_0_80_43 ();
 DECAPx2_ASAP7_75t_R FILLER_0_80_51 ();
 FILLER_ASAP7_75t_R FILLER_0_80_77 ();
 DECAPx1_ASAP7_75t_R FILLER_0_80_89 ();
 FILLER_ASAP7_75t_R FILLER_0_80_98 ();
 FILLER_ASAP7_75t_R FILLER_0_80_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_110 ();
 FILLER_ASAP7_75t_R FILLER_0_80_135 ();
 FILLER_ASAP7_75t_R FILLER_0_80_143 ();
 FILLER_ASAP7_75t_R FILLER_0_80_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_153 ();
 DECAPx2_ASAP7_75t_R FILLER_0_80_164 ();
 FILLER_ASAP7_75t_R FILLER_0_80_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_172 ();
 FILLER_ASAP7_75t_R FILLER_0_80_183 ();
 DECAPx4_ASAP7_75t_R FILLER_0_80_193 ();
 FILLER_ASAP7_75t_R FILLER_0_80_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_205 ();
 FILLER_ASAP7_75t_R FILLER_0_80_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_215 ();
 FILLER_ASAP7_75t_R FILLER_0_80_226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_238 ();
 DECAPx2_ASAP7_75t_R FILLER_0_80_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_266 ();
 DECAPx1_ASAP7_75t_R FILLER_0_80_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_274 ();
 FILLER_ASAP7_75t_R FILLER_0_80_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_283 ();
 DECAPx1_ASAP7_75t_R FILLER_0_80_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_294 ();
 FILLER_ASAP7_75t_R FILLER_0_80_298 ();
 FILLER_ASAP7_75t_R FILLER_0_80_306 ();
 FILLER_ASAP7_75t_R FILLER_0_80_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_313 ();
 FILLER_ASAP7_75t_R FILLER_0_80_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_321 ();
 DECAPx2_ASAP7_75t_R FILLER_0_80_328 ();
 FILLER_ASAP7_75t_R FILLER_0_80_337 ();
 FILLER_ASAP7_75t_R FILLER_0_80_354 ();
 FILLER_ASAP7_75t_R FILLER_0_80_364 ();
 FILLER_ASAP7_75t_R FILLER_0_80_372 ();
 FILLER_ASAP7_75t_R FILLER_0_80_380 ();
 FILLER_ASAP7_75t_R FILLER_0_80_389 ();
 DECAPx2_ASAP7_75t_R FILLER_0_80_396 ();
 DECAPx1_ASAP7_75t_R FILLER_0_80_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_413 ();
 DECAPx2_ASAP7_75t_R FILLER_0_80_420 ();
 FILLER_ASAP7_75t_R FILLER_0_80_426 ();
 DECAPx2_ASAP7_75t_R FILLER_0_80_438 ();
 DECAPx2_ASAP7_75t_R FILLER_0_80_456 ();
 DECAPx6_ASAP7_75t_R FILLER_0_80_464 ();
 DECAPx2_ASAP7_75t_R FILLER_0_80_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_484 ();
 FILLER_ASAP7_75t_R FILLER_0_80_488 ();
 DECAPx6_ASAP7_75t_R FILLER_0_80_496 ();
 DECAPx2_ASAP7_75t_R FILLER_0_80_510 ();
 DECAPx6_ASAP7_75t_R FILLER_0_80_522 ();
 DECAPx1_ASAP7_75t_R FILLER_0_80_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_540 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_547 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_591 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_642 ();
 DECAPx4_ASAP7_75t_R FILLER_0_80_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_674 ();
 FILLER_ASAP7_75t_R FILLER_0_80_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_682 ();
 DECAPx2_ASAP7_75t_R FILLER_0_80_689 ();
 FILLER_ASAP7_75t_R FILLER_0_80_700 ();
 FILLER_ASAP7_75t_R FILLER_0_80_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_709 ();
 FILLER_ASAP7_75t_R FILLER_0_80_715 ();
 DECAPx2_ASAP7_75t_R FILLER_0_80_723 ();
 FILLER_ASAP7_75t_R FILLER_0_80_729 ();
 FILLER_ASAP7_75t_R FILLER_0_80_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_740 ();
 DECAPx1_ASAP7_75t_R FILLER_0_80_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_751 ();
 DECAPx2_ASAP7_75t_R FILLER_0_80_759 ();
 FILLER_ASAP7_75t_R FILLER_0_80_765 ();
 DECAPx1_ASAP7_75t_R FILLER_0_80_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_781 ();
 FILLER_ASAP7_75t_R FILLER_0_80_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_790 ();
 DECAPx6_ASAP7_75t_R FILLER_0_80_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_812 ();
 DECAPx1_ASAP7_75t_R FILLER_0_80_819 ();
 FILLER_ASAP7_75t_R FILLER_0_80_829 ();
 DECAPx2_ASAP7_75t_R FILLER_0_80_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_843 ();
 FILLER_ASAP7_75t_R FILLER_0_80_850 ();
 DECAPx2_ASAP7_75t_R FILLER_0_80_858 ();
 DECAPx4_ASAP7_75t_R FILLER_0_80_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_885 ();
 FILLER_ASAP7_75t_R FILLER_0_80_893 ();
 DECAPx2_ASAP7_75t_R FILLER_0_80_906 ();
 FILLER_ASAP7_75t_R FILLER_0_80_912 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_920 ();
 DECAPx1_ASAP7_75t_R FILLER_0_80_942 ();
 FILLER_ASAP7_75t_R FILLER_0_80_958 ();
 FILLER_ASAP7_75t_R FILLER_0_80_966 ();
 FILLER_ASAP7_75t_R FILLER_0_80_978 ();
 DECAPx1_ASAP7_75t_R FILLER_0_80_985 ();
 DECAPx2_ASAP7_75t_R FILLER_0_80_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_1001 ();
 FILLER_ASAP7_75t_R FILLER_0_80_1012 ();
 DECAPx2_ASAP7_75t_R FILLER_0_80_1021 ();
 FILLER_ASAP7_75t_R FILLER_0_80_1027 ();
 FILLER_ASAP7_75t_R FILLER_0_80_1039 ();
 FILLER_ASAP7_75t_R FILLER_0_80_1051 ();
 FILLER_ASAP7_75t_R FILLER_0_80_1058 ();
 FILLER_ASAP7_75t_R FILLER_0_80_1065 ();
 FILLER_ASAP7_75t_R FILLER_0_80_1077 ();
 DECAPx1_ASAP7_75t_R FILLER_0_80_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_0_80_1100 ();
 DECAPx2_ASAP7_75t_R FILLER_0_80_1124 ();
 FILLER_ASAP7_75t_R FILLER_0_80_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_1140 ();
 DECAPx4_ASAP7_75t_R FILLER_0_80_1153 ();
 FILLER_ASAP7_75t_R FILLER_0_80_1163 ();
 DECAPx1_ASAP7_75t_R FILLER_0_80_1171 ();
 FILLER_ASAP7_75t_R FILLER_0_80_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_1180 ();
 DECAPx2_ASAP7_75t_R FILLER_0_80_1187 ();
 FILLER_ASAP7_75t_R FILLER_0_80_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_1206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_1338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_1360 ();
 DECAPx1_ASAP7_75t_R FILLER_0_81_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_28 ();
 DECAPx1_ASAP7_75t_R FILLER_0_81_40 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_54 ();
 DECAPx1_ASAP7_75t_R FILLER_0_81_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_80 ();
 FILLER_ASAP7_75t_R FILLER_0_81_88 ();
 DECAPx1_ASAP7_75t_R FILLER_0_81_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_100 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_114 ();
 FILLER_ASAP7_75t_R FILLER_0_81_121 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_133 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_145 ();
 FILLER_ASAP7_75t_R FILLER_0_81_157 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_179 ();
 FILLER_ASAP7_75t_R FILLER_0_81_187 ();
 DECAPx4_ASAP7_75t_R FILLER_0_81_201 ();
 FILLER_ASAP7_75t_R FILLER_0_81_211 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_219 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_241 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_257 ();
 FILLER_ASAP7_75t_R FILLER_0_81_263 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_277 ();
 DECAPx6_ASAP7_75t_R FILLER_0_81_284 ();
 FILLER_ASAP7_75t_R FILLER_0_81_298 ();
 DECAPx1_ASAP7_75t_R FILLER_0_81_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_310 ();
 DECAPx4_ASAP7_75t_R FILLER_0_81_317 ();
 FILLER_ASAP7_75t_R FILLER_0_81_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_329 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_340 ();
 FILLER_ASAP7_75t_R FILLER_0_81_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_348 ();
 FILLER_ASAP7_75t_R FILLER_0_81_359 ();
 DECAPx4_ASAP7_75t_R FILLER_0_81_367 ();
 FILLER_ASAP7_75t_R FILLER_0_81_377 ();
 FILLER_ASAP7_75t_R FILLER_0_81_386 ();
 FILLER_ASAP7_75t_R FILLER_0_81_396 ();
 FILLER_ASAP7_75t_R FILLER_0_81_406 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_414 ();
 FILLER_ASAP7_75t_R FILLER_0_81_420 ();
 FILLER_ASAP7_75t_R FILLER_0_81_427 ();
 FILLER_ASAP7_75t_R FILLER_0_81_434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_468 ();
 FILLER_ASAP7_75t_R FILLER_0_81_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_492 ();
 FILLER_ASAP7_75t_R FILLER_0_81_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_502 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_519 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_532 ();
 FILLER_ASAP7_75t_R FILLER_0_81_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_545 ();
 FILLER_ASAP7_75t_R FILLER_0_81_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_554 ();
 FILLER_ASAP7_75t_R FILLER_0_81_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_563 ();
 FILLER_ASAP7_75t_R FILLER_0_81_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_588 ();
 DECAPx1_ASAP7_75t_R FILLER_0_81_600 ();
 FILLER_ASAP7_75t_R FILLER_0_81_610 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_617 ();
 FILLER_ASAP7_75t_R FILLER_0_81_629 ();
 FILLER_ASAP7_75t_R FILLER_0_81_637 ();
 DECAPx6_ASAP7_75t_R FILLER_0_81_645 ();
 FILLER_ASAP7_75t_R FILLER_0_81_659 ();
 FILLER_ASAP7_75t_R FILLER_0_81_667 ();
 FILLER_ASAP7_75t_R FILLER_0_81_675 ();
 FILLER_ASAP7_75t_R FILLER_0_81_683 ();
 FILLER_ASAP7_75t_R FILLER_0_81_691 ();
 DECAPx1_ASAP7_75t_R FILLER_0_81_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_703 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_714 ();
 FILLER_ASAP7_75t_R FILLER_0_81_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_730 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_739 ();
 FILLER_ASAP7_75t_R FILLER_0_81_745 ();
 DECAPx6_ASAP7_75t_R FILLER_0_81_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_781 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_788 ();
 DECAPx6_ASAP7_75t_R FILLER_0_81_810 ();
 DECAPx4_ASAP7_75t_R FILLER_0_81_834 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_850 ();
 FILLER_ASAP7_75t_R FILLER_0_81_856 ();
 FILLER_ASAP7_75t_R FILLER_0_81_868 ();
 FILLER_ASAP7_75t_R FILLER_0_81_877 ();
 FILLER_ASAP7_75t_R FILLER_0_81_885 ();
 DECAPx6_ASAP7_75t_R FILLER_0_81_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_908 ();
 FILLER_ASAP7_75t_R FILLER_0_81_915 ();
 FILLER_ASAP7_75t_R FILLER_0_81_923 ();
 DECAPx6_ASAP7_75t_R FILLER_0_81_927 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_941 ();
 FILLER_ASAP7_75t_R FILLER_0_81_950 ();
 FILLER_ASAP7_75t_R FILLER_0_81_957 ();
 FILLER_ASAP7_75t_R FILLER_0_81_967 ();
 FILLER_ASAP7_75t_R FILLER_0_81_975 ();
 FILLER_ASAP7_75t_R FILLER_0_81_983 ();
 FILLER_ASAP7_75t_R FILLER_0_81_991 ();
 FILLER_ASAP7_75t_R FILLER_0_81_999 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_1001 ();
 FILLER_ASAP7_75t_R FILLER_0_81_1012 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_1020 ();
 FILLER_ASAP7_75t_R FILLER_0_81_1034 ();
 FILLER_ASAP7_75t_R FILLER_0_81_1046 ();
 DECAPx1_ASAP7_75t_R FILLER_0_81_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_1062 ();
 FILLER_ASAP7_75t_R FILLER_0_81_1071 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_1083 ();
 FILLER_ASAP7_75t_R FILLER_0_81_1089 ();
 DECAPx6_ASAP7_75t_R FILLER_0_81_1098 ();
 FILLER_ASAP7_75t_R FILLER_0_81_1115 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_1128 ();
 FILLER_ASAP7_75t_R FILLER_0_81_1135 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_1153 ();
 FILLER_ASAP7_75t_R FILLER_0_81_1160 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_1172 ();
 FILLER_ASAP7_75t_R FILLER_0_81_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_1180 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_1192 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_1198 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_1227 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_1293 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_1315 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_1337 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_1359 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_82_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_13 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_29 ();
 FILLER_ASAP7_75t_R FILLER_0_82_41 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_49 ();
 DECAPx2_ASAP7_75t_R FILLER_0_82_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_77 ();
 DECAPx6_ASAP7_75t_R FILLER_0_82_84 ();
 FILLER_ASAP7_75t_R FILLER_0_82_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_106 ();
 FILLER_ASAP7_75t_R FILLER_0_82_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_115 ();
 FILLER_ASAP7_75t_R FILLER_0_82_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_128 ();
 FILLER_ASAP7_75t_R FILLER_0_82_139 ();
 DECAPx2_ASAP7_75t_R FILLER_0_82_147 ();
 FILLER_ASAP7_75t_R FILLER_0_82_153 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_166 ();
 FILLER_ASAP7_75t_R FILLER_0_82_170 ();
 FILLER_ASAP7_75t_R FILLER_0_82_178 ();
 FILLER_ASAP7_75t_R FILLER_0_82_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_190 ();
 DECAPx6_ASAP7_75t_R FILLER_0_82_201 ();
 FILLER_ASAP7_75t_R FILLER_0_82_215 ();
 FILLER_ASAP7_75t_R FILLER_0_82_237 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_250 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_261 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_272 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_284 ();
 FILLER_ASAP7_75t_R FILLER_0_82_308 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_321 ();
 DECAPx4_ASAP7_75t_R FILLER_0_82_343 ();
 DECAPx2_ASAP7_75t_R FILLER_0_82_358 ();
 FILLER_ASAP7_75t_R FILLER_0_82_364 ();
 DECAPx4_ASAP7_75t_R FILLER_0_82_373 ();
 FILLER_ASAP7_75t_R FILLER_0_82_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_385 ();
 DECAPx6_ASAP7_75t_R FILLER_0_82_392 ();
 FILLER_ASAP7_75t_R FILLER_0_82_412 ();
 FILLER_ASAP7_75t_R FILLER_0_82_421 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_433 ();
 DECAPx2_ASAP7_75t_R FILLER_0_82_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_461 ();
 DECAPx4_ASAP7_75t_R FILLER_0_82_464 ();
 FILLER_ASAP7_75t_R FILLER_0_82_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_476 ();
 DECAPx4_ASAP7_75t_R FILLER_0_82_483 ();
 FILLER_ASAP7_75t_R FILLER_0_82_513 ();
 FILLER_ASAP7_75t_R FILLER_0_82_525 ();
 DECAPx2_ASAP7_75t_R FILLER_0_82_547 ();
 DECAPx2_ASAP7_75t_R FILLER_0_82_563 ();
 FILLER_ASAP7_75t_R FILLER_0_82_569 ();
 FILLER_ASAP7_75t_R FILLER_0_82_577 ();
 FILLER_ASAP7_75t_R FILLER_0_82_590 ();
 DECAPx2_ASAP7_75t_R FILLER_0_82_598 ();
 FILLER_ASAP7_75t_R FILLER_0_82_604 ();
 FILLER_ASAP7_75t_R FILLER_0_82_617 ();
 DECAPx2_ASAP7_75t_R FILLER_0_82_625 ();
 FILLER_ASAP7_75t_R FILLER_0_82_631 ();
 FILLER_ASAP7_75t_R FILLER_0_82_639 ();
 DECAPx6_ASAP7_75t_R FILLER_0_82_647 ();
 FILLER_ASAP7_75t_R FILLER_0_82_661 ();
 DECAPx2_ASAP7_75t_R FILLER_0_82_674 ();
 FILLER_ASAP7_75t_R FILLER_0_82_680 ();
 FILLER_ASAP7_75t_R FILLER_0_82_690 ();
 FILLER_ASAP7_75t_R FILLER_0_82_698 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_710 ();
 FILLER_ASAP7_75t_R FILLER_0_82_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_722 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_729 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_739 ();
 DECAPx2_ASAP7_75t_R FILLER_0_82_749 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_761 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_776 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_791 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_806 ();
 FILLER_ASAP7_75t_R FILLER_0_82_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_817 ();
 DECAPx6_ASAP7_75t_R FILLER_0_82_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_841 ();
 DECAPx4_ASAP7_75t_R FILLER_0_82_848 ();
 FILLER_ASAP7_75t_R FILLER_0_82_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_860 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_873 ();
 FILLER_ASAP7_75t_R FILLER_0_82_883 ();
 DECAPx2_ASAP7_75t_R FILLER_0_82_891 ();
 FILLER_ASAP7_75t_R FILLER_0_82_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_899 ();
 FILLER_ASAP7_75t_R FILLER_0_82_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_915 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_937 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_941 ();
 DECAPx2_ASAP7_75t_R FILLER_0_82_948 ();
 DECAPx2_ASAP7_75t_R FILLER_0_82_974 ();
 FILLER_ASAP7_75t_R FILLER_0_82_986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_82_994 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_1000 ();
 FILLER_ASAP7_75t_R FILLER_0_82_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_1013 ();
 FILLER_ASAP7_75t_R FILLER_0_82_1021 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_1029 ();
 FILLER_ASAP7_75t_R FILLER_0_82_1043 ();
 FILLER_ASAP7_75t_R FILLER_0_82_1055 ();
 FILLER_ASAP7_75t_R FILLER_0_82_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_1065 ();
 FILLER_ASAP7_75t_R FILLER_0_82_1071 ();
 DECAPx2_ASAP7_75t_R FILLER_0_82_1083 ();
 FILLER_ASAP7_75t_R FILLER_0_82_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_1091 ();
 DECAPx4_ASAP7_75t_R FILLER_0_82_1095 ();
 FILLER_ASAP7_75t_R FILLER_0_82_1111 ();
 DECAPx2_ASAP7_75t_R FILLER_0_82_1119 ();
 FILLER_ASAP7_75t_R FILLER_0_82_1131 ();
 FILLER_ASAP7_75t_R FILLER_0_82_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_1141 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_1147 ();
 DECAPx6_ASAP7_75t_R FILLER_0_82_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_1170 ();
 DECAPx4_ASAP7_75t_R FILLER_0_82_1179 ();
 FILLER_ASAP7_75t_R FILLER_0_82_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_1204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_1226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_1270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_1336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_1358 ();
 FILLER_ASAP7_75t_R FILLER_0_82_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_83_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_15 ();
 FILLER_ASAP7_75t_R FILLER_0_83_19 ();
 DECAPx1_ASAP7_75t_R FILLER_0_83_24 ();
 DECAPx6_ASAP7_75t_R FILLER_0_83_34 ();
 DECAPx1_ASAP7_75t_R FILLER_0_83_48 ();
 FILLER_ASAP7_75t_R FILLER_0_83_62 ();
 DECAPx4_ASAP7_75t_R FILLER_0_83_76 ();
 FILLER_ASAP7_75t_R FILLER_0_83_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_95 ();
 FILLER_ASAP7_75t_R FILLER_0_83_103 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_117 ();
 FILLER_ASAP7_75t_R FILLER_0_83_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_130 ();
 FILLER_ASAP7_75t_R FILLER_0_83_137 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_156 ();
 DECAPx4_ASAP7_75t_R FILLER_0_83_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_177 ();
 DECAPx6_ASAP7_75t_R FILLER_0_83_202 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_224 ();
 FILLER_ASAP7_75t_R FILLER_0_83_242 ();
 DECAPx6_ASAP7_75t_R FILLER_0_83_264 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_284 ();
 FILLER_ASAP7_75t_R FILLER_0_83_291 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_302 ();
 FILLER_ASAP7_75t_R FILLER_0_83_308 ();
 FILLER_ASAP7_75t_R FILLER_0_83_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_318 ();
 DECAPx1_ASAP7_75t_R FILLER_0_83_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_329 ();
 DECAPx6_ASAP7_75t_R FILLER_0_83_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_350 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_363 ();
 FILLER_ASAP7_75t_R FILLER_0_83_370 ();
 FILLER_ASAP7_75t_R FILLER_0_83_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_381 ();
 DECAPx4_ASAP7_75t_R FILLER_0_83_392 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_414 ();
 DECAPx1_ASAP7_75t_R FILLER_0_83_423 ();
 DECAPx1_ASAP7_75t_R FILLER_0_83_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_437 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_444 ();
 DECAPx6_ASAP7_75t_R FILLER_0_83_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_480 ();
 DECAPx4_ASAP7_75t_R FILLER_0_83_487 ();
 FILLER_ASAP7_75t_R FILLER_0_83_500 ();
 DECAPx6_ASAP7_75t_R FILLER_0_83_508 ();
 FILLER_ASAP7_75t_R FILLER_0_83_522 ();
 DECAPx4_ASAP7_75t_R FILLER_0_83_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_540 ();
 DECAPx4_ASAP7_75t_R FILLER_0_83_552 ();
 FILLER_ASAP7_75t_R FILLER_0_83_562 ();
 DECAPx4_ASAP7_75t_R FILLER_0_83_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_586 ();
 FILLER_ASAP7_75t_R FILLER_0_83_592 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_597 ();
 FILLER_ASAP7_75t_R FILLER_0_83_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_605 ();
 DECAPx1_ASAP7_75t_R FILLER_0_83_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_616 ();
 FILLER_ASAP7_75t_R FILLER_0_83_620 ();
 DECAPx1_ASAP7_75t_R FILLER_0_83_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_632 ();
 FILLER_ASAP7_75t_R FILLER_0_83_639 ();
 DECAPx4_ASAP7_75t_R FILLER_0_83_644 ();
 FILLER_ASAP7_75t_R FILLER_0_83_654 ();
 FILLER_ASAP7_75t_R FILLER_0_83_662 ();
 FILLER_ASAP7_75t_R FILLER_0_83_670 ();
 FILLER_ASAP7_75t_R FILLER_0_83_678 ();
 FILLER_ASAP7_75t_R FILLER_0_83_690 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_702 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_716 ();
 FILLER_ASAP7_75t_R FILLER_0_83_729 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_741 ();
 FILLER_ASAP7_75t_R FILLER_0_83_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_749 ();
 DECAPx4_ASAP7_75t_R FILLER_0_83_757 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_773 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_787 ();
 FILLER_ASAP7_75t_R FILLER_0_83_798 ();
 FILLER_ASAP7_75t_R FILLER_0_83_814 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_822 ();
 FILLER_ASAP7_75t_R FILLER_0_83_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_830 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_837 ();
 FILLER_ASAP7_75t_R FILLER_0_83_843 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_851 ();
 FILLER_ASAP7_75t_R FILLER_0_83_857 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_869 ();
 FILLER_ASAP7_75t_R FILLER_0_83_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_893 ();
 FILLER_ASAP7_75t_R FILLER_0_83_906 ();
 FILLER_ASAP7_75t_R FILLER_0_83_914 ();
 FILLER_ASAP7_75t_R FILLER_0_83_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_924 ();
 DECAPx6_ASAP7_75t_R FILLER_0_83_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_941 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_962 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_990 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_994 ();
 FILLER_ASAP7_75t_R FILLER_0_83_1000 ();
 FILLER_ASAP7_75t_R FILLER_0_83_1012 ();
 FILLER_ASAP7_75t_R FILLER_0_83_1022 ();
 FILLER_ASAP7_75t_R FILLER_0_83_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_1032 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_1049 ();
 FILLER_ASAP7_75t_R FILLER_0_83_1058 ();
 FILLER_ASAP7_75t_R FILLER_0_83_1063 ();
 FILLER_ASAP7_75t_R FILLER_0_83_1069 ();
 FILLER_ASAP7_75t_R FILLER_0_83_1076 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_1092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_1098 ();
 DECAPx1_ASAP7_75t_R FILLER_0_83_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_1124 ();
 DECAPx1_ASAP7_75t_R FILLER_0_83_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_1135 ();
 DECAPx6_ASAP7_75t_R FILLER_0_83_1141 ();
 FILLER_ASAP7_75t_R FILLER_0_83_1161 ();
 DECAPx1_ASAP7_75t_R FILLER_0_83_1183 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_1251 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_1273 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_1295 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_1317 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_1339 ();
 DECAPx6_ASAP7_75t_R FILLER_0_83_1361 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_84_2 ();
 FILLER_ASAP7_75t_R FILLER_0_84_7 ();
 FILLER_ASAP7_75t_R FILLER_0_84_20 ();
 DECAPx6_ASAP7_75t_R FILLER_0_84_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_46 ();
 FILLER_ASAP7_75t_R FILLER_0_84_53 ();
 DECAPx1_ASAP7_75t_R FILLER_0_84_61 ();
 DECAPx1_ASAP7_75t_R FILLER_0_84_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_75 ();
 FILLER_ASAP7_75t_R FILLER_0_84_83 ();
 DECAPx1_ASAP7_75t_R FILLER_0_84_95 ();
 DECAPx1_ASAP7_75t_R FILLER_0_84_106 ();
 DECAPx2_ASAP7_75t_R FILLER_0_84_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_122 ();
 DECAPx2_ASAP7_75t_R FILLER_0_84_133 ();
 FILLER_ASAP7_75t_R FILLER_0_84_150 ();
 FILLER_ASAP7_75t_R FILLER_0_84_157 ();
 DECAPx1_ASAP7_75t_R FILLER_0_84_165 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_180 ();
 DECAPx2_ASAP7_75t_R FILLER_0_84_202 ();
 FILLER_ASAP7_75t_R FILLER_0_84_208 ();
 DECAPx6_ASAP7_75t_R FILLER_0_84_220 ();
 DECAPx1_ASAP7_75t_R FILLER_0_84_234 ();
 DECAPx1_ASAP7_75t_R FILLER_0_84_248 ();
 DECAPx1_ASAP7_75t_R FILLER_0_84_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_259 ();
 DECAPx2_ASAP7_75t_R FILLER_0_84_266 ();
 FILLER_ASAP7_75t_R FILLER_0_84_272 ();
 FILLER_ASAP7_75t_R FILLER_0_84_280 ();
 FILLER_ASAP7_75t_R FILLER_0_84_288 ();
 DECAPx1_ASAP7_75t_R FILLER_0_84_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_302 ();
 FILLER_ASAP7_75t_R FILLER_0_84_311 ();
 FILLER_ASAP7_75t_R FILLER_0_84_316 ();
 FILLER_ASAP7_75t_R FILLER_0_84_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_326 ();
 FILLER_ASAP7_75t_R FILLER_0_84_333 ();
 DECAPx2_ASAP7_75t_R FILLER_0_84_338 ();
 FILLER_ASAP7_75t_R FILLER_0_84_350 ();
 FILLER_ASAP7_75t_R FILLER_0_84_358 ();
 DECAPx6_ASAP7_75t_R FILLER_0_84_367 ();
 DECAPx1_ASAP7_75t_R FILLER_0_84_381 ();
 FILLER_ASAP7_75t_R FILLER_0_84_391 ();
 FILLER_ASAP7_75t_R FILLER_0_84_396 ();
 FILLER_ASAP7_75t_R FILLER_0_84_404 ();
 FILLER_ASAP7_75t_R FILLER_0_84_414 ();
 DECAPx1_ASAP7_75t_R FILLER_0_84_422 ();
 DECAPx2_ASAP7_75t_R FILLER_0_84_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_438 ();
 FILLER_ASAP7_75t_R FILLER_0_84_448 ();
 FILLER_ASAP7_75t_R FILLER_0_84_460 ();
 DECAPx4_ASAP7_75t_R FILLER_0_84_464 ();
 FILLER_ASAP7_75t_R FILLER_0_84_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_476 ();
 DECAPx6_ASAP7_75t_R FILLER_0_84_483 ();
 FILLER_ASAP7_75t_R FILLER_0_84_497 ();
 DECAPx1_ASAP7_75t_R FILLER_0_84_505 ();
 DECAPx2_ASAP7_75t_R FILLER_0_84_515 ();
 DECAPx4_ASAP7_75t_R FILLER_0_84_527 ();
 FILLER_ASAP7_75t_R FILLER_0_84_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_539 ();
 FILLER_ASAP7_75t_R FILLER_0_84_546 ();
 DECAPx4_ASAP7_75t_R FILLER_0_84_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_564 ();
 DECAPx6_ASAP7_75t_R FILLER_0_84_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_582 ();
 FILLER_ASAP7_75t_R FILLER_0_84_591 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_599 ();
 FILLER_ASAP7_75t_R FILLER_0_84_631 ();
 DECAPx4_ASAP7_75t_R FILLER_0_84_639 ();
 FILLER_ASAP7_75t_R FILLER_0_84_654 ();
 FILLER_ASAP7_75t_R FILLER_0_84_666 ();
 FILLER_ASAP7_75t_R FILLER_0_84_678 ();
 FILLER_ASAP7_75t_R FILLER_0_84_688 ();
 FILLER_ASAP7_75t_R FILLER_0_84_700 ();
 FILLER_ASAP7_75t_R FILLER_0_84_712 ();
 FILLER_ASAP7_75t_R FILLER_0_84_724 ();
 FILLER_ASAP7_75t_R FILLER_0_84_736 ();
 FILLER_ASAP7_75t_R FILLER_0_84_743 ();
 FILLER_ASAP7_75t_R FILLER_0_84_750 ();
 DECAPx2_ASAP7_75t_R FILLER_0_84_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_761 ();
 FILLER_ASAP7_75t_R FILLER_0_84_768 ();
 FILLER_ASAP7_75t_R FILLER_0_84_777 ();
 FILLER_ASAP7_75t_R FILLER_0_84_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_787 ();
 DECAPx2_ASAP7_75t_R FILLER_0_84_798 ();
 DECAPx1_ASAP7_75t_R FILLER_0_84_815 ();
 DECAPx2_ASAP7_75t_R FILLER_0_84_828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_84_845 ();
 DECAPx2_ASAP7_75t_R FILLER_0_84_857 ();
 FILLER_ASAP7_75t_R FILLER_0_84_869 ();
 DECAPx2_ASAP7_75t_R FILLER_0_84_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_882 ();
 FILLER_ASAP7_75t_R FILLER_0_84_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_891 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_918 ();
 DECAPx2_ASAP7_75t_R FILLER_0_84_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_946 ();
 DECAPx2_ASAP7_75t_R FILLER_0_84_957 ();
 FILLER_ASAP7_75t_R FILLER_0_84_963 ();
 FILLER_ASAP7_75t_R FILLER_0_84_972 ();
 DECAPx2_ASAP7_75t_R FILLER_0_84_980 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_986 ();
 FILLER_ASAP7_75t_R FILLER_0_84_997 ();
 DECAPx6_ASAP7_75t_R FILLER_0_84_1004 ();
 DECAPx2_ASAP7_75t_R FILLER_0_84_1024 ();
 FILLER_ASAP7_75t_R FILLER_0_84_1030 ();
 FILLER_ASAP7_75t_R FILLER_0_84_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_1044 ();
 FILLER_ASAP7_75t_R FILLER_0_84_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_0_84_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_1068 ();
 DECAPx2_ASAP7_75t_R FILLER_0_84_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_1085 ();
 FILLER_ASAP7_75t_R FILLER_0_84_1093 ();
 DECAPx4_ASAP7_75t_R FILLER_0_84_1102 ();
 FILLER_ASAP7_75t_R FILLER_0_84_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_1114 ();
 DECAPx4_ASAP7_75t_R FILLER_0_84_1121 ();
 FILLER_ASAP7_75t_R FILLER_0_84_1141 ();
 DECAPx6_ASAP7_75t_R FILLER_0_84_1153 ();
 FILLER_ASAP7_75t_R FILLER_0_84_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_1169 ();
 FILLER_ASAP7_75t_R FILLER_0_84_1176 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_1178 ();
 DECAPx1_ASAP7_75t_R FILLER_0_84_1185 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_1189 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_1240 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_1262 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_1284 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_1306 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_1328 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_1350 ();
 DECAPx4_ASAP7_75t_R FILLER_0_84_1372 ();
 FILLER_ASAP7_75t_R FILLER_0_85_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_4 ();
 FILLER_ASAP7_75t_R FILLER_0_85_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_12 ();
 FILLER_ASAP7_75t_R FILLER_0_85_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_21 ();
 DECAPx1_ASAP7_75t_R FILLER_0_85_28 ();
 FILLER_ASAP7_75t_R FILLER_0_85_48 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_83 ();
 FILLER_ASAP7_75t_R FILLER_0_85_90 ();
 DECAPx2_ASAP7_75t_R FILLER_0_85_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_104 ();
 DECAPx1_ASAP7_75t_R FILLER_0_85_117 ();
 FILLER_ASAP7_75t_R FILLER_0_85_127 ();
 FILLER_ASAP7_75t_R FILLER_0_85_137 ();
 DECAPx2_ASAP7_75t_R FILLER_0_85_144 ();
 FILLER_ASAP7_75t_R FILLER_0_85_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_152 ();
 FILLER_ASAP7_75t_R FILLER_0_85_159 ();
 FILLER_ASAP7_75t_R FILLER_0_85_168 ();
 FILLER_ASAP7_75t_R FILLER_0_85_180 ();
 DECAPx2_ASAP7_75t_R FILLER_0_85_190 ();
 FILLER_ASAP7_75t_R FILLER_0_85_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_198 ();
 FILLER_ASAP7_75t_R FILLER_0_85_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_207 ();
 FILLER_ASAP7_75t_R FILLER_0_85_213 ();
 FILLER_ASAP7_75t_R FILLER_0_85_225 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_237 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_259 ();
 DECAPx1_ASAP7_75t_R FILLER_0_85_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_285 ();
 DECAPx2_ASAP7_75t_R FILLER_0_85_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_300 ();
 DECAPx2_ASAP7_75t_R FILLER_0_85_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_313 ();
 DECAPx2_ASAP7_75t_R FILLER_0_85_321 ();
 FILLER_ASAP7_75t_R FILLER_0_85_327 ();
 FILLER_ASAP7_75t_R FILLER_0_85_337 ();
 DECAPx2_ASAP7_75t_R FILLER_0_85_344 ();
 FILLER_ASAP7_75t_R FILLER_0_85_350 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_358 ();
 DECAPx1_ASAP7_75t_R FILLER_0_85_380 ();
 DECAPx1_ASAP7_75t_R FILLER_0_85_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_396 ();
 DECAPx2_ASAP7_75t_R FILLER_0_85_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_410 ();
 DECAPx2_ASAP7_75t_R FILLER_0_85_417 ();
 FILLER_ASAP7_75t_R FILLER_0_85_429 ();
 FILLER_ASAP7_75t_R FILLER_0_85_437 ();
 DECAPx6_ASAP7_75t_R FILLER_0_85_445 ();
 FILLER_ASAP7_75t_R FILLER_0_85_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_461 ();
 FILLER_ASAP7_75t_R FILLER_0_85_482 ();
 DECAPx2_ASAP7_75t_R FILLER_0_85_491 ();
 FILLER_ASAP7_75t_R FILLER_0_85_504 ();
 FILLER_ASAP7_75t_R FILLER_0_85_513 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_521 ();
 DECAPx6_ASAP7_75t_R FILLER_0_85_549 ();
 DECAPx1_ASAP7_75t_R FILLER_0_85_563 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_574 ();
 FILLER_ASAP7_75t_R FILLER_0_85_602 ();
 DECAPx6_ASAP7_75t_R FILLER_0_85_610 ();
 DECAPx2_ASAP7_75t_R FILLER_0_85_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_630 ();
 DECAPx4_ASAP7_75t_R FILLER_0_85_638 ();
 FILLER_ASAP7_75t_R FILLER_0_85_648 ();
 FILLER_ASAP7_75t_R FILLER_0_85_655 ();
 FILLER_ASAP7_75t_R FILLER_0_85_662 ();
 FILLER_ASAP7_75t_R FILLER_0_85_674 ();
 FILLER_ASAP7_75t_R FILLER_0_85_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_688 ();
 FILLER_ASAP7_75t_R FILLER_0_85_694 ();
 FILLER_ASAP7_75t_R FILLER_0_85_706 ();
 FILLER_ASAP7_75t_R FILLER_0_85_718 ();
 FILLER_ASAP7_75t_R FILLER_0_85_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_732 ();
 FILLER_ASAP7_75t_R FILLER_0_85_743 ();
 DECAPx4_ASAP7_75t_R FILLER_0_85_757 ();
 DECAPx6_ASAP7_75t_R FILLER_0_85_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_789 ();
 FILLER_ASAP7_75t_R FILLER_0_85_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_802 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_809 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_831 ();
 DECAPx2_ASAP7_75t_R FILLER_0_85_853 ();
 FILLER_ASAP7_75t_R FILLER_0_85_859 ();
 DECAPx2_ASAP7_75t_R FILLER_0_85_871 ();
 FILLER_ASAP7_75t_R FILLER_0_85_885 ();
 DECAPx4_ASAP7_75t_R FILLER_0_85_893 ();
 DECAPx6_ASAP7_75t_R FILLER_0_85_909 ();
 FILLER_ASAP7_75t_R FILLER_0_85_923 ();
 DECAPx4_ASAP7_75t_R FILLER_0_85_927 ();
 FILLER_ASAP7_75t_R FILLER_0_85_937 ();
 DECAPx2_ASAP7_75t_R FILLER_0_85_951 ();
 FILLER_ASAP7_75t_R FILLER_0_85_967 ();
 DECAPx4_ASAP7_75t_R FILLER_0_85_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_987 ();
 DECAPx4_ASAP7_75t_R FILLER_0_85_994 ();
 FILLER_ASAP7_75t_R FILLER_0_85_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_1006 ();
 FILLER_ASAP7_75t_R FILLER_0_85_1010 ();
 FILLER_ASAP7_75t_R FILLER_0_85_1018 ();
 FILLER_ASAP7_75t_R FILLER_0_85_1026 ();
 DECAPx2_ASAP7_75t_R FILLER_0_85_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_1040 ();
 FILLER_ASAP7_75t_R FILLER_0_85_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_1055 ();
 FILLER_ASAP7_75t_R FILLER_0_85_1066 ();
 DECAPx2_ASAP7_75t_R FILLER_0_85_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_1079 ();
 FILLER_ASAP7_75t_R FILLER_0_85_1092 ();
 FILLER_ASAP7_75t_R FILLER_0_85_1105 ();
 FILLER_ASAP7_75t_R FILLER_0_85_1113 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_1121 ();
 DECAPx1_ASAP7_75t_R FILLER_0_85_1143 ();
 DECAPx1_ASAP7_75t_R FILLER_0_85_1155 ();
 DECAPx4_ASAP7_75t_R FILLER_0_85_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_1175 ();
 DECAPx1_ASAP7_75t_R FILLER_0_85_1182 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_85_1193 ();
 FILLER_ASAP7_75t_R FILLER_0_85_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_1231 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_1319 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_1341 ();
 DECAPx6_ASAP7_75t_R FILLER_0_85_1363 ();
 DECAPx1_ASAP7_75t_R FILLER_0_85_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_86_2 ();
 FILLER_ASAP7_75t_R FILLER_0_86_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_11 ();
 FILLER_ASAP7_75t_R FILLER_0_86_22 ();
 DECAPx1_ASAP7_75t_R FILLER_0_86_32 ();
 DECAPx2_ASAP7_75t_R FILLER_0_86_42 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_54 ();
 DECAPx6_ASAP7_75t_R FILLER_0_86_76 ();
 DECAPx2_ASAP7_75t_R FILLER_0_86_90 ();
 DECAPx4_ASAP7_75t_R FILLER_0_86_104 ();
 FILLER_ASAP7_75t_R FILLER_0_86_114 ();
 FILLER_ASAP7_75t_R FILLER_0_86_121 ();
 FILLER_ASAP7_75t_R FILLER_0_86_128 ();
 FILLER_ASAP7_75t_R FILLER_0_86_140 ();
 DECAPx2_ASAP7_75t_R FILLER_0_86_148 ();
 FILLER_ASAP7_75t_R FILLER_0_86_154 ();
 DECAPx2_ASAP7_75t_R FILLER_0_86_166 ();
 FILLER_ASAP7_75t_R FILLER_0_86_192 ();
 DECAPx2_ASAP7_75t_R FILLER_0_86_201 ();
 FILLER_ASAP7_75t_R FILLER_0_86_207 ();
 FILLER_ASAP7_75t_R FILLER_0_86_215 ();
 FILLER_ASAP7_75t_R FILLER_0_86_223 ();
 FILLER_ASAP7_75t_R FILLER_0_86_233 ();
 DECAPx1_ASAP7_75t_R FILLER_0_86_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_247 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_254 ();
 FILLER_ASAP7_75t_R FILLER_0_86_282 ();
 DECAPx4_ASAP7_75t_R FILLER_0_86_292 ();
 FILLER_ASAP7_75t_R FILLER_0_86_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_319 ();
 DECAPx4_ASAP7_75t_R FILLER_0_86_341 ();
 DECAPx6_ASAP7_75t_R FILLER_0_86_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_371 ();
 FILLER_ASAP7_75t_R FILLER_0_86_378 ();
 FILLER_ASAP7_75t_R FILLER_0_86_386 ();
 FILLER_ASAP7_75t_R FILLER_0_86_393 ();
 DECAPx6_ASAP7_75t_R FILLER_0_86_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_412 ();
 DECAPx2_ASAP7_75t_R FILLER_0_86_423 ();
 FILLER_ASAP7_75t_R FILLER_0_86_435 ();
 FILLER_ASAP7_75t_R FILLER_0_86_443 ();
 FILLER_ASAP7_75t_R FILLER_0_86_452 ();
 FILLER_ASAP7_75t_R FILLER_0_86_460 ();
 DECAPx2_ASAP7_75t_R FILLER_0_86_464 ();
 FILLER_ASAP7_75t_R FILLER_0_86_476 ();
 DECAPx1_ASAP7_75t_R FILLER_0_86_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_485 ();
 DECAPx4_ASAP7_75t_R FILLER_0_86_492 ();
 FILLER_ASAP7_75t_R FILLER_0_86_502 ();
 DECAPx1_ASAP7_75t_R FILLER_0_86_510 ();
 FILLER_ASAP7_75t_R FILLER_0_86_525 ();
 DECAPx2_ASAP7_75t_R FILLER_0_86_537 ();
 FILLER_ASAP7_75t_R FILLER_0_86_543 ();
 FILLER_ASAP7_75t_R FILLER_0_86_551 ();
 DECAPx2_ASAP7_75t_R FILLER_0_86_559 ();
 DECAPx1_ASAP7_75t_R FILLER_0_86_576 ();
 FILLER_ASAP7_75t_R FILLER_0_86_586 ();
 DECAPx2_ASAP7_75t_R FILLER_0_86_599 ();
 FILLER_ASAP7_75t_R FILLER_0_86_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_607 ();
 FILLER_ASAP7_75t_R FILLER_0_86_619 ();
 FILLER_ASAP7_75t_R FILLER_0_86_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_633 ();
 FILLER_ASAP7_75t_R FILLER_0_86_640 ();
 DECAPx1_ASAP7_75t_R FILLER_0_86_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_652 ();
 FILLER_ASAP7_75t_R FILLER_0_86_658 ();
 FILLER_ASAP7_75t_R FILLER_0_86_665 ();
 FILLER_ASAP7_75t_R FILLER_0_86_677 ();
 FILLER_ASAP7_75t_R FILLER_0_86_689 ();
 DECAPx1_ASAP7_75t_R FILLER_0_86_696 ();
 FILLER_ASAP7_75t_R FILLER_0_86_706 ();
 FILLER_ASAP7_75t_R FILLER_0_86_718 ();
 DECAPx1_ASAP7_75t_R FILLER_0_86_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_734 ();
 FILLER_ASAP7_75t_R FILLER_0_86_741 ();
 DECAPx2_ASAP7_75t_R FILLER_0_86_755 ();
 FILLER_ASAP7_75t_R FILLER_0_86_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_763 ();
 DECAPx6_ASAP7_75t_R FILLER_0_86_774 ();
 FILLER_ASAP7_75t_R FILLER_0_86_788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_795 ();
 DECAPx2_ASAP7_75t_R FILLER_0_86_817 ();
 FILLER_ASAP7_75t_R FILLER_0_86_823 ();
 DECAPx2_ASAP7_75t_R FILLER_0_86_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_839 ();
 DECAPx2_ASAP7_75t_R FILLER_0_86_846 ();
 FILLER_ASAP7_75t_R FILLER_0_86_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_860 ();
 DECAPx1_ASAP7_75t_R FILLER_0_86_867 ();
 DECAPx4_ASAP7_75t_R FILLER_0_86_891 ();
 FILLER_ASAP7_75t_R FILLER_0_86_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_903 ();
 FILLER_ASAP7_75t_R FILLER_0_86_911 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_919 ();
 FILLER_ASAP7_75t_R FILLER_0_86_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_943 ();
 DECAPx4_ASAP7_75t_R FILLER_0_86_956 ();
 FILLER_ASAP7_75t_R FILLER_0_86_966 ();
 DECAPx1_ASAP7_75t_R FILLER_0_86_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_976 ();
 FILLER_ASAP7_75t_R FILLER_0_86_984 ();
 FILLER_ASAP7_75t_R FILLER_0_86_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_995 ();
 DECAPx1_ASAP7_75t_R FILLER_0_86_1004 ();
 FILLER_ASAP7_75t_R FILLER_0_86_1013 ();
 DECAPx1_ASAP7_75t_R FILLER_0_86_1026 ();
 FILLER_ASAP7_75t_R FILLER_0_86_1040 ();
 DECAPx1_ASAP7_75t_R FILLER_0_86_1050 ();
 DECAPx1_ASAP7_75t_R FILLER_0_86_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_1065 ();
 FILLER_ASAP7_75t_R FILLER_0_86_1076 ();
 DECAPx1_ASAP7_75t_R FILLER_0_86_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_1087 ();
 FILLER_ASAP7_75t_R FILLER_0_86_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_1121 ();
 FILLER_ASAP7_75t_R FILLER_0_86_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_1145 ();
 DECAPx6_ASAP7_75t_R FILLER_0_86_1157 ();
 FILLER_ASAP7_75t_R FILLER_0_86_1171 ();
 FILLER_ASAP7_75t_R FILLER_0_86_1179 ();
 FILLER_ASAP7_75t_R FILLER_0_86_1187 ();
 FILLER_ASAP7_75t_R FILLER_0_86_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_1203 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_1269 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_1313 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_1335 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_86_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_87_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_87_9 ();
 DECAPx1_ASAP7_75t_R FILLER_0_87_25 ();
 FILLER_ASAP7_75t_R FILLER_0_87_35 ();
 FILLER_ASAP7_75t_R FILLER_0_87_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_45 ();
 FILLER_ASAP7_75t_R FILLER_0_87_52 ();
 DECAPx6_ASAP7_75t_R FILLER_0_87_57 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_77 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_86 ();
 FILLER_ASAP7_75t_R FILLER_0_87_92 ();
 FILLER_ASAP7_75t_R FILLER_0_87_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_102 ();
 DECAPx1_ASAP7_75t_R FILLER_0_87_113 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_133 ();
 FILLER_ASAP7_75t_R FILLER_0_87_140 ();
 DECAPx1_ASAP7_75t_R FILLER_0_87_148 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_166 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_170 ();
 FILLER_ASAP7_75t_R FILLER_0_87_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_178 ();
 DECAPx1_ASAP7_75t_R FILLER_0_87_189 ();
 FILLER_ASAP7_75t_R FILLER_0_87_199 ();
 FILLER_ASAP7_75t_R FILLER_0_87_211 ();
 DECAPx1_ASAP7_75t_R FILLER_0_87_219 ();
 FILLER_ASAP7_75t_R FILLER_0_87_233 ();
 FILLER_ASAP7_75t_R FILLER_0_87_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_256 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_278 ();
 DECAPx4_ASAP7_75t_R FILLER_0_87_290 ();
 FILLER_ASAP7_75t_R FILLER_0_87_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_302 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_310 ();
 DECAPx1_ASAP7_75t_R FILLER_0_87_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_326 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_333 ();
 FILLER_ASAP7_75t_R FILLER_0_87_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_347 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_356 ();
 FILLER_ASAP7_75t_R FILLER_0_87_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_380 ();
 DECAPx1_ASAP7_75t_R FILLER_0_87_387 ();
 DECAPx1_ASAP7_75t_R FILLER_0_87_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_398 ();
 FILLER_ASAP7_75t_R FILLER_0_87_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_408 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_415 ();
 FILLER_ASAP7_75t_R FILLER_0_87_437 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_445 ();
 DECAPx1_ASAP7_75t_R FILLER_0_87_467 ();
 FILLER_ASAP7_75t_R FILLER_0_87_477 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_489 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_511 ();
 FILLER_ASAP7_75t_R FILLER_0_87_517 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_535 ();
 FILLER_ASAP7_75t_R FILLER_0_87_542 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_561 ();
 FILLER_ASAP7_75t_R FILLER_0_87_570 ();
 DECAPx1_ASAP7_75t_R FILLER_0_87_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_582 ();
 DECAPx1_ASAP7_75t_R FILLER_0_87_589 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_599 ();
 DECAPx1_ASAP7_75t_R FILLER_0_87_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_615 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_622 ();
 FILLER_ASAP7_75t_R FILLER_0_87_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_630 ();
 DECAPx1_ASAP7_75t_R FILLER_0_87_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_641 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_655 ();
 FILLER_ASAP7_75t_R FILLER_0_87_662 ();
 FILLER_ASAP7_75t_R FILLER_0_87_670 ();
 FILLER_ASAP7_75t_R FILLER_0_87_682 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_696 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_707 ();
 FILLER_ASAP7_75t_R FILLER_0_87_723 ();
 FILLER_ASAP7_75t_R FILLER_0_87_735 ();
 DECAPx6_ASAP7_75t_R FILLER_0_87_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_757 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_770 ();
 FILLER_ASAP7_75t_R FILLER_0_87_777 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_785 ();
 DECAPx1_ASAP7_75t_R FILLER_0_87_798 ();
 FILLER_ASAP7_75t_R FILLER_0_87_809 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_818 ();
 FILLER_ASAP7_75t_R FILLER_0_87_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_826 ();
 DECAPx1_ASAP7_75t_R FILLER_0_87_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_841 ();
 DECAPx4_ASAP7_75t_R FILLER_0_87_852 ();
 FILLER_ASAP7_75t_R FILLER_0_87_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_864 ();
 DECAPx6_ASAP7_75t_R FILLER_0_87_870 ();
 FILLER_ASAP7_75t_R FILLER_0_87_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_886 ();
 FILLER_ASAP7_75t_R FILLER_0_87_893 ();
 FILLER_ASAP7_75t_R FILLER_0_87_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_907 ();
 DECAPx4_ASAP7_75t_R FILLER_0_87_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_924 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_927 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_955 ();
 DECAPx6_ASAP7_75t_R FILLER_0_87_962 ();
 FILLER_ASAP7_75t_R FILLER_0_87_976 ();
 FILLER_ASAP7_75t_R FILLER_0_87_990 ();
 DECAPx6_ASAP7_75t_R FILLER_0_87_998 ();
 FILLER_ASAP7_75t_R FILLER_0_87_1012 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_1026 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_1047 ();
 FILLER_ASAP7_75t_R FILLER_0_87_1053 ();
 FILLER_ASAP7_75t_R FILLER_0_87_1061 ();
 FILLER_ASAP7_75t_R FILLER_0_87_1073 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_1109 ();
 FILLER_ASAP7_75t_R FILLER_0_87_1116 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_1130 ();
 FILLER_ASAP7_75t_R FILLER_0_87_1138 ();
 DECAPx6_ASAP7_75t_R FILLER_0_87_1150 ();
 FILLER_ASAP7_75t_R FILLER_0_87_1164 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_1172 ();
 FILLER_ASAP7_75t_R FILLER_0_87_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_1180 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_1187 ();
 FILLER_ASAP7_75t_R FILLER_0_87_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_1195 ();
 FILLER_ASAP7_75t_R FILLER_0_87_1202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_1251 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_1273 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_1295 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_1317 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_1339 ();
 DECAPx6_ASAP7_75t_R FILLER_0_87_1361 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_88_2 ();
 FILLER_ASAP7_75t_R FILLER_0_88_9 ();
 FILLER_ASAP7_75t_R FILLER_0_88_16 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_22 ();
 FILLER_ASAP7_75t_R FILLER_0_88_34 ();
 FILLER_ASAP7_75t_R FILLER_0_88_42 ();
 FILLER_ASAP7_75t_R FILLER_0_88_50 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_58 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_77 ();
 DECAPx6_ASAP7_75t_R FILLER_0_88_84 ();
 DECAPx1_ASAP7_75t_R FILLER_0_88_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_102 ();
 FILLER_ASAP7_75t_R FILLER_0_88_110 ();
 FILLER_ASAP7_75t_R FILLER_0_88_132 ();
 FILLER_ASAP7_75t_R FILLER_0_88_140 ();
 FILLER_ASAP7_75t_R FILLER_0_88_146 ();
 FILLER_ASAP7_75t_R FILLER_0_88_160 ();
 DECAPx6_ASAP7_75t_R FILLER_0_88_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_181 ();
 DECAPx1_ASAP7_75t_R FILLER_0_88_202 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_216 ();
 FILLER_ASAP7_75t_R FILLER_0_88_230 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_238 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_260 ();
 FILLER_ASAP7_75t_R FILLER_0_88_272 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_280 ();
 FILLER_ASAP7_75t_R FILLER_0_88_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_288 ();
 FILLER_ASAP7_75t_R FILLER_0_88_295 ();
 DECAPx1_ASAP7_75t_R FILLER_0_88_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_307 ();
 FILLER_ASAP7_75t_R FILLER_0_88_314 ();
 DECAPx1_ASAP7_75t_R FILLER_0_88_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_327 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_336 ();
 FILLER_ASAP7_75t_R FILLER_0_88_348 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_356 ();
 FILLER_ASAP7_75t_R FILLER_0_88_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_370 ();
 DECAPx1_ASAP7_75t_R FILLER_0_88_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_381 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_394 ();
 FILLER_ASAP7_75t_R FILLER_0_88_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_403 ();
 FILLER_ASAP7_75t_R FILLER_0_88_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_409 ();
 FILLER_ASAP7_75t_R FILLER_0_88_416 ();
 FILLER_ASAP7_75t_R FILLER_0_88_424 ();
 FILLER_ASAP7_75t_R FILLER_0_88_434 ();
 FILLER_ASAP7_75t_R FILLER_0_88_460 ();
 DECAPx1_ASAP7_75t_R FILLER_0_88_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_468 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_475 ();
 FILLER_ASAP7_75t_R FILLER_0_88_487 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_501 ();
 DECAPx1_ASAP7_75t_R FILLER_0_88_505 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_515 ();
 FILLER_ASAP7_75t_R FILLER_0_88_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_523 ();
 FILLER_ASAP7_75t_R FILLER_0_88_530 ();
 DECAPx4_ASAP7_75t_R FILLER_0_88_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_545 ();
 DECAPx4_ASAP7_75t_R FILLER_0_88_554 ();
 FILLER_ASAP7_75t_R FILLER_0_88_564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_574 ();
 DECAPx1_ASAP7_75t_R FILLER_0_88_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_600 ();
 DECAPx4_ASAP7_75t_R FILLER_0_88_607 ();
 FILLER_ASAP7_75t_R FILLER_0_88_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_619 ();
 DECAPx1_ASAP7_75t_R FILLER_0_88_625 ();
 FILLER_ASAP7_75t_R FILLER_0_88_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_638 ();
 DECAPx4_ASAP7_75t_R FILLER_0_88_645 ();
 FILLER_ASAP7_75t_R FILLER_0_88_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_657 ();
 FILLER_ASAP7_75t_R FILLER_0_88_664 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_676 ();
 FILLER_ASAP7_75t_R FILLER_0_88_682 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_694 ();
 FILLER_ASAP7_75t_R FILLER_0_88_700 ();
 FILLER_ASAP7_75t_R FILLER_0_88_712 ();
 FILLER_ASAP7_75t_R FILLER_0_88_724 ();
 FILLER_ASAP7_75t_R FILLER_0_88_734 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_742 ();
 FILLER_ASAP7_75t_R FILLER_0_88_764 ();
 DECAPx1_ASAP7_75t_R FILLER_0_88_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_777 ();
 FILLER_ASAP7_75t_R FILLER_0_88_789 ();
 DECAPx4_ASAP7_75t_R FILLER_0_88_802 ();
 DECAPx1_ASAP7_75t_R FILLER_0_88_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_826 ();
 FILLER_ASAP7_75t_R FILLER_0_88_833 ();
 DECAPx1_ASAP7_75t_R FILLER_0_88_841 ();
 DECAPx1_ASAP7_75t_R FILLER_0_88_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_855 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_862 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_878 ();
 DECAPx1_ASAP7_75t_R FILLER_0_88_887 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_897 ();
 DECAPx1_ASAP7_75t_R FILLER_0_88_909 ();
 FILLER_ASAP7_75t_R FILLER_0_88_919 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_927 ();
 DECAPx1_ASAP7_75t_R FILLER_0_88_949 ();
 FILLER_ASAP7_75t_R FILLER_0_88_959 ();
 DECAPx4_ASAP7_75t_R FILLER_0_88_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_977 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_984 ();
 FILLER_ASAP7_75t_R FILLER_0_88_990 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_1000 ();
 DECAPx4_ASAP7_75t_R FILLER_0_88_1022 ();
 FILLER_ASAP7_75t_R FILLER_0_88_1032 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_1050 ();
 DECAPx1_ASAP7_75t_R FILLER_0_88_1061 ();
 FILLER_ASAP7_75t_R FILLER_0_88_1075 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_1082 ();
 FILLER_ASAP7_75t_R FILLER_0_88_1088 ();
 FILLER_ASAP7_75t_R FILLER_0_88_1097 ();
 FILLER_ASAP7_75t_R FILLER_0_88_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_1108 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_1137 ();
 FILLER_ASAP7_75t_R FILLER_0_88_1144 ();
 FILLER_ASAP7_75t_R FILLER_0_88_1157 ();
 DECAPx4_ASAP7_75t_R FILLER_0_88_1169 ();
 FILLER_ASAP7_75t_R FILLER_0_88_1185 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_1215 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_1259 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_1281 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_1303 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_1325 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_1347 ();
 DECAPx4_ASAP7_75t_R FILLER_0_88_1369 ();
 FILLER_ASAP7_75t_R FILLER_0_88_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_89_2 ();
 FILLER_ASAP7_75t_R FILLER_0_89_9 ();
 FILLER_ASAP7_75t_R FILLER_0_89_16 ();
 FILLER_ASAP7_75t_R FILLER_0_89_23 ();
 FILLER_ASAP7_75t_R FILLER_0_89_28 ();
 DECAPx1_ASAP7_75t_R FILLER_0_89_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_40 ();
 FILLER_ASAP7_75t_R FILLER_0_89_47 ();
 FILLER_ASAP7_75t_R FILLER_0_89_55 ();
 FILLER_ASAP7_75t_R FILLER_0_89_63 ();
 DECAPx2_ASAP7_75t_R FILLER_0_89_71 ();
 FILLER_ASAP7_75t_R FILLER_0_89_83 ();
 FILLER_ASAP7_75t_R FILLER_0_89_91 ();
 FILLER_ASAP7_75t_R FILLER_0_89_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_102 ();
 FILLER_ASAP7_75t_R FILLER_0_89_109 ();
 FILLER_ASAP7_75t_R FILLER_0_89_118 ();
 DECAPx1_ASAP7_75t_R FILLER_0_89_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_134 ();
 FILLER_ASAP7_75t_R FILLER_0_89_145 ();
 FILLER_ASAP7_75t_R FILLER_0_89_154 ();
 DECAPx1_ASAP7_75t_R FILLER_0_89_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_166 ();
 DECAPx6_ASAP7_75t_R FILLER_0_89_174 ();
 DECAPx2_ASAP7_75t_R FILLER_0_89_188 ();
 DECAPx6_ASAP7_75t_R FILLER_0_89_200 ();
 FILLER_ASAP7_75t_R FILLER_0_89_234 ();
 FILLER_ASAP7_75t_R FILLER_0_89_246 ();
 DECAPx6_ASAP7_75t_R FILLER_0_89_253 ();
 DECAPx2_ASAP7_75t_R FILLER_0_89_267 ();
 DECAPx2_ASAP7_75t_R FILLER_0_89_293 ();
 DECAPx2_ASAP7_75t_R FILLER_0_89_305 ();
 FILLER_ASAP7_75t_R FILLER_0_89_311 ();
 DECAPx6_ASAP7_75t_R FILLER_0_89_319 ();
 DECAPx2_ASAP7_75t_R FILLER_0_89_339 ();
 FILLER_ASAP7_75t_R FILLER_0_89_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_347 ();
 DECAPx6_ASAP7_75t_R FILLER_0_89_351 ();
 DECAPx6_ASAP7_75t_R FILLER_0_89_371 ();
 DECAPx2_ASAP7_75t_R FILLER_0_89_385 ();
 FILLER_ASAP7_75t_R FILLER_0_89_401 ();
 DECAPx6_ASAP7_75t_R FILLER_0_89_423 ();
 FILLER_ASAP7_75t_R FILLER_0_89_443 ();
 DECAPx2_ASAP7_75t_R FILLER_0_89_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_462 ();
 DECAPx1_ASAP7_75t_R FILLER_0_89_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_488 ();
 DECAPx2_ASAP7_75t_R FILLER_0_89_495 ();
 DECAPx1_ASAP7_75t_R FILLER_0_89_507 ();
 DECAPx2_ASAP7_75t_R FILLER_0_89_517 ();
 FILLER_ASAP7_75t_R FILLER_0_89_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_532 ();
 FILLER_ASAP7_75t_R FILLER_0_89_544 ();
 DECAPx2_ASAP7_75t_R FILLER_0_89_556 ();
 FILLER_ASAP7_75t_R FILLER_0_89_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_564 ();
 FILLER_ASAP7_75t_R FILLER_0_89_577 ();
 FILLER_ASAP7_75t_R FILLER_0_89_591 ();
 FILLER_ASAP7_75t_R FILLER_0_89_599 ();
 FILLER_ASAP7_75t_R FILLER_0_89_607 ();
 FILLER_ASAP7_75t_R FILLER_0_89_616 ();
 DECAPx1_ASAP7_75t_R FILLER_0_89_626 ();
 FILLER_ASAP7_75t_R FILLER_0_89_635 ();
 DECAPx1_ASAP7_75t_R FILLER_0_89_652 ();
 FILLER_ASAP7_75t_R FILLER_0_89_666 ();
 DECAPx2_ASAP7_75t_R FILLER_0_89_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_684 ();
 DECAPx1_ASAP7_75t_R FILLER_0_89_695 ();
 FILLER_ASAP7_75t_R FILLER_0_89_705 ();
 FILLER_ASAP7_75t_R FILLER_0_89_713 ();
 FILLER_ASAP7_75t_R FILLER_0_89_723 ();
 FILLER_ASAP7_75t_R FILLER_0_89_733 ();
 FILLER_ASAP7_75t_R FILLER_0_89_741 ();
 DECAPx6_ASAP7_75t_R FILLER_0_89_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_763 ();
 DECAPx1_ASAP7_75t_R FILLER_0_89_774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_807 ();
 DECAPx6_ASAP7_75t_R FILLER_0_89_811 ();
 DECAPx1_ASAP7_75t_R FILLER_0_89_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_829 ();
 FILLER_ASAP7_75t_R FILLER_0_89_840 ();
 FILLER_ASAP7_75t_R FILLER_0_89_848 ();
 FILLER_ASAP7_75t_R FILLER_0_89_856 ();
 FILLER_ASAP7_75t_R FILLER_0_89_865 ();
 FILLER_ASAP7_75t_R FILLER_0_89_873 ();
 FILLER_ASAP7_75t_R FILLER_0_89_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_883 ();
 FILLER_ASAP7_75t_R FILLER_0_89_890 ();
 FILLER_ASAP7_75t_R FILLER_0_89_898 ();
 DECAPx1_ASAP7_75t_R FILLER_0_89_905 ();
 FILLER_ASAP7_75t_R FILLER_0_89_915 ();
 FILLER_ASAP7_75t_R FILLER_0_89_923 ();
 DECAPx6_ASAP7_75t_R FILLER_0_89_927 ();
 FILLER_ASAP7_75t_R FILLER_0_89_953 ();
 FILLER_ASAP7_75t_R FILLER_0_89_967 ();
 FILLER_ASAP7_75t_R FILLER_0_89_975 ();
 FILLER_ASAP7_75t_R FILLER_0_89_985 ();
 FILLER_ASAP7_75t_R FILLER_0_89_999 ();
 FILLER_ASAP7_75t_R FILLER_0_89_1013 ();
 DECAPx1_ASAP7_75t_R FILLER_0_89_1021 ();
 FILLER_ASAP7_75t_R FILLER_0_89_1031 ();
 DECAPx1_ASAP7_75t_R FILLER_0_89_1043 ();
 FILLER_ASAP7_75t_R FILLER_0_89_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_0_89_1062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_89_1076 ();
 FILLER_ASAP7_75t_R FILLER_0_89_1092 ();
 FILLER_ASAP7_75t_R FILLER_0_89_1105 ();
 DECAPx1_ASAP7_75t_R FILLER_0_89_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_1123 ();
 FILLER_ASAP7_75t_R FILLER_0_89_1136 ();
 DECAPx6_ASAP7_75t_R FILLER_0_89_1144 ();
 FILLER_ASAP7_75t_R FILLER_0_89_1168 ();
 FILLER_ASAP7_75t_R FILLER_0_89_1180 ();
 FILLER_ASAP7_75t_R FILLER_0_89_1188 ();
 FILLER_ASAP7_75t_R FILLER_0_89_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_1333 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_1355 ();
 DECAPx1_ASAP7_75t_R FILLER_0_89_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_1381 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_6 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_12 ();
 DECAPx2_ASAP7_75t_R FILLER_0_90_21 ();
 FILLER_ASAP7_75t_R FILLER_0_90_27 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_35 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_53 ();
 FILLER_ASAP7_75t_R FILLER_0_90_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_62 ();
 DECAPx6_ASAP7_75t_R FILLER_0_90_69 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_83 ();
 FILLER_ASAP7_75t_R FILLER_0_90_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_96 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_105 ();
 DECAPx2_ASAP7_75t_R FILLER_0_90_117 ();
 DECAPx2_ASAP7_75t_R FILLER_0_90_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_135 ();
 FILLER_ASAP7_75t_R FILLER_0_90_146 ();
 DECAPx2_ASAP7_75t_R FILLER_0_90_153 ();
 FILLER_ASAP7_75t_R FILLER_0_90_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_168 ();
 FILLER_ASAP7_75t_R FILLER_0_90_175 ();
 DECAPx4_ASAP7_75t_R FILLER_0_90_183 ();
 FILLER_ASAP7_75t_R FILLER_0_90_193 ();
 FILLER_ASAP7_75t_R FILLER_0_90_203 ();
 DECAPx2_ASAP7_75t_R FILLER_0_90_213 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_231 ();
 FILLER_ASAP7_75t_R FILLER_0_90_242 ();
 DECAPx6_ASAP7_75t_R FILLER_0_90_255 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_273 ();
 FILLER_ASAP7_75t_R FILLER_0_90_280 ();
 FILLER_ASAP7_75t_R FILLER_0_90_288 ();
 FILLER_ASAP7_75t_R FILLER_0_90_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_299 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_308 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_330 ();
 DECAPx6_ASAP7_75t_R FILLER_0_90_340 ();
 FILLER_ASAP7_75t_R FILLER_0_90_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_356 ();
 FILLER_ASAP7_75t_R FILLER_0_90_363 ();
 DECAPx6_ASAP7_75t_R FILLER_0_90_373 ();
 FILLER_ASAP7_75t_R FILLER_0_90_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_389 ();
 FILLER_ASAP7_75t_R FILLER_0_90_396 ();
 FILLER_ASAP7_75t_R FILLER_0_90_404 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_412 ();
 DECAPx4_ASAP7_75t_R FILLER_0_90_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_432 ();
 FILLER_ASAP7_75t_R FILLER_0_90_439 ();
 FILLER_ASAP7_75t_R FILLER_0_90_444 ();
 DECAPx2_ASAP7_75t_R FILLER_0_90_454 ();
 FILLER_ASAP7_75t_R FILLER_0_90_460 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_464 ();
 FILLER_ASAP7_75t_R FILLER_0_90_488 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_496 ();
 DECAPx2_ASAP7_75t_R FILLER_0_90_506 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_522 ();
 DECAPx2_ASAP7_75t_R FILLER_0_90_530 ();
 DECAPx2_ASAP7_75t_R FILLER_0_90_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_545 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_556 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_567 ();
 FILLER_ASAP7_75t_R FILLER_0_90_581 ();
 FILLER_ASAP7_75t_R FILLER_0_90_588 ();
 FILLER_ASAP7_75t_R FILLER_0_90_602 ();
 FILLER_ASAP7_75t_R FILLER_0_90_609 ();
 FILLER_ASAP7_75t_R FILLER_0_90_617 ();
 FILLER_ASAP7_75t_R FILLER_0_90_625 ();
 FILLER_ASAP7_75t_R FILLER_0_90_633 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_643 ();
 DECAPx2_ASAP7_75t_R FILLER_0_90_655 ();
 FILLER_ASAP7_75t_R FILLER_0_90_661 ();
 FILLER_ASAP7_75t_R FILLER_0_90_673 ();
 FILLER_ASAP7_75t_R FILLER_0_90_680 ();
 FILLER_ASAP7_75t_R FILLER_0_90_692 ();
 DECAPx2_ASAP7_75t_R FILLER_0_90_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_705 ();
 DECAPx4_ASAP7_75t_R FILLER_0_90_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_726 ();
 DECAPx2_ASAP7_75t_R FILLER_0_90_737 ();
 FILLER_ASAP7_75t_R FILLER_0_90_743 ();
 DECAPx2_ASAP7_75t_R FILLER_0_90_752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_90_778 ();
 FILLER_ASAP7_75t_R FILLER_0_90_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_786 ();
 FILLER_ASAP7_75t_R FILLER_0_90_793 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_803 ();
 DECAPx2_ASAP7_75t_R FILLER_0_90_813 ();
 FILLER_ASAP7_75t_R FILLER_0_90_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_821 ();
 DECAPx6_ASAP7_75t_R FILLER_0_90_842 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_856 ();
 DECAPx6_ASAP7_75t_R FILLER_0_90_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_880 ();
 DECAPx2_ASAP7_75t_R FILLER_0_90_887 ();
 FILLER_ASAP7_75t_R FILLER_0_90_899 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_916 ();
 FILLER_ASAP7_75t_R FILLER_0_90_923 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_931 ();
 FILLER_ASAP7_75t_R FILLER_0_90_953 ();
 FILLER_ASAP7_75t_R FILLER_0_90_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_963 ();
 FILLER_ASAP7_75t_R FILLER_0_90_970 ();
 FILLER_ASAP7_75t_R FILLER_0_90_977 ();
 DECAPx4_ASAP7_75t_R FILLER_0_90_982 ();
 FILLER_ASAP7_75t_R FILLER_0_90_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_1003 ();
 DECAPx4_ASAP7_75t_R FILLER_0_90_1025 ();
 FILLER_ASAP7_75t_R FILLER_0_90_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_1037 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_1048 ();
 FILLER_ASAP7_75t_R FILLER_0_90_1058 ();
 DECAPx2_ASAP7_75t_R FILLER_0_90_1066 ();
 DECAPx6_ASAP7_75t_R FILLER_0_90_1080 ();
 DECAPx4_ASAP7_75t_R FILLER_0_90_1100 ();
 DECAPx2_ASAP7_75t_R FILLER_0_90_1116 ();
 FILLER_ASAP7_75t_R FILLER_0_90_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_1124 ();
 FILLER_ASAP7_75t_R FILLER_0_90_1131 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_1143 ();
 DECAPx2_ASAP7_75t_R FILLER_0_90_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_1160 ();
 FILLER_ASAP7_75t_R FILLER_0_90_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_1169 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_1181 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_1191 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_1255 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_1277 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_1299 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_1321 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_1343 ();
 DECAPx6_ASAP7_75t_R FILLER_0_90_1365 ();
 FILLER_ASAP7_75t_R FILLER_0_90_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_91_2 ();
 FILLER_ASAP7_75t_R FILLER_0_91_9 ();
 DECAPx1_ASAP7_75t_R FILLER_0_91_16 ();
 FILLER_ASAP7_75t_R FILLER_0_91_25 ();
 FILLER_ASAP7_75t_R FILLER_0_91_33 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_41 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_63 ();
 FILLER_ASAP7_75t_R FILLER_0_91_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_71 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_78 ();
 FILLER_ASAP7_75t_R FILLER_0_91_84 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_112 ();
 FILLER_ASAP7_75t_R FILLER_0_91_119 ();
 DECAPx1_ASAP7_75t_R FILLER_0_91_127 ();
 FILLER_ASAP7_75t_R FILLER_0_91_141 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_153 ();
 FILLER_ASAP7_75t_R FILLER_0_91_159 ();
 FILLER_ASAP7_75t_R FILLER_0_91_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_169 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_177 ();
 FILLER_ASAP7_75t_R FILLER_0_91_183 ();
 FILLER_ASAP7_75t_R FILLER_0_91_195 ();
 FILLER_ASAP7_75t_R FILLER_0_91_217 ();
 FILLER_ASAP7_75t_R FILLER_0_91_229 ();
 FILLER_ASAP7_75t_R FILLER_0_91_251 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_263 ();
 FILLER_ASAP7_75t_R FILLER_0_91_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_287 ();
 DECAPx6_ASAP7_75t_R FILLER_0_91_294 ();
 DECAPx1_ASAP7_75t_R FILLER_0_91_308 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_318 ();
 FILLER_ASAP7_75t_R FILLER_0_91_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_326 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_333 ();
 FILLER_ASAP7_75t_R FILLER_0_91_339 ();
 FILLER_ASAP7_75t_R FILLER_0_91_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_363 ();
 DECAPx4_ASAP7_75t_R FILLER_0_91_370 ();
 FILLER_ASAP7_75t_R FILLER_0_91_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_382 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_392 ();
 FILLER_ASAP7_75t_R FILLER_0_91_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_401 ();
 FILLER_ASAP7_75t_R FILLER_0_91_408 ();
 FILLER_ASAP7_75t_R FILLER_0_91_416 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_446 ();
 FILLER_ASAP7_75t_R FILLER_0_91_469 ();
 FILLER_ASAP7_75t_R FILLER_0_91_477 ();
 DECAPx1_ASAP7_75t_R FILLER_0_91_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_489 ();
 FILLER_ASAP7_75t_R FILLER_0_91_496 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_503 ();
 DECAPx1_ASAP7_75t_R FILLER_0_91_519 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_523 ();
 DECAPx1_ASAP7_75t_R FILLER_0_91_531 ();
 FILLER_ASAP7_75t_R FILLER_0_91_540 ();
 DECAPx4_ASAP7_75t_R FILLER_0_91_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_559 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_570 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_587 ();
 FILLER_ASAP7_75t_R FILLER_0_91_593 ();
 FILLER_ASAP7_75t_R FILLER_0_91_601 ();
 FILLER_ASAP7_75t_R FILLER_0_91_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_611 ();
 DECAPx1_ASAP7_75t_R FILLER_0_91_622 ();
 DECAPx1_ASAP7_75t_R FILLER_0_91_636 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_653 ();
 FILLER_ASAP7_75t_R FILLER_0_91_659 ();
 FILLER_ASAP7_75t_R FILLER_0_91_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_668 ();
 FILLER_ASAP7_75t_R FILLER_0_91_677 ();
 DECAPx4_ASAP7_75t_R FILLER_0_91_687 ();
 FILLER_ASAP7_75t_R FILLER_0_91_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_699 ();
 DECAPx4_ASAP7_75t_R FILLER_0_91_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_713 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_720 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_733 ();
 FILLER_ASAP7_75t_R FILLER_0_91_739 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_747 ();
 DECAPx1_ASAP7_75t_R FILLER_0_91_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_777 ();
 DECAPx1_ASAP7_75t_R FILLER_0_91_784 ();
 DECAPx1_ASAP7_75t_R FILLER_0_91_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_800 ();
 DECAPx1_ASAP7_75t_R FILLER_0_91_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_811 ();
 FILLER_ASAP7_75t_R FILLER_0_91_823 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_831 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_843 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_865 ();
 DECAPx1_ASAP7_75t_R FILLER_0_91_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_891 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_911 ();
 FILLER_ASAP7_75t_R FILLER_0_91_923 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_927 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_949 ();
 FILLER_ASAP7_75t_R FILLER_0_91_966 ();
 DECAPx1_ASAP7_75t_R FILLER_0_91_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_980 ();
 FILLER_ASAP7_75t_R FILLER_0_91_987 ();
 DECAPx6_ASAP7_75t_R FILLER_0_91_996 ();
 FILLER_ASAP7_75t_R FILLER_0_91_1010 ();
 DECAPx4_ASAP7_75t_R FILLER_0_91_1019 ();
 FILLER_ASAP7_75t_R FILLER_0_91_1029 ();
 FILLER_ASAP7_75t_R FILLER_0_91_1051 ();
 FILLER_ASAP7_75t_R FILLER_0_91_1063 ();
 DECAPx4_ASAP7_75t_R FILLER_0_91_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_1089 ();
 DECAPx4_ASAP7_75t_R FILLER_0_91_1100 ();
 FILLER_ASAP7_75t_R FILLER_0_91_1110 ();
 DECAPx1_ASAP7_75t_R FILLER_0_91_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_1122 ();
 FILLER_ASAP7_75t_R FILLER_0_91_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_1131 ();
 DECAPx1_ASAP7_75t_R FILLER_0_91_1138 ();
 DECAPx4_ASAP7_75t_R FILLER_0_91_1148 ();
 FILLER_ASAP7_75t_R FILLER_0_91_1158 ();
 DECAPx1_ASAP7_75t_R FILLER_0_91_1164 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_1180 ();
 FILLER_ASAP7_75t_R FILLER_0_91_1187 ();
 DECAPx4_ASAP7_75t_R FILLER_0_91_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_1211 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_1255 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_1277 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_1299 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_1321 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_1343 ();
 DECAPx6_ASAP7_75t_R FILLER_0_91_1365 ();
 FILLER_ASAP7_75t_R FILLER_0_91_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_92_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_92_9 ();
 FILLER_ASAP7_75t_R FILLER_0_92_34 ();
 DECAPx6_ASAP7_75t_R FILLER_0_92_42 ();
 DECAPx2_ASAP7_75t_R FILLER_0_92_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_62 ();
 DECAPx4_ASAP7_75t_R FILLER_0_92_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_79 ();
 FILLER_ASAP7_75t_R FILLER_0_92_90 ();
 FILLER_ASAP7_75t_R FILLER_0_92_102 ();
 FILLER_ASAP7_75t_R FILLER_0_92_114 ();
 FILLER_ASAP7_75t_R FILLER_0_92_136 ();
 DECAPx4_ASAP7_75t_R FILLER_0_92_148 ();
 DECAPx2_ASAP7_75t_R FILLER_0_92_168 ();
 FILLER_ASAP7_75t_R FILLER_0_92_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_176 ();
 DECAPx6_ASAP7_75t_R FILLER_0_92_183 ();
 FILLER_ASAP7_75t_R FILLER_0_92_197 ();
 FILLER_ASAP7_75t_R FILLER_0_92_205 ();
 DECAPx6_ASAP7_75t_R FILLER_0_92_213 ();
 DECAPx1_ASAP7_75t_R FILLER_0_92_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_231 ();
 DECAPx2_ASAP7_75t_R FILLER_0_92_242 ();
 FILLER_ASAP7_75t_R FILLER_0_92_248 ();
 DECAPx2_ASAP7_75t_R FILLER_0_92_256 ();
 DECAPx6_ASAP7_75t_R FILLER_0_92_270 ();
 DECAPx1_ASAP7_75t_R FILLER_0_92_284 ();
 FILLER_ASAP7_75t_R FILLER_0_92_296 ();
 FILLER_ASAP7_75t_R FILLER_0_92_320 ();
 FILLER_ASAP7_75t_R FILLER_0_92_328 ();
 DECAPx1_ASAP7_75t_R FILLER_0_92_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_341 ();
 FILLER_ASAP7_75t_R FILLER_0_92_362 ();
 DECAPx1_ASAP7_75t_R FILLER_0_92_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_374 ();
 FILLER_ASAP7_75t_R FILLER_0_92_381 ();
 FILLER_ASAP7_75t_R FILLER_0_92_388 ();
 DECAPx2_ASAP7_75t_R FILLER_0_92_393 ();
 FILLER_ASAP7_75t_R FILLER_0_92_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_401 ();
 DECAPx6_ASAP7_75t_R FILLER_0_92_410 ();
 FILLER_ASAP7_75t_R FILLER_0_92_424 ();
 DECAPx4_ASAP7_75t_R FILLER_0_92_429 ();
 DECAPx6_ASAP7_75t_R FILLER_0_92_446 ();
 FILLER_ASAP7_75t_R FILLER_0_92_460 ();
 DECAPx6_ASAP7_75t_R FILLER_0_92_464 ();
 FILLER_ASAP7_75t_R FILLER_0_92_478 ();
 DECAPx1_ASAP7_75t_R FILLER_0_92_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_487 ();
 FILLER_ASAP7_75t_R FILLER_0_92_494 ();
 DECAPx2_ASAP7_75t_R FILLER_0_92_516 ();
 FILLER_ASAP7_75t_R FILLER_0_92_522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_527 ();
 DECAPx6_ASAP7_75t_R FILLER_0_92_549 ();
 DECAPx2_ASAP7_75t_R FILLER_0_92_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_569 ();
 FILLER_ASAP7_75t_R FILLER_0_92_580 ();
 DECAPx2_ASAP7_75t_R FILLER_0_92_592 ();
 FILLER_ASAP7_75t_R FILLER_0_92_603 ();
 DECAPx2_ASAP7_75t_R FILLER_0_92_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_621 ();
 FILLER_ASAP7_75t_R FILLER_0_92_632 ();
 DECAPx1_ASAP7_75t_R FILLER_0_92_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_648 ();
 FILLER_ASAP7_75t_R FILLER_0_92_657 ();
 FILLER_ASAP7_75t_R FILLER_0_92_665 ();
 FILLER_ASAP7_75t_R FILLER_0_92_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_675 ();
 DECAPx4_ASAP7_75t_R FILLER_0_92_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_697 ();
 FILLER_ASAP7_75t_R FILLER_0_92_703 ();
 DECAPx1_ASAP7_75t_R FILLER_0_92_711 ();
 DECAPx2_ASAP7_75t_R FILLER_0_92_722 ();
 DECAPx4_ASAP7_75t_R FILLER_0_92_738 ();
 DECAPx2_ASAP7_75t_R FILLER_0_92_758 ();
 FILLER_ASAP7_75t_R FILLER_0_92_770 ();
 DECAPx2_ASAP7_75t_R FILLER_0_92_777 ();
 FILLER_ASAP7_75t_R FILLER_0_92_793 ();
 FILLER_ASAP7_75t_R FILLER_0_92_805 ();
 DECAPx1_ASAP7_75t_R FILLER_0_92_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_816 ();
 DECAPx4_ASAP7_75t_R FILLER_0_92_823 ();
 FILLER_ASAP7_75t_R FILLER_0_92_833 ();
 DECAPx2_ASAP7_75t_R FILLER_0_92_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_851 ();
 DECAPx1_ASAP7_75t_R FILLER_0_92_858 ();
 FILLER_ASAP7_75t_R FILLER_0_92_868 ();
 DECAPx4_ASAP7_75t_R FILLER_0_92_876 ();
 FILLER_ASAP7_75t_R FILLER_0_92_886 ();
 DECAPx2_ASAP7_75t_R FILLER_0_92_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_905 ();
 DECAPx2_ASAP7_75t_R FILLER_0_92_916 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_922 ();
 DECAPx4_ASAP7_75t_R FILLER_0_92_945 ();
 FILLER_ASAP7_75t_R FILLER_0_92_961 ();
 DECAPx6_ASAP7_75t_R FILLER_0_92_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_983 ();
 DECAPx6_ASAP7_75t_R FILLER_0_92_994 ();
 DECAPx6_ASAP7_75t_R FILLER_0_92_1014 ();
 DECAPx2_ASAP7_75t_R FILLER_0_92_1028 ();
 DECAPx1_ASAP7_75t_R FILLER_0_92_1044 ();
 FILLER_ASAP7_75t_R FILLER_0_92_1054 ();
 DECAPx2_ASAP7_75t_R FILLER_0_92_1062 ();
 DECAPx4_ASAP7_75t_R FILLER_0_92_1073 ();
 FILLER_ASAP7_75t_R FILLER_0_92_1083 ();
 FILLER_ASAP7_75t_R FILLER_0_92_1091 ();
 DECAPx2_ASAP7_75t_R FILLER_0_92_1101 ();
 DECAPx2_ASAP7_75t_R FILLER_0_92_1113 ();
 FILLER_ASAP7_75t_R FILLER_0_92_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_1134 ();
 DECAPx1_ASAP7_75t_R FILLER_0_92_1156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_1166 ();
 FILLER_ASAP7_75t_R FILLER_0_92_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_1196 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_1240 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_1262 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_1284 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_1306 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_1328 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_1350 ();
 DECAPx4_ASAP7_75t_R FILLER_0_92_1372 ();
 FILLER_ASAP7_75t_R FILLER_0_93_2 ();
 FILLER_ASAP7_75t_R FILLER_0_93_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_11 ();
 FILLER_ASAP7_75t_R FILLER_0_93_15 ();
 DECAPx2_ASAP7_75t_R FILLER_0_93_23 ();
 FILLER_ASAP7_75t_R FILLER_0_93_29 ();
 FILLER_ASAP7_75t_R FILLER_0_93_51 ();
 FILLER_ASAP7_75t_R FILLER_0_93_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_65 ();
 FILLER_ASAP7_75t_R FILLER_0_93_72 ();
 DECAPx2_ASAP7_75t_R FILLER_0_93_84 ();
 FILLER_ASAP7_75t_R FILLER_0_93_90 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_102 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_116 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_127 ();
 FILLER_ASAP7_75t_R FILLER_0_93_138 ();
 DECAPx4_ASAP7_75t_R FILLER_0_93_150 ();
 FILLER_ASAP7_75t_R FILLER_0_93_166 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_175 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_186 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_214 ();
 FILLER_ASAP7_75t_R FILLER_0_93_221 ();
 FILLER_ASAP7_75t_R FILLER_0_93_233 ();
 FILLER_ASAP7_75t_R FILLER_0_93_240 ();
 FILLER_ASAP7_75t_R FILLER_0_93_252 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_259 ();
 DECAPx2_ASAP7_75t_R FILLER_0_93_281 ();
 FILLER_ASAP7_75t_R FILLER_0_93_287 ();
 FILLER_ASAP7_75t_R FILLER_0_93_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_299 ();
 FILLER_ASAP7_75t_R FILLER_0_93_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_316 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_323 ();
 DECAPx2_ASAP7_75t_R FILLER_0_93_333 ();
 FILLER_ASAP7_75t_R FILLER_0_93_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_341 ();
 FILLER_ASAP7_75t_R FILLER_0_93_350 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_358 ();
 DECAPx4_ASAP7_75t_R FILLER_0_93_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_390 ();
 DECAPx2_ASAP7_75t_R FILLER_0_93_398 ();
 FILLER_ASAP7_75t_R FILLER_0_93_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_406 ();
 DECAPx2_ASAP7_75t_R FILLER_0_93_410 ();
 FILLER_ASAP7_75t_R FILLER_0_93_422 ();
 FILLER_ASAP7_75t_R FILLER_0_93_432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_440 ();
 DECAPx6_ASAP7_75t_R FILLER_0_93_462 ();
 DECAPx2_ASAP7_75t_R FILLER_0_93_476 ();
 DECAPx2_ASAP7_75t_R FILLER_0_93_488 ();
 FILLER_ASAP7_75t_R FILLER_0_93_494 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_516 ();
 FILLER_ASAP7_75t_R FILLER_0_93_526 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_537 ();
 DECAPx6_ASAP7_75t_R FILLER_0_93_544 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_558 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_562 ();
 FILLER_ASAP7_75t_R FILLER_0_93_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_572 ();
 DECAPx6_ASAP7_75t_R FILLER_0_93_579 ();
 FILLER_ASAP7_75t_R FILLER_0_93_593 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_601 ();
 FILLER_ASAP7_75t_R FILLER_0_93_611 ();
 FILLER_ASAP7_75t_R FILLER_0_93_620 ();
 FILLER_ASAP7_75t_R FILLER_0_93_632 ();
 FILLER_ASAP7_75t_R FILLER_0_93_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_646 ();
 DECAPx2_ASAP7_75t_R FILLER_0_93_657 ();
 FILLER_ASAP7_75t_R FILLER_0_93_669 ();
 FILLER_ASAP7_75t_R FILLER_0_93_679 ();
 DECAPx2_ASAP7_75t_R FILLER_0_93_693 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_705 ();
 FILLER_ASAP7_75t_R FILLER_0_93_719 ();
 FILLER_ASAP7_75t_R FILLER_0_93_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_93_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_741 ();
 FILLER_ASAP7_75t_R FILLER_0_93_762 ();
 FILLER_ASAP7_75t_R FILLER_0_93_772 ();
 FILLER_ASAP7_75t_R FILLER_0_93_780 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_788 ();
 FILLER_ASAP7_75t_R FILLER_0_93_802 ();
 FILLER_ASAP7_75t_R FILLER_0_93_810 ();
 FILLER_ASAP7_75t_R FILLER_0_93_818 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_830 ();
 DECAPx2_ASAP7_75t_R FILLER_0_93_836 ();
 FILLER_ASAP7_75t_R FILLER_0_93_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_844 ();
 FILLER_ASAP7_75t_R FILLER_0_93_851 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_865 ();
 FILLER_ASAP7_75t_R FILLER_0_93_872 ();
 FILLER_ASAP7_75t_R FILLER_0_93_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_882 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_889 ();
 FILLER_ASAP7_75t_R FILLER_0_93_899 ();
 DECAPx2_ASAP7_75t_R FILLER_0_93_907 ();
 FILLER_ASAP7_75t_R FILLER_0_93_913 ();
 FILLER_ASAP7_75t_R FILLER_0_93_923 ();
 FILLER_ASAP7_75t_R FILLER_0_93_927 ();
 DECAPx2_ASAP7_75t_R FILLER_0_93_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_941 ();
 FILLER_ASAP7_75t_R FILLER_0_93_948 ();
 FILLER_ASAP7_75t_R FILLER_0_93_960 ();
 DECAPx6_ASAP7_75t_R FILLER_0_93_970 ();
 DECAPx2_ASAP7_75t_R FILLER_0_93_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_990 ();
 DECAPx6_ASAP7_75t_R FILLER_0_93_1007 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_1025 ();
 DECAPx6_ASAP7_75t_R FILLER_0_93_1033 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_1047 ();
 DECAPx6_ASAP7_75t_R FILLER_0_93_1054 ();
 FILLER_ASAP7_75t_R FILLER_0_93_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_0_93_1082 ();
 FILLER_ASAP7_75t_R FILLER_0_93_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_1090 ();
 DECAPx2_ASAP7_75t_R FILLER_0_93_1097 ();
 FILLER_ASAP7_75t_R FILLER_0_93_1109 ();
 FILLER_ASAP7_75t_R FILLER_0_93_1117 ();
 FILLER_ASAP7_75t_R FILLER_0_93_1125 ();
 FILLER_ASAP7_75t_R FILLER_0_93_1133 ();
 DECAPx6_ASAP7_75t_R FILLER_0_93_1141 ();
 FILLER_ASAP7_75t_R FILLER_0_93_1155 ();
 FILLER_ASAP7_75t_R FILLER_0_93_1163 ();
 DECAPx4_ASAP7_75t_R FILLER_0_93_1171 ();
 FILLER_ASAP7_75t_R FILLER_0_93_1187 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_1197 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_1207 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_1251 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_1273 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_1295 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_1317 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_1339 ();
 DECAPx6_ASAP7_75t_R FILLER_0_93_1361 ();
 DECAPx2_ASAP7_75t_R FILLER_0_93_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_94_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_94_9 ();
 FILLER_ASAP7_75t_R FILLER_0_94_15 ();
 DECAPx2_ASAP7_75t_R FILLER_0_94_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_28 ();
 DECAPx1_ASAP7_75t_R FILLER_0_94_35 ();
 DECAPx1_ASAP7_75t_R FILLER_0_94_45 ();
 DECAPx2_ASAP7_75t_R FILLER_0_94_55 ();
 FILLER_ASAP7_75t_R FILLER_0_94_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_69 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_76 ();
 DECAPx2_ASAP7_75t_R FILLER_0_94_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_104 ();
 DECAPx2_ASAP7_75t_R FILLER_0_94_115 ();
 DECAPx2_ASAP7_75t_R FILLER_0_94_127 ();
 FILLER_ASAP7_75t_R FILLER_0_94_133 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_145 ();
 DECAPx6_ASAP7_75t_R FILLER_0_94_167 ();
 FILLER_ASAP7_75t_R FILLER_0_94_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_183 ();
 FILLER_ASAP7_75t_R FILLER_0_94_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_196 ();
 DECAPx2_ASAP7_75t_R FILLER_0_94_203 ();
 FILLER_ASAP7_75t_R FILLER_0_94_209 ();
 FILLER_ASAP7_75t_R FILLER_0_94_221 ();
 FILLER_ASAP7_75t_R FILLER_0_94_230 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_242 ();
 DECAPx6_ASAP7_75t_R FILLER_0_94_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_278 ();
 FILLER_ASAP7_75t_R FILLER_0_94_289 ();
 FILLER_ASAP7_75t_R FILLER_0_94_299 ();
 FILLER_ASAP7_75t_R FILLER_0_94_311 ();
 FILLER_ASAP7_75t_R FILLER_0_94_319 ();
 FILLER_ASAP7_75t_R FILLER_0_94_327 ();
 FILLER_ASAP7_75t_R FILLER_0_94_339 ();
 FILLER_ASAP7_75t_R FILLER_0_94_347 ();
 DECAPx1_ASAP7_75t_R FILLER_0_94_352 ();
 FILLER_ASAP7_75t_R FILLER_0_94_366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_380 ();
 DECAPx1_ASAP7_75t_R FILLER_0_94_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_406 ();
 FILLER_ASAP7_75t_R FILLER_0_94_413 ();
 DECAPx2_ASAP7_75t_R FILLER_0_94_421 ();
 FILLER_ASAP7_75t_R FILLER_0_94_433 ();
 DECAPx2_ASAP7_75t_R FILLER_0_94_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_449 ();
 FILLER_ASAP7_75t_R FILLER_0_94_460 ();
 FILLER_ASAP7_75t_R FILLER_0_94_464 ();
 DECAPx1_ASAP7_75t_R FILLER_0_94_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_476 ();
 FILLER_ASAP7_75t_R FILLER_0_94_483 ();
 FILLER_ASAP7_75t_R FILLER_0_94_496 ();
 DECAPx1_ASAP7_75t_R FILLER_0_94_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_508 ();
 DECAPx1_ASAP7_75t_R FILLER_0_94_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_516 ();
 FILLER_ASAP7_75t_R FILLER_0_94_523 ();
 DECAPx1_ASAP7_75t_R FILLER_0_94_531 ();
 DECAPx1_ASAP7_75t_R FILLER_0_94_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_546 ();
 FILLER_ASAP7_75t_R FILLER_0_94_553 ();
 FILLER_ASAP7_75t_R FILLER_0_94_562 ();
 DECAPx4_ASAP7_75t_R FILLER_0_94_575 ();
 DECAPx2_ASAP7_75t_R FILLER_0_94_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_597 ();
 DECAPx2_ASAP7_75t_R FILLER_0_94_604 ();
 FILLER_ASAP7_75t_R FILLER_0_94_615 ();
 FILLER_ASAP7_75t_R FILLER_0_94_629 ();
 FILLER_ASAP7_75t_R FILLER_0_94_641 ();
 DECAPx4_ASAP7_75t_R FILLER_0_94_653 ();
 FILLER_ASAP7_75t_R FILLER_0_94_663 ();
 FILLER_ASAP7_75t_R FILLER_0_94_675 ();
 FILLER_ASAP7_75t_R FILLER_0_94_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_685 ();
 FILLER_ASAP7_75t_R FILLER_0_94_696 ();
 DECAPx1_ASAP7_75t_R FILLER_0_94_704 ();
 FILLER_ASAP7_75t_R FILLER_0_94_718 ();
 FILLER_ASAP7_75t_R FILLER_0_94_727 ();
 FILLER_ASAP7_75t_R FILLER_0_94_747 ();
 FILLER_ASAP7_75t_R FILLER_0_94_759 ();
 DECAPx1_ASAP7_75t_R FILLER_0_94_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_773 ();
 FILLER_ASAP7_75t_R FILLER_0_94_781 ();
 DECAPx2_ASAP7_75t_R FILLER_0_94_789 ();
 FILLER_ASAP7_75t_R FILLER_0_94_805 ();
 DECAPx1_ASAP7_75t_R FILLER_0_94_815 ();
 DECAPx1_ASAP7_75t_R FILLER_0_94_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_828 ();
 FILLER_ASAP7_75t_R FILLER_0_94_839 ();
 DECAPx6_ASAP7_75t_R FILLER_0_94_849 ();
 FILLER_ASAP7_75t_R FILLER_0_94_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_871 ();
 DECAPx2_ASAP7_75t_R FILLER_0_94_877 ();
 FILLER_ASAP7_75t_R FILLER_0_94_889 ();
 FILLER_ASAP7_75t_R FILLER_0_94_897 ();
 FILLER_ASAP7_75t_R FILLER_0_94_905 ();
 FILLER_ASAP7_75t_R FILLER_0_94_913 ();
 DECAPx6_ASAP7_75t_R FILLER_0_94_921 ();
 DECAPx2_ASAP7_75t_R FILLER_0_94_935 ();
 FILLER_ASAP7_75t_R FILLER_0_94_947 ();
 FILLER_ASAP7_75t_R FILLER_0_94_959 ();
 FILLER_ASAP7_75t_R FILLER_0_94_967 ();
 FILLER_ASAP7_75t_R FILLER_0_94_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_977 ();
 DECAPx2_ASAP7_75t_R FILLER_0_94_984 ();
 DECAPx4_ASAP7_75t_R FILLER_0_94_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_1006 ();
 DECAPx4_ASAP7_75t_R FILLER_0_94_1018 ();
 FILLER_ASAP7_75t_R FILLER_0_94_1034 ();
 DECAPx1_ASAP7_75t_R FILLER_0_94_1042 ();
 DECAPx2_ASAP7_75t_R FILLER_0_94_1056 ();
 FILLER_ASAP7_75t_R FILLER_0_94_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_1064 ();
 FILLER_ASAP7_75t_R FILLER_0_94_1071 ();
 FILLER_ASAP7_75t_R FILLER_0_94_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_1081 ();
 FILLER_ASAP7_75t_R FILLER_0_94_1088 ();
 DECAPx4_ASAP7_75t_R FILLER_0_94_1097 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_1107 ();
 DECAPx4_ASAP7_75t_R FILLER_0_94_1114 ();
 FILLER_ASAP7_75t_R FILLER_0_94_1124 ();
 DECAPx6_ASAP7_75t_R FILLER_0_94_1136 ();
 FILLER_ASAP7_75t_R FILLER_0_94_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_1152 ();
 FILLER_ASAP7_75t_R FILLER_0_94_1159 ();
 DECAPx2_ASAP7_75t_R FILLER_0_94_1167 ();
 FILLER_ASAP7_75t_R FILLER_0_94_1183 ();
 FILLER_ASAP7_75t_R FILLER_0_94_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_1209 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_1231 ();
 FILLER_ASAP7_75t_R FILLER_0_94_1253 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_1255 ();
 DECAPx1_ASAP7_75t_R FILLER_0_94_1262 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_1266 ();
 FILLER_ASAP7_75t_R FILLER_0_94_1270 ();
 DECAPx6_ASAP7_75t_R FILLER_0_94_1278 ();
 DECAPx2_ASAP7_75t_R FILLER_0_94_1292 ();
 FILLER_ASAP7_75t_R FILLER_0_94_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_1312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_1334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_1356 ();
 DECAPx1_ASAP7_75t_R FILLER_0_94_1378 ();
 FILLER_ASAP7_75t_R FILLER_0_95_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_95_9 ();
 DECAPx1_ASAP7_75t_R FILLER_0_95_33 ();
 FILLER_ASAP7_75t_R FILLER_0_95_43 ();
 DECAPx1_ASAP7_75t_R FILLER_0_95_50 ();
 DECAPx6_ASAP7_75t_R FILLER_0_95_60 ();
 DECAPx1_ASAP7_75t_R FILLER_0_95_74 ();
 FILLER_ASAP7_75t_R FILLER_0_95_88 ();
 DECAPx1_ASAP7_75t_R FILLER_0_95_97 ();
 FILLER_ASAP7_75t_R FILLER_0_95_119 ();
 FILLER_ASAP7_75t_R FILLER_0_95_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_129 ();
 FILLER_ASAP7_75t_R FILLER_0_95_136 ();
 DECAPx6_ASAP7_75t_R FILLER_0_95_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_158 ();
 FILLER_ASAP7_75t_R FILLER_0_95_165 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_178 ();
 FILLER_ASAP7_75t_R FILLER_0_95_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_202 ();
 FILLER_ASAP7_75t_R FILLER_0_95_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_211 ();
 FILLER_ASAP7_75t_R FILLER_0_95_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_219 ();
 FILLER_ASAP7_75t_R FILLER_0_95_227 ();
 DECAPx6_ASAP7_75t_R FILLER_0_95_234 ();
 FILLER_ASAP7_75t_R FILLER_0_95_248 ();
 FILLER_ASAP7_75t_R FILLER_0_95_270 ();
 FILLER_ASAP7_75t_R FILLER_0_95_276 ();
 FILLER_ASAP7_75t_R FILLER_0_95_288 ();
 FILLER_ASAP7_75t_R FILLER_0_95_300 ();
 FILLER_ASAP7_75t_R FILLER_0_95_309 ();
 FILLER_ASAP7_75t_R FILLER_0_95_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_318 ();
 DECAPx6_ASAP7_75t_R FILLER_0_95_325 ();
 DECAPx1_ASAP7_75t_R FILLER_0_95_339 ();
 DECAPx4_ASAP7_75t_R FILLER_0_95_349 ();
 FILLER_ASAP7_75t_R FILLER_0_95_359 ();
 FILLER_ASAP7_75t_R FILLER_0_95_367 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_379 ();
 FILLER_ASAP7_75t_R FILLER_0_95_385 ();
 FILLER_ASAP7_75t_R FILLER_0_95_393 ();
 DECAPx1_ASAP7_75t_R FILLER_0_95_401 ();
 FILLER_ASAP7_75t_R FILLER_0_95_412 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_420 ();
 FILLER_ASAP7_75t_R FILLER_0_95_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_434 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_448 ();
 FILLER_ASAP7_75t_R FILLER_0_95_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_457 ();
 FILLER_ASAP7_75t_R FILLER_0_95_461 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_475 ();
 FILLER_ASAP7_75t_R FILLER_0_95_486 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_491 ();
 FILLER_ASAP7_75t_R FILLER_0_95_497 ();
 FILLER_ASAP7_75t_R FILLER_0_95_504 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_517 ();
 FILLER_ASAP7_75t_R FILLER_0_95_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_526 ();
 DECAPx1_ASAP7_75t_R FILLER_0_95_535 ();
 FILLER_ASAP7_75t_R FILLER_0_95_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_547 ();
 FILLER_ASAP7_75t_R FILLER_0_95_554 ();
 DECAPx1_ASAP7_75t_R FILLER_0_95_560 ();
 FILLER_ASAP7_75t_R FILLER_0_95_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_576 ();
 FILLER_ASAP7_75t_R FILLER_0_95_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_585 ();
 FILLER_ASAP7_75t_R FILLER_0_95_594 ();
 DECAPx4_ASAP7_75t_R FILLER_0_95_607 ();
 FILLER_ASAP7_75t_R FILLER_0_95_620 ();
 DECAPx1_ASAP7_75t_R FILLER_0_95_628 ();
 FILLER_ASAP7_75t_R FILLER_0_95_642 ();
 DECAPx4_ASAP7_75t_R FILLER_0_95_654 ();
 FILLER_ASAP7_75t_R FILLER_0_95_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_666 ();
 FILLER_ASAP7_75t_R FILLER_0_95_672 ();
 FILLER_ASAP7_75t_R FILLER_0_95_684 ();
 FILLER_ASAP7_75t_R FILLER_0_95_696 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_724 ();
 FILLER_ASAP7_75t_R FILLER_0_95_732 ();
 FILLER_ASAP7_75t_R FILLER_0_95_739 ();
 FILLER_ASAP7_75t_R FILLER_0_95_746 ();
 FILLER_ASAP7_75t_R FILLER_0_95_752 ();
 DECAPx4_ASAP7_75t_R FILLER_0_95_760 ();
 FILLER_ASAP7_75t_R FILLER_0_95_770 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_788 ();
 FILLER_ASAP7_75t_R FILLER_0_95_795 ();
 DECAPx1_ASAP7_75t_R FILLER_0_95_804 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_820 ();
 FILLER_ASAP7_75t_R FILLER_0_95_836 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_844 ();
 FILLER_ASAP7_75t_R FILLER_0_95_850 ();
 DECAPx1_ASAP7_75t_R FILLER_0_95_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_866 ();
 FILLER_ASAP7_75t_R FILLER_0_95_877 ();
 FILLER_ASAP7_75t_R FILLER_0_95_885 ();
 DECAPx1_ASAP7_75t_R FILLER_0_95_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_897 ();
 FILLER_ASAP7_75t_R FILLER_0_95_908 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_916 ();
 FILLER_ASAP7_75t_R FILLER_0_95_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_924 ();
 DECAPx6_ASAP7_75t_R FILLER_0_95_927 ();
 DECAPx1_ASAP7_75t_R FILLER_0_95_941 ();
 DECAPx4_ASAP7_75t_R FILLER_0_95_948 ();
 FILLER_ASAP7_75t_R FILLER_0_95_958 ();
 FILLER_ASAP7_75t_R FILLER_0_95_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_973 ();
 FILLER_ASAP7_75t_R FILLER_0_95_980 ();
 FILLER_ASAP7_75t_R FILLER_0_95_988 ();
 FILLER_ASAP7_75t_R FILLER_0_95_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_998 ();
 FILLER_ASAP7_75t_R FILLER_0_95_1005 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_1014 ();
 DECAPx6_ASAP7_75t_R FILLER_0_95_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_1050 ();
 FILLER_ASAP7_75t_R FILLER_0_95_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_1059 ();
 FILLER_ASAP7_75t_R FILLER_0_95_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_1068 ();
 FILLER_ASAP7_75t_R FILLER_0_95_1075 ();
 DECAPx6_ASAP7_75t_R FILLER_0_95_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_1101 ();
 FILLER_ASAP7_75t_R FILLER_0_95_1108 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_1116 ();
 FILLER_ASAP7_75t_R FILLER_0_95_1144 ();
 DECAPx4_ASAP7_75t_R FILLER_0_95_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_1162 ();
 DECAPx6_ASAP7_75t_R FILLER_0_95_1169 ();
 FILLER_ASAP7_75t_R FILLER_0_95_1189 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_1197 ();
 FILLER_ASAP7_75t_R FILLER_0_95_1203 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_1211 ();
 FILLER_ASAP7_75t_R FILLER_0_95_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_1219 ();
 FILLER_ASAP7_75t_R FILLER_0_95_1226 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_1228 ();
 FILLER_ASAP7_75t_R FILLER_0_95_1236 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_1244 ();
 FILLER_ASAP7_75t_R FILLER_0_95_1250 ();
 FILLER_ASAP7_75t_R FILLER_0_95_1259 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_1268 ();
 FILLER_ASAP7_75t_R FILLER_0_95_1274 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_1282 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_1294 ();
 FILLER_ASAP7_75t_R FILLER_0_95_1300 ();
 FILLER_ASAP7_75t_R FILLER_0_95_1308 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_1321 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_1343 ();
 DECAPx6_ASAP7_75t_R FILLER_0_95_1365 ();
 FILLER_ASAP7_75t_R FILLER_0_95_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_96_2 ();
 FILLER_ASAP7_75t_R FILLER_0_96_9 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_20 ();
 FILLER_ASAP7_75t_R FILLER_0_96_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_28 ();
 FILLER_ASAP7_75t_R FILLER_0_96_32 ();
 FILLER_ASAP7_75t_R FILLER_0_96_40 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_48 ();
 FILLER_ASAP7_75t_R FILLER_0_96_60 ();
 DECAPx2_ASAP7_75t_R FILLER_0_96_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_80 ();
 FILLER_ASAP7_75t_R FILLER_0_96_86 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_94 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_105 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_119 ();
 DECAPx2_ASAP7_75t_R FILLER_0_96_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_136 ();
 FILLER_ASAP7_75t_R FILLER_0_96_145 ();
 FILLER_ASAP7_75t_R FILLER_0_96_153 ();
 FILLER_ASAP7_75t_R FILLER_0_96_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_169 ();
 DECAPx6_ASAP7_75t_R FILLER_0_96_176 ();
 FILLER_ASAP7_75t_R FILLER_0_96_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_192 ();
 FILLER_ASAP7_75t_R FILLER_0_96_209 ();
 FILLER_ASAP7_75t_R FILLER_0_96_217 ();
 FILLER_ASAP7_75t_R FILLER_0_96_225 ();
 FILLER_ASAP7_75t_R FILLER_0_96_233 ();
 FILLER_ASAP7_75t_R FILLER_0_96_245 ();
 DECAPx4_ASAP7_75t_R FILLER_0_96_253 ();
 FILLER_ASAP7_75t_R FILLER_0_96_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_265 ();
 DECAPx6_ASAP7_75t_R FILLER_0_96_269 ();
 FILLER_ASAP7_75t_R FILLER_0_96_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_285 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_296 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_307 ();
 FILLER_ASAP7_75t_R FILLER_0_96_317 ();
 DECAPx6_ASAP7_75t_R FILLER_0_96_326 ();
 FILLER_ASAP7_75t_R FILLER_0_96_346 ();
 FILLER_ASAP7_75t_R FILLER_0_96_358 ();
 FILLER_ASAP7_75t_R FILLER_0_96_370 ();
 FILLER_ASAP7_75t_R FILLER_0_96_378 ();
 FILLER_ASAP7_75t_R FILLER_0_96_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_389 ();
 FILLER_ASAP7_75t_R FILLER_0_96_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_406 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_450 ();
 DECAPx2_ASAP7_75t_R FILLER_0_96_454 ();
 FILLER_ASAP7_75t_R FILLER_0_96_460 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_492 ();
 FILLER_ASAP7_75t_R FILLER_0_96_520 ();
 FILLER_ASAP7_75t_R FILLER_0_96_532 ();
 FILLER_ASAP7_75t_R FILLER_0_96_541 ();
 FILLER_ASAP7_75t_R FILLER_0_96_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_551 ();
 FILLER_ASAP7_75t_R FILLER_0_96_557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_96_570 ();
 FILLER_ASAP7_75t_R FILLER_0_96_576 ();
 FILLER_ASAP7_75t_R FILLER_0_96_584 ();
 FILLER_ASAP7_75t_R FILLER_0_96_592 ();
 FILLER_ASAP7_75t_R FILLER_0_96_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_604 ();
 FILLER_ASAP7_75t_R FILLER_0_96_611 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_633 ();
 FILLER_ASAP7_75t_R FILLER_0_96_643 ();
 DECAPx4_ASAP7_75t_R FILLER_0_96_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_660 ();
 FILLER_ASAP7_75t_R FILLER_0_96_666 ();
 DECAPx2_ASAP7_75t_R FILLER_0_96_689 ();
 FILLER_ASAP7_75t_R FILLER_0_96_695 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_717 ();
 FILLER_ASAP7_75t_R FILLER_0_96_727 ();
 FILLER_ASAP7_75t_R FILLER_0_96_737 ();
 FILLER_ASAP7_75t_R FILLER_0_96_745 ();
 FILLER_ASAP7_75t_R FILLER_0_96_753 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_759 ();
 FILLER_ASAP7_75t_R FILLER_0_96_781 ();
 FILLER_ASAP7_75t_R FILLER_0_96_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_797 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_808 ();
 FILLER_ASAP7_75t_R FILLER_0_96_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_824 ();
 FILLER_ASAP7_75t_R FILLER_0_96_832 ();
 FILLER_ASAP7_75t_R FILLER_0_96_840 ();
 FILLER_ASAP7_75t_R FILLER_0_96_848 ();
 FILLER_ASAP7_75t_R FILLER_0_96_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_862 ();
 FILLER_ASAP7_75t_R FILLER_0_96_868 ();
 FILLER_ASAP7_75t_R FILLER_0_96_878 ();
 FILLER_ASAP7_75t_R FILLER_0_96_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_890 ();
 FILLER_ASAP7_75t_R FILLER_0_96_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_903 ();
 DECAPx2_ASAP7_75t_R FILLER_0_96_910 ();
 FILLER_ASAP7_75t_R FILLER_0_96_916 ();
 FILLER_ASAP7_75t_R FILLER_0_96_924 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_932 ();
 FILLER_ASAP7_75t_R FILLER_0_96_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_956 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_963 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_989 ();
 FILLER_ASAP7_75t_R FILLER_0_96_1000 ();
 DECAPx6_ASAP7_75t_R FILLER_0_96_1005 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_1019 ();
 FILLER_ASAP7_75t_R FILLER_0_96_1043 ();
 FILLER_ASAP7_75t_R FILLER_0_96_1051 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_1060 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_1064 ();
 DECAPx6_ASAP7_75t_R FILLER_0_96_1071 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_1085 ();
 DECAPx2_ASAP7_75t_R FILLER_0_96_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_1101 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_1117 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_1121 ();
 FILLER_ASAP7_75t_R FILLER_0_96_1131 ();
 FILLER_ASAP7_75t_R FILLER_0_96_1140 ();
 DECAPx6_ASAP7_75t_R FILLER_0_96_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_1166 ();
 FILLER_ASAP7_75t_R FILLER_0_96_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_1175 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_1182 ();
 DECAPx6_ASAP7_75t_R FILLER_0_96_1204 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_1218 ();
 FILLER_ASAP7_75t_R FILLER_0_96_1228 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_1236 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_1240 ();
 FILLER_ASAP7_75t_R FILLER_0_96_1261 ();
 FILLER_ASAP7_75t_R FILLER_0_96_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_1271 ();
 FILLER_ASAP7_75t_R FILLER_0_96_1278 ();
 DECAPx2_ASAP7_75t_R FILLER_0_96_1286 ();
 FILLER_ASAP7_75t_R FILLER_0_96_1292 ();
 FILLER_ASAP7_75t_R FILLER_0_96_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_1315 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_1337 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_1359 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_97_2 ();
 FILLER_ASAP7_75t_R FILLER_0_97_10 ();
 FILLER_ASAP7_75t_R FILLER_0_97_18 ();
 DECAPx1_ASAP7_75t_R FILLER_0_97_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_29 ();
 FILLER_ASAP7_75t_R FILLER_0_97_36 ();
 DECAPx2_ASAP7_75t_R FILLER_0_97_44 ();
 FILLER_ASAP7_75t_R FILLER_0_97_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_52 ();
 DECAPx6_ASAP7_75t_R FILLER_0_97_59 ();
 FILLER_ASAP7_75t_R FILLER_0_97_79 ();
 DECAPx2_ASAP7_75t_R FILLER_0_97_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_99 ();
 FILLER_ASAP7_75t_R FILLER_0_97_108 ();
 FILLER_ASAP7_75t_R FILLER_0_97_117 ();
 DECAPx2_ASAP7_75t_R FILLER_0_97_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_131 ();
 FILLER_ASAP7_75t_R FILLER_0_97_142 ();
 FILLER_ASAP7_75t_R FILLER_0_97_154 ();
 DECAPx4_ASAP7_75t_R FILLER_0_97_163 ();
 FILLER_ASAP7_75t_R FILLER_0_97_179 ();
 DECAPx1_ASAP7_75t_R FILLER_0_97_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_189 ();
 DECAPx4_ASAP7_75t_R FILLER_0_97_196 ();
 DECAPx1_ASAP7_75t_R FILLER_0_97_212 ();
 DECAPx2_ASAP7_75t_R FILLER_0_97_224 ();
 FILLER_ASAP7_75t_R FILLER_0_97_230 ();
 DECAPx6_ASAP7_75t_R FILLER_0_97_242 ();
 DECAPx1_ASAP7_75t_R FILLER_0_97_256 ();
 FILLER_ASAP7_75t_R FILLER_0_97_263 ();
 DECAPx6_ASAP7_75t_R FILLER_0_97_273 ();
 DECAPx1_ASAP7_75t_R FILLER_0_97_287 ();
 FILLER_ASAP7_75t_R FILLER_0_97_301 ();
 FILLER_ASAP7_75t_R FILLER_0_97_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_319 ();
 DECAPx2_ASAP7_75t_R FILLER_0_97_326 ();
 FILLER_ASAP7_75t_R FILLER_0_97_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_334 ();
 DECAPx2_ASAP7_75t_R FILLER_0_97_345 ();
 FILLER_ASAP7_75t_R FILLER_0_97_351 ();
 FILLER_ASAP7_75t_R FILLER_0_97_365 ();
 FILLER_ASAP7_75t_R FILLER_0_97_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_375 ();
 DECAPx1_ASAP7_75t_R FILLER_0_97_386 ();
 DECAPx1_ASAP7_75t_R FILLER_0_97_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_400 ();
 DECAPx2_ASAP7_75t_R FILLER_0_97_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_417 ();
 DECAPx1_ASAP7_75t_R FILLER_0_97_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_425 ();
 DECAPx4_ASAP7_75t_R FILLER_0_97_432 ();
 FILLER_ASAP7_75t_R FILLER_0_97_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_454 ();
 DECAPx4_ASAP7_75t_R FILLER_0_97_476 ();
 FILLER_ASAP7_75t_R FILLER_0_97_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_488 ();
 FILLER_ASAP7_75t_R FILLER_0_97_492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_97_500 ();
 FILLER_ASAP7_75t_R FILLER_0_97_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_512 ();
 FILLER_ASAP7_75t_R FILLER_0_97_519 ();
 FILLER_ASAP7_75t_R FILLER_0_97_531 ();
 FILLER_ASAP7_75t_R FILLER_0_97_539 ();
 DECAPx2_ASAP7_75t_R FILLER_0_97_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_553 ();
 DECAPx2_ASAP7_75t_R FILLER_0_97_561 ();
 FILLER_ASAP7_75t_R FILLER_0_97_573 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_581 ();
 FILLER_ASAP7_75t_R FILLER_0_97_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_605 ();
 DECAPx6_ASAP7_75t_R FILLER_0_97_612 ();
 DECAPx2_ASAP7_75t_R FILLER_0_97_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_638 ();
 DECAPx2_ASAP7_75t_R FILLER_0_97_649 ();
 FILLER_ASAP7_75t_R FILLER_0_97_655 ();
 FILLER_ASAP7_75t_R FILLER_0_97_660 ();
 FILLER_ASAP7_75t_R FILLER_0_97_667 ();
 FILLER_ASAP7_75t_R FILLER_0_97_687 ();
 FILLER_ASAP7_75t_R FILLER_0_97_701 ();
 DECAPx2_ASAP7_75t_R FILLER_0_97_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_719 ();
 FILLER_ASAP7_75t_R FILLER_0_97_727 ();
 FILLER_ASAP7_75t_R FILLER_0_97_735 ();
 FILLER_ASAP7_75t_R FILLER_0_97_742 ();
 DECAPx2_ASAP7_75t_R FILLER_0_97_749 ();
 FILLER_ASAP7_75t_R FILLER_0_97_755 ();
 FILLER_ASAP7_75t_R FILLER_0_97_767 ();
 FILLER_ASAP7_75t_R FILLER_0_97_789 ();
 FILLER_ASAP7_75t_R FILLER_0_97_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_799 ();
 FILLER_ASAP7_75t_R FILLER_0_97_806 ();
 FILLER_ASAP7_75t_R FILLER_0_97_814 ();
 FILLER_ASAP7_75t_R FILLER_0_97_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_838 ();
 DECAPx2_ASAP7_75t_R FILLER_0_97_849 ();
 FILLER_ASAP7_75t_R FILLER_0_97_879 ();
 DECAPx2_ASAP7_75t_R FILLER_0_97_891 ();
 FILLER_ASAP7_75t_R FILLER_0_97_897 ();
 DECAPx6_ASAP7_75t_R FILLER_0_97_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_924 ();
 DECAPx6_ASAP7_75t_R FILLER_0_97_927 ();
 DECAPx2_ASAP7_75t_R FILLER_0_97_941 ();
 FILLER_ASAP7_75t_R FILLER_0_97_957 ();
 DECAPx2_ASAP7_75t_R FILLER_0_97_965 ();
 FILLER_ASAP7_75t_R FILLER_0_97_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_983 ();
 DECAPx2_ASAP7_75t_R FILLER_0_97_990 ();
 FILLER_ASAP7_75t_R FILLER_0_97_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_998 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_1007 ();
 DECAPx4_ASAP7_75t_R FILLER_0_97_1014 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1024 ();
 DECAPx4_ASAP7_75t_R FILLER_0_97_1036 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1046 ();
 DECAPx1_ASAP7_75t_R FILLER_0_97_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_1058 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1065 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_1075 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_0_97_1090 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1104 ();
 DECAPx1_ASAP7_75t_R FILLER_0_97_1112 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1122 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1130 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_1157 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1164 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1172 ();
 DECAPx6_ASAP7_75t_R FILLER_0_97_1180 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_1196 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1207 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1219 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1227 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1235 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1244 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1252 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1260 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1268 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1276 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1284 ();
 DECAPx2_ASAP7_75t_R FILLER_0_97_1291 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_1305 ();
 DECAPx4_ASAP7_75t_R FILLER_0_97_1327 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1337 ();
 FILLER_ASAP7_75t_R FILLER_0_97_1345 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_1350 ();
 DECAPx4_ASAP7_75t_R FILLER_0_97_1372 ();
 FILLER_ASAP7_75t_R FILLER_0_98_2 ();
 FILLER_ASAP7_75t_R FILLER_0_98_25 ();
 FILLER_ASAP7_75t_R FILLER_0_98_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_32 ();
 FILLER_ASAP7_75t_R FILLER_0_98_43 ();
 DECAPx1_ASAP7_75t_R FILLER_0_98_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_54 ();
 DECAPx4_ASAP7_75t_R FILLER_0_98_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_88 ();
 FILLER_ASAP7_75t_R FILLER_0_98_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_112 ();
 FILLER_ASAP7_75t_R FILLER_0_98_119 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_131 ();
 FILLER_ASAP7_75t_R FILLER_0_98_153 ();
 DECAPx2_ASAP7_75t_R FILLER_0_98_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_173 ();
 FILLER_ASAP7_75t_R FILLER_0_98_180 ();
 DECAPx2_ASAP7_75t_R FILLER_0_98_192 ();
 DECAPx2_ASAP7_75t_R FILLER_0_98_204 ();
 FILLER_ASAP7_75t_R FILLER_0_98_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_212 ();
 FILLER_ASAP7_75t_R FILLER_0_98_218 ();
 DECAPx1_ASAP7_75t_R FILLER_0_98_228 ();
 FILLER_ASAP7_75t_R FILLER_0_98_242 ();
 DECAPx1_ASAP7_75t_R FILLER_0_98_254 ();
 FILLER_ASAP7_75t_R FILLER_0_98_269 ();
 DECAPx6_ASAP7_75t_R FILLER_0_98_277 ();
 DECAPx1_ASAP7_75t_R FILLER_0_98_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_295 ();
 FILLER_ASAP7_75t_R FILLER_0_98_305 ();
 FILLER_ASAP7_75t_R FILLER_0_98_312 ();
 DECAPx1_ASAP7_75t_R FILLER_0_98_317 ();
 FILLER_ASAP7_75t_R FILLER_0_98_328 ();
 DECAPx4_ASAP7_75t_R FILLER_0_98_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_346 ();
 FILLER_ASAP7_75t_R FILLER_0_98_352 ();
 FILLER_ASAP7_75t_R FILLER_0_98_378 ();
 DECAPx2_ASAP7_75t_R FILLER_0_98_383 ();
 DECAPx6_ASAP7_75t_R FILLER_0_98_395 ();
 DECAPx2_ASAP7_75t_R FILLER_0_98_409 ();
 DECAPx2_ASAP7_75t_R FILLER_0_98_421 ();
 FILLER_ASAP7_75t_R FILLER_0_98_427 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_436 ();
 DECAPx1_ASAP7_75t_R FILLER_0_98_458 ();
 FILLER_ASAP7_75t_R FILLER_0_98_464 ();
 FILLER_ASAP7_75t_R FILLER_0_98_469 ();
 FILLER_ASAP7_75t_R FILLER_0_98_491 ();
 FILLER_ASAP7_75t_R FILLER_0_98_499 ();
 DECAPx2_ASAP7_75t_R FILLER_0_98_507 ();
 DECAPx1_ASAP7_75t_R FILLER_0_98_519 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_523 ();
 DECAPx2_ASAP7_75t_R FILLER_0_98_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_540 ();
 FILLER_ASAP7_75t_R FILLER_0_98_549 ();
 FILLER_ASAP7_75t_R FILLER_0_98_556 ();
 FILLER_ASAP7_75t_R FILLER_0_98_564 ();
 DECAPx6_ASAP7_75t_R FILLER_0_98_572 ();
 FILLER_ASAP7_75t_R FILLER_0_98_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_588 ();
 FILLER_ASAP7_75t_R FILLER_0_98_595 ();
 DECAPx1_ASAP7_75t_R FILLER_0_98_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_607 ();
 FILLER_ASAP7_75t_R FILLER_0_98_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_617 ();
 FILLER_ASAP7_75t_R FILLER_0_98_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_630 ();
 FILLER_ASAP7_75t_R FILLER_0_98_637 ();
 DECAPx4_ASAP7_75t_R FILLER_0_98_645 ();
 FILLER_ASAP7_75t_R FILLER_0_98_655 ();
 FILLER_ASAP7_75t_R FILLER_0_98_662 ();
 FILLER_ASAP7_75t_R FILLER_0_98_674 ();
 DECAPx1_ASAP7_75t_R FILLER_0_98_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_700 ();
 FILLER_ASAP7_75t_R FILLER_0_98_707 ();
 FILLER_ASAP7_75t_R FILLER_0_98_715 ();
 DECAPx1_ASAP7_75t_R FILLER_0_98_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_727 ();
 FILLER_ASAP7_75t_R FILLER_0_98_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_735 ();
 DECAPx1_ASAP7_75t_R FILLER_0_98_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_750 ();
 DECAPx1_ASAP7_75t_R FILLER_0_98_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_761 ();
 FILLER_ASAP7_75t_R FILLER_0_98_772 ();
 DECAPx2_ASAP7_75t_R FILLER_0_98_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_787 ();
 DECAPx2_ASAP7_75t_R FILLER_0_98_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_800 ();
 FILLER_ASAP7_75t_R FILLER_0_98_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_813 ();
 FILLER_ASAP7_75t_R FILLER_0_98_820 ();
 DECAPx2_ASAP7_75t_R FILLER_0_98_832 ();
 FILLER_ASAP7_75t_R FILLER_0_98_838 ();
 DECAPx2_ASAP7_75t_R FILLER_0_98_850 ();
 FILLER_ASAP7_75t_R FILLER_0_98_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_858 ();
 FILLER_ASAP7_75t_R FILLER_0_98_863 ();
 DECAPx6_ASAP7_75t_R FILLER_0_98_872 ();
 DECAPx6_ASAP7_75t_R FILLER_0_98_897 ();
 DECAPx2_ASAP7_75t_R FILLER_0_98_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_917 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_924 ();
 FILLER_ASAP7_75t_R FILLER_0_98_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_948 ();
 DECAPx2_ASAP7_75t_R FILLER_0_98_955 ();
 FILLER_ASAP7_75t_R FILLER_0_98_981 ();
 DECAPx2_ASAP7_75t_R FILLER_0_98_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_999 ();
 FILLER_ASAP7_75t_R FILLER_0_98_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_1009 ();
 DECAPx1_ASAP7_75t_R FILLER_0_98_1021 ();
 FILLER_ASAP7_75t_R FILLER_0_98_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_1047 ();
 DECAPx1_ASAP7_75t_R FILLER_0_98_1054 ();
 FILLER_ASAP7_75t_R FILLER_0_98_1068 ();
 DECAPx2_ASAP7_75t_R FILLER_0_98_1076 ();
 FILLER_ASAP7_75t_R FILLER_0_98_1082 ();
 DECAPx6_ASAP7_75t_R FILLER_0_98_1089 ();
 DECAPx2_ASAP7_75t_R FILLER_0_98_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_1115 ();
 FILLER_ASAP7_75t_R FILLER_0_98_1121 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_1129 ();
 FILLER_ASAP7_75t_R FILLER_0_98_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_1153 ();
 DECAPx1_ASAP7_75t_R FILLER_0_98_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_1175 ();
 FILLER_ASAP7_75t_R FILLER_0_98_1197 ();
 FILLER_ASAP7_75t_R FILLER_0_98_1219 ();
 DECAPx2_ASAP7_75t_R FILLER_0_98_1241 ();
 FILLER_ASAP7_75t_R FILLER_0_98_1247 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_1249 ();
 DECAPx2_ASAP7_75t_R FILLER_0_98_1260 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_1266 ();
 FILLER_ASAP7_75t_R FILLER_0_98_1273 ();
 FILLER_ASAP7_75t_R FILLER_0_98_1281 ();
 DECAPx4_ASAP7_75t_R FILLER_0_98_1291 ();
 FILLER_ASAP7_75t_R FILLER_0_98_1301 ();
 FILLER_ASAP7_75t_R FILLER_0_98_1309 ();
 FILLER_ASAP7_75t_R FILLER_0_98_1321 ();
 FILLER_ASAP7_75t_R FILLER_0_98_1329 ();
 FILLER_ASAP7_75t_R FILLER_0_98_1337 ();
 FILLER_ASAP7_75t_R FILLER_0_98_1345 ();
 FILLER_ASAP7_75t_R FILLER_0_98_1353 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_1358 ();
 FILLER_ASAP7_75t_R FILLER_0_98_1380 ();
 DECAPx2_ASAP7_75t_R FILLER_0_99_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_13 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_27 ();
 FILLER_ASAP7_75t_R FILLER_0_99_38 ();
 DECAPx4_ASAP7_75t_R FILLER_0_99_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_58 ();
 DECAPx6_ASAP7_75t_R FILLER_0_99_65 ();
 FILLER_ASAP7_75t_R FILLER_0_99_79 ();
 DECAPx2_ASAP7_75t_R FILLER_0_99_87 ();
 FILLER_ASAP7_75t_R FILLER_0_99_99 ();
 FILLER_ASAP7_75t_R FILLER_0_99_107 ();
 DECAPx4_ASAP7_75t_R FILLER_0_99_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_125 ();
 DECAPx2_ASAP7_75t_R FILLER_0_99_134 ();
 FILLER_ASAP7_75t_R FILLER_0_99_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_142 ();
 DECAPx4_ASAP7_75t_R FILLER_0_99_148 ();
 DECAPx4_ASAP7_75t_R FILLER_0_99_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_173 ();
 FILLER_ASAP7_75t_R FILLER_0_99_181 ();
 DECAPx2_ASAP7_75t_R FILLER_0_99_189 ();
 FILLER_ASAP7_75t_R FILLER_0_99_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_197 ();
 FILLER_ASAP7_75t_R FILLER_0_99_205 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_213 ();
 DECAPx2_ASAP7_75t_R FILLER_0_99_223 ();
 FILLER_ASAP7_75t_R FILLER_0_99_229 ();
 FILLER_ASAP7_75t_R FILLER_0_99_241 ();
 DECAPx6_ASAP7_75t_R FILLER_0_99_253 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_267 ();
 DECAPx6_ASAP7_75t_R FILLER_0_99_292 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_306 ();
 DECAPx2_ASAP7_75t_R FILLER_0_99_317 ();
 FILLER_ASAP7_75t_R FILLER_0_99_323 ();
 DECAPx6_ASAP7_75t_R FILLER_0_99_331 ();
 FILLER_ASAP7_75t_R FILLER_0_99_345 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_354 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_372 ();
 FILLER_ASAP7_75t_R FILLER_0_99_379 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_387 ();
 DECAPx4_ASAP7_75t_R FILLER_0_99_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_408 ();
 DECAPx2_ASAP7_75t_R FILLER_0_99_412 ();
 FILLER_ASAP7_75t_R FILLER_0_99_424 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_432 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_447 ();
 FILLER_ASAP7_75t_R FILLER_0_99_457 ();
 FILLER_ASAP7_75t_R FILLER_0_99_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_464 ();
 DECAPx2_ASAP7_75t_R FILLER_0_99_471 ();
 FILLER_ASAP7_75t_R FILLER_0_99_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_479 ();
 DECAPx2_ASAP7_75t_R FILLER_0_99_490 ();
 DECAPx6_ASAP7_75t_R FILLER_0_99_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_516 ();
 FILLER_ASAP7_75t_R FILLER_0_99_522 ();
 FILLER_ASAP7_75t_R FILLER_0_99_534 ();
 FILLER_ASAP7_75t_R FILLER_0_99_547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_559 ();
 FILLER_ASAP7_75t_R FILLER_0_99_566 ();
 DECAPx6_ASAP7_75t_R FILLER_0_99_574 ();
 FILLER_ASAP7_75t_R FILLER_0_99_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_596 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_607 ();
 FILLER_ASAP7_75t_R FILLER_0_99_614 ();
 FILLER_ASAP7_75t_R FILLER_0_99_619 ();
 FILLER_ASAP7_75t_R FILLER_0_99_627 ();
 FILLER_ASAP7_75t_R FILLER_0_99_635 ();
 DECAPx4_ASAP7_75t_R FILLER_0_99_643 ();
 FILLER_ASAP7_75t_R FILLER_0_99_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_655 ();
 FILLER_ASAP7_75t_R FILLER_0_99_661 ();
 FILLER_ASAP7_75t_R FILLER_0_99_673 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_683 ();
 FILLER_ASAP7_75t_R FILLER_0_99_697 ();
 FILLER_ASAP7_75t_R FILLER_0_99_706 ();
 FILLER_ASAP7_75t_R FILLER_0_99_714 ();
 FILLER_ASAP7_75t_R FILLER_0_99_721 ();
 FILLER_ASAP7_75t_R FILLER_0_99_733 ();
 FILLER_ASAP7_75t_R FILLER_0_99_747 ();
 FILLER_ASAP7_75t_R FILLER_0_99_755 ();
 FILLER_ASAP7_75t_R FILLER_0_99_762 ();
 FILLER_ASAP7_75t_R FILLER_0_99_770 ();
 DECAPx2_ASAP7_75t_R FILLER_0_99_778 ();
 FILLER_ASAP7_75t_R FILLER_0_99_784 ();
 FILLER_ASAP7_75t_R FILLER_0_99_796 ();
 FILLER_ASAP7_75t_R FILLER_0_99_803 ();
 FILLER_ASAP7_75t_R FILLER_0_99_811 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_822 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_843 ();
 DECAPx2_ASAP7_75t_R FILLER_0_99_857 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_869 ();
 DECAPx2_ASAP7_75t_R FILLER_0_99_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_99_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_903 ();
 DECAPx2_ASAP7_75t_R FILLER_0_99_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_916 ();
 FILLER_ASAP7_75t_R FILLER_0_99_923 ();
 FILLER_ASAP7_75t_R FILLER_0_99_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_929 ();
 DECAPx2_ASAP7_75t_R FILLER_0_99_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_942 ();
 FILLER_ASAP7_75t_R FILLER_0_99_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_948 ();
 FILLER_ASAP7_75t_R FILLER_0_99_955 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_963 ();
 FILLER_ASAP7_75t_R FILLER_0_99_978 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_990 ();
 DECAPx4_ASAP7_75t_R FILLER_0_99_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_1007 ();
 FILLER_ASAP7_75t_R FILLER_0_99_1014 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_1023 ();
 FILLER_ASAP7_75t_R FILLER_0_99_1032 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_1044 ();
 DECAPx2_ASAP7_75t_R FILLER_0_99_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_1057 ();
 DECAPx6_ASAP7_75t_R FILLER_0_99_1064 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_0_99_1093 ();
 FILLER_ASAP7_75t_R FILLER_0_99_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_1101 ();
 DECAPx4_ASAP7_75t_R FILLER_0_99_1108 ();
 FILLER_ASAP7_75t_R FILLER_0_99_1118 ();
 FILLER_ASAP7_75t_R FILLER_0_99_1126 ();
 DECAPx4_ASAP7_75t_R FILLER_0_99_1134 ();
 FILLER_ASAP7_75t_R FILLER_0_99_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_1146 ();
 FILLER_ASAP7_75t_R FILLER_0_99_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_1155 ();
 DECAPx4_ASAP7_75t_R FILLER_0_99_1163 ();
 FILLER_ASAP7_75t_R FILLER_0_99_1179 ();
 FILLER_ASAP7_75t_R FILLER_0_99_1187 ();
 DECAPx6_ASAP7_75t_R FILLER_0_99_1209 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_1223 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_1233 ();
 DECAPx2_ASAP7_75t_R FILLER_0_99_1247 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_1253 ();
 FILLER_ASAP7_75t_R FILLER_0_99_1274 ();
 FILLER_ASAP7_75t_R FILLER_0_99_1290 ();
 FILLER_ASAP7_75t_R FILLER_0_99_1298 ();
 DECAPx2_ASAP7_75t_R FILLER_0_99_1306 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_1312 ();
 FILLER_ASAP7_75t_R FILLER_0_99_1323 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_1325 ();
 DECAPx2_ASAP7_75t_R FILLER_0_99_1332 ();
 FILLER_ASAP7_75t_R FILLER_0_99_1338 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_1340 ();
 FILLER_ASAP7_75t_R FILLER_0_99_1347 ();
 DECAPx6_ASAP7_75t_R FILLER_0_99_1352 ();
 DECAPx2_ASAP7_75t_R FILLER_0_99_1366 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_1372 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_1378 ();
 DECAPx2_ASAP7_75t_R FILLER_0_100_2 ();
 FILLER_ASAP7_75t_R FILLER_0_100_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_100_50 ();
 FILLER_ASAP7_75t_R FILLER_0_100_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_66 ();
 FILLER_ASAP7_75t_R FILLER_0_100_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_75 ();
 DECAPx6_ASAP7_75t_R FILLER_0_100_82 ();
 DECAPx1_ASAP7_75t_R FILLER_0_100_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_111 ();
 DECAPx4_ASAP7_75t_R FILLER_0_100_120 ();
 FILLER_ASAP7_75t_R FILLER_0_100_130 ();
 FILLER_ASAP7_75t_R FILLER_0_100_139 ();
 FILLER_ASAP7_75t_R FILLER_0_100_148 ();
 DECAPx1_ASAP7_75t_R FILLER_0_100_160 ();
 DECAPx2_ASAP7_75t_R FILLER_0_100_170 ();
 FILLER_ASAP7_75t_R FILLER_0_100_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_178 ();
 DECAPx1_ASAP7_75t_R FILLER_0_100_185 ();
 DECAPx1_ASAP7_75t_R FILLER_0_100_196 ();
 DECAPx1_ASAP7_75t_R FILLER_0_100_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_215 ();
 DECAPx1_ASAP7_75t_R FILLER_0_100_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_230 ();
 DECAPx1_ASAP7_75t_R FILLER_0_100_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_245 ();
 FILLER_ASAP7_75t_R FILLER_0_100_256 ();
 FILLER_ASAP7_75t_R FILLER_0_100_265 ();
 DECAPx1_ASAP7_75t_R FILLER_0_100_277 ();
 DECAPx4_ASAP7_75t_R FILLER_0_100_291 ();
 DECAPx4_ASAP7_75t_R FILLER_0_100_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_317 ();
 FILLER_ASAP7_75t_R FILLER_0_100_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_323 ();
 FILLER_ASAP7_75t_R FILLER_0_100_344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_100_352 ();
 DECAPx1_ASAP7_75t_R FILLER_0_100_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_370 ();
 DECAPx1_ASAP7_75t_R FILLER_0_100_379 ();
 FILLER_ASAP7_75t_R FILLER_0_100_389 ();
 DECAPx4_ASAP7_75t_R FILLER_0_100_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_407 ();
 DECAPx4_ASAP7_75t_R FILLER_0_100_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_425 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_434 ();
 DECAPx2_ASAP7_75t_R FILLER_0_100_456 ();
 DECAPx4_ASAP7_75t_R FILLER_0_100_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_474 ();
 FILLER_ASAP7_75t_R FILLER_0_100_481 ();
 FILLER_ASAP7_75t_R FILLER_0_100_486 ();
 FILLER_ASAP7_75t_R FILLER_0_100_494 ();
 FILLER_ASAP7_75t_R FILLER_0_100_502 ();
 DECAPx1_ASAP7_75t_R FILLER_0_100_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_514 ();
 FILLER_ASAP7_75t_R FILLER_0_100_520 ();
 FILLER_ASAP7_75t_R FILLER_0_100_527 ();
 DECAPx2_ASAP7_75t_R FILLER_0_100_534 ();
 FILLER_ASAP7_75t_R FILLER_0_100_546 ();
 FILLER_ASAP7_75t_R FILLER_0_100_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_555 ();
 FILLER_ASAP7_75t_R FILLER_0_100_561 ();
 FILLER_ASAP7_75t_R FILLER_0_100_568 ();
 DECAPx4_ASAP7_75t_R FILLER_0_100_573 ();
 FILLER_ASAP7_75t_R FILLER_0_100_590 ();
 FILLER_ASAP7_75t_R FILLER_0_100_602 ();
 FILLER_ASAP7_75t_R FILLER_0_100_610 ();
 DECAPx1_ASAP7_75t_R FILLER_0_100_617 ();
 FILLER_ASAP7_75t_R FILLER_0_100_626 ();
 FILLER_ASAP7_75t_R FILLER_0_100_634 ();
 FILLER_ASAP7_75t_R FILLER_0_100_641 ();
 FILLER_ASAP7_75t_R FILLER_0_100_649 ();
 FILLER_ASAP7_75t_R FILLER_0_100_655 ();
 FILLER_ASAP7_75t_R FILLER_0_100_662 ();
 FILLER_ASAP7_75t_R FILLER_0_100_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_676 ();
 FILLER_ASAP7_75t_R FILLER_0_100_683 ();
 FILLER_ASAP7_75t_R FILLER_0_100_709 ();
 FILLER_ASAP7_75t_R FILLER_0_100_716 ();
 FILLER_ASAP7_75t_R FILLER_0_100_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_100_736 ();
 FILLER_ASAP7_75t_R FILLER_0_100_752 ();
 DECAPx1_ASAP7_75t_R FILLER_0_100_759 ();
 DECAPx4_ASAP7_75t_R FILLER_0_100_773 ();
 FILLER_ASAP7_75t_R FILLER_0_100_783 ();
 DECAPx6_ASAP7_75t_R FILLER_0_100_792 ();
 FILLER_ASAP7_75t_R FILLER_0_100_816 ();
 DECAPx1_ASAP7_75t_R FILLER_0_100_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_825 ();
 FILLER_ASAP7_75t_R FILLER_0_100_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_834 ();
 FILLER_ASAP7_75t_R FILLER_0_100_845 ();
 DECAPx1_ASAP7_75t_R FILLER_0_100_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_857 ();
 FILLER_ASAP7_75t_R FILLER_0_100_869 ();
 DECAPx2_ASAP7_75t_R FILLER_0_100_877 ();
 FILLER_ASAP7_75t_R FILLER_0_100_883 ();
 FILLER_ASAP7_75t_R FILLER_0_100_891 ();
 FILLER_ASAP7_75t_R FILLER_0_100_896 ();
 FILLER_ASAP7_75t_R FILLER_0_100_904 ();
 FILLER_ASAP7_75t_R FILLER_0_100_912 ();
 FILLER_ASAP7_75t_R FILLER_0_100_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_922 ();
 DECAPx6_ASAP7_75t_R FILLER_0_100_929 ();
 FILLER_ASAP7_75t_R FILLER_0_100_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_945 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_957 ();
 DECAPx2_ASAP7_75t_R FILLER_0_100_979 ();
 FILLER_ASAP7_75t_R FILLER_0_100_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_987 ();
 FILLER_ASAP7_75t_R FILLER_0_100_994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_1002 ();
 DECAPx2_ASAP7_75t_R FILLER_0_100_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_1030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_1041 ();
 DECAPx2_ASAP7_75t_R FILLER_0_100_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_1069 ();
 DECAPx1_ASAP7_75t_R FILLER_0_100_1076 ();
 DECAPx4_ASAP7_75t_R FILLER_0_100_1084 ();
 FILLER_ASAP7_75t_R FILLER_0_100_1100 ();
 DECAPx4_ASAP7_75t_R FILLER_0_100_1108 ();
 FILLER_ASAP7_75t_R FILLER_0_100_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_1120 ();
 FILLER_ASAP7_75t_R FILLER_0_100_1128 ();
 FILLER_ASAP7_75t_R FILLER_0_100_1141 ();
 FILLER_ASAP7_75t_R FILLER_0_100_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_1151 ();
 DECAPx4_ASAP7_75t_R FILLER_0_100_1158 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_1168 ();
 DECAPx6_ASAP7_75t_R FILLER_0_100_1179 ();
 FILLER_ASAP7_75t_R FILLER_0_100_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_1201 ();
 DECAPx6_ASAP7_75t_R FILLER_0_100_1208 ();
 FILLER_ASAP7_75t_R FILLER_0_100_1229 ();
 FILLER_ASAP7_75t_R FILLER_0_100_1236 ();
 FILLER_ASAP7_75t_R FILLER_0_100_1245 ();
 DECAPx2_ASAP7_75t_R FILLER_0_100_1253 ();
 FILLER_ASAP7_75t_R FILLER_0_100_1265 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_1267 ();
 FILLER_ASAP7_75t_R FILLER_0_100_1275 ();
 DECAPx1_ASAP7_75t_R FILLER_0_100_1283 ();
 FILLER_ASAP7_75t_R FILLER_0_100_1311 ();
 FILLER_ASAP7_75t_R FILLER_0_100_1319 ();
 DECAPx1_ASAP7_75t_R FILLER_0_100_1327 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_1331 ();
 DECAPx6_ASAP7_75t_R FILLER_0_100_1338 ();
 DECAPx1_ASAP7_75t_R FILLER_0_100_1352 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_1356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_1360 ();
 FILLER_ASAP7_75t_R FILLER_0_101_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_4 ();
 FILLER_ASAP7_75t_R FILLER_0_101_8 ();
 FILLER_ASAP7_75t_R FILLER_0_101_16 ();
 DECAPx2_ASAP7_75t_R FILLER_0_101_28 ();
 FILLER_ASAP7_75t_R FILLER_0_101_34 ();
 FILLER_ASAP7_75t_R FILLER_0_101_44 ();
 FILLER_ASAP7_75t_R FILLER_0_101_51 ();
 DECAPx4_ASAP7_75t_R FILLER_0_101_64 ();
 FILLER_ASAP7_75t_R FILLER_0_101_74 ();
 DECAPx4_ASAP7_75t_R FILLER_0_101_87 ();
 FILLER_ASAP7_75t_R FILLER_0_101_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_99 ();
 FILLER_ASAP7_75t_R FILLER_0_101_106 ();
 FILLER_ASAP7_75t_R FILLER_0_101_118 ();
 DECAPx2_ASAP7_75t_R FILLER_0_101_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_129 ();
 FILLER_ASAP7_75t_R FILLER_0_101_137 ();
 DECAPx1_ASAP7_75t_R FILLER_0_101_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_149 ();
 FILLER_ASAP7_75t_R FILLER_0_101_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_158 ();
 DECAPx1_ASAP7_75t_R FILLER_0_101_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_169 ();
 DECAPx4_ASAP7_75t_R FILLER_0_101_185 ();
 DECAPx4_ASAP7_75t_R FILLER_0_101_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_215 ();
 DECAPx1_ASAP7_75t_R FILLER_0_101_222 ();
 DECAPx6_ASAP7_75t_R FILLER_0_101_232 ();
 DECAPx1_ASAP7_75t_R FILLER_0_101_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_250 ();
 FILLER_ASAP7_75t_R FILLER_0_101_261 ();
 FILLER_ASAP7_75t_R FILLER_0_101_273 ();
 FILLER_ASAP7_75t_R FILLER_0_101_279 ();
 DECAPx4_ASAP7_75t_R FILLER_0_101_284 ();
 FILLER_ASAP7_75t_R FILLER_0_101_308 ();
 FILLER_ASAP7_75t_R FILLER_0_101_316 ();
 FILLER_ASAP7_75t_R FILLER_0_101_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_326 ();
 FILLER_ASAP7_75t_R FILLER_0_101_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_335 ();
 FILLER_ASAP7_75t_R FILLER_0_101_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_366 ();
 FILLER_ASAP7_75t_R FILLER_0_101_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_375 ();
 DECAPx1_ASAP7_75t_R FILLER_0_101_385 ();
 FILLER_ASAP7_75t_R FILLER_0_101_395 ();
 FILLER_ASAP7_75t_R FILLER_0_101_408 ();
 FILLER_ASAP7_75t_R FILLER_0_101_418 ();
 DECAPx1_ASAP7_75t_R FILLER_0_101_426 ();
 FILLER_ASAP7_75t_R FILLER_0_101_436 ();
 DECAPx2_ASAP7_75t_R FILLER_0_101_458 ();
 FILLER_ASAP7_75t_R FILLER_0_101_464 ();
 FILLER_ASAP7_75t_R FILLER_0_101_472 ();
 DECAPx6_ASAP7_75t_R FILLER_0_101_480 ();
 DECAPx1_ASAP7_75t_R FILLER_0_101_494 ();
 DECAPx6_ASAP7_75t_R FILLER_0_101_503 ();
 DECAPx1_ASAP7_75t_R FILLER_0_101_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_521 ();
 FILLER_ASAP7_75t_R FILLER_0_101_528 ();
 DECAPx1_ASAP7_75t_R FILLER_0_101_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_540 ();
 FILLER_ASAP7_75t_R FILLER_0_101_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_551 ();
 DECAPx1_ASAP7_75t_R FILLER_0_101_558 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_562 ();
 DECAPx2_ASAP7_75t_R FILLER_0_101_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_575 ();
 FILLER_ASAP7_75t_R FILLER_0_101_582 ();
 FILLER_ASAP7_75t_R FILLER_0_101_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_592 ();
 DECAPx2_ASAP7_75t_R FILLER_0_101_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_606 ();
 FILLER_ASAP7_75t_R FILLER_0_101_617 ();
 DECAPx2_ASAP7_75t_R FILLER_0_101_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_633 ();
 FILLER_ASAP7_75t_R FILLER_0_101_640 ();
 FILLER_ASAP7_75t_R FILLER_0_101_652 ();
 DECAPx2_ASAP7_75t_R FILLER_0_101_659 ();
 FILLER_ASAP7_75t_R FILLER_0_101_670 ();
 FILLER_ASAP7_75t_R FILLER_0_101_678 ();
 FILLER_ASAP7_75t_R FILLER_0_101_690 ();
 FILLER_ASAP7_75t_R FILLER_0_101_702 ();
 FILLER_ASAP7_75t_R FILLER_0_101_714 ();
 FILLER_ASAP7_75t_R FILLER_0_101_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_726 ();
 DECAPx2_ASAP7_75t_R FILLER_0_101_733 ();
 FILLER_ASAP7_75t_R FILLER_0_101_739 ();
 FILLER_ASAP7_75t_R FILLER_0_101_747 ();
 FILLER_ASAP7_75t_R FILLER_0_101_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_757 ();
 FILLER_ASAP7_75t_R FILLER_0_101_778 ();
 DECAPx6_ASAP7_75t_R FILLER_0_101_788 ();
 FILLER_ASAP7_75t_R FILLER_0_101_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_804 ();
 FILLER_ASAP7_75t_R FILLER_0_101_811 ();
 FILLER_ASAP7_75t_R FILLER_0_101_819 ();
 DECAPx2_ASAP7_75t_R FILLER_0_101_824 ();
 FILLER_ASAP7_75t_R FILLER_0_101_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_832 ();
 FILLER_ASAP7_75t_R FILLER_0_101_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_841 ();
 DECAPx4_ASAP7_75t_R FILLER_0_101_848 ();
 FILLER_ASAP7_75t_R FILLER_0_101_858 ();
 FILLER_ASAP7_75t_R FILLER_0_101_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_872 ();
 FILLER_ASAP7_75t_R FILLER_0_101_883 ();
 DECAPx6_ASAP7_75t_R FILLER_0_101_895 ();
 DECAPx4_ASAP7_75t_R FILLER_0_101_915 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_927 ();
 FILLER_ASAP7_75t_R FILLER_0_101_949 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_957 ();
 DECAPx6_ASAP7_75t_R FILLER_0_101_979 ();
 DECAPx1_ASAP7_75t_R FILLER_0_101_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_997 ();
 DECAPx1_ASAP7_75t_R FILLER_0_101_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_1013 ();
 FILLER_ASAP7_75t_R FILLER_0_101_1020 ();
 FILLER_ASAP7_75t_R FILLER_0_101_1029 ();
 DECAPx6_ASAP7_75t_R FILLER_0_101_1037 ();
 DECAPx1_ASAP7_75t_R FILLER_0_101_1051 ();
 DECAPx2_ASAP7_75t_R FILLER_0_101_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_1068 ();
 FILLER_ASAP7_75t_R FILLER_0_101_1075 ();
 DECAPx1_ASAP7_75t_R FILLER_0_101_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_1087 ();
 DECAPx4_ASAP7_75t_R FILLER_0_101_1094 ();
 DECAPx4_ASAP7_75t_R FILLER_0_101_1110 ();
 FILLER_ASAP7_75t_R FILLER_0_101_1126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_1156 ();
 DECAPx4_ASAP7_75t_R FILLER_0_101_1178 ();
 DECAPx2_ASAP7_75t_R FILLER_0_101_1195 ();
 FILLER_ASAP7_75t_R FILLER_0_101_1201 ();
 DECAPx4_ASAP7_75t_R FILLER_0_101_1211 ();
 FILLER_ASAP7_75t_R FILLER_0_101_1221 ();
 FILLER_ASAP7_75t_R FILLER_0_101_1229 ();
 FILLER_ASAP7_75t_R FILLER_0_101_1237 ();
 FILLER_ASAP7_75t_R FILLER_0_101_1245 ();
 DECAPx4_ASAP7_75t_R FILLER_0_101_1252 ();
 FILLER_ASAP7_75t_R FILLER_0_101_1268 ();
 FILLER_ASAP7_75t_R FILLER_0_101_1276 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_1283 ();
 DECAPx6_ASAP7_75t_R FILLER_0_101_1305 ();
 FILLER_ASAP7_75t_R FILLER_0_101_1319 ();
 DECAPx2_ASAP7_75t_R FILLER_0_101_1324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_1336 ();
 FILLER_ASAP7_75t_R FILLER_0_101_1358 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_1360 ();
 DECAPx6_ASAP7_75t_R FILLER_0_101_1366 ();
 FILLER_ASAP7_75t_R FILLER_0_101_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_102_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_9 ();
 FILLER_ASAP7_75t_R FILLER_0_102_20 ();
 DECAPx1_ASAP7_75t_R FILLER_0_102_32 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_48 ();
 DECAPx1_ASAP7_75t_R FILLER_0_102_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_59 ();
 FILLER_ASAP7_75t_R FILLER_0_102_63 ();
 FILLER_ASAP7_75t_R FILLER_0_102_71 ();
 FILLER_ASAP7_75t_R FILLER_0_102_80 ();
 FILLER_ASAP7_75t_R FILLER_0_102_88 ();
 DECAPx1_ASAP7_75t_R FILLER_0_102_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_100 ();
 DECAPx6_ASAP7_75t_R FILLER_0_102_107 ();
 FILLER_ASAP7_75t_R FILLER_0_102_121 ();
 DECAPx4_ASAP7_75t_R FILLER_0_102_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_139 ();
 DECAPx4_ASAP7_75t_R FILLER_0_102_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_156 ();
 FILLER_ASAP7_75t_R FILLER_0_102_163 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_172 ();
 FILLER_ASAP7_75t_R FILLER_0_102_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_180 ();
 DECAPx1_ASAP7_75t_R FILLER_0_102_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_205 ();
 FILLER_ASAP7_75t_R FILLER_0_102_209 ();
 FILLER_ASAP7_75t_R FILLER_0_102_217 ();
 FILLER_ASAP7_75t_R FILLER_0_102_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_228 ();
 FILLER_ASAP7_75t_R FILLER_0_102_239 ();
 FILLER_ASAP7_75t_R FILLER_0_102_251 ();
 FILLER_ASAP7_75t_R FILLER_0_102_263 ();
 FILLER_ASAP7_75t_R FILLER_0_102_269 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_281 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_303 ();
 FILLER_ASAP7_75t_R FILLER_0_102_319 ();
 FILLER_ASAP7_75t_R FILLER_0_102_328 ();
 DECAPx1_ASAP7_75t_R FILLER_0_102_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_340 ();
 DECAPx4_ASAP7_75t_R FILLER_0_102_346 ();
 FILLER_ASAP7_75t_R FILLER_0_102_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_363 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_370 ();
 FILLER_ASAP7_75t_R FILLER_0_102_376 ();
 DECAPx1_ASAP7_75t_R FILLER_0_102_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_388 ();
 FILLER_ASAP7_75t_R FILLER_0_102_395 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_402 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_420 ();
 FILLER_ASAP7_75t_R FILLER_0_102_427 ();
 FILLER_ASAP7_75t_R FILLER_0_102_438 ();
 FILLER_ASAP7_75t_R FILLER_0_102_446 ();
 DECAPx1_ASAP7_75t_R FILLER_0_102_458 ();
 FILLER_ASAP7_75t_R FILLER_0_102_464 ();
 FILLER_ASAP7_75t_R FILLER_0_102_469 ();
 FILLER_ASAP7_75t_R FILLER_0_102_482 ();
 DECAPx1_ASAP7_75t_R FILLER_0_102_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_494 ();
 DECAPx6_ASAP7_75t_R FILLER_0_102_501 ();
 FILLER_ASAP7_75t_R FILLER_0_102_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_517 ();
 DECAPx1_ASAP7_75t_R FILLER_0_102_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_528 ();
 FILLER_ASAP7_75t_R FILLER_0_102_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_537 ();
 FILLER_ASAP7_75t_R FILLER_0_102_544 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_552 ();
 FILLER_ASAP7_75t_R FILLER_0_102_558 ();
 FILLER_ASAP7_75t_R FILLER_0_102_571 ();
 DECAPx1_ASAP7_75t_R FILLER_0_102_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_583 ();
 FILLER_ASAP7_75t_R FILLER_0_102_594 ();
 FILLER_ASAP7_75t_R FILLER_0_102_602 ();
 FILLER_ASAP7_75t_R FILLER_0_102_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_616 ();
 FILLER_ASAP7_75t_R FILLER_0_102_627 ();
 FILLER_ASAP7_75t_R FILLER_0_102_635 ();
 FILLER_ASAP7_75t_R FILLER_0_102_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_645 ();
 FILLER_ASAP7_75t_R FILLER_0_102_651 ();
 FILLER_ASAP7_75t_R FILLER_0_102_658 ();
 FILLER_ASAP7_75t_R FILLER_0_102_670 ();
 FILLER_ASAP7_75t_R FILLER_0_102_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_692 ();
 FILLER_ASAP7_75t_R FILLER_0_102_699 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_711 ();
 FILLER_ASAP7_75t_R FILLER_0_102_725 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_741 ();
 FILLER_ASAP7_75t_R FILLER_0_102_750 ();
 DECAPx1_ASAP7_75t_R FILLER_0_102_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_762 ();
 DECAPx1_ASAP7_75t_R FILLER_0_102_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_777 ();
 DECAPx4_ASAP7_75t_R FILLER_0_102_788 ();
 FILLER_ASAP7_75t_R FILLER_0_102_798 ();
 FILLER_ASAP7_75t_R FILLER_0_102_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_812 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_818 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_830 ();
 FILLER_ASAP7_75t_R FILLER_0_102_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_838 ();
 DECAPx4_ASAP7_75t_R FILLER_0_102_845 ();
 FILLER_ASAP7_75t_R FILLER_0_102_861 ();
 DECAPx4_ASAP7_75t_R FILLER_0_102_869 ();
 FILLER_ASAP7_75t_R FILLER_0_102_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_881 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_888 ();
 FILLER_ASAP7_75t_R FILLER_0_102_901 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_909 ();
 DECAPx6_ASAP7_75t_R FILLER_0_102_931 ();
 FILLER_ASAP7_75t_R FILLER_0_102_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_947 ();
 FILLER_ASAP7_75t_R FILLER_0_102_954 ();
 DECAPx6_ASAP7_75t_R FILLER_0_102_962 ();
 FILLER_ASAP7_75t_R FILLER_0_102_986 ();
 DECAPx1_ASAP7_75t_R FILLER_0_102_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_1008 ();
 FILLER_ASAP7_75t_R FILLER_0_102_1015 ();
 FILLER_ASAP7_75t_R FILLER_0_102_1023 ();
 FILLER_ASAP7_75t_R FILLER_0_102_1031 ();
 FILLER_ASAP7_75t_R FILLER_0_102_1039 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_1053 ();
 DECAPx6_ASAP7_75t_R FILLER_0_102_1061 ();
 DECAPx1_ASAP7_75t_R FILLER_0_102_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_1079 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_1086 ();
 DECAPx6_ASAP7_75t_R FILLER_0_102_1108 ();
 FILLER_ASAP7_75t_R FILLER_0_102_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_1129 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_1151 ();
 FILLER_ASAP7_75t_R FILLER_0_102_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_1159 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_1169 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_1176 ();
 FILLER_ASAP7_75t_R FILLER_0_102_1182 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_1196 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_1223 ();
 DECAPx1_ASAP7_75t_R FILLER_0_102_1230 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_1234 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_1255 ();
 FILLER_ASAP7_75t_R FILLER_0_102_1261 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_1273 ();
 FILLER_ASAP7_75t_R FILLER_0_102_1279 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_1297 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_1303 ();
 FILLER_ASAP7_75t_R FILLER_0_102_1314 ();
 FILLER_ASAP7_75t_R FILLER_0_102_1324 ();
 FILLER_ASAP7_75t_R FILLER_0_102_1332 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_1334 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_1341 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_1347 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_1351 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_102_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_103_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_4 ();
 FILLER_ASAP7_75t_R FILLER_0_103_11 ();
 FILLER_ASAP7_75t_R FILLER_0_103_18 ();
 FILLER_ASAP7_75t_R FILLER_0_103_25 ();
 DECAPx2_ASAP7_75t_R FILLER_0_103_33 ();
 DECAPx1_ASAP7_75t_R FILLER_0_103_50 ();
 FILLER_ASAP7_75t_R FILLER_0_103_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_68 ();
 DECAPx4_ASAP7_75t_R FILLER_0_103_75 ();
 FILLER_ASAP7_75t_R FILLER_0_103_88 ();
 DECAPx1_ASAP7_75t_R FILLER_0_103_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_102 ();
 DECAPx1_ASAP7_75t_R FILLER_0_103_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_117 ();
 DECAPx6_ASAP7_75t_R FILLER_0_103_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_144 ();
 FILLER_ASAP7_75t_R FILLER_0_103_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_153 ();
 FILLER_ASAP7_75t_R FILLER_0_103_160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_172 ();
 DECAPx2_ASAP7_75t_R FILLER_0_103_194 ();
 FILLER_ASAP7_75t_R FILLER_0_103_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_202 ();
 FILLER_ASAP7_75t_R FILLER_0_103_223 ();
 FILLER_ASAP7_75t_R FILLER_0_103_235 ();
 FILLER_ASAP7_75t_R FILLER_0_103_247 ();
 DECAPx1_ASAP7_75t_R FILLER_0_103_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_259 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_270 ();
 DECAPx4_ASAP7_75t_R FILLER_0_103_292 ();
 FILLER_ASAP7_75t_R FILLER_0_103_302 ();
 DECAPx4_ASAP7_75t_R FILLER_0_103_307 ();
 FILLER_ASAP7_75t_R FILLER_0_103_317 ();
 FILLER_ASAP7_75t_R FILLER_0_103_327 ();
 FILLER_ASAP7_75t_R FILLER_0_103_332 ();
 DECAPx4_ASAP7_75t_R FILLER_0_103_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_350 ();
 FILLER_ASAP7_75t_R FILLER_0_103_361 ();
 FILLER_ASAP7_75t_R FILLER_0_103_369 ();
 FILLER_ASAP7_75t_R FILLER_0_103_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_379 ();
 DECAPx2_ASAP7_75t_R FILLER_0_103_390 ();
 DECAPx6_ASAP7_75t_R FILLER_0_103_402 ();
 DECAPx1_ASAP7_75t_R FILLER_0_103_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_420 ();
 FILLER_ASAP7_75t_R FILLER_0_103_427 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_435 ();
 DECAPx2_ASAP7_75t_R FILLER_0_103_457 ();
 FILLER_ASAP7_75t_R FILLER_0_103_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_465 ();
 FILLER_ASAP7_75t_R FILLER_0_103_476 ();
 FILLER_ASAP7_75t_R FILLER_0_103_484 ();
 FILLER_ASAP7_75t_R FILLER_0_103_492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_103_500 ();
 FILLER_ASAP7_75t_R FILLER_0_103_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_526 ();
 DECAPx1_ASAP7_75t_R FILLER_0_103_537 ();
 FILLER_ASAP7_75t_R FILLER_0_103_551 ();
 DECAPx2_ASAP7_75t_R FILLER_0_103_559 ();
 FILLER_ASAP7_75t_R FILLER_0_103_565 ();
 DECAPx1_ASAP7_75t_R FILLER_0_103_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_577 ();
 FILLER_ASAP7_75t_R FILLER_0_103_584 ();
 FILLER_ASAP7_75t_R FILLER_0_103_592 ();
 FILLER_ASAP7_75t_R FILLER_0_103_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_608 ();
 FILLER_ASAP7_75t_R FILLER_0_103_615 ();
 FILLER_ASAP7_75t_R FILLER_0_103_632 ();
 DECAPx1_ASAP7_75t_R FILLER_0_103_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_644 ();
 FILLER_ASAP7_75t_R FILLER_0_103_650 ();
 FILLER_ASAP7_75t_R FILLER_0_103_657 ();
 FILLER_ASAP7_75t_R FILLER_0_103_665 ();
 FILLER_ASAP7_75t_R FILLER_0_103_677 ();
 FILLER_ASAP7_75t_R FILLER_0_103_689 ();
 FILLER_ASAP7_75t_R FILLER_0_103_701 ();
 FILLER_ASAP7_75t_R FILLER_0_103_713 ();
 FILLER_ASAP7_75t_R FILLER_0_103_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_727 ();
 FILLER_ASAP7_75t_R FILLER_0_103_734 ();
 FILLER_ASAP7_75t_R FILLER_0_103_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_741 ();
 FILLER_ASAP7_75t_R FILLER_0_103_748 ();
 FILLER_ASAP7_75t_R FILLER_0_103_755 ();
 FILLER_ASAP7_75t_R FILLER_0_103_777 ();
 FILLER_ASAP7_75t_R FILLER_0_103_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_786 ();
 DECAPx1_ASAP7_75t_R FILLER_0_103_793 ();
 DECAPx2_ASAP7_75t_R FILLER_0_103_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_810 ();
 DECAPx4_ASAP7_75t_R FILLER_0_103_817 ();
 DECAPx2_ASAP7_75t_R FILLER_0_103_833 ();
 DECAPx4_ASAP7_75t_R FILLER_0_103_847 ();
 FILLER_ASAP7_75t_R FILLER_0_103_867 ();
 FILLER_ASAP7_75t_R FILLER_0_103_875 ();
 DECAPx2_ASAP7_75t_R FILLER_0_103_884 ();
 FILLER_ASAP7_75t_R FILLER_0_103_890 ();
 DECAPx4_ASAP7_75t_R FILLER_0_103_895 ();
 DECAPx4_ASAP7_75t_R FILLER_0_103_913 ();
 FILLER_ASAP7_75t_R FILLER_0_103_923 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_927 ();
 FILLER_ASAP7_75t_R FILLER_0_103_955 ();
 FILLER_ASAP7_75t_R FILLER_0_103_965 ();
 FILLER_ASAP7_75t_R FILLER_0_103_973 ();
 FILLER_ASAP7_75t_R FILLER_0_103_981 ();
 DECAPx2_ASAP7_75t_R FILLER_0_103_989 ();
 FILLER_ASAP7_75t_R FILLER_0_103_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_997 ();
 FILLER_ASAP7_75t_R FILLER_0_103_1004 ();
 FILLER_ASAP7_75t_R FILLER_0_103_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_1014 ();
 FILLER_ASAP7_75t_R FILLER_0_103_1025 ();
 DECAPx1_ASAP7_75t_R FILLER_0_103_1033 ();
 DECAPx2_ASAP7_75t_R FILLER_0_103_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_1053 ();
 DECAPx4_ASAP7_75t_R FILLER_0_103_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_1090 ();
 DECAPx2_ASAP7_75t_R FILLER_0_103_1112 ();
 DECAPx6_ASAP7_75t_R FILLER_0_103_1124 ();
 FILLER_ASAP7_75t_R FILLER_0_103_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_1146 ();
 DECAPx1_ASAP7_75t_R FILLER_0_103_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_1172 ();
 FILLER_ASAP7_75t_R FILLER_0_103_1179 ();
 DECAPx1_ASAP7_75t_R FILLER_0_103_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_1193 ();
 DECAPx1_ASAP7_75t_R FILLER_0_103_1199 ();
 DECAPx4_ASAP7_75t_R FILLER_0_103_1213 ();
 FILLER_ASAP7_75t_R FILLER_0_103_1223 ();
 FILLER_ASAP7_75t_R FILLER_0_103_1231 ();
 DECAPx6_ASAP7_75t_R FILLER_0_103_1239 ();
 FILLER_ASAP7_75t_R FILLER_0_103_1253 ();
 FILLER_ASAP7_75t_R FILLER_0_103_1262 ();
 DECAPx4_ASAP7_75t_R FILLER_0_103_1274 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_1284 ();
 DECAPx1_ASAP7_75t_R FILLER_0_103_1293 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_1297 ();
 DECAPx1_ASAP7_75t_R FILLER_0_103_1304 ();
 FILLER_ASAP7_75t_R FILLER_0_103_1314 ();
 DECAPx4_ASAP7_75t_R FILLER_0_103_1322 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_1332 ();
 DECAPx6_ASAP7_75t_R FILLER_0_103_1339 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_1353 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_1359 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_104_2 ();
 FILLER_ASAP7_75t_R FILLER_0_104_9 ();
 DECAPx2_ASAP7_75t_R FILLER_0_104_17 ();
 FILLER_ASAP7_75t_R FILLER_0_104_23 ();
 FILLER_ASAP7_75t_R FILLER_0_104_53 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_61 ();
 DECAPx6_ASAP7_75t_R FILLER_0_104_83 ();
 FILLER_ASAP7_75t_R FILLER_0_104_97 ();
 FILLER_ASAP7_75t_R FILLER_0_104_109 ();
 FILLER_ASAP7_75t_R FILLER_0_104_121 ();
 DECAPx4_ASAP7_75t_R FILLER_0_104_133 ();
 FILLER_ASAP7_75t_R FILLER_0_104_143 ();
 DECAPx6_ASAP7_75t_R FILLER_0_104_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_179 ();
 FILLER_ASAP7_75t_R FILLER_0_104_200 ();
 FILLER_ASAP7_75t_R FILLER_0_104_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_210 ();
 FILLER_ASAP7_75t_R FILLER_0_104_218 ();
 FILLER_ASAP7_75t_R FILLER_0_104_230 ();
 FILLER_ASAP7_75t_R FILLER_0_104_242 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_254 ();
 DECAPx1_ASAP7_75t_R FILLER_0_104_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_280 ();
 FILLER_ASAP7_75t_R FILLER_0_104_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_304 ();
 DECAPx1_ASAP7_75t_R FILLER_0_104_311 ();
 FILLER_ASAP7_75t_R FILLER_0_104_320 ();
 DECAPx1_ASAP7_75t_R FILLER_0_104_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_336 ();
 FILLER_ASAP7_75t_R FILLER_0_104_340 ();
 FILLER_ASAP7_75t_R FILLER_0_104_352 ();
 FILLER_ASAP7_75t_R FILLER_0_104_360 ();
 FILLER_ASAP7_75t_R FILLER_0_104_369 ();
 DECAPx1_ASAP7_75t_R FILLER_0_104_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_381 ();
 FILLER_ASAP7_75t_R FILLER_0_104_389 ();
 FILLER_ASAP7_75t_R FILLER_0_104_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_402 ();
 DECAPx4_ASAP7_75t_R FILLER_0_104_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_420 ();
 FILLER_ASAP7_75t_R FILLER_0_104_431 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_461 ();
 FILLER_ASAP7_75t_R FILLER_0_104_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_472 ();
 FILLER_ASAP7_75t_R FILLER_0_104_494 ();
 DECAPx2_ASAP7_75t_R FILLER_0_104_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_508 ();
 FILLER_ASAP7_75t_R FILLER_0_104_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_517 ();
 FILLER_ASAP7_75t_R FILLER_0_104_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_530 ();
 FILLER_ASAP7_75t_R FILLER_0_104_537 ();
 FILLER_ASAP7_75t_R FILLER_0_104_549 ();
 DECAPx1_ASAP7_75t_R FILLER_0_104_561 ();
 FILLER_ASAP7_75t_R FILLER_0_104_571 ();
 DECAPx1_ASAP7_75t_R FILLER_0_104_578 ();
 FILLER_ASAP7_75t_R FILLER_0_104_588 ();
 FILLER_ASAP7_75t_R FILLER_0_104_596 ();
 FILLER_ASAP7_75t_R FILLER_0_104_608 ();
 FILLER_ASAP7_75t_R FILLER_0_104_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_622 ();
 FILLER_ASAP7_75t_R FILLER_0_104_633 ();
 FILLER_ASAP7_75t_R FILLER_0_104_645 ();
 FILLER_ASAP7_75t_R FILLER_0_104_657 ();
 FILLER_ASAP7_75t_R FILLER_0_104_664 ();
 FILLER_ASAP7_75t_R FILLER_0_104_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_678 ();
 FILLER_ASAP7_75t_R FILLER_0_104_689 ();
 FILLER_ASAP7_75t_R FILLER_0_104_696 ();
 FILLER_ASAP7_75t_R FILLER_0_104_708 ();
 DECAPx1_ASAP7_75t_R FILLER_0_104_720 ();
 FILLER_ASAP7_75t_R FILLER_0_104_732 ();
 DECAPx2_ASAP7_75t_R FILLER_0_104_743 ();
 FILLER_ASAP7_75t_R FILLER_0_104_749 ();
 FILLER_ASAP7_75t_R FILLER_0_104_767 ();
 DECAPx4_ASAP7_75t_R FILLER_0_104_775 ();
 FILLER_ASAP7_75t_R FILLER_0_104_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_787 ();
 DECAPx6_ASAP7_75t_R FILLER_0_104_796 ();
 FILLER_ASAP7_75t_R FILLER_0_104_810 ();
 FILLER_ASAP7_75t_R FILLER_0_104_818 ();
 DECAPx2_ASAP7_75t_R FILLER_0_104_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_836 ();
 DECAPx6_ASAP7_75t_R FILLER_0_104_848 ();
 FILLER_ASAP7_75t_R FILLER_0_104_868 ();
 DECAPx4_ASAP7_75t_R FILLER_0_104_876 ();
 DECAPx2_ASAP7_75t_R FILLER_0_104_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_900 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_911 ();
 DECAPx4_ASAP7_75t_R FILLER_0_104_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_943 ();
 FILLER_ASAP7_75t_R FILLER_0_104_947 ();
 DECAPx6_ASAP7_75t_R FILLER_0_104_955 ();
 FILLER_ASAP7_75t_R FILLER_0_104_969 ();
 FILLER_ASAP7_75t_R FILLER_0_104_977 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_1004 ();
 DECAPx2_ASAP7_75t_R FILLER_0_104_1011 ();
 FILLER_ASAP7_75t_R FILLER_0_104_1027 ();
 DECAPx1_ASAP7_75t_R FILLER_0_104_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_1039 ();
 FILLER_ASAP7_75t_R FILLER_0_104_1046 ();
 DECAPx1_ASAP7_75t_R FILLER_0_104_1054 ();
 DECAPx6_ASAP7_75t_R FILLER_0_104_1064 ();
 FILLER_ASAP7_75t_R FILLER_0_104_1084 ();
 FILLER_ASAP7_75t_R FILLER_0_104_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_1094 ();
 DECAPx4_ASAP7_75t_R FILLER_0_104_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_1111 ();
 FILLER_ASAP7_75t_R FILLER_0_104_1118 ();
 FILLER_ASAP7_75t_R FILLER_0_104_1126 ();
 DECAPx2_ASAP7_75t_R FILLER_0_104_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_1140 ();
 DECAPx2_ASAP7_75t_R FILLER_0_104_1151 ();
 FILLER_ASAP7_75t_R FILLER_0_104_1168 ();
 DECAPx2_ASAP7_75t_R FILLER_0_104_1176 ();
 FILLER_ASAP7_75t_R FILLER_0_104_1182 ();
 DECAPx1_ASAP7_75t_R FILLER_0_104_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_1194 ();
 FILLER_ASAP7_75t_R FILLER_0_104_1202 ();
 FILLER_ASAP7_75t_R FILLER_0_104_1212 ();
 DECAPx4_ASAP7_75t_R FILLER_0_104_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_1229 ();
 FILLER_ASAP7_75t_R FILLER_0_104_1237 ();
 DECAPx4_ASAP7_75t_R FILLER_0_104_1245 ();
 DECAPx1_ASAP7_75t_R FILLER_0_104_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_0_104_1272 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_1278 ();
 FILLER_ASAP7_75t_R FILLER_0_104_1299 ();
 FILLER_ASAP7_75t_R FILLER_0_104_1307 ();
 DECAPx6_ASAP7_75t_R FILLER_0_104_1315 ();
 FILLER_ASAP7_75t_R FILLER_0_104_1335 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_104_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_105_2 ();
 FILLER_ASAP7_75t_R FILLER_0_105_25 ();
 FILLER_ASAP7_75t_R FILLER_0_105_32 ();
 DECAPx1_ASAP7_75t_R FILLER_0_105_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_43 ();
 FILLER_ASAP7_75t_R FILLER_0_105_50 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_58 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_80 ();
 FILLER_ASAP7_75t_R FILLER_0_105_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_104 ();
 FILLER_ASAP7_75t_R FILLER_0_105_115 ();
 FILLER_ASAP7_75t_R FILLER_0_105_123 ();
 DECAPx4_ASAP7_75t_R FILLER_0_105_131 ();
 FILLER_ASAP7_75t_R FILLER_0_105_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_143 ();
 FILLER_ASAP7_75t_R FILLER_0_105_152 ();
 DECAPx2_ASAP7_75t_R FILLER_0_105_164 ();
 FILLER_ASAP7_75t_R FILLER_0_105_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_172 ();
 DECAPx2_ASAP7_75t_R FILLER_0_105_179 ();
 DECAPx4_ASAP7_75t_R FILLER_0_105_195 ();
 FILLER_ASAP7_75t_R FILLER_0_105_205 ();
 DECAPx1_ASAP7_75t_R FILLER_0_105_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_221 ();
 DECAPx4_ASAP7_75t_R FILLER_0_105_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_242 ();
 FILLER_ASAP7_75t_R FILLER_0_105_253 ();
 DECAPx2_ASAP7_75t_R FILLER_0_105_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_267 ();
 FILLER_ASAP7_75t_R FILLER_0_105_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_281 ();
 DECAPx2_ASAP7_75t_R FILLER_0_105_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_294 ();
 DECAPx2_ASAP7_75t_R FILLER_0_105_302 ();
 FILLER_ASAP7_75t_R FILLER_0_105_314 ();
 FILLER_ASAP7_75t_R FILLER_0_105_326 ();
 FILLER_ASAP7_75t_R FILLER_0_105_336 ();
 DECAPx1_ASAP7_75t_R FILLER_0_105_344 ();
 FILLER_ASAP7_75t_R FILLER_0_105_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_358 ();
 FILLER_ASAP7_75t_R FILLER_0_105_362 ();
 FILLER_ASAP7_75t_R FILLER_0_105_370 ();
 FILLER_ASAP7_75t_R FILLER_0_105_378 ();
 FILLER_ASAP7_75t_R FILLER_0_105_386 ();
 FILLER_ASAP7_75t_R FILLER_0_105_394 ();
 DECAPx4_ASAP7_75t_R FILLER_0_105_403 ();
 FILLER_ASAP7_75t_R FILLER_0_105_413 ();
 FILLER_ASAP7_75t_R FILLER_0_105_418 ();
 FILLER_ASAP7_75t_R FILLER_0_105_426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_431 ();
 FILLER_ASAP7_75t_R FILLER_0_105_459 ();
 DECAPx2_ASAP7_75t_R FILLER_0_105_467 ();
 FILLER_ASAP7_75t_R FILLER_0_105_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_475 ();
 DECAPx6_ASAP7_75t_R FILLER_0_105_482 ();
 FILLER_ASAP7_75t_R FILLER_0_105_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_498 ();
 DECAPx1_ASAP7_75t_R FILLER_0_105_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_519 ();
 FILLER_ASAP7_75t_R FILLER_0_105_525 ();
 FILLER_ASAP7_75t_R FILLER_0_105_534 ();
 FILLER_ASAP7_75t_R FILLER_0_105_546 ();
 FILLER_ASAP7_75t_R FILLER_0_105_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_555 ();
 DECAPx1_ASAP7_75t_R FILLER_0_105_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_570 ();
 FILLER_ASAP7_75t_R FILLER_0_105_577 ();
 FILLER_ASAP7_75t_R FILLER_0_105_585 ();
 FILLER_ASAP7_75t_R FILLER_0_105_597 ();
 FILLER_ASAP7_75t_R FILLER_0_105_609 ();
 FILLER_ASAP7_75t_R FILLER_0_105_621 ();
 FILLER_ASAP7_75t_R FILLER_0_105_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_635 ();
 FILLER_ASAP7_75t_R FILLER_0_105_643 ();
 FILLER_ASAP7_75t_R FILLER_0_105_651 ();
 FILLER_ASAP7_75t_R FILLER_0_105_663 ();
 FILLER_ASAP7_75t_R FILLER_0_105_669 ();
 FILLER_ASAP7_75t_R FILLER_0_105_677 ();
 DECAPx1_ASAP7_75t_R FILLER_0_105_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_693 ();
 FILLER_ASAP7_75t_R FILLER_0_105_704 ();
 FILLER_ASAP7_75t_R FILLER_0_105_711 ();
 FILLER_ASAP7_75t_R FILLER_0_105_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_725 ();
 FILLER_ASAP7_75t_R FILLER_0_105_729 ();
 DECAPx2_ASAP7_75t_R FILLER_0_105_749 ();
 FILLER_ASAP7_75t_R FILLER_0_105_755 ();
 FILLER_ASAP7_75t_R FILLER_0_105_767 ();
 DECAPx1_ASAP7_75t_R FILLER_0_105_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_783 ();
 DECAPx2_ASAP7_75t_R FILLER_0_105_794 ();
 FILLER_ASAP7_75t_R FILLER_0_105_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_802 ();
 DECAPx4_ASAP7_75t_R FILLER_0_105_825 ();
 FILLER_ASAP7_75t_R FILLER_0_105_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_843 ();
 DECAPx2_ASAP7_75t_R FILLER_0_105_850 ();
 FILLER_ASAP7_75t_R FILLER_0_105_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_858 ();
 DECAPx4_ASAP7_75t_R FILLER_0_105_871 ();
 FILLER_ASAP7_75t_R FILLER_0_105_881 ();
 FILLER_ASAP7_75t_R FILLER_0_105_888 ();
 DECAPx4_ASAP7_75t_R FILLER_0_105_902 ();
 DECAPx1_ASAP7_75t_R FILLER_0_105_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_924 ();
 DECAPx6_ASAP7_75t_R FILLER_0_105_927 ();
 DECAPx1_ASAP7_75t_R FILLER_0_105_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_945 ();
 FILLER_ASAP7_75t_R FILLER_0_105_967 ();
 FILLER_ASAP7_75t_R FILLER_0_105_974 ();
 FILLER_ASAP7_75t_R FILLER_0_105_982 ();
 DECAPx4_ASAP7_75t_R FILLER_0_105_990 ();
 FILLER_ASAP7_75t_R FILLER_0_105_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_1002 ();
 DECAPx6_ASAP7_75t_R FILLER_0_105_1009 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_1029 ();
 DECAPx6_ASAP7_75t_R FILLER_0_105_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_1071 ();
 DECAPx2_ASAP7_75t_R FILLER_0_105_1077 ();
 FILLER_ASAP7_75t_R FILLER_0_105_1088 ();
 FILLER_ASAP7_75t_R FILLER_0_105_1096 ();
 DECAPx2_ASAP7_75t_R FILLER_0_105_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_1110 ();
 FILLER_ASAP7_75t_R FILLER_0_105_1117 ();
 FILLER_ASAP7_75t_R FILLER_0_105_1130 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_1138 ();
 FILLER_ASAP7_75t_R FILLER_0_105_1160 ();
 DECAPx4_ASAP7_75t_R FILLER_0_105_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_1178 ();
 FILLER_ASAP7_75t_R FILLER_0_105_1185 ();
 DECAPx4_ASAP7_75t_R FILLER_0_105_1209 ();
 FILLER_ASAP7_75t_R FILLER_0_105_1219 ();
 FILLER_ASAP7_75t_R FILLER_0_105_1227 ();
 FILLER_ASAP7_75t_R FILLER_0_105_1235 ();
 DECAPx2_ASAP7_75t_R FILLER_0_105_1243 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_1249 ();
 DECAPx1_ASAP7_75t_R FILLER_0_105_1260 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_1264 ();
 DECAPx6_ASAP7_75t_R FILLER_0_105_1270 ();
 DECAPx1_ASAP7_75t_R FILLER_0_105_1287 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_1291 ();
 FILLER_ASAP7_75t_R FILLER_0_105_1298 ();
 FILLER_ASAP7_75t_R FILLER_0_105_1306 ();
 FILLER_ASAP7_75t_R FILLER_0_105_1314 ();
 FILLER_ASAP7_75t_R FILLER_0_105_1322 ();
 DECAPx1_ASAP7_75t_R FILLER_0_105_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_1341 ();
 DECAPx6_ASAP7_75t_R FILLER_0_105_1363 ();
 FILLER_ASAP7_75t_R FILLER_0_105_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_106_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_106_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_13 ();
 FILLER_ASAP7_75t_R FILLER_0_106_19 ();
 FILLER_ASAP7_75t_R FILLER_0_106_29 ();
 FILLER_ASAP7_75t_R FILLER_0_106_47 ();
 FILLER_ASAP7_75t_R FILLER_0_106_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_54 ();
 FILLER_ASAP7_75t_R FILLER_0_106_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_63 ();
 FILLER_ASAP7_75t_R FILLER_0_106_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_72 ();
 FILLER_ASAP7_75t_R FILLER_0_106_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_85 ();
 DECAPx1_ASAP7_75t_R FILLER_0_106_92 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_104 ();
 DECAPx6_ASAP7_75t_R FILLER_0_106_132 ();
 FILLER_ASAP7_75t_R FILLER_0_106_146 ();
 FILLER_ASAP7_75t_R FILLER_0_106_158 ();
 FILLER_ASAP7_75t_R FILLER_0_106_164 ();
 DECAPx6_ASAP7_75t_R FILLER_0_106_178 ();
 DECAPx1_ASAP7_75t_R FILLER_0_106_192 ();
 FILLER_ASAP7_75t_R FILLER_0_106_202 ();
 FILLER_ASAP7_75t_R FILLER_0_106_210 ();
 FILLER_ASAP7_75t_R FILLER_0_106_220 ();
 DECAPx1_ASAP7_75t_R FILLER_0_106_227 ();
 FILLER_ASAP7_75t_R FILLER_0_106_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_237 ();
 FILLER_ASAP7_75t_R FILLER_0_106_244 ();
 FILLER_ASAP7_75t_R FILLER_0_106_252 ();
 DECAPx6_ASAP7_75t_R FILLER_0_106_260 ();
 FILLER_ASAP7_75t_R FILLER_0_106_277 ();
 FILLER_ASAP7_75t_R FILLER_0_106_282 ();
 DECAPx2_ASAP7_75t_R FILLER_0_106_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_298 ();
 FILLER_ASAP7_75t_R FILLER_0_106_309 ();
 DECAPx1_ASAP7_75t_R FILLER_0_106_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_325 ();
 DECAPx2_ASAP7_75t_R FILLER_0_106_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_352 ();
 FILLER_ASAP7_75t_R FILLER_0_106_363 ();
 FILLER_ASAP7_75t_R FILLER_0_106_370 ();
 FILLER_ASAP7_75t_R FILLER_0_106_379 ();
 DECAPx2_ASAP7_75t_R FILLER_0_106_391 ();
 FILLER_ASAP7_75t_R FILLER_0_106_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_399 ();
 FILLER_ASAP7_75t_R FILLER_0_106_410 ();
 DECAPx4_ASAP7_75t_R FILLER_0_106_418 ();
 FILLER_ASAP7_75t_R FILLER_0_106_428 ();
 DECAPx6_ASAP7_75t_R FILLER_0_106_438 ();
 FILLER_ASAP7_75t_R FILLER_0_106_452 ();
 FILLER_ASAP7_75t_R FILLER_0_106_460 ();
 FILLER_ASAP7_75t_R FILLER_0_106_464 ();
 DECAPx1_ASAP7_75t_R FILLER_0_106_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_477 ();
 FILLER_ASAP7_75t_R FILLER_0_106_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_486 ();
 FILLER_ASAP7_75t_R FILLER_0_106_493 ();
 FILLER_ASAP7_75t_R FILLER_0_106_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_503 ();
 FILLER_ASAP7_75t_R FILLER_0_106_510 ();
 FILLER_ASAP7_75t_R FILLER_0_106_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_520 ();
 FILLER_ASAP7_75t_R FILLER_0_106_529 ();
 FILLER_ASAP7_75t_R FILLER_0_106_539 ();
 FILLER_ASAP7_75t_R FILLER_0_106_551 ();
 FILLER_ASAP7_75t_R FILLER_0_106_563 ();
 FILLER_ASAP7_75t_R FILLER_0_106_570 ();
 FILLER_ASAP7_75t_R FILLER_0_106_582 ();
 FILLER_ASAP7_75t_R FILLER_0_106_589 ();
 FILLER_ASAP7_75t_R FILLER_0_106_601 ();
 DECAPx1_ASAP7_75t_R FILLER_0_106_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_617 ();
 DECAPx2_ASAP7_75t_R FILLER_0_106_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_634 ();
 DECAPx2_ASAP7_75t_R FILLER_0_106_659 ();
 FILLER_ASAP7_75t_R FILLER_0_106_671 ();
 FILLER_ASAP7_75t_R FILLER_0_106_683 ();
 FILLER_ASAP7_75t_R FILLER_0_106_695 ();
 FILLER_ASAP7_75t_R FILLER_0_106_707 ();
 FILLER_ASAP7_75t_R FILLER_0_106_717 ();
 FILLER_ASAP7_75t_R FILLER_0_106_729 ();
 FILLER_ASAP7_75t_R FILLER_0_106_743 ();
 FILLER_ASAP7_75t_R FILLER_0_106_767 ();
 FILLER_ASAP7_75t_R FILLER_0_106_775 ();
 DECAPx4_ASAP7_75t_R FILLER_0_106_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_807 ();
 DECAPx2_ASAP7_75t_R FILLER_0_106_815 ();
 FILLER_ASAP7_75t_R FILLER_0_106_843 ();
 DECAPx2_ASAP7_75t_R FILLER_0_106_852 ();
 FILLER_ASAP7_75t_R FILLER_0_106_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_860 ();
 DECAPx4_ASAP7_75t_R FILLER_0_106_871 ();
 FILLER_ASAP7_75t_R FILLER_0_106_888 ();
 DECAPx1_ASAP7_75t_R FILLER_0_106_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_904 ();
 FILLER_ASAP7_75t_R FILLER_0_106_929 ();
 FILLER_ASAP7_75t_R FILLER_0_106_937 ();
 DECAPx6_ASAP7_75t_R FILLER_0_106_943 ();
 DECAPx2_ASAP7_75t_R FILLER_0_106_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_963 ();
 FILLER_ASAP7_75t_R FILLER_0_106_967 ();
 FILLER_ASAP7_75t_R FILLER_0_106_975 ();
 FILLER_ASAP7_75t_R FILLER_0_106_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_985 ();
 DECAPx1_ASAP7_75t_R FILLER_0_106_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_996 ();
 DECAPx2_ASAP7_75t_R FILLER_0_106_1017 ();
 FILLER_ASAP7_75t_R FILLER_0_106_1023 ();
 DECAPx6_ASAP7_75t_R FILLER_0_106_1033 ();
 DECAPx2_ASAP7_75t_R FILLER_0_106_1047 ();
 FILLER_ASAP7_75t_R FILLER_0_106_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_1061 ();
 FILLER_ASAP7_75t_R FILLER_0_106_1072 ();
 DECAPx2_ASAP7_75t_R FILLER_0_106_1080 ();
 DECAPx1_ASAP7_75t_R FILLER_0_106_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_1096 ();
 DECAPx2_ASAP7_75t_R FILLER_0_106_1103 ();
 DECAPx1_ASAP7_75t_R FILLER_0_106_1115 ();
 FILLER_ASAP7_75t_R FILLER_0_106_1125 ();
 FILLER_ASAP7_75t_R FILLER_0_106_1133 ();
 DECAPx6_ASAP7_75t_R FILLER_0_106_1140 ();
 DECAPx1_ASAP7_75t_R FILLER_0_106_1154 ();
 FILLER_ASAP7_75t_R FILLER_0_106_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_1166 ();
 FILLER_ASAP7_75t_R FILLER_0_106_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_1177 ();
 DECAPx1_ASAP7_75t_R FILLER_0_106_1185 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_1189 ();
 DECAPx2_ASAP7_75t_R FILLER_0_106_1196 ();
 FILLER_ASAP7_75t_R FILLER_0_106_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_1204 ();
 FILLER_ASAP7_75t_R FILLER_0_106_1211 ();
 DECAPx2_ASAP7_75t_R FILLER_0_106_1219 ();
 FILLER_ASAP7_75t_R FILLER_0_106_1235 ();
 DECAPx2_ASAP7_75t_R FILLER_0_106_1248 ();
 FILLER_ASAP7_75t_R FILLER_0_106_1257 ();
 FILLER_ASAP7_75t_R FILLER_0_106_1265 ();
 FILLER_ASAP7_75t_R FILLER_0_106_1273 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_1281 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_1303 ();
 DECAPx2_ASAP7_75t_R FILLER_0_106_1310 ();
 DECAPx2_ASAP7_75t_R FILLER_0_106_1322 ();
 FILLER_ASAP7_75t_R FILLER_0_106_1334 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_1336 ();
 FILLER_ASAP7_75t_R FILLER_0_106_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_106_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_107_2 ();
 FILLER_ASAP7_75t_R FILLER_0_107_9 ();
 FILLER_ASAP7_75t_R FILLER_0_107_16 ();
 FILLER_ASAP7_75t_R FILLER_0_107_21 ();
 FILLER_ASAP7_75t_R FILLER_0_107_29 ();
 FILLER_ASAP7_75t_R FILLER_0_107_36 ();
 FILLER_ASAP7_75t_R FILLER_0_107_44 ();
 DECAPx1_ASAP7_75t_R FILLER_0_107_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_55 ();
 DECAPx2_ASAP7_75t_R FILLER_0_107_62 ();
 FILLER_ASAP7_75t_R FILLER_0_107_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_70 ();
 DECAPx2_ASAP7_75t_R FILLER_0_107_82 ();
 DECAPx2_ASAP7_75t_R FILLER_0_107_94 ();
 DECAPx1_ASAP7_75t_R FILLER_0_107_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_112 ();
 DECAPx2_ASAP7_75t_R FILLER_0_107_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_129 ();
 FILLER_ASAP7_75t_R FILLER_0_107_140 ();
 FILLER_ASAP7_75t_R FILLER_0_107_146 ();
 FILLER_ASAP7_75t_R FILLER_0_107_154 ();
 FILLER_ASAP7_75t_R FILLER_0_107_162 ();
 FILLER_ASAP7_75t_R FILLER_0_107_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_171 ();
 FILLER_ASAP7_75t_R FILLER_0_107_178 ();
 FILLER_ASAP7_75t_R FILLER_0_107_186 ();
 FILLER_ASAP7_75t_R FILLER_0_107_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_198 ();
 FILLER_ASAP7_75t_R FILLER_0_107_204 ();
 DECAPx1_ASAP7_75t_R FILLER_0_107_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_230 ();
 DECAPx4_ASAP7_75t_R FILLER_0_107_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_247 ();
 DECAPx6_ASAP7_75t_R FILLER_0_107_268 ();
 DECAPx2_ASAP7_75t_R FILLER_0_107_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_288 ();
 DECAPx2_ASAP7_75t_R FILLER_0_107_299 ();
 FILLER_ASAP7_75t_R FILLER_0_107_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_328 ();
 DECAPx6_ASAP7_75t_R FILLER_0_107_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_348 ();
 FILLER_ASAP7_75t_R FILLER_0_107_355 ();
 FILLER_ASAP7_75t_R FILLER_0_107_367 ();
 DECAPx1_ASAP7_75t_R FILLER_0_107_374 ();
 FILLER_ASAP7_75t_R FILLER_0_107_390 ();
 FILLER_ASAP7_75t_R FILLER_0_107_402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_414 ();
 DECAPx2_ASAP7_75t_R FILLER_0_107_436 ();
 DECAPx1_ASAP7_75t_R FILLER_0_107_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_452 ();
 FILLER_ASAP7_75t_R FILLER_0_107_473 ();
 FILLER_ASAP7_75t_R FILLER_0_107_483 ();
 FILLER_ASAP7_75t_R FILLER_0_107_488 ();
 FILLER_ASAP7_75t_R FILLER_0_107_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_498 ();
 DECAPx2_ASAP7_75t_R FILLER_0_107_505 ();
 FILLER_ASAP7_75t_R FILLER_0_107_517 ();
 FILLER_ASAP7_75t_R FILLER_0_107_525 ();
 FILLER_ASAP7_75t_R FILLER_0_107_537 ();
 DECAPx1_ASAP7_75t_R FILLER_0_107_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_553 ();
 DECAPx1_ASAP7_75t_R FILLER_0_107_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_568 ();
 FILLER_ASAP7_75t_R FILLER_0_107_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_581 ();
 DECAPx1_ASAP7_75t_R FILLER_0_107_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_596 ();
 FILLER_ASAP7_75t_R FILLER_0_107_607 ();
 FILLER_ASAP7_75t_R FILLER_0_107_615 ();
 DECAPx1_ASAP7_75t_R FILLER_0_107_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_631 ();
 DECAPx1_ASAP7_75t_R FILLER_0_107_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_658 ();
 FILLER_ASAP7_75t_R FILLER_0_107_669 ();
 DECAPx1_ASAP7_75t_R FILLER_0_107_681 ();
 FILLER_ASAP7_75t_R FILLER_0_107_695 ();
 FILLER_ASAP7_75t_R FILLER_0_107_707 ();
 FILLER_ASAP7_75t_R FILLER_0_107_715 ();
 DECAPx1_ASAP7_75t_R FILLER_0_107_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_731 ();
 FILLER_ASAP7_75t_R FILLER_0_107_743 ();
 FILLER_ASAP7_75t_R FILLER_0_107_755 ();
 FILLER_ASAP7_75t_R FILLER_0_107_767 ();
 FILLER_ASAP7_75t_R FILLER_0_107_779 ();
 DECAPx2_ASAP7_75t_R FILLER_0_107_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_797 ();
 FILLER_ASAP7_75t_R FILLER_0_107_805 ();
 FILLER_ASAP7_75t_R FILLER_0_107_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_815 ();
 FILLER_ASAP7_75t_R FILLER_0_107_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_828 ();
 FILLER_ASAP7_75t_R FILLER_0_107_839 ();
 DECAPx1_ASAP7_75t_R FILLER_0_107_853 ();
 DECAPx2_ASAP7_75t_R FILLER_0_107_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_872 ();
 FILLER_ASAP7_75t_R FILLER_0_107_883 ();
 FILLER_ASAP7_75t_R FILLER_0_107_892 ();
 FILLER_ASAP7_75t_R FILLER_0_107_897 ();
 DECAPx2_ASAP7_75t_R FILLER_0_107_919 ();
 DECAPx6_ASAP7_75t_R FILLER_0_107_927 ();
 DECAPx2_ASAP7_75t_R FILLER_0_107_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_947 ();
 FILLER_ASAP7_75t_R FILLER_0_107_960 ();
 DECAPx2_ASAP7_75t_R FILLER_0_107_982 ();
 DECAPx2_ASAP7_75t_R FILLER_0_107_994 ();
 FILLER_ASAP7_75t_R FILLER_0_107_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_1002 ();
 DECAPx6_ASAP7_75t_R FILLER_0_107_1011 ();
 FILLER_ASAP7_75t_R FILLER_0_107_1032 ();
 DECAPx2_ASAP7_75t_R FILLER_0_107_1040 ();
 FILLER_ASAP7_75t_R FILLER_0_107_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_1048 ();
 FILLER_ASAP7_75t_R FILLER_0_107_1055 ();
 FILLER_ASAP7_75t_R FILLER_0_107_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_1067 ();
 FILLER_ASAP7_75t_R FILLER_0_107_1074 ();
 FILLER_ASAP7_75t_R FILLER_0_107_1082 ();
 DECAPx4_ASAP7_75t_R FILLER_0_107_1104 ();
 FILLER_ASAP7_75t_R FILLER_0_107_1114 ();
 FILLER_ASAP7_75t_R FILLER_0_107_1122 ();
 FILLER_ASAP7_75t_R FILLER_0_107_1130 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_1135 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_1179 ();
 DECAPx4_ASAP7_75t_R FILLER_0_107_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_1201 ();
 FILLER_ASAP7_75t_R FILLER_0_107_1208 ();
 FILLER_ASAP7_75t_R FILLER_0_107_1216 ();
 FILLER_ASAP7_75t_R FILLER_0_107_1224 ();
 FILLER_ASAP7_75t_R FILLER_0_107_1232 ();
 FILLER_ASAP7_75t_R FILLER_0_107_1240 ();
 FILLER_ASAP7_75t_R FILLER_0_107_1248 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_1250 ();
 DECAPx2_ASAP7_75t_R FILLER_0_107_1257 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_1263 ();
 DECAPx1_ASAP7_75t_R FILLER_0_107_1271 ();
 DECAPx6_ASAP7_75t_R FILLER_0_107_1281 ();
 DECAPx1_ASAP7_75t_R FILLER_0_107_1295 ();
 DECAPx1_ASAP7_75t_R FILLER_0_107_1319 ();
 DECAPx1_ASAP7_75t_R FILLER_0_107_1330 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_1334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_1345 ();
 FILLER_ASAP7_75t_R FILLER_0_107_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_107_1380 ();
 DECAPx1_ASAP7_75t_R FILLER_0_108_2 ();
 FILLER_ASAP7_75t_R FILLER_0_108_11 ();
 FILLER_ASAP7_75t_R FILLER_0_108_18 ();
 FILLER_ASAP7_75t_R FILLER_0_108_23 ();
 FILLER_ASAP7_75t_R FILLER_0_108_33 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_40 ();
 DECAPx6_ASAP7_75t_R FILLER_0_108_62 ();
 DECAPx2_ASAP7_75t_R FILLER_0_108_76 ();
 FILLER_ASAP7_75t_R FILLER_0_108_88 ();
 DECAPx2_ASAP7_75t_R FILLER_0_108_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_102 ();
 DECAPx1_ASAP7_75t_R FILLER_0_108_123 ();
 DECAPx4_ASAP7_75t_R FILLER_0_108_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_147 ();
 FILLER_ASAP7_75t_R FILLER_0_108_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_170 ();
 DECAPx4_ASAP7_75t_R FILLER_0_108_177 ();
 FILLER_ASAP7_75t_R FILLER_0_108_197 ();
 DECAPx2_ASAP7_75t_R FILLER_0_108_206 ();
 DECAPx2_ASAP7_75t_R FILLER_0_108_222 ();
 FILLER_ASAP7_75t_R FILLER_0_108_228 ();
 FILLER_ASAP7_75t_R FILLER_0_108_241 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_249 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_293 ();
 DECAPx2_ASAP7_75t_R FILLER_0_108_312 ();
 FILLER_ASAP7_75t_R FILLER_0_108_324 ();
 DECAPx1_ASAP7_75t_R FILLER_0_108_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_335 ();
 DECAPx4_ASAP7_75t_R FILLER_0_108_346 ();
 FILLER_ASAP7_75t_R FILLER_0_108_356 ();
 DECAPx2_ASAP7_75t_R FILLER_0_108_368 ();
 FILLER_ASAP7_75t_R FILLER_0_108_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_376 ();
 FILLER_ASAP7_75t_R FILLER_0_108_383 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_412 ();
 DECAPx4_ASAP7_75t_R FILLER_0_108_434 ();
 DECAPx1_ASAP7_75t_R FILLER_0_108_450 ();
 FILLER_ASAP7_75t_R FILLER_0_108_460 ();
 FILLER_ASAP7_75t_R FILLER_0_108_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_494 ();
 FILLER_ASAP7_75t_R FILLER_0_108_498 ();
 FILLER_ASAP7_75t_R FILLER_0_108_514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_108_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_531 ();
 FILLER_ASAP7_75t_R FILLER_0_108_542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_108_554 ();
 FILLER_ASAP7_75t_R FILLER_0_108_568 ();
 DECAPx1_ASAP7_75t_R FILLER_0_108_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_580 ();
 FILLER_ASAP7_75t_R FILLER_0_108_591 ();
 FILLER_ASAP7_75t_R FILLER_0_108_603 ();
 DECAPx2_ASAP7_75t_R FILLER_0_108_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_621 ();
 FILLER_ASAP7_75t_R FILLER_0_108_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_634 ();
 FILLER_ASAP7_75t_R FILLER_0_108_641 ();
 FILLER_ASAP7_75t_R FILLER_0_108_653 ();
 FILLER_ASAP7_75t_R FILLER_0_108_665 ();
 FILLER_ASAP7_75t_R FILLER_0_108_671 ();
 FILLER_ASAP7_75t_R FILLER_0_108_680 ();
 FILLER_ASAP7_75t_R FILLER_0_108_692 ();
 FILLER_ASAP7_75t_R FILLER_0_108_704 ();
 DECAPx1_ASAP7_75t_R FILLER_0_108_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_718 ();
 FILLER_ASAP7_75t_R FILLER_0_108_729 ();
 FILLER_ASAP7_75t_R FILLER_0_108_737 ();
 FILLER_ASAP7_75t_R FILLER_0_108_757 ();
 DECAPx1_ASAP7_75t_R FILLER_0_108_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_769 ();
 FILLER_ASAP7_75t_R FILLER_0_108_780 ();
 FILLER_ASAP7_75t_R FILLER_0_108_792 ();
 FILLER_ASAP7_75t_R FILLER_0_108_799 ();
 FILLER_ASAP7_75t_R FILLER_0_108_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_808 ();
 DECAPx1_ASAP7_75t_R FILLER_0_108_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_820 ();
 DECAPx6_ASAP7_75t_R FILLER_0_108_826 ();
 FILLER_ASAP7_75t_R FILLER_0_108_840 ();
 DECAPx2_ASAP7_75t_R FILLER_0_108_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_855 ();
 FILLER_ASAP7_75t_R FILLER_0_108_860 ();
 DECAPx2_ASAP7_75t_R FILLER_0_108_868 ();
 FILLER_ASAP7_75t_R FILLER_0_108_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_876 ();
 FILLER_ASAP7_75t_R FILLER_0_108_885 ();
 DECAPx2_ASAP7_75t_R FILLER_0_108_894 ();
 FILLER_ASAP7_75t_R FILLER_0_108_900 ();
 DECAPx1_ASAP7_75t_R FILLER_0_108_912 ();
 FILLER_ASAP7_75t_R FILLER_0_108_937 ();
 DECAPx2_ASAP7_75t_R FILLER_0_108_942 ();
 DECAPx2_ASAP7_75t_R FILLER_0_108_954 ();
 FILLER_ASAP7_75t_R FILLER_0_108_960 ();
 DECAPx1_ASAP7_75t_R FILLER_0_108_968 ();
 FILLER_ASAP7_75t_R FILLER_0_108_978 ();
 DECAPx1_ASAP7_75t_R FILLER_0_108_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_990 ();
 FILLER_ASAP7_75t_R FILLER_0_108_1001 ();
 DECAPx4_ASAP7_75t_R FILLER_0_108_1009 ();
 FILLER_ASAP7_75t_R FILLER_0_108_1019 ();
 FILLER_ASAP7_75t_R FILLER_0_108_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_1029 ();
 DECAPx1_ASAP7_75t_R FILLER_0_108_1036 ();
 FILLER_ASAP7_75t_R FILLER_0_108_1051 ();
 DECAPx2_ASAP7_75t_R FILLER_0_108_1059 ();
 FILLER_ASAP7_75t_R FILLER_0_108_1065 ();
 FILLER_ASAP7_75t_R FILLER_0_108_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_0_108_1079 ();
 FILLER_ASAP7_75t_R FILLER_0_108_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_1087 ();
 FILLER_ASAP7_75t_R FILLER_0_108_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_1105 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_1127 ();
 FILLER_ASAP7_75t_R FILLER_0_108_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_1151 ();
 FILLER_ASAP7_75t_R FILLER_0_108_1155 ();
 FILLER_ASAP7_75t_R FILLER_0_108_1163 ();
 FILLER_ASAP7_75t_R FILLER_0_108_1171 ();
 FILLER_ASAP7_75t_R FILLER_0_108_1179 ();
 DECAPx1_ASAP7_75t_R FILLER_0_108_1187 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_1201 ();
 DECAPx4_ASAP7_75t_R FILLER_0_108_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_1239 ();
 DECAPx6_ASAP7_75t_R FILLER_0_108_1261 ();
 FILLER_ASAP7_75t_R FILLER_0_108_1275 ();
 FILLER_ASAP7_75t_R FILLER_0_108_1297 ();
 FILLER_ASAP7_75t_R FILLER_0_108_1309 ();
 FILLER_ASAP7_75t_R FILLER_0_108_1331 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_1333 ();
 FILLER_ASAP7_75t_R FILLER_0_108_1340 ();
 DECAPx4_ASAP7_75t_R FILLER_0_108_1352 ();
 FILLER_ASAP7_75t_R FILLER_0_108_1365 ();
 DECAPx1_ASAP7_75t_R FILLER_0_108_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_108_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_109_2 ();
 FILLER_ASAP7_75t_R FILLER_0_109_25 ();
 DECAPx2_ASAP7_75t_R FILLER_0_109_33 ();
 FILLER_ASAP7_75t_R FILLER_0_109_39 ();
 DECAPx4_ASAP7_75t_R FILLER_0_109_47 ();
 DECAPx6_ASAP7_75t_R FILLER_0_109_67 ();
 FILLER_ASAP7_75t_R FILLER_0_109_92 ();
 DECAPx6_ASAP7_75t_R FILLER_0_109_100 ();
 DECAPx2_ASAP7_75t_R FILLER_0_109_120 ();
 DECAPx2_ASAP7_75t_R FILLER_0_109_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_142 ();
 DECAPx2_ASAP7_75t_R FILLER_0_109_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_157 ();
 FILLER_ASAP7_75t_R FILLER_0_109_164 ();
 FILLER_ASAP7_75t_R FILLER_0_109_172 ();
 DECAPx2_ASAP7_75t_R FILLER_0_109_179 ();
 FILLER_ASAP7_75t_R FILLER_0_109_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_187 ();
 DECAPx2_ASAP7_75t_R FILLER_0_109_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_202 ();
 DECAPx2_ASAP7_75t_R FILLER_0_109_209 ();
 DECAPx4_ASAP7_75t_R FILLER_0_109_221 ();
 DECAPx2_ASAP7_75t_R FILLER_0_109_241 ();
 DECAPx4_ASAP7_75t_R FILLER_0_109_258 ();
 FILLER_ASAP7_75t_R FILLER_0_109_268 ();
 DECAPx1_ASAP7_75t_R FILLER_0_109_291 ();
 DECAPx2_ASAP7_75t_R FILLER_0_109_300 ();
 FILLER_ASAP7_75t_R FILLER_0_109_310 ();
 FILLER_ASAP7_75t_R FILLER_0_109_333 ();
 FILLER_ASAP7_75t_R FILLER_0_109_341 ();
 FILLER_ASAP7_75t_R FILLER_0_109_348 ();
 DECAPx4_ASAP7_75t_R FILLER_0_109_353 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_369 ();
 DECAPx2_ASAP7_75t_R FILLER_0_109_391 ();
 FILLER_ASAP7_75t_R FILLER_0_109_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_399 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_403 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_425 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_447 ();
 DECAPx6_ASAP7_75t_R FILLER_0_109_469 ();
 FILLER_ASAP7_75t_R FILLER_0_109_483 ();
 FILLER_ASAP7_75t_R FILLER_0_109_491 ();
 DECAPx4_ASAP7_75t_R FILLER_0_109_500 ();
 FILLER_ASAP7_75t_R FILLER_0_109_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_512 ();
 FILLER_ASAP7_75t_R FILLER_0_109_519 ();
 FILLER_ASAP7_75t_R FILLER_0_109_530 ();
 FILLER_ASAP7_75t_R FILLER_0_109_542 ();
 FILLER_ASAP7_75t_R FILLER_0_109_558 ();
 FILLER_ASAP7_75t_R FILLER_0_109_568 ();
 DECAPx1_ASAP7_75t_R FILLER_0_109_577 ();
 FILLER_ASAP7_75t_R FILLER_0_109_587 ();
 FILLER_ASAP7_75t_R FILLER_0_109_596 ();
 FILLER_ASAP7_75t_R FILLER_0_109_606 ();
 FILLER_ASAP7_75t_R FILLER_0_109_615 ();
 FILLER_ASAP7_75t_R FILLER_0_109_622 ();
 DECAPx1_ASAP7_75t_R FILLER_0_109_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_638 ();
 FILLER_ASAP7_75t_R FILLER_0_109_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_651 ();
 FILLER_ASAP7_75t_R FILLER_0_109_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_664 ();
 FILLER_ASAP7_75t_R FILLER_0_109_670 ();
 FILLER_ASAP7_75t_R FILLER_0_109_682 ();
 FILLER_ASAP7_75t_R FILLER_0_109_694 ();
 FILLER_ASAP7_75t_R FILLER_0_109_706 ();
 FILLER_ASAP7_75t_R FILLER_0_109_716 ();
 DECAPx1_ASAP7_75t_R FILLER_0_109_728 ();
 FILLER_ASAP7_75t_R FILLER_0_109_742 ();
 FILLER_ASAP7_75t_R FILLER_0_109_754 ();
 DECAPx1_ASAP7_75t_R FILLER_0_109_764 ();
 FILLER_ASAP7_75t_R FILLER_0_109_788 ();
 FILLER_ASAP7_75t_R FILLER_0_109_796 ();
 FILLER_ASAP7_75t_R FILLER_0_109_804 ();
 DECAPx2_ASAP7_75t_R FILLER_0_109_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_822 ();
 FILLER_ASAP7_75t_R FILLER_0_109_831 ();
 DECAPx2_ASAP7_75t_R FILLER_0_109_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_849 ();
 FILLER_ASAP7_75t_R FILLER_0_109_860 ();
 DECAPx4_ASAP7_75t_R FILLER_0_109_868 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_884 ();
 DECAPx4_ASAP7_75t_R FILLER_0_109_906 ();
 FILLER_ASAP7_75t_R FILLER_0_109_916 ();
 DECAPx1_ASAP7_75t_R FILLER_0_109_921 ();
 DECAPx6_ASAP7_75t_R FILLER_0_109_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_941 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_953 ();
 FILLER_ASAP7_75t_R FILLER_0_109_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_977 ();
 FILLER_ASAP7_75t_R FILLER_0_109_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_986 ();
 FILLER_ASAP7_75t_R FILLER_0_109_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_995 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_1002 ();
 DECAPx2_ASAP7_75t_R FILLER_0_109_1024 ();
 FILLER_ASAP7_75t_R FILLER_0_109_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_1032 ();
 DECAPx6_ASAP7_75t_R FILLER_0_109_1039 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_1053 ();
 DECAPx2_ASAP7_75t_R FILLER_0_109_1059 ();
 FILLER_ASAP7_75t_R FILLER_0_109_1071 ();
 DECAPx6_ASAP7_75t_R FILLER_0_109_1079 ();
 FILLER_ASAP7_75t_R FILLER_0_109_1093 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_1095 ();
 DECAPx4_ASAP7_75t_R FILLER_0_109_1102 ();
 FILLER_ASAP7_75t_R FILLER_0_109_1112 ();
 FILLER_ASAP7_75t_R FILLER_0_109_1135 ();
 DECAPx4_ASAP7_75t_R FILLER_0_109_1147 ();
 FILLER_ASAP7_75t_R FILLER_0_109_1157 ();
 FILLER_ASAP7_75t_R FILLER_0_109_1162 ();
 FILLER_ASAP7_75t_R FILLER_0_109_1174 ();
 FILLER_ASAP7_75t_R FILLER_0_109_1182 ();
 DECAPx1_ASAP7_75t_R FILLER_0_109_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_1194 ();
 FILLER_ASAP7_75t_R FILLER_0_109_1201 ();
 DECAPx2_ASAP7_75t_R FILLER_0_109_1209 ();
 FILLER_ASAP7_75t_R FILLER_0_109_1215 ();
 DECAPx4_ASAP7_75t_R FILLER_0_109_1228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_1249 ();
 DECAPx2_ASAP7_75t_R FILLER_0_109_1271 ();
 FILLER_ASAP7_75t_R FILLER_0_109_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_1292 ();
 FILLER_ASAP7_75t_R FILLER_0_109_1314 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_1316 ();
 DECAPx6_ASAP7_75t_R FILLER_0_109_1325 ();
 FILLER_ASAP7_75t_R FILLER_0_109_1339 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_1341 ();
 DECAPx4_ASAP7_75t_R FILLER_0_109_1345 ();
 FILLER_ASAP7_75t_R FILLER_0_109_1355 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_109_1363 ();
 FILLER_ASAP7_75t_R FILLER_0_109_1370 ();
 DECAPx1_ASAP7_75t_R FILLER_0_109_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_110_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_4 ();
 FILLER_ASAP7_75t_R FILLER_0_110_11 ();
 FILLER_ASAP7_75t_R FILLER_0_110_18 ();
 FILLER_ASAP7_75t_R FILLER_0_110_25 ();
 DECAPx2_ASAP7_75t_R FILLER_0_110_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_39 ();
 DECAPx1_ASAP7_75t_R FILLER_0_110_46 ();
 FILLER_ASAP7_75t_R FILLER_0_110_56 ();
 DECAPx6_ASAP7_75t_R FILLER_0_110_64 ();
 DECAPx1_ASAP7_75t_R FILLER_0_110_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_82 ();
 DECAPx6_ASAP7_75t_R FILLER_0_110_89 ();
 FILLER_ASAP7_75t_R FILLER_0_110_109 ();
 FILLER_ASAP7_75t_R FILLER_0_110_118 ();
 DECAPx1_ASAP7_75t_R FILLER_0_110_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_130 ();
 FILLER_ASAP7_75t_R FILLER_0_110_141 ();
 FILLER_ASAP7_75t_R FILLER_0_110_151 ();
 FILLER_ASAP7_75t_R FILLER_0_110_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_158 ();
 FILLER_ASAP7_75t_R FILLER_0_110_165 ();
 FILLER_ASAP7_75t_R FILLER_0_110_174 ();
 DECAPx1_ASAP7_75t_R FILLER_0_110_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_186 ();
 FILLER_ASAP7_75t_R FILLER_0_110_197 ();
 FILLER_ASAP7_75t_R FILLER_0_110_205 ();
 DECAPx4_ASAP7_75t_R FILLER_0_110_212 ();
 FILLER_ASAP7_75t_R FILLER_0_110_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_224 ();
 FILLER_ASAP7_75t_R FILLER_0_110_232 ();
 FILLER_ASAP7_75t_R FILLER_0_110_244 ();
 DECAPx1_ASAP7_75t_R FILLER_0_110_252 ();
 DECAPx4_ASAP7_75t_R FILLER_0_110_262 ();
 DECAPx4_ASAP7_75t_R FILLER_0_110_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_288 ();
 FILLER_ASAP7_75t_R FILLER_0_110_292 ();
 FILLER_ASAP7_75t_R FILLER_0_110_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_306 ();
 FILLER_ASAP7_75t_R FILLER_0_110_310 ();
 FILLER_ASAP7_75t_R FILLER_0_110_318 ();
 FILLER_ASAP7_75t_R FILLER_0_110_325 ();
 DECAPx6_ASAP7_75t_R FILLER_0_110_330 ();
 FILLER_ASAP7_75t_R FILLER_0_110_348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_356 ();
 DECAPx1_ASAP7_75t_R FILLER_0_110_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_382 ();
 DECAPx1_ASAP7_75t_R FILLER_0_110_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_399 ();
 DECAPx1_ASAP7_75t_R FILLER_0_110_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_412 ();
 FILLER_ASAP7_75t_R FILLER_0_110_434 ();
 DECAPx2_ASAP7_75t_R FILLER_0_110_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_453 ();
 FILLER_ASAP7_75t_R FILLER_0_110_460 ();
 FILLER_ASAP7_75t_R FILLER_0_110_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_476 ();
 DECAPx4_ASAP7_75t_R FILLER_0_110_498 ();
 DECAPx6_ASAP7_75t_R FILLER_0_110_518 ();
 DECAPx2_ASAP7_75t_R FILLER_0_110_540 ();
 FILLER_ASAP7_75t_R FILLER_0_110_556 ();
 FILLER_ASAP7_75t_R FILLER_0_110_576 ();
 DECAPx2_ASAP7_75t_R FILLER_0_110_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_595 ();
 DECAPx2_ASAP7_75t_R FILLER_0_110_608 ();
 FILLER_ASAP7_75t_R FILLER_0_110_620 ();
 FILLER_ASAP7_75t_R FILLER_0_110_628 ();
 FILLER_ASAP7_75t_R FILLER_0_110_640 ();
 DECAPx2_ASAP7_75t_R FILLER_0_110_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_658 ();
 FILLER_ASAP7_75t_R FILLER_0_110_664 ();
 FILLER_ASAP7_75t_R FILLER_0_110_671 ();
 FILLER_ASAP7_75t_R FILLER_0_110_683 ();
 FILLER_ASAP7_75t_R FILLER_0_110_695 ();
 FILLER_ASAP7_75t_R FILLER_0_110_707 ();
 FILLER_ASAP7_75t_R FILLER_0_110_715 ();
 FILLER_ASAP7_75t_R FILLER_0_110_727 ();
 FILLER_ASAP7_75t_R FILLER_0_110_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_741 ();
 FILLER_ASAP7_75t_R FILLER_0_110_752 ();
 FILLER_ASAP7_75t_R FILLER_0_110_762 ();
 FILLER_ASAP7_75t_R FILLER_0_110_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_769 ();
 DECAPx2_ASAP7_75t_R FILLER_0_110_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_786 ();
 FILLER_ASAP7_75t_R FILLER_0_110_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_799 ();
 FILLER_ASAP7_75t_R FILLER_0_110_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_812 ();
 FILLER_ASAP7_75t_R FILLER_0_110_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_821 ();
 DECAPx1_ASAP7_75t_R FILLER_0_110_833 ();
 DECAPx6_ASAP7_75t_R FILLER_0_110_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_857 ();
 FILLER_ASAP7_75t_R FILLER_0_110_863 ();
 DECAPx1_ASAP7_75t_R FILLER_0_110_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_877 ();
 FILLER_ASAP7_75t_R FILLER_0_110_888 ();
 FILLER_ASAP7_75t_R FILLER_0_110_914 ();
 DECAPx6_ASAP7_75t_R FILLER_0_110_928 ();
 DECAPx2_ASAP7_75t_R FILLER_0_110_942 ();
 FILLER_ASAP7_75t_R FILLER_0_110_954 ();
 FILLER_ASAP7_75t_R FILLER_0_110_959 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_967 ();
 DECAPx6_ASAP7_75t_R FILLER_0_110_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_1003 ();
 FILLER_ASAP7_75t_R FILLER_0_110_1024 ();
 DECAPx4_ASAP7_75t_R FILLER_0_110_1036 ();
 DECAPx6_ASAP7_75t_R FILLER_0_110_1052 ();
 FILLER_ASAP7_75t_R FILLER_0_110_1066 ();
 FILLER_ASAP7_75t_R FILLER_0_110_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_1082 ();
 DECAPx4_ASAP7_75t_R FILLER_0_110_1104 ();
 FILLER_ASAP7_75t_R FILLER_0_110_1114 ();
 DECAPx4_ASAP7_75t_R FILLER_0_110_1119 ();
 FILLER_ASAP7_75t_R FILLER_0_110_1129 ();
 FILLER_ASAP7_75t_R FILLER_0_110_1151 ();
 FILLER_ASAP7_75t_R FILLER_0_110_1159 ();
 DECAPx2_ASAP7_75t_R FILLER_0_110_1167 ();
 FILLER_ASAP7_75t_R FILLER_0_110_1173 ();
 FILLER_ASAP7_75t_R FILLER_0_110_1183 ();
 DECAPx1_ASAP7_75t_R FILLER_0_110_1193 ();
 FILLER_ASAP7_75t_R FILLER_0_110_1203 ();
 DECAPx2_ASAP7_75t_R FILLER_0_110_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_1217 ();
 DECAPx2_ASAP7_75t_R FILLER_0_110_1224 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_1230 ();
 FILLER_ASAP7_75t_R FILLER_0_110_1237 ();
 DECAPx6_ASAP7_75t_R FILLER_0_110_1245 ();
 DECAPx1_ASAP7_75t_R FILLER_0_110_1259 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_1273 ();
 FILLER_ASAP7_75t_R FILLER_0_110_1295 ();
 DECAPx2_ASAP7_75t_R FILLER_0_110_1303 ();
 FILLER_ASAP7_75t_R FILLER_0_110_1315 ();
 FILLER_ASAP7_75t_R FILLER_0_110_1323 ();
 FILLER_ASAP7_75t_R FILLER_0_110_1333 ();
 DECAPx4_ASAP7_75t_R FILLER_0_110_1341 ();
 FILLER_ASAP7_75t_R FILLER_0_110_1351 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_1353 ();
 FILLER_ASAP7_75t_R FILLER_0_110_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_110_1380 ();
 DECAPx2_ASAP7_75t_R FILLER_0_111_2 ();
 FILLER_ASAP7_75t_R FILLER_0_111_13 ();
 FILLER_ASAP7_75t_R FILLER_0_111_18 ();
 DECAPx1_ASAP7_75t_R FILLER_0_111_25 ();
 FILLER_ASAP7_75t_R FILLER_0_111_35 ();
 FILLER_ASAP7_75t_R FILLER_0_111_48 ();
 FILLER_ASAP7_75t_R FILLER_0_111_56 ();
 FILLER_ASAP7_75t_R FILLER_0_111_64 ();
 FILLER_ASAP7_75t_R FILLER_0_111_82 ();
 DECAPx1_ASAP7_75t_R FILLER_0_111_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_94 ();
 FILLER_ASAP7_75t_R FILLER_0_111_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_102 ();
 DECAPx2_ASAP7_75t_R FILLER_0_111_111 ();
 FILLER_ASAP7_75t_R FILLER_0_111_117 ();
 FILLER_ASAP7_75t_R FILLER_0_111_129 ();
 FILLER_ASAP7_75t_R FILLER_0_111_141 ();
 DECAPx2_ASAP7_75t_R FILLER_0_111_149 ();
 FILLER_ASAP7_75t_R FILLER_0_111_161 ();
 DECAPx2_ASAP7_75t_R FILLER_0_111_168 ();
 FILLER_ASAP7_75t_R FILLER_0_111_174 ();
 FILLER_ASAP7_75t_R FILLER_0_111_181 ();
 DECAPx2_ASAP7_75t_R FILLER_0_111_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_195 ();
 FILLER_ASAP7_75t_R FILLER_0_111_204 ();
 FILLER_ASAP7_75t_R FILLER_0_111_212 ();
 FILLER_ASAP7_75t_R FILLER_0_111_220 ();
 DECAPx6_ASAP7_75t_R FILLER_0_111_228 ();
 DECAPx2_ASAP7_75t_R FILLER_0_111_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_248 ();
 DECAPx6_ASAP7_75t_R FILLER_0_111_255 ();
 DECAPx4_ASAP7_75t_R FILLER_0_111_281 ();
 FILLER_ASAP7_75t_R FILLER_0_111_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_293 ();
 DECAPx2_ASAP7_75t_R FILLER_0_111_300 ();
 FILLER_ASAP7_75t_R FILLER_0_111_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_308 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_315 ();
 DECAPx4_ASAP7_75t_R FILLER_0_111_337 ();
 FILLER_ASAP7_75t_R FILLER_0_111_347 ();
 FILLER_ASAP7_75t_R FILLER_0_111_370 ();
 DECAPx1_ASAP7_75t_R FILLER_0_111_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_380 ();
 DECAPx1_ASAP7_75t_R FILLER_0_111_393 ();
 FILLER_ASAP7_75t_R FILLER_0_111_400 ();
 DECAPx1_ASAP7_75t_R FILLER_0_111_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_440 ();
 FILLER_ASAP7_75t_R FILLER_0_111_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_449 ();
 FILLER_ASAP7_75t_R FILLER_0_111_458 ();
 FILLER_ASAP7_75t_R FILLER_0_111_466 ();
 DECAPx2_ASAP7_75t_R FILLER_0_111_478 ();
 FILLER_ASAP7_75t_R FILLER_0_111_484 ();
 DECAPx1_ASAP7_75t_R FILLER_0_111_492 ();
 FILLER_ASAP7_75t_R FILLER_0_111_516 ();
 DECAPx1_ASAP7_75t_R FILLER_0_111_528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_111_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_543 ();
 DECAPx2_ASAP7_75t_R FILLER_0_111_549 ();
 FILLER_ASAP7_75t_R FILLER_0_111_560 ();
 FILLER_ASAP7_75t_R FILLER_0_111_574 ();
 DECAPx6_ASAP7_75t_R FILLER_0_111_583 ();
 DECAPx1_ASAP7_75t_R FILLER_0_111_597 ();
 FILLER_ASAP7_75t_R FILLER_0_111_607 ();
 FILLER_ASAP7_75t_R FILLER_0_111_619 ();
 DECAPx1_ASAP7_75t_R FILLER_0_111_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_635 ();
 FILLER_ASAP7_75t_R FILLER_0_111_646 ();
 DECAPx2_ASAP7_75t_R FILLER_0_111_653 ();
 FILLER_ASAP7_75t_R FILLER_0_111_664 ();
 FILLER_ASAP7_75t_R FILLER_0_111_671 ();
 DECAPx1_ASAP7_75t_R FILLER_0_111_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_687 ();
 FILLER_ASAP7_75t_R FILLER_0_111_698 ();
 DECAPx2_ASAP7_75t_R FILLER_0_111_710 ();
 FILLER_ASAP7_75t_R FILLER_0_111_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_728 ();
 FILLER_ASAP7_75t_R FILLER_0_111_734 ();
 FILLER_ASAP7_75t_R FILLER_0_111_746 ();
 DECAPx2_ASAP7_75t_R FILLER_0_111_758 ();
 FILLER_ASAP7_75t_R FILLER_0_111_774 ();
 FILLER_ASAP7_75t_R FILLER_0_111_782 ();
 DECAPx1_ASAP7_75t_R FILLER_0_111_792 ();
 FILLER_ASAP7_75t_R FILLER_0_111_806 ();
 FILLER_ASAP7_75t_R FILLER_0_111_818 ();
 FILLER_ASAP7_75t_R FILLER_0_111_830 ();
 DECAPx6_ASAP7_75t_R FILLER_0_111_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_852 ();
 FILLER_ASAP7_75t_R FILLER_0_111_863 ();
 FILLER_ASAP7_75t_R FILLER_0_111_875 ();
 DECAPx6_ASAP7_75t_R FILLER_0_111_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_903 ();
 FILLER_ASAP7_75t_R FILLER_0_111_909 ();
 DECAPx2_ASAP7_75t_R FILLER_0_111_917 ();
 FILLER_ASAP7_75t_R FILLER_0_111_923 ();
 DECAPx1_ASAP7_75t_R FILLER_0_111_927 ();
 DECAPx2_ASAP7_75t_R FILLER_0_111_937 ();
 FILLER_ASAP7_75t_R FILLER_0_111_943 ();
 FILLER_ASAP7_75t_R FILLER_0_111_948 ();
 FILLER_ASAP7_75t_R FILLER_0_111_960 ();
 FILLER_ASAP7_75t_R FILLER_0_111_972 ();
 FILLER_ASAP7_75t_R FILLER_0_111_1012 ();
 DECAPx4_ASAP7_75t_R FILLER_0_111_1017 ();
 FILLER_ASAP7_75t_R FILLER_0_111_1027 ();
 DECAPx2_ASAP7_75t_R FILLER_0_111_1032 ();
 FILLER_ASAP7_75t_R FILLER_0_111_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_1040 ();
 DECAPx2_ASAP7_75t_R FILLER_0_111_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_1057 ();
 FILLER_ASAP7_75t_R FILLER_0_111_1079 ();
 DECAPx2_ASAP7_75t_R FILLER_0_111_1087 ();
 FILLER_ASAP7_75t_R FILLER_0_111_1093 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_1101 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_1123 ();
 DECAPx2_ASAP7_75t_R FILLER_0_111_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_1151 ();
 DECAPx4_ASAP7_75t_R FILLER_0_111_1164 ();
 FILLER_ASAP7_75t_R FILLER_0_111_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_1176 ();
 FILLER_ASAP7_75t_R FILLER_0_111_1187 ();
 FILLER_ASAP7_75t_R FILLER_0_111_1195 ();
 FILLER_ASAP7_75t_R FILLER_0_111_1203 ();
 DECAPx2_ASAP7_75t_R FILLER_0_111_1211 ();
 DECAPx4_ASAP7_75t_R FILLER_0_111_1223 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_1233 ();
 FILLER_ASAP7_75t_R FILLER_0_111_1240 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_1242 ();
 FILLER_ASAP7_75t_R FILLER_0_111_1253 ();
 FILLER_ASAP7_75t_R FILLER_0_111_1275 ();
 DECAPx4_ASAP7_75t_R FILLER_0_111_1283 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_1293 ();
 FILLER_ASAP7_75t_R FILLER_0_111_1304 ();
 DECAPx4_ASAP7_75t_R FILLER_0_111_1313 ();
 DECAPx2_ASAP7_75t_R FILLER_0_111_1329 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_1335 ();
 DECAPx1_ASAP7_75t_R FILLER_0_111_1343 ();
 DECAPx1_ASAP7_75t_R FILLER_0_111_1368 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_1372 ();
 FILLER_ASAP7_75t_R FILLER_0_111_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_112_2 ();
 FILLER_ASAP7_75t_R FILLER_0_112_9 ();
 FILLER_ASAP7_75t_R FILLER_0_112_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_16 ();
 FILLER_ASAP7_75t_R FILLER_0_112_23 ();
 FILLER_ASAP7_75t_R FILLER_0_112_30 ();
 FILLER_ASAP7_75t_R FILLER_0_112_38 ();
 DECAPx2_ASAP7_75t_R FILLER_0_112_46 ();
 FILLER_ASAP7_75t_R FILLER_0_112_52 ();
 FILLER_ASAP7_75t_R FILLER_0_112_65 ();
 DECAPx2_ASAP7_75t_R FILLER_0_112_73 ();
 FILLER_ASAP7_75t_R FILLER_0_112_87 ();
 DECAPx1_ASAP7_75t_R FILLER_0_112_99 ();
 FILLER_ASAP7_75t_R FILLER_0_112_111 ();
 DECAPx2_ASAP7_75t_R FILLER_0_112_119 ();
 FILLER_ASAP7_75t_R FILLER_0_112_125 ();
 FILLER_ASAP7_75t_R FILLER_0_112_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_139 ();
 FILLER_ASAP7_75t_R FILLER_0_112_150 ();
 DECAPx2_ASAP7_75t_R FILLER_0_112_158 ();
 FILLER_ASAP7_75t_R FILLER_0_112_164 ();
 DECAPx4_ASAP7_75t_R FILLER_0_112_172 ();
 FILLER_ASAP7_75t_R FILLER_0_112_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_184 ();
 FILLER_ASAP7_75t_R FILLER_0_112_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_193 ();
 DECAPx2_ASAP7_75t_R FILLER_0_112_200 ();
 FILLER_ASAP7_75t_R FILLER_0_112_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_208 ();
 FILLER_ASAP7_75t_R FILLER_0_112_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_217 ();
 FILLER_ASAP7_75t_R FILLER_0_112_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_226 ();
 DECAPx6_ASAP7_75t_R FILLER_0_112_235 ();
 DECAPx1_ASAP7_75t_R FILLER_0_112_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_263 ();
 FILLER_ASAP7_75t_R FILLER_0_112_267 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_299 ();
 DECAPx2_ASAP7_75t_R FILLER_0_112_321 ();
 FILLER_ASAP7_75t_R FILLER_0_112_333 ();
 DECAPx1_ASAP7_75t_R FILLER_0_112_347 ();
 DECAPx6_ASAP7_75t_R FILLER_0_112_354 ();
 FILLER_ASAP7_75t_R FILLER_0_112_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_370 ();
 FILLER_ASAP7_75t_R FILLER_0_112_383 ();
 DECAPx1_ASAP7_75t_R FILLER_0_112_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_401 ();
 FILLER_ASAP7_75t_R FILLER_0_112_408 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_438 ();
 DECAPx2_ASAP7_75t_R FILLER_0_112_445 ();
 FILLER_ASAP7_75t_R FILLER_0_112_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_453 ();
 FILLER_ASAP7_75t_R FILLER_0_112_460 ();
 DECAPx1_ASAP7_75t_R FILLER_0_112_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_468 ();
 DECAPx1_ASAP7_75t_R FILLER_0_112_476 ();
 FILLER_ASAP7_75t_R FILLER_0_112_500 ();
 FILLER_ASAP7_75t_R FILLER_0_112_508 ();
 FILLER_ASAP7_75t_R FILLER_0_112_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_518 ();
 FILLER_ASAP7_75t_R FILLER_0_112_526 ();
 FILLER_ASAP7_75t_R FILLER_0_112_538 ();
 FILLER_ASAP7_75t_R FILLER_0_112_552 ();
 FILLER_ASAP7_75t_R FILLER_0_112_562 ();
 DECAPx2_ASAP7_75t_R FILLER_0_112_569 ();
 FILLER_ASAP7_75t_R FILLER_0_112_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_577 ();
 DECAPx4_ASAP7_75t_R FILLER_0_112_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_594 ();
 FILLER_ASAP7_75t_R FILLER_0_112_601 ();
 DECAPx1_ASAP7_75t_R FILLER_0_112_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_613 ();
 FILLER_ASAP7_75t_R FILLER_0_112_624 ();
 DECAPx2_ASAP7_75t_R FILLER_0_112_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_642 ();
 FILLER_ASAP7_75t_R FILLER_0_112_653 ();
 FILLER_ASAP7_75t_R FILLER_0_112_661 ();
 FILLER_ASAP7_75t_R FILLER_0_112_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_670 ();
 FILLER_ASAP7_75t_R FILLER_0_112_681 ();
 DECAPx2_ASAP7_75t_R FILLER_0_112_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_699 ();
 DECAPx1_ASAP7_75t_R FILLER_0_112_710 ();
 FILLER_ASAP7_75t_R FILLER_0_112_719 ();
 FILLER_ASAP7_75t_R FILLER_0_112_727 ();
 FILLER_ASAP7_75t_R FILLER_0_112_734 ();
 FILLER_ASAP7_75t_R FILLER_0_112_741 ();
 FILLER_ASAP7_75t_R FILLER_0_112_753 ();
 FILLER_ASAP7_75t_R FILLER_0_112_765 ();
 DECAPx2_ASAP7_75t_R FILLER_0_112_777 ();
 FILLER_ASAP7_75t_R FILLER_0_112_783 ();
 DECAPx2_ASAP7_75t_R FILLER_0_112_795 ();
 FILLER_ASAP7_75t_R FILLER_0_112_811 ();
 DECAPx2_ASAP7_75t_R FILLER_0_112_823 ();
 FILLER_ASAP7_75t_R FILLER_0_112_829 ();
 FILLER_ASAP7_75t_R FILLER_0_112_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_844 ();
 FILLER_ASAP7_75t_R FILLER_0_112_855 ();
 FILLER_ASAP7_75t_R FILLER_0_112_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_865 ();
 FILLER_ASAP7_75t_R FILLER_0_112_876 ();
 DECAPx1_ASAP7_75t_R FILLER_0_112_883 ();
 DECAPx2_ASAP7_75t_R FILLER_0_112_925 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_931 ();
 FILLER_ASAP7_75t_R FILLER_0_112_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_940 ();
 FILLER_ASAP7_75t_R FILLER_0_112_963 ();
 FILLER_ASAP7_75t_R FILLER_0_112_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_970 ();
 DECAPx4_ASAP7_75t_R FILLER_0_112_974 ();
 FILLER_ASAP7_75t_R FILLER_0_112_984 ();
 DECAPx1_ASAP7_75t_R FILLER_0_112_1006 ();
 DECAPx1_ASAP7_75t_R FILLER_0_112_1016 ();
 DECAPx2_ASAP7_75t_R FILLER_0_112_1030 ();
 FILLER_ASAP7_75t_R FILLER_0_112_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_1038 ();
 FILLER_ASAP7_75t_R FILLER_0_112_1047 ();
 DECAPx2_ASAP7_75t_R FILLER_0_112_1070 ();
 FILLER_ASAP7_75t_R FILLER_0_112_1076 ();
 FILLER_ASAP7_75t_R FILLER_0_112_1088 ();
 FILLER_ASAP7_75t_R FILLER_0_112_1093 ();
 DECAPx4_ASAP7_75t_R FILLER_0_112_1107 ();
 FILLER_ASAP7_75t_R FILLER_0_112_1123 ();
 FILLER_ASAP7_75t_R FILLER_0_112_1131 ();
 DECAPx1_ASAP7_75t_R FILLER_0_112_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_1140 ();
 DECAPx1_ASAP7_75t_R FILLER_0_112_1151 ();
 FILLER_ASAP7_75t_R FILLER_0_112_1161 ();
 DECAPx2_ASAP7_75t_R FILLER_0_112_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_1177 ();
 FILLER_ASAP7_75t_R FILLER_0_112_1181 ();
 FILLER_ASAP7_75t_R FILLER_0_112_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_1191 ();
 DECAPx4_ASAP7_75t_R FILLER_0_112_1198 ();
 FILLER_ASAP7_75t_R FILLER_0_112_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_1210 ();
 FILLER_ASAP7_75t_R FILLER_0_112_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_1225 ();
 FILLER_ASAP7_75t_R FILLER_0_112_1247 ();
 DECAPx2_ASAP7_75t_R FILLER_0_112_1259 ();
 FILLER_ASAP7_75t_R FILLER_0_112_1265 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_1267 ();
 FILLER_ASAP7_75t_R FILLER_0_112_1274 ();
 DECAPx2_ASAP7_75t_R FILLER_0_112_1287 ();
 FILLER_ASAP7_75t_R FILLER_0_112_1293 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_1295 ();
 DECAPx1_ASAP7_75t_R FILLER_0_112_1302 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_1306 ();
 FILLER_ASAP7_75t_R FILLER_0_112_1313 ();
 FILLER_ASAP7_75t_R FILLER_0_112_1326 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_1328 ();
 FILLER_ASAP7_75t_R FILLER_0_112_1349 ();
 FILLER_ASAP7_75t_R FILLER_0_112_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_112_1365 ();
 FILLER_ASAP7_75t_R FILLER_0_112_1370 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_1372 ();
 FILLER_ASAP7_75t_R FILLER_0_112_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_113_2 ();
 FILLER_ASAP7_75t_R FILLER_0_113_9 ();
 DECAPx1_ASAP7_75t_R FILLER_0_113_16 ();
 FILLER_ASAP7_75t_R FILLER_0_113_25 ();
 FILLER_ASAP7_75t_R FILLER_0_113_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_34 ();
 DECAPx1_ASAP7_75t_R FILLER_0_113_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_45 ();
 DECAPx2_ASAP7_75t_R FILLER_0_113_52 ();
 FILLER_ASAP7_75t_R FILLER_0_113_58 ();
 DECAPx6_ASAP7_75t_R FILLER_0_113_63 ();
 DECAPx2_ASAP7_75t_R FILLER_0_113_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_83 ();
 FILLER_ASAP7_75t_R FILLER_0_113_94 ();
 FILLER_ASAP7_75t_R FILLER_0_113_101 ();
 FILLER_ASAP7_75t_R FILLER_0_113_110 ();
 FILLER_ASAP7_75t_R FILLER_0_113_118 ();
 FILLER_ASAP7_75t_R FILLER_0_113_130 ();
 FILLER_ASAP7_75t_R FILLER_0_113_142 ();
 DECAPx2_ASAP7_75t_R FILLER_0_113_150 ();
 FILLER_ASAP7_75t_R FILLER_0_113_166 ();
 DECAPx4_ASAP7_75t_R FILLER_0_113_174 ();
 FILLER_ASAP7_75t_R FILLER_0_113_184 ();
 DECAPx2_ASAP7_75t_R FILLER_0_113_192 ();
 FILLER_ASAP7_75t_R FILLER_0_113_198 ();
 DECAPx4_ASAP7_75t_R FILLER_0_113_212 ();
 DECAPx2_ASAP7_75t_R FILLER_0_113_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_231 ();
 DECAPx2_ASAP7_75t_R FILLER_0_113_238 ();
 FILLER_ASAP7_75t_R FILLER_0_113_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_246 ();
 DECAPx6_ASAP7_75t_R FILLER_0_113_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_267 ();
 DECAPx1_ASAP7_75t_R FILLER_0_113_274 ();
 FILLER_ASAP7_75t_R FILLER_0_113_299 ();
 FILLER_ASAP7_75t_R FILLER_0_113_307 ();
 FILLER_ASAP7_75t_R FILLER_0_113_314 ();
 DECAPx1_ASAP7_75t_R FILLER_0_113_321 ();
 DECAPx2_ASAP7_75t_R FILLER_0_113_346 ();
 FILLER_ASAP7_75t_R FILLER_0_113_352 ();
 DECAPx1_ASAP7_75t_R FILLER_0_113_364 ();
 FILLER_ASAP7_75t_R FILLER_0_113_374 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_404 ();
 DECAPx6_ASAP7_75t_R FILLER_0_113_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_440 ();
 DECAPx1_ASAP7_75t_R FILLER_0_113_448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_113_458 ();
 DECAPx1_ASAP7_75t_R FILLER_0_113_470 ();
 DECAPx2_ASAP7_75t_R FILLER_0_113_480 ();
 DECAPx2_ASAP7_75t_R FILLER_0_113_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_502 ();
 FILLER_ASAP7_75t_R FILLER_0_113_507 ();
 FILLER_ASAP7_75t_R FILLER_0_113_514 ();
 FILLER_ASAP7_75t_R FILLER_0_113_522 ();
 FILLER_ASAP7_75t_R FILLER_0_113_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_532 ();
 FILLER_ASAP7_75t_R FILLER_0_113_538 ();
 FILLER_ASAP7_75t_R FILLER_0_113_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_560 ();
 DECAPx1_ASAP7_75t_R FILLER_0_113_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_586 ();
 DECAPx1_ASAP7_75t_R FILLER_0_113_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_601 ();
 FILLER_ASAP7_75t_R FILLER_0_113_608 ();
 FILLER_ASAP7_75t_R FILLER_0_113_620 ();
 FILLER_ASAP7_75t_R FILLER_0_113_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_634 ();
 FILLER_ASAP7_75t_R FILLER_0_113_639 ();
 DECAPx1_ASAP7_75t_R FILLER_0_113_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_655 ();
 DECAPx1_ASAP7_75t_R FILLER_0_113_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_670 ();
 FILLER_ASAP7_75t_R FILLER_0_113_676 ();
 DECAPx1_ASAP7_75t_R FILLER_0_113_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_692 ();
 FILLER_ASAP7_75t_R FILLER_0_113_698 ();
 FILLER_ASAP7_75t_R FILLER_0_113_705 ();
 FILLER_ASAP7_75t_R FILLER_0_113_745 ();
 FILLER_ASAP7_75t_R FILLER_0_113_757 ();
 DECAPx2_ASAP7_75t_R FILLER_0_113_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_775 ();
 DECAPx2_ASAP7_75t_R FILLER_0_113_786 ();
 FILLER_ASAP7_75t_R FILLER_0_113_792 ();
 FILLER_ASAP7_75t_R FILLER_0_113_804 ();
 DECAPx1_ASAP7_75t_R FILLER_0_113_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_830 ();
 DECAPx2_ASAP7_75t_R FILLER_0_113_837 ();
 DECAPx1_ASAP7_75t_R FILLER_0_113_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_852 ();
 FILLER_ASAP7_75t_R FILLER_0_113_861 ();
 FILLER_ASAP7_75t_R FILLER_0_113_868 ();
 FILLER_ASAP7_75t_R FILLER_0_113_875 ();
 DECAPx1_ASAP7_75t_R FILLER_0_113_915 ();
 FILLER_ASAP7_75t_R FILLER_0_113_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_924 ();
 FILLER_ASAP7_75t_R FILLER_0_113_927 ();
 FILLER_ASAP7_75t_R FILLER_0_113_937 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_945 ();
 DECAPx2_ASAP7_75t_R FILLER_0_113_967 ();
 FILLER_ASAP7_75t_R FILLER_0_113_973 ();
 DECAPx2_ASAP7_75t_R FILLER_0_113_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_987 ();
 FILLER_ASAP7_75t_R FILLER_0_113_998 ();
 DECAPx2_ASAP7_75t_R FILLER_0_113_1006 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1012 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_1022 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1033 ();
 DECAPx2_ASAP7_75t_R FILLER_0_113_1043 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1049 ();
 DECAPx2_ASAP7_75t_R FILLER_0_113_1054 ();
 DECAPx4_ASAP7_75t_R FILLER_0_113_1063 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1081 ();
 DECAPx6_ASAP7_75t_R FILLER_0_113_1089 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_1105 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_1116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_1143 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1150 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1158 ();
 DECAPx2_ASAP7_75t_R FILLER_0_113_1166 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1172 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1177 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1185 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1193 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1201 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1209 ();
 DECAPx6_ASAP7_75t_R FILLER_0_113_1217 ();
 DECAPx1_ASAP7_75t_R FILLER_0_113_1237 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_1241 ();
 DECAPx1_ASAP7_75t_R FILLER_0_113_1248 ();
 DECAPx1_ASAP7_75t_R FILLER_0_113_1262 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_1266 ();
 DECAPx1_ASAP7_75t_R FILLER_0_113_1273 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_1277 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1284 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_1286 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1293 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1303 ();
 DECAPx6_ASAP7_75t_R FILLER_0_113_1315 ();
 DECAPx2_ASAP7_75t_R FILLER_0_113_1329 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_1335 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1341 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1348 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1356 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1361 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1368 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1375 ();
 FILLER_ASAP7_75t_R FILLER_0_113_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_114_2 ();
 FILLER_ASAP7_75t_R FILLER_0_114_9 ();
 DECAPx1_ASAP7_75t_R FILLER_0_114_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_20 ();
 FILLER_ASAP7_75t_R FILLER_0_114_26 ();
 DECAPx1_ASAP7_75t_R FILLER_0_114_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_35 ();
 FILLER_ASAP7_75t_R FILLER_0_114_42 ();
 DECAPx2_ASAP7_75t_R FILLER_0_114_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_57 ();
 DECAPx2_ASAP7_75t_R FILLER_0_114_70 ();
 FILLER_ASAP7_75t_R FILLER_0_114_82 ();
 FILLER_ASAP7_75t_R FILLER_0_114_90 ();
 FILLER_ASAP7_75t_R FILLER_0_114_98 ();
 FILLER_ASAP7_75t_R FILLER_0_114_106 ();
 FILLER_ASAP7_75t_R FILLER_0_114_118 ();
 FILLER_ASAP7_75t_R FILLER_0_114_130 ();
 FILLER_ASAP7_75t_R FILLER_0_114_142 ();
 FILLER_ASAP7_75t_R FILLER_0_114_152 ();
 FILLER_ASAP7_75t_R FILLER_0_114_160 ();
 DECAPx1_ASAP7_75t_R FILLER_0_114_168 ();
 FILLER_ASAP7_75t_R FILLER_0_114_177 ();
 FILLER_ASAP7_75t_R FILLER_0_114_185 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_193 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_215 ();
 DECAPx4_ASAP7_75t_R FILLER_0_114_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_247 ();
 FILLER_ASAP7_75t_R FILLER_0_114_251 ();
 DECAPx1_ASAP7_75t_R FILLER_0_114_259 ();
 DECAPx4_ASAP7_75t_R FILLER_0_114_269 ();
 FILLER_ASAP7_75t_R FILLER_0_114_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_281 ();
 FILLER_ASAP7_75t_R FILLER_0_114_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_296 ();
 DECAPx2_ASAP7_75t_R FILLER_0_114_300 ();
 FILLER_ASAP7_75t_R FILLER_0_114_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_308 ();
 DECAPx4_ASAP7_75t_R FILLER_0_114_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_322 ();
 FILLER_ASAP7_75t_R FILLER_0_114_329 ();
 DECAPx2_ASAP7_75t_R FILLER_0_114_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_340 ();
 DECAPx4_ASAP7_75t_R FILLER_0_114_347 ();
 FILLER_ASAP7_75t_R FILLER_0_114_357 ();
 FILLER_ASAP7_75t_R FILLER_0_114_365 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_375 ();
 DECAPx6_ASAP7_75t_R FILLER_0_114_407 ();
 DECAPx1_ASAP7_75t_R FILLER_0_114_421 ();
 DECAPx2_ASAP7_75t_R FILLER_0_114_436 ();
 FILLER_ASAP7_75t_R FILLER_0_114_442 ();
 FILLER_ASAP7_75t_R FILLER_0_114_451 ();
 FILLER_ASAP7_75t_R FILLER_0_114_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_461 ();
 FILLER_ASAP7_75t_R FILLER_0_114_464 ();
 FILLER_ASAP7_75t_R FILLER_0_114_474 ();
 DECAPx2_ASAP7_75t_R FILLER_0_114_486 ();
 DECAPx1_ASAP7_75t_R FILLER_0_114_498 ();
 DECAPx1_ASAP7_75t_R FILLER_0_114_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_516 ();
 FILLER_ASAP7_75t_R FILLER_0_114_523 ();
 DECAPx6_ASAP7_75t_R FILLER_0_114_530 ();
 FILLER_ASAP7_75t_R FILLER_0_114_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_546 ();
 DECAPx4_ASAP7_75t_R FILLER_0_114_553 ();
 DECAPx2_ASAP7_75t_R FILLER_0_114_568 ();
 FILLER_ASAP7_75t_R FILLER_0_114_574 ();
 FILLER_ASAP7_75t_R FILLER_0_114_582 ();
 DECAPx4_ASAP7_75t_R FILLER_0_114_590 ();
 FILLER_ASAP7_75t_R FILLER_0_114_600 ();
 FILLER_ASAP7_75t_R FILLER_0_114_607 ();
 FILLER_ASAP7_75t_R FILLER_0_114_615 ();
 FILLER_ASAP7_75t_R FILLER_0_114_627 ();
 FILLER_ASAP7_75t_R FILLER_0_114_639 ();
 FILLER_ASAP7_75t_R FILLER_0_114_651 ();
 FILLER_ASAP7_75t_R FILLER_0_114_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_665 ();
 DECAPx2_ASAP7_75t_R FILLER_0_114_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_682 ();
 FILLER_ASAP7_75t_R FILLER_0_114_689 ();
 FILLER_ASAP7_75t_R FILLER_0_114_695 ();
 FILLER_ASAP7_75t_R FILLER_0_114_707 ();
 FILLER_ASAP7_75t_R FILLER_0_114_719 ();
 FILLER_ASAP7_75t_R FILLER_0_114_739 ();
 FILLER_ASAP7_75t_R FILLER_0_114_751 ();
 FILLER_ASAP7_75t_R FILLER_0_114_763 ();
 DECAPx2_ASAP7_75t_R FILLER_0_114_775 ();
 FILLER_ASAP7_75t_R FILLER_0_114_791 ();
 FILLER_ASAP7_75t_R FILLER_0_114_803 ();
 FILLER_ASAP7_75t_R FILLER_0_114_810 ();
 FILLER_ASAP7_75t_R FILLER_0_114_822 ();
 FILLER_ASAP7_75t_R FILLER_0_114_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_831 ();
 DECAPx1_ASAP7_75t_R FILLER_0_114_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_842 ();
 DECAPx1_ASAP7_75t_R FILLER_0_114_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_867 ();
 DECAPx2_ASAP7_75t_R FILLER_0_114_892 ();
 FILLER_ASAP7_75t_R FILLER_0_114_919 ();
 FILLER_ASAP7_75t_R FILLER_0_114_927 ();
 FILLER_ASAP7_75t_R FILLER_0_114_950 ();
 FILLER_ASAP7_75t_R FILLER_0_114_973 ();
 FILLER_ASAP7_75t_R FILLER_0_114_978 ();
 DECAPx6_ASAP7_75t_R FILLER_0_114_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_997 ();
 DECAPx2_ASAP7_75t_R FILLER_0_114_1008 ();
 FILLER_ASAP7_75t_R FILLER_0_114_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_1016 ();
 FILLER_ASAP7_75t_R FILLER_0_114_1023 ();
 DECAPx2_ASAP7_75t_R FILLER_0_114_1037 ();
 FILLER_ASAP7_75t_R FILLER_0_114_1043 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_1048 ();
 DECAPx4_ASAP7_75t_R FILLER_0_114_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_1080 ();
 DECAPx4_ASAP7_75t_R FILLER_0_114_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_1097 ();
 FILLER_ASAP7_75t_R FILLER_0_114_1106 ();
 DECAPx1_ASAP7_75t_R FILLER_0_114_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_1122 ();
 DECAPx6_ASAP7_75t_R FILLER_0_114_1131 ();
 FILLER_ASAP7_75t_R FILLER_0_114_1150 ();
 DECAPx1_ASAP7_75t_R FILLER_0_114_1164 ();
 FILLER_ASAP7_75t_R FILLER_0_114_1178 ();
 FILLER_ASAP7_75t_R FILLER_0_114_1190 ();
 FILLER_ASAP7_75t_R FILLER_0_114_1199 ();
 FILLER_ASAP7_75t_R FILLER_0_114_1207 ();
 DECAPx2_ASAP7_75t_R FILLER_0_114_1215 ();
 FILLER_ASAP7_75t_R FILLER_0_114_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_1223 ();
 FILLER_ASAP7_75t_R FILLER_0_114_1234 ();
 FILLER_ASAP7_75t_R FILLER_0_114_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_0_114_1272 ();
 DECAPx1_ASAP7_75t_R FILLER_0_114_1286 ();
 FILLER_ASAP7_75t_R FILLER_0_114_1297 ();
 DECAPx2_ASAP7_75t_R FILLER_0_114_1305 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_1311 ();
 DECAPx4_ASAP7_75t_R FILLER_0_114_1318 ();
 FILLER_ASAP7_75t_R FILLER_0_114_1328 ();
 FILLER_ASAP7_75t_R FILLER_0_114_1336 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_1338 ();
 FILLER_ASAP7_75t_R FILLER_0_114_1342 ();
 FILLER_ASAP7_75t_R FILLER_0_114_1349 ();
 FILLER_ASAP7_75t_R FILLER_0_114_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_114_1380 ();
 DECAPx1_ASAP7_75t_R FILLER_0_115_2 ();
 FILLER_ASAP7_75t_R FILLER_0_115_11 ();
 DECAPx2_ASAP7_75t_R FILLER_0_115_18 ();
 DECAPx2_ASAP7_75t_R FILLER_0_115_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_36 ();
 DECAPx4_ASAP7_75t_R FILLER_0_115_43 ();
 FILLER_ASAP7_75t_R FILLER_0_115_53 ();
 FILLER_ASAP7_75t_R FILLER_0_115_60 ();
 FILLER_ASAP7_75t_R FILLER_0_115_67 ();
 DECAPx2_ASAP7_75t_R FILLER_0_115_75 ();
 FILLER_ASAP7_75t_R FILLER_0_115_81 ();
 FILLER_ASAP7_75t_R FILLER_0_115_90 ();
 FILLER_ASAP7_75t_R FILLER_0_115_98 ();
 FILLER_ASAP7_75t_R FILLER_0_115_108 ();
 FILLER_ASAP7_75t_R FILLER_0_115_120 ();
 FILLER_ASAP7_75t_R FILLER_0_115_132 ();
 DECAPx1_ASAP7_75t_R FILLER_0_115_148 ();
 FILLER_ASAP7_75t_R FILLER_0_115_158 ();
 FILLER_ASAP7_75t_R FILLER_0_115_166 ();
 FILLER_ASAP7_75t_R FILLER_0_115_174 ();
 FILLER_ASAP7_75t_R FILLER_0_115_181 ();
 FILLER_ASAP7_75t_R FILLER_0_115_188 ();
 DECAPx6_ASAP7_75t_R FILLER_0_115_196 ();
 FILLER_ASAP7_75t_R FILLER_0_115_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_212 ();
 FILLER_ASAP7_75t_R FILLER_0_115_219 ();
 DECAPx2_ASAP7_75t_R FILLER_0_115_227 ();
 FILLER_ASAP7_75t_R FILLER_0_115_233 ();
 FILLER_ASAP7_75t_R FILLER_0_115_241 ();
 FILLER_ASAP7_75t_R FILLER_0_115_254 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_266 ();
 DECAPx4_ASAP7_75t_R FILLER_0_115_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_319 ();
 DECAPx4_ASAP7_75t_R FILLER_0_115_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_333 ();
 FILLER_ASAP7_75t_R FILLER_0_115_355 ();
 DECAPx4_ASAP7_75t_R FILLER_0_115_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_388 ();
 DECAPx2_ASAP7_75t_R FILLER_0_115_397 ();
 FILLER_ASAP7_75t_R FILLER_0_115_415 ();
 DECAPx4_ASAP7_75t_R FILLER_0_115_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_439 ();
 DECAPx1_ASAP7_75t_R FILLER_0_115_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_450 ();
 FILLER_ASAP7_75t_R FILLER_0_115_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_463 ();
 FILLER_ASAP7_75t_R FILLER_0_115_470 ();
 DECAPx2_ASAP7_75t_R FILLER_0_115_477 ();
 FILLER_ASAP7_75t_R FILLER_0_115_483 ();
 FILLER_ASAP7_75t_R FILLER_0_115_505 ();
 FILLER_ASAP7_75t_R FILLER_0_115_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_519 ();
 FILLER_ASAP7_75t_R FILLER_0_115_529 ();
 DECAPx2_ASAP7_75t_R FILLER_0_115_536 ();
 FILLER_ASAP7_75t_R FILLER_0_115_548 ();
 DECAPx2_ASAP7_75t_R FILLER_0_115_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_561 ();
 DECAPx1_ASAP7_75t_R FILLER_0_115_574 ();
 FILLER_ASAP7_75t_R FILLER_0_115_584 ();
 FILLER_ASAP7_75t_R FILLER_0_115_593 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_595 ();
 FILLER_ASAP7_75t_R FILLER_0_115_602 ();
 DECAPx1_ASAP7_75t_R FILLER_0_115_615 ();
 DECAPx1_ASAP7_75t_R FILLER_0_115_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_633 ();
 FILLER_ASAP7_75t_R FILLER_0_115_639 ();
 FILLER_ASAP7_75t_R FILLER_0_115_651 ();
 DECAPx1_ASAP7_75t_R FILLER_0_115_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_667 ();
 FILLER_ASAP7_75t_R FILLER_0_115_678 ();
 FILLER_ASAP7_75t_R FILLER_0_115_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_704 ();
 FILLER_ASAP7_75t_R FILLER_0_115_715 ();
 FILLER_ASAP7_75t_R FILLER_0_115_735 ();
 FILLER_ASAP7_75t_R FILLER_0_115_759 ();
 FILLER_ASAP7_75t_R FILLER_0_115_767 ();
 FILLER_ASAP7_75t_R FILLER_0_115_774 ();
 FILLER_ASAP7_75t_R FILLER_0_115_782 ();
 FILLER_ASAP7_75t_R FILLER_0_115_789 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_796 ();
 DECAPx6_ASAP7_75t_R FILLER_0_115_818 ();
 FILLER_ASAP7_75t_R FILLER_0_115_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_834 ();
 DECAPx1_ASAP7_75t_R FILLER_0_115_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_851 ();
 DECAPx2_ASAP7_75t_R FILLER_0_115_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_868 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_874 ();
 DECAPx6_ASAP7_75t_R FILLER_0_115_896 ();
 DECAPx1_ASAP7_75t_R FILLER_0_115_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_914 ();
 FILLER_ASAP7_75t_R FILLER_0_115_923 ();
 DECAPx2_ASAP7_75t_R FILLER_0_115_927 ();
 FILLER_ASAP7_75t_R FILLER_0_115_941 ();
 DECAPx1_ASAP7_75t_R FILLER_0_115_946 ();
 DECAPx2_ASAP7_75t_R FILLER_0_115_957 ();
 FILLER_ASAP7_75t_R FILLER_0_115_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_965 ();
 FILLER_ASAP7_75t_R FILLER_0_115_972 ();
 DECAPx2_ASAP7_75t_R FILLER_0_115_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_991 ();
 DECAPx1_ASAP7_75t_R FILLER_0_115_1012 ();
 FILLER_ASAP7_75t_R FILLER_0_115_1021 ();
 DECAPx1_ASAP7_75t_R FILLER_0_115_1029 ();
 FILLER_ASAP7_75t_R FILLER_0_115_1041 ();
 FILLER_ASAP7_75t_R FILLER_0_115_1053 ();
 DECAPx4_ASAP7_75t_R FILLER_0_115_1060 ();
 FILLER_ASAP7_75t_R FILLER_0_115_1070 ();
 FILLER_ASAP7_75t_R FILLER_0_115_1082 ();
 FILLER_ASAP7_75t_R FILLER_0_115_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_1106 ();
 DECAPx2_ASAP7_75t_R FILLER_0_115_1128 ();
 FILLER_ASAP7_75t_R FILLER_0_115_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_1142 ();
 FILLER_ASAP7_75t_R FILLER_0_115_1155 ();
 FILLER_ASAP7_75t_R FILLER_0_115_1167 ();
 FILLER_ASAP7_75t_R FILLER_0_115_1179 ();
 DECAPx2_ASAP7_75t_R FILLER_0_115_1191 ();
 FILLER_ASAP7_75t_R FILLER_0_115_1197 ();
 DECAPx1_ASAP7_75t_R FILLER_0_115_1209 ();
 FILLER_ASAP7_75t_R FILLER_0_115_1219 ();
 FILLER_ASAP7_75t_R FILLER_0_115_1227 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_1229 ();
 DECAPx1_ASAP7_75t_R FILLER_0_115_1236 ();
 FILLER_ASAP7_75t_R FILLER_0_115_1246 ();
 DECAPx1_ASAP7_75t_R FILLER_0_115_1255 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_1259 ();
 FILLER_ASAP7_75t_R FILLER_0_115_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_0_115_1280 ();
 FILLER_ASAP7_75t_R FILLER_0_115_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_1288 ();
 FILLER_ASAP7_75t_R FILLER_0_115_1299 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_1301 ();
 DECAPx1_ASAP7_75t_R FILLER_0_115_1309 ();
 FILLER_ASAP7_75t_R FILLER_0_115_1323 ();
 FILLER_ASAP7_75t_R FILLER_0_115_1345 ();
 FILLER_ASAP7_75t_R FILLER_0_115_1368 ();
 DECAPx2_ASAP7_75t_R FILLER_0_115_1376 ();
 FILLER_ASAP7_75t_R FILLER_0_116_2 ();
 FILLER_ASAP7_75t_R FILLER_0_116_26 ();
 FILLER_ASAP7_75t_R FILLER_0_116_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_41 ();
 DECAPx2_ASAP7_75t_R FILLER_0_116_48 ();
 FILLER_ASAP7_75t_R FILLER_0_116_66 ();
 FILLER_ASAP7_75t_R FILLER_0_116_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_78 ();
 DECAPx1_ASAP7_75t_R FILLER_0_116_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_103 ();
 FILLER_ASAP7_75t_R FILLER_0_116_111 ();
 FILLER_ASAP7_75t_R FILLER_0_116_123 ();
 FILLER_ASAP7_75t_R FILLER_0_116_135 ();
 FILLER_ASAP7_75t_R FILLER_0_116_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_149 ();
 DECAPx1_ASAP7_75t_R FILLER_0_116_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_165 ();
 FILLER_ASAP7_75t_R FILLER_0_116_172 ();
 DECAPx1_ASAP7_75t_R FILLER_0_116_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_184 ();
 DECAPx1_ASAP7_75t_R FILLER_0_116_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_200 ();
 FILLER_ASAP7_75t_R FILLER_0_116_217 ();
 FILLER_ASAP7_75t_R FILLER_0_116_230 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_238 ();
 DECAPx4_ASAP7_75t_R FILLER_0_116_260 ();
 DECAPx4_ASAP7_75t_R FILLER_0_116_276 ();
 DECAPx6_ASAP7_75t_R FILLER_0_116_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_304 ();
 FILLER_ASAP7_75t_R FILLER_0_116_308 ();
 FILLER_ASAP7_75t_R FILLER_0_116_321 ();
 FILLER_ASAP7_75t_R FILLER_0_116_326 ();
 FILLER_ASAP7_75t_R FILLER_0_116_331 ();
 DECAPx1_ASAP7_75t_R FILLER_0_116_339 ();
 DECAPx1_ASAP7_75t_R FILLER_0_116_355 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_362 ();
 FILLER_ASAP7_75t_R FILLER_0_116_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_386 ();
 DECAPx4_ASAP7_75t_R FILLER_0_116_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_403 ();
 DECAPx2_ASAP7_75t_R FILLER_0_116_415 ();
 FILLER_ASAP7_75t_R FILLER_0_116_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_423 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_434 ();
 DECAPx2_ASAP7_75t_R FILLER_0_116_456 ();
 DECAPx1_ASAP7_75t_R FILLER_0_116_464 ();
 DECAPx4_ASAP7_75t_R FILLER_0_116_474 ();
 DECAPx4_ASAP7_75t_R FILLER_0_116_490 ();
 FILLER_ASAP7_75t_R FILLER_0_116_506 ();
 DECAPx1_ASAP7_75t_R FILLER_0_116_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_518 ();
 FILLER_ASAP7_75t_R FILLER_0_116_525 ();
 FILLER_ASAP7_75t_R FILLER_0_116_534 ();
 FILLER_ASAP7_75t_R FILLER_0_116_542 ();
 FILLER_ASAP7_75t_R FILLER_0_116_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_552 ();
 FILLER_ASAP7_75t_R FILLER_0_116_559 ();
 FILLER_ASAP7_75t_R FILLER_0_116_573 ();
 FILLER_ASAP7_75t_R FILLER_0_116_581 ();
 FILLER_ASAP7_75t_R FILLER_0_116_589 ();
 DECAPx1_ASAP7_75t_R FILLER_0_116_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_600 ();
 FILLER_ASAP7_75t_R FILLER_0_116_607 ();
 DECAPx1_ASAP7_75t_R FILLER_0_116_612 ();
 FILLER_ASAP7_75t_R FILLER_0_116_621 ();
 DECAPx2_ASAP7_75t_R FILLER_0_116_633 ();
 FILLER_ASAP7_75t_R FILLER_0_116_644 ();
 FILLER_ASAP7_75t_R FILLER_0_116_651 ();
 DECAPx2_ASAP7_75t_R FILLER_0_116_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_669 ();
 FILLER_ASAP7_75t_R FILLER_0_116_676 ();
 DECAPx4_ASAP7_75t_R FILLER_0_116_682 ();
 FILLER_ASAP7_75t_R FILLER_0_116_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_694 ();
 FILLER_ASAP7_75t_R FILLER_0_116_698 ();
 FILLER_ASAP7_75t_R FILLER_0_116_704 ();
 FILLER_ASAP7_75t_R FILLER_0_116_728 ();
 FILLER_ASAP7_75t_R FILLER_0_116_752 ();
 FILLER_ASAP7_75t_R FILLER_0_116_764 ();
 FILLER_ASAP7_75t_R FILLER_0_116_776 ();
 DECAPx6_ASAP7_75t_R FILLER_0_116_783 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_809 ();
 DECAPx2_ASAP7_75t_R FILLER_0_116_831 ();
 FILLER_ASAP7_75t_R FILLER_0_116_837 ();
 DECAPx6_ASAP7_75t_R FILLER_0_116_857 ();
 FILLER_ASAP7_75t_R FILLER_0_116_892 ();
 FILLER_ASAP7_75t_R FILLER_0_116_900 ();
 DECAPx2_ASAP7_75t_R FILLER_0_116_908 ();
 FILLER_ASAP7_75t_R FILLER_0_116_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_916 ();
 DECAPx1_ASAP7_75t_R FILLER_0_116_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_924 ();
 DECAPx2_ASAP7_75t_R FILLER_0_116_931 ();
 FILLER_ASAP7_75t_R FILLER_0_116_945 ();
 DECAPx1_ASAP7_75t_R FILLER_0_116_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_954 ();
 DECAPx1_ASAP7_75t_R FILLER_0_116_966 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_970 ();
 FILLER_ASAP7_75t_R FILLER_0_116_979 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_981 ();
 DECAPx1_ASAP7_75t_R FILLER_0_116_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_989 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_1002 ();
 DECAPx4_ASAP7_75t_R FILLER_0_116_1030 ();
 FILLER_ASAP7_75t_R FILLER_0_116_1060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_1072 ();
 DECAPx1_ASAP7_75t_R FILLER_0_116_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_1104 ();
 DECAPx4_ASAP7_75t_R FILLER_0_116_1126 ();
 FILLER_ASAP7_75t_R FILLER_0_116_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_1138 ();
 FILLER_ASAP7_75t_R FILLER_0_116_1144 ();
 FILLER_ASAP7_75t_R FILLER_0_116_1156 ();
 FILLER_ASAP7_75t_R FILLER_0_116_1168 ();
 FILLER_ASAP7_75t_R FILLER_0_116_1180 ();
 FILLER_ASAP7_75t_R FILLER_0_116_1192 ();
 DECAPx1_ASAP7_75t_R FILLER_0_116_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_1203 ();
 DECAPx6_ASAP7_75t_R FILLER_0_116_1209 ();
 DECAPx1_ASAP7_75t_R FILLER_0_116_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_1233 ();
 DECAPx2_ASAP7_75t_R FILLER_0_116_1269 ();
 DECAPx1_ASAP7_75t_R FILLER_0_116_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_1286 ();
 FILLER_ASAP7_75t_R FILLER_0_116_1292 ();
 FILLER_ASAP7_75t_R FILLER_0_116_1300 ();
 FILLER_ASAP7_75t_R FILLER_0_116_1307 ();
 DECAPx1_ASAP7_75t_R FILLER_0_116_1314 ();
 FILLER_ASAP7_75t_R FILLER_0_116_1324 ();
 FILLER_ASAP7_75t_R FILLER_0_116_1329 ();
 FILLER_ASAP7_75t_R FILLER_0_116_1361 ();
 FILLER_ASAP7_75t_R FILLER_0_116_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_116_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_117_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_117_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_13 ();
 FILLER_ASAP7_75t_R FILLER_0_117_20 ();
 FILLER_ASAP7_75t_R FILLER_0_117_28 ();
 DECAPx2_ASAP7_75t_R FILLER_0_117_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_42 ();
 FILLER_ASAP7_75t_R FILLER_0_117_49 ();
 DECAPx2_ASAP7_75t_R FILLER_0_117_57 ();
 FILLER_ASAP7_75t_R FILLER_0_117_63 ();
 FILLER_ASAP7_75t_R FILLER_0_117_70 ();
 FILLER_ASAP7_75t_R FILLER_0_117_77 ();
 FILLER_ASAP7_75t_R FILLER_0_117_85 ();
 FILLER_ASAP7_75t_R FILLER_0_117_93 ();
 FILLER_ASAP7_75t_R FILLER_0_117_101 ();
 DECAPx2_ASAP7_75t_R FILLER_0_117_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_129 ();
 FILLER_ASAP7_75t_R FILLER_0_117_148 ();
 FILLER_ASAP7_75t_R FILLER_0_117_160 ();
 DECAPx2_ASAP7_75t_R FILLER_0_117_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_175 ();
 DECAPx2_ASAP7_75t_R FILLER_0_117_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_188 ();
 DECAPx4_ASAP7_75t_R FILLER_0_117_195 ();
 FILLER_ASAP7_75t_R FILLER_0_117_205 ();
 DECAPx1_ASAP7_75t_R FILLER_0_117_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_217 ();
 DECAPx1_ASAP7_75t_R FILLER_0_117_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_228 ();
 DECAPx1_ASAP7_75t_R FILLER_0_117_235 ();
 DECAPx2_ASAP7_75t_R FILLER_0_117_245 ();
 FILLER_ASAP7_75t_R FILLER_0_117_251 ();
 FILLER_ASAP7_75t_R FILLER_0_117_259 ();
 FILLER_ASAP7_75t_R FILLER_0_117_264 ();
 FILLER_ASAP7_75t_R FILLER_0_117_272 ();
 DECAPx1_ASAP7_75t_R FILLER_0_117_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_286 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_292 ();
 DECAPx2_ASAP7_75t_R FILLER_0_117_314 ();
 DECAPx1_ASAP7_75t_R FILLER_0_117_328 ();
 FILLER_ASAP7_75t_R FILLER_0_117_344 ();
 DECAPx4_ASAP7_75t_R FILLER_0_117_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_368 ();
 DECAPx2_ASAP7_75t_R FILLER_0_117_380 ();
 FILLER_ASAP7_75t_R FILLER_0_117_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_388 ();
 DECAPx4_ASAP7_75t_R FILLER_0_117_397 ();
 DECAPx6_ASAP7_75t_R FILLER_0_117_419 ();
 FILLER_ASAP7_75t_R FILLER_0_117_433 ();
 FILLER_ASAP7_75t_R FILLER_0_117_438 ();
 FILLER_ASAP7_75t_R FILLER_0_117_446 ();
 DECAPx6_ASAP7_75t_R FILLER_0_117_451 ();
 DECAPx2_ASAP7_75t_R FILLER_0_117_471 ();
 FILLER_ASAP7_75t_R FILLER_0_117_477 ();
 FILLER_ASAP7_75t_R FILLER_0_117_485 ();
 FILLER_ASAP7_75t_R FILLER_0_117_493 ();
 FILLER_ASAP7_75t_R FILLER_0_117_498 ();
 FILLER_ASAP7_75t_R FILLER_0_117_505 ();
 FILLER_ASAP7_75t_R FILLER_0_117_513 ();
 DECAPx1_ASAP7_75t_R FILLER_0_117_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_530 ();
 DECAPx2_ASAP7_75t_R FILLER_0_117_538 ();
 DECAPx4_ASAP7_75t_R FILLER_0_117_550 ();
 FILLER_ASAP7_75t_R FILLER_0_117_563 ();
 DECAPx6_ASAP7_75t_R FILLER_0_117_572 ();
 DECAPx2_ASAP7_75t_R FILLER_0_117_586 ();
 FILLER_ASAP7_75t_R FILLER_0_117_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_117_606 ();
 FILLER_ASAP7_75t_R FILLER_0_117_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_614 ();
 DECAPx2_ASAP7_75t_R FILLER_0_117_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_627 ();
 DECAPx2_ASAP7_75t_R FILLER_0_117_638 ();
 FILLER_ASAP7_75t_R FILLER_0_117_644 ();
 FILLER_ASAP7_75t_R FILLER_0_117_656 ();
 DECAPx1_ASAP7_75t_R FILLER_0_117_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_667 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_678 ();
 DECAPx4_ASAP7_75t_R FILLER_0_117_700 ();
 FILLER_ASAP7_75t_R FILLER_0_117_710 ();
 FILLER_ASAP7_75t_R FILLER_0_117_733 ();
 FILLER_ASAP7_75t_R FILLER_0_117_738 ();
 DECAPx6_ASAP7_75t_R FILLER_0_117_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_757 ();
 FILLER_ASAP7_75t_R FILLER_0_117_768 ();
 FILLER_ASAP7_75t_R FILLER_0_117_776 ();
 FILLER_ASAP7_75t_R FILLER_0_117_784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_792 ();
 FILLER_ASAP7_75t_R FILLER_0_117_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_816 ();
 FILLER_ASAP7_75t_R FILLER_0_117_829 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_837 ();
 DECAPx2_ASAP7_75t_R FILLER_0_117_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_865 ();
 FILLER_ASAP7_75t_R FILLER_0_117_872 ();
 DECAPx2_ASAP7_75t_R FILLER_0_117_880 ();
 FILLER_ASAP7_75t_R FILLER_0_117_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_888 ();
 FILLER_ASAP7_75t_R FILLER_0_117_892 ();
 DECAPx4_ASAP7_75t_R FILLER_0_117_915 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_927 ();
 DECAPx2_ASAP7_75t_R FILLER_0_117_949 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_961 ();
 DECAPx1_ASAP7_75t_R FILLER_0_117_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_987 ();
 DECAPx2_ASAP7_75t_R FILLER_0_117_1009 ();
 DECAPx6_ASAP7_75t_R FILLER_0_117_1027 ();
 DECAPx1_ASAP7_75t_R FILLER_0_117_1041 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_0_117_1077 ();
 FILLER_ASAP7_75t_R FILLER_0_117_1083 ();
 FILLER_ASAP7_75t_R FILLER_0_117_1097 ();
 FILLER_ASAP7_75t_R FILLER_0_117_1105 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_1107 ();
 FILLER_ASAP7_75t_R FILLER_0_117_1114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_1124 ();
 FILLER_ASAP7_75t_R FILLER_0_117_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_1148 ();
 FILLER_ASAP7_75t_R FILLER_0_117_1155 ();
 FILLER_ASAP7_75t_R FILLER_0_117_1163 ();
 FILLER_ASAP7_75t_R FILLER_0_117_1170 ();
 FILLER_ASAP7_75t_R FILLER_0_117_1182 ();
 FILLER_ASAP7_75t_R FILLER_0_117_1192 ();
 FILLER_ASAP7_75t_R FILLER_0_117_1202 ();
 DECAPx4_ASAP7_75t_R FILLER_0_117_1207 ();
 FILLER_ASAP7_75t_R FILLER_0_117_1227 ();
 FILLER_ASAP7_75t_R FILLER_0_117_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_1246 ();
 FILLER_ASAP7_75t_R FILLER_0_117_1268 ();
 FILLER_ASAP7_75t_R FILLER_0_117_1276 ();
 DECAPx2_ASAP7_75t_R FILLER_0_117_1284 ();
 DECAPx2_ASAP7_75t_R FILLER_0_117_1302 ();
 FILLER_ASAP7_75t_R FILLER_0_117_1308 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_1310 ();
 FILLER_ASAP7_75t_R FILLER_0_117_1316 ();
 FILLER_ASAP7_75t_R FILLER_0_117_1325 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_1327 ();
 FILLER_ASAP7_75t_R FILLER_0_117_1334 ();
 FILLER_ASAP7_75t_R FILLER_0_117_1339 ();
 FILLER_ASAP7_75t_R FILLER_0_117_1363 ();
 FILLER_ASAP7_75t_R FILLER_0_117_1371 ();
 DECAPx1_ASAP7_75t_R FILLER_0_117_1378 ();
 FILLER_ASAP7_75t_R FILLER_0_118_2 ();
 FILLER_ASAP7_75t_R FILLER_0_118_9 ();
 FILLER_ASAP7_75t_R FILLER_0_118_16 ();
 FILLER_ASAP7_75t_R FILLER_0_118_23 ();
 FILLER_ASAP7_75t_R FILLER_0_118_31 ();
 FILLER_ASAP7_75t_R FILLER_0_118_36 ();
 DECAPx2_ASAP7_75t_R FILLER_0_118_44 ();
 FILLER_ASAP7_75t_R FILLER_0_118_50 ();
 FILLER_ASAP7_75t_R FILLER_0_118_58 ();
 FILLER_ASAP7_75t_R FILLER_0_118_66 ();
 DECAPx1_ASAP7_75t_R FILLER_0_118_79 ();
 FILLER_ASAP7_75t_R FILLER_0_118_94 ();
 FILLER_ASAP7_75t_R FILLER_0_118_101 ();
 FILLER_ASAP7_75t_R FILLER_0_118_109 ();
 FILLER_ASAP7_75t_R FILLER_0_118_117 ();
 FILLER_ASAP7_75t_R FILLER_0_118_129 ();
 FILLER_ASAP7_75t_R FILLER_0_118_149 ();
 DECAPx2_ASAP7_75t_R FILLER_0_118_161 ();
 FILLER_ASAP7_75t_R FILLER_0_118_173 ();
 FILLER_ASAP7_75t_R FILLER_0_118_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_183 ();
 DECAPx2_ASAP7_75t_R FILLER_0_118_190 ();
 FILLER_ASAP7_75t_R FILLER_0_118_196 ();
 FILLER_ASAP7_75t_R FILLER_0_118_204 ();
 DECAPx2_ASAP7_75t_R FILLER_0_118_212 ();
 FILLER_ASAP7_75t_R FILLER_0_118_218 ();
 DECAPx6_ASAP7_75t_R FILLER_0_118_236 ();
 FILLER_ASAP7_75t_R FILLER_0_118_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_252 ();
 FILLER_ASAP7_75t_R FILLER_0_118_263 ();
 FILLER_ASAP7_75t_R FILLER_0_118_271 ();
 DECAPx2_ASAP7_75t_R FILLER_0_118_281 ();
 FILLER_ASAP7_75t_R FILLER_0_118_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_289 ();
 DECAPx1_ASAP7_75t_R FILLER_0_118_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_306 ();
 FILLER_ASAP7_75t_R FILLER_0_118_313 ();
 DECAPx2_ASAP7_75t_R FILLER_0_118_325 ();
 FILLER_ASAP7_75t_R FILLER_0_118_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_333 ();
 DECAPx2_ASAP7_75t_R FILLER_0_118_346 ();
 DECAPx6_ASAP7_75t_R FILLER_0_118_358 ();
 DECAPx1_ASAP7_75t_R FILLER_0_118_372 ();
 DECAPx6_ASAP7_75t_R FILLER_0_118_388 ();
 FILLER_ASAP7_75t_R FILLER_0_118_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_404 ();
 DECAPx2_ASAP7_75t_R FILLER_0_118_417 ();
 FILLER_ASAP7_75t_R FILLER_0_118_423 ();
 FILLER_ASAP7_75t_R FILLER_0_118_431 ();
 FILLER_ASAP7_75t_R FILLER_0_118_439 ();
 DECAPx6_ASAP7_75t_R FILLER_0_118_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_486 ();
 DECAPx4_ASAP7_75t_R FILLER_0_118_507 ();
 FILLER_ASAP7_75t_R FILLER_0_118_524 ();
 FILLER_ASAP7_75t_R FILLER_0_118_532 ();
 FILLER_ASAP7_75t_R FILLER_0_118_544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_551 ();
 DECAPx4_ASAP7_75t_R FILLER_0_118_573 ();
 FILLER_ASAP7_75t_R FILLER_0_118_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_585 ();
 DECAPx2_ASAP7_75t_R FILLER_0_118_598 ();
 FILLER_ASAP7_75t_R FILLER_0_118_604 ();
 FILLER_ASAP7_75t_R FILLER_0_118_616 ();
 DECAPx2_ASAP7_75t_R FILLER_0_118_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_630 ();
 FILLER_ASAP7_75t_R FILLER_0_118_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_641 ();
 DECAPx1_ASAP7_75t_R FILLER_0_118_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_677 ();
 FILLER_ASAP7_75t_R FILLER_0_118_705 ();
 FILLER_ASAP7_75t_R FILLER_0_118_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_715 ();
 DECAPx1_ASAP7_75t_R FILLER_0_118_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_726 ();
 FILLER_ASAP7_75t_R FILLER_0_118_730 ();
 FILLER_ASAP7_75t_R FILLER_0_118_742 ();
 DECAPx1_ASAP7_75t_R FILLER_0_118_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_751 ();
 DECAPx2_ASAP7_75t_R FILLER_0_118_758 ();
 FILLER_ASAP7_75t_R FILLER_0_118_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_766 ();
 DECAPx2_ASAP7_75t_R FILLER_0_118_773 ();
 DECAPx2_ASAP7_75t_R FILLER_0_118_789 ();
 DECAPx6_ASAP7_75t_R FILLER_0_118_802 ();
 FILLER_ASAP7_75t_R FILLER_0_118_816 ();
 DECAPx4_ASAP7_75t_R FILLER_0_118_830 ();
 FILLER_ASAP7_75t_R FILLER_0_118_840 ();
 FILLER_ASAP7_75t_R FILLER_0_118_848 ();
 DECAPx1_ASAP7_75t_R FILLER_0_118_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_860 ();
 DECAPx1_ASAP7_75t_R FILLER_0_118_872 ();
 DECAPx2_ASAP7_75t_R FILLER_0_118_886 ();
 FILLER_ASAP7_75t_R FILLER_0_118_892 ();
 FILLER_ASAP7_75t_R FILLER_0_118_897 ();
 FILLER_ASAP7_75t_R FILLER_0_118_904 ();
 DECAPx4_ASAP7_75t_R FILLER_0_118_909 ();
 FILLER_ASAP7_75t_R FILLER_0_118_919 ();
 FILLER_ASAP7_75t_R FILLER_0_118_931 ();
 DECAPx2_ASAP7_75t_R FILLER_0_118_954 ();
 FILLER_ASAP7_75t_R FILLER_0_118_960 ();
 FILLER_ASAP7_75t_R FILLER_0_118_982 ();
 DECAPx4_ASAP7_75t_R FILLER_0_118_988 ();
 FILLER_ASAP7_75t_R FILLER_0_118_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_1000 ();
 FILLER_ASAP7_75t_R FILLER_0_118_1004 ();
 FILLER_ASAP7_75t_R FILLER_0_118_1016 ();
 FILLER_ASAP7_75t_R FILLER_0_118_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_1032 ();
 DECAPx1_ASAP7_75t_R FILLER_0_118_1045 ();
 DECAPx1_ASAP7_75t_R FILLER_0_118_1059 ();
 DECAPx1_ASAP7_75t_R FILLER_0_118_1084 ();
 FILLER_ASAP7_75t_R FILLER_0_118_1100 ();
 FILLER_ASAP7_75t_R FILLER_0_118_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_1144 ();
 FILLER_ASAP7_75t_R FILLER_0_118_1155 ();
 DECAPx2_ASAP7_75t_R FILLER_0_118_1165 ();
 FILLER_ASAP7_75t_R FILLER_0_118_1181 ();
 FILLER_ASAP7_75t_R FILLER_0_118_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_1193 ();
 DECAPx2_ASAP7_75t_R FILLER_0_118_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_1211 ();
 FILLER_ASAP7_75t_R FILLER_0_118_1224 ();
 DECAPx4_ASAP7_75t_R FILLER_0_118_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_0_118_1272 ();
 FILLER_ASAP7_75t_R FILLER_0_118_1292 ();
 DECAPx6_ASAP7_75t_R FILLER_0_118_1299 ();
 FILLER_ASAP7_75t_R FILLER_0_118_1318 ();
 FILLER_ASAP7_75t_R FILLER_0_118_1332 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_1334 ();
 FILLER_ASAP7_75t_R FILLER_0_118_1340 ();
 DECAPx1_ASAP7_75t_R FILLER_0_118_1364 ();
 FILLER_ASAP7_75t_R FILLER_0_118_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_118_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_119_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_119_9 ();
 FILLER_ASAP7_75t_R FILLER_0_119_20 ();
 DECAPx2_ASAP7_75t_R FILLER_0_119_28 ();
 FILLER_ASAP7_75t_R FILLER_0_119_40 ();
 DECAPx2_ASAP7_75t_R FILLER_0_119_48 ();
 FILLER_ASAP7_75t_R FILLER_0_119_54 ();
 DECAPx4_ASAP7_75t_R FILLER_0_119_62 ();
 FILLER_ASAP7_75t_R FILLER_0_119_78 ();
 FILLER_ASAP7_75t_R FILLER_0_119_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_88 ();
 FILLER_ASAP7_75t_R FILLER_0_119_94 ();
 DECAPx2_ASAP7_75t_R FILLER_0_119_112 ();
 FILLER_ASAP7_75t_R FILLER_0_119_118 ();
 FILLER_ASAP7_75t_R FILLER_0_119_130 ();
 FILLER_ASAP7_75t_R FILLER_0_119_150 ();
 FILLER_ASAP7_75t_R FILLER_0_119_170 ();
 FILLER_ASAP7_75t_R FILLER_0_119_177 ();
 DECAPx1_ASAP7_75t_R FILLER_0_119_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_189 ();
 FILLER_ASAP7_75t_R FILLER_0_119_195 ();
 FILLER_ASAP7_75t_R FILLER_0_119_203 ();
 FILLER_ASAP7_75t_R FILLER_0_119_216 ();
 FILLER_ASAP7_75t_R FILLER_0_119_234 ();
 FILLER_ASAP7_75t_R FILLER_0_119_242 ();
 DECAPx2_ASAP7_75t_R FILLER_0_119_250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_277 ();
 DECAPx2_ASAP7_75t_R FILLER_0_119_299 ();
 FILLER_ASAP7_75t_R FILLER_0_119_305 ();
 DECAPx1_ASAP7_75t_R FILLER_0_119_328 ();
 DECAPx2_ASAP7_75t_R FILLER_0_119_344 ();
 DECAPx4_ASAP7_75t_R FILLER_0_119_371 ();
 FILLER_ASAP7_75t_R FILLER_0_119_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_383 ();
 DECAPx4_ASAP7_75t_R FILLER_0_119_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_402 ();
 DECAPx4_ASAP7_75t_R FILLER_0_119_415 ();
 FILLER_ASAP7_75t_R FILLER_0_119_428 ();
 DECAPx1_ASAP7_75t_R FILLER_0_119_436 ();
 FILLER_ASAP7_75t_R FILLER_0_119_451 ();
 DECAPx6_ASAP7_75t_R FILLER_0_119_459 ();
 FILLER_ASAP7_75t_R FILLER_0_119_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_475 ();
 FILLER_ASAP7_75t_R FILLER_0_119_482 ();
 DECAPx4_ASAP7_75t_R FILLER_0_119_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_500 ();
 FILLER_ASAP7_75t_R FILLER_0_119_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_508 ();
 FILLER_ASAP7_75t_R FILLER_0_119_515 ();
 FILLER_ASAP7_75t_R FILLER_0_119_523 ();
 FILLER_ASAP7_75t_R FILLER_0_119_531 ();
 DECAPx1_ASAP7_75t_R FILLER_0_119_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_547 ();
 DECAPx6_ASAP7_75t_R FILLER_0_119_554 ();
 DECAPx2_ASAP7_75t_R FILLER_0_119_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_574 ();
 FILLER_ASAP7_75t_R FILLER_0_119_582 ();
 FILLER_ASAP7_75t_R FILLER_0_119_590 ();
 DECAPx6_ASAP7_75t_R FILLER_0_119_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_614 ();
 FILLER_ASAP7_75t_R FILLER_0_119_621 ();
 FILLER_ASAP7_75t_R FILLER_0_119_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_631 ();
 FILLER_ASAP7_75t_R FILLER_0_119_638 ();
 FILLER_ASAP7_75t_R FILLER_0_119_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_650 ();
 FILLER_ASAP7_75t_R FILLER_0_119_657 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_708 ();
 FILLER_ASAP7_75t_R FILLER_0_119_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_717 ();
 FILLER_ASAP7_75t_R FILLER_0_119_724 ();
 FILLER_ASAP7_75t_R FILLER_0_119_729 ();
 FILLER_ASAP7_75t_R FILLER_0_119_736 ();
 DECAPx1_ASAP7_75t_R FILLER_0_119_746 ();
 DECAPx1_ASAP7_75t_R FILLER_0_119_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_760 ();
 FILLER_ASAP7_75t_R FILLER_0_119_764 ();
 FILLER_ASAP7_75t_R FILLER_0_119_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_786 ();
 DECAPx2_ASAP7_75t_R FILLER_0_119_813 ();
 FILLER_ASAP7_75t_R FILLER_0_119_819 ();
 FILLER_ASAP7_75t_R FILLER_0_119_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_829 ();
 FILLER_ASAP7_75t_R FILLER_0_119_836 ();
 DECAPx1_ASAP7_75t_R FILLER_0_119_844 ();
 FILLER_ASAP7_75t_R FILLER_0_119_854 ();
 FILLER_ASAP7_75t_R FILLER_0_119_862 ();
 FILLER_ASAP7_75t_R FILLER_0_119_870 ();
 DECAPx4_ASAP7_75t_R FILLER_0_119_878 ();
 FILLER_ASAP7_75t_R FILLER_0_119_888 ();
 DECAPx6_ASAP7_75t_R FILLER_0_119_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_924 ();
 DECAPx2_ASAP7_75t_R FILLER_0_119_927 ();
 FILLER_ASAP7_75t_R FILLER_0_119_933 ();
 DECAPx4_ASAP7_75t_R FILLER_0_119_938 ();
 FILLER_ASAP7_75t_R FILLER_0_119_958 ();
 DECAPx1_ASAP7_75t_R FILLER_0_119_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_972 ();
 FILLER_ASAP7_75t_R FILLER_0_119_981 ();
 DECAPx6_ASAP7_75t_R FILLER_0_119_991 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1005 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1018 ();
 DECAPx1_ASAP7_75t_R FILLER_0_119_1027 ();
 DECAPx1_ASAP7_75t_R FILLER_0_119_1042 ();
 DECAPx1_ASAP7_75t_R FILLER_0_119_1054 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1064 ();
 DECAPx6_ASAP7_75t_R FILLER_0_119_1069 ();
 DECAPx1_ASAP7_75t_R FILLER_0_119_1083 ();
 DECAPx2_ASAP7_75t_R FILLER_0_119_1099 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1105 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1111 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1119 ();
 DECAPx1_ASAP7_75t_R FILLER_0_119_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_1137 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1148 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1160 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1170 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_1180 ();
 DECAPx1_ASAP7_75t_R FILLER_0_119_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_1195 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1204 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1212 ();
 DECAPx2_ASAP7_75t_R FILLER_0_119_1220 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1226 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1235 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1243 ();
 DECAPx4_ASAP7_75t_R FILLER_0_119_1251 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1261 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1271 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1284 ();
 DECAPx2_ASAP7_75t_R FILLER_0_119_1292 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_1298 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1309 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1319 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1327 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1335 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1343 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1350 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1374 ();
 FILLER_ASAP7_75t_R FILLER_0_119_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_120_2 ();
 FILLER_ASAP7_75t_R FILLER_0_120_9 ();
 FILLER_ASAP7_75t_R FILLER_0_120_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_18 ();
 FILLER_ASAP7_75t_R FILLER_0_120_24 ();
 FILLER_ASAP7_75t_R FILLER_0_120_29 ();
 FILLER_ASAP7_75t_R FILLER_0_120_37 ();
 FILLER_ASAP7_75t_R FILLER_0_120_45 ();
 DECAPx6_ASAP7_75t_R FILLER_0_120_50 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_70 ();
 FILLER_ASAP7_75t_R FILLER_0_120_81 ();
 FILLER_ASAP7_75t_R FILLER_0_120_89 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_97 ();
 FILLER_ASAP7_75t_R FILLER_0_120_103 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_111 ();
 FILLER_ASAP7_75t_R FILLER_0_120_117 ();
 FILLER_ASAP7_75t_R FILLER_0_120_124 ();
 FILLER_ASAP7_75t_R FILLER_0_120_136 ();
 FILLER_ASAP7_75t_R FILLER_0_120_148 ();
 FILLER_ASAP7_75t_R FILLER_0_120_160 ();
 DECAPx1_ASAP7_75t_R FILLER_0_120_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_172 ();
 FILLER_ASAP7_75t_R FILLER_0_120_179 ();
 FILLER_ASAP7_75t_R FILLER_0_120_187 ();
 FILLER_ASAP7_75t_R FILLER_0_120_195 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_203 ();
 FILLER_ASAP7_75t_R FILLER_0_120_214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_226 ();
 FILLER_ASAP7_75t_R FILLER_0_120_232 ();
 FILLER_ASAP7_75t_R FILLER_0_120_239 ();
 FILLER_ASAP7_75t_R FILLER_0_120_247 ();
 DECAPx6_ASAP7_75t_R FILLER_0_120_254 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_274 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_278 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_300 ();
 FILLER_ASAP7_75t_R FILLER_0_120_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_308 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_312 ();
 FILLER_ASAP7_75t_R FILLER_0_120_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_336 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_343 ();
 FILLER_ASAP7_75t_R FILLER_0_120_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_351 ();
 FILLER_ASAP7_75t_R FILLER_0_120_355 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_360 ();
 FILLER_ASAP7_75t_R FILLER_0_120_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_368 ();
 DECAPx1_ASAP7_75t_R FILLER_0_120_375 ();
 FILLER_ASAP7_75t_R FILLER_0_120_382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_405 ();
 DECAPx1_ASAP7_75t_R FILLER_0_120_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_431 ();
 FILLER_ASAP7_75t_R FILLER_0_120_438 ();
 DECAPx1_ASAP7_75t_R FILLER_0_120_450 ();
 FILLER_ASAP7_75t_R FILLER_0_120_460 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_470 ();
 FILLER_ASAP7_75t_R FILLER_0_120_477 ();
 DECAPx4_ASAP7_75t_R FILLER_0_120_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_495 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_501 ();
 FILLER_ASAP7_75t_R FILLER_0_120_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_509 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_531 ();
 DECAPx1_ASAP7_75t_R FILLER_0_120_538 ();
 FILLER_ASAP7_75t_R FILLER_0_120_548 ();
 FILLER_ASAP7_75t_R FILLER_0_120_556 ();
 DECAPx4_ASAP7_75t_R FILLER_0_120_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_574 ();
 FILLER_ASAP7_75t_R FILLER_0_120_581 ();
 DECAPx1_ASAP7_75t_R FILLER_0_120_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_593 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_600 ();
 FILLER_ASAP7_75t_R FILLER_0_120_606 ();
 DECAPx1_ASAP7_75t_R FILLER_0_120_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_623 ();
 FILLER_ASAP7_75t_R FILLER_0_120_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_632 ();
 FILLER_ASAP7_75t_R FILLER_0_120_636 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_644 ();
 FILLER_ASAP7_75t_R FILLER_0_120_650 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_662 ();
 DECAPx1_ASAP7_75t_R FILLER_0_120_684 ();
 DECAPx4_ASAP7_75t_R FILLER_0_120_698 ();
 FILLER_ASAP7_75t_R FILLER_0_120_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_710 ();
 FILLER_ASAP7_75t_R FILLER_0_120_717 ();
 DECAPx1_ASAP7_75t_R FILLER_0_120_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_731 ();
 FILLER_ASAP7_75t_R FILLER_0_120_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_740 ();
 FILLER_ASAP7_75t_R FILLER_0_120_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_753 ();
 FILLER_ASAP7_75t_R FILLER_0_120_760 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_769 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_781 ();
 DECAPx1_ASAP7_75t_R FILLER_0_120_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_807 ();
 DECAPx1_ASAP7_75t_R FILLER_0_120_813 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_833 ();
 FILLER_ASAP7_75t_R FILLER_0_120_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_841 ();
 DECAPx4_ASAP7_75t_R FILLER_0_120_848 ();
 FILLER_ASAP7_75t_R FILLER_0_120_858 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_866 ();
 FILLER_ASAP7_75t_R FILLER_0_120_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_874 ();
 FILLER_ASAP7_75t_R FILLER_0_120_881 ();
 FILLER_ASAP7_75t_R FILLER_0_120_889 ();
 FILLER_ASAP7_75t_R FILLER_0_120_897 ();
 FILLER_ASAP7_75t_R FILLER_0_120_905 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_917 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_945 ();
 FILLER_ASAP7_75t_R FILLER_0_120_967 ();
 FILLER_ASAP7_75t_R FILLER_0_120_972 ();
 FILLER_ASAP7_75t_R FILLER_0_120_984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_990 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_1012 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_1030 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1052 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_1070 ();
 DECAPx6_ASAP7_75t_R FILLER_0_120_1092 ();
 DECAPx1_ASAP7_75t_R FILLER_0_120_1106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_1116 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_1138 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1144 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1151 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1165 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_1179 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1194 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1204 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_1218 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1226 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_1234 ();
 DECAPx4_ASAP7_75t_R FILLER_0_120_1250 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1260 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1268 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1275 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1288 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1296 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1304 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1309 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1317 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1331 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1338 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1345 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1352 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1359 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_1361 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1367 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1374 ();
 FILLER_ASAP7_75t_R FILLER_0_120_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_121_2 ();
 FILLER_ASAP7_75t_R FILLER_0_121_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_28 ();
 DECAPx1_ASAP7_75t_R FILLER_0_121_32 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_42 ();
 DECAPx6_ASAP7_75t_R FILLER_0_121_64 ();
 DECAPx1_ASAP7_75t_R FILLER_0_121_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_82 ();
 FILLER_ASAP7_75t_R FILLER_0_121_89 ();
 DECAPx2_ASAP7_75t_R FILLER_0_121_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_103 ();
 FILLER_ASAP7_75t_R FILLER_0_121_110 ();
 DECAPx2_ASAP7_75t_R FILLER_0_121_119 ();
 FILLER_ASAP7_75t_R FILLER_0_121_135 ();
 FILLER_ASAP7_75t_R FILLER_0_121_141 ();
 FILLER_ASAP7_75t_R FILLER_0_121_153 ();
 FILLER_ASAP7_75t_R FILLER_0_121_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_163 ();
 DECAPx4_ASAP7_75t_R FILLER_0_121_170 ();
 FILLER_ASAP7_75t_R FILLER_0_121_186 ();
 FILLER_ASAP7_75t_R FILLER_0_121_194 ();
 FILLER_ASAP7_75t_R FILLER_0_121_203 ();
 DECAPx2_ASAP7_75t_R FILLER_0_121_210 ();
 FILLER_ASAP7_75t_R FILLER_0_121_216 ();
 FILLER_ASAP7_75t_R FILLER_0_121_240 ();
 FILLER_ASAP7_75t_R FILLER_0_121_245 ();
 FILLER_ASAP7_75t_R FILLER_0_121_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_260 ();
 DECAPx1_ASAP7_75t_R FILLER_0_121_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_273 ();
 DECAPx2_ASAP7_75t_R FILLER_0_121_282 ();
 FILLER_ASAP7_75t_R FILLER_0_121_299 ();
 DECAPx2_ASAP7_75t_R FILLER_0_121_322 ();
 DECAPx2_ASAP7_75t_R FILLER_0_121_349 ();
 DECAPx1_ASAP7_75t_R FILLER_0_121_358 ();
 FILLER_ASAP7_75t_R FILLER_0_121_383 ();
 DECAPx6_ASAP7_75t_R FILLER_0_121_406 ();
 DECAPx2_ASAP7_75t_R FILLER_0_121_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_426 ();
 FILLER_ASAP7_75t_R FILLER_0_121_430 ();
 DECAPx4_ASAP7_75t_R FILLER_0_121_442 ();
 FILLER_ASAP7_75t_R FILLER_0_121_472 ();
 DECAPx2_ASAP7_75t_R FILLER_0_121_480 ();
 DECAPx1_ASAP7_75t_R FILLER_0_121_492 ();
 DECAPx1_ASAP7_75t_R FILLER_0_121_502 ();
 FILLER_ASAP7_75t_R FILLER_0_121_528 ();
 DECAPx1_ASAP7_75t_R FILLER_0_121_538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_548 ();
 DECAPx1_ASAP7_75t_R FILLER_0_121_570 ();
 DECAPx2_ASAP7_75t_R FILLER_0_121_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_586 ();
 FILLER_ASAP7_75t_R FILLER_0_121_593 ();
 FILLER_ASAP7_75t_R FILLER_0_121_605 ();
 DECAPx4_ASAP7_75t_R FILLER_0_121_613 ();
 FILLER_ASAP7_75t_R FILLER_0_121_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_625 ();
 FILLER_ASAP7_75t_R FILLER_0_121_634 ();
 DECAPx1_ASAP7_75t_R FILLER_0_121_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_647 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_658 ();
 DECAPx4_ASAP7_75t_R FILLER_0_121_680 ();
 DECAPx4_ASAP7_75t_R FILLER_0_121_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_706 ();
 DECAPx6_ASAP7_75t_R FILLER_0_121_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_729 ();
 DECAPx2_ASAP7_75t_R FILLER_0_121_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_742 ();
 FILLER_ASAP7_75t_R FILLER_0_121_749 ();
 DECAPx6_ASAP7_75t_R FILLER_0_121_757 ();
 DECAPx2_ASAP7_75t_R FILLER_0_121_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_777 ();
 FILLER_ASAP7_75t_R FILLER_0_121_784 ();
 FILLER_ASAP7_75t_R FILLER_0_121_792 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_805 ();
 DECAPx2_ASAP7_75t_R FILLER_0_121_827 ();
 FILLER_ASAP7_75t_R FILLER_0_121_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_835 ();
 DECAPx2_ASAP7_75t_R FILLER_0_121_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_848 ();
 FILLER_ASAP7_75t_R FILLER_0_121_854 ();
 DECAPx2_ASAP7_75t_R FILLER_0_121_862 ();
 FILLER_ASAP7_75t_R FILLER_0_121_874 ();
 DECAPx6_ASAP7_75t_R FILLER_0_121_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_896 ();
 FILLER_ASAP7_75t_R FILLER_0_121_903 ();
 DECAPx6_ASAP7_75t_R FILLER_0_121_911 ();
 DECAPx4_ASAP7_75t_R FILLER_0_121_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_937 ();
 FILLER_ASAP7_75t_R FILLER_0_121_950 ();
 DECAPx4_ASAP7_75t_R FILLER_0_121_962 ();
 FILLER_ASAP7_75t_R FILLER_0_121_972 ();
 DECAPx2_ASAP7_75t_R FILLER_0_121_984 ();
 DECAPx2_ASAP7_75t_R FILLER_0_121_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_1015 ();
 DECAPx1_ASAP7_75t_R FILLER_0_121_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_1041 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_1050 ();
 FILLER_ASAP7_75t_R FILLER_0_121_1072 ();
 FILLER_ASAP7_75t_R FILLER_0_121_1082 ();
 FILLER_ASAP7_75t_R FILLER_0_121_1092 ();
 DECAPx6_ASAP7_75t_R FILLER_0_121_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_1112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_1119 ();
 DECAPx2_ASAP7_75t_R FILLER_0_121_1141 ();
 FILLER_ASAP7_75t_R FILLER_0_121_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_1149 ();
 DECAPx1_ASAP7_75t_R FILLER_0_121_1160 ();
 FILLER_ASAP7_75t_R FILLER_0_121_1168 ();
 DECAPx2_ASAP7_75t_R FILLER_0_121_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_1196 ();
 FILLER_ASAP7_75t_R FILLER_0_121_1207 ();
 FILLER_ASAP7_75t_R FILLER_0_121_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_1214 ();
 FILLER_ASAP7_75t_R FILLER_0_121_1225 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_1227 ();
 FILLER_ASAP7_75t_R FILLER_0_121_1234 ();
 DECAPx4_ASAP7_75t_R FILLER_0_121_1242 ();
 FILLER_ASAP7_75t_R FILLER_0_121_1258 ();
 DECAPx1_ASAP7_75t_R FILLER_0_121_1266 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_1270 ();
 DECAPx6_ASAP7_75t_R FILLER_0_121_1277 ();
 FILLER_ASAP7_75t_R FILLER_0_121_1291 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_1293 ();
 DECAPx4_ASAP7_75t_R FILLER_0_121_1300 ();
 FILLER_ASAP7_75t_R FILLER_0_121_1317 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_1319 ();
 FILLER_ASAP7_75t_R FILLER_0_121_1323 ();
 DECAPx1_ASAP7_75t_R FILLER_0_121_1347 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_1351 ();
 FILLER_ASAP7_75t_R FILLER_0_121_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_121_1364 ();
 DECAPx1_ASAP7_75t_R FILLER_0_121_1371 ();
 FILLER_ASAP7_75t_R FILLER_0_121_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_122_2 ();
 FILLER_ASAP7_75t_R FILLER_0_122_9 ();
 FILLER_ASAP7_75t_R FILLER_0_122_16 ();
 FILLER_ASAP7_75t_R FILLER_0_122_23 ();
 FILLER_ASAP7_75t_R FILLER_0_122_30 ();
 DECAPx1_ASAP7_75t_R FILLER_0_122_35 ();
 FILLER_ASAP7_75t_R FILLER_0_122_50 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_55 ();
 DECAPx4_ASAP7_75t_R FILLER_0_122_77 ();
 DECAPx4_ASAP7_75t_R FILLER_0_122_93 ();
 FILLER_ASAP7_75t_R FILLER_0_122_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_105 ();
 DECAPx2_ASAP7_75t_R FILLER_0_122_116 ();
 FILLER_ASAP7_75t_R FILLER_0_122_122 ();
 DECAPx1_ASAP7_75t_R FILLER_0_122_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_122_145 ();
 FILLER_ASAP7_75t_R FILLER_0_122_157 ();
 FILLER_ASAP7_75t_R FILLER_0_122_164 ();
 FILLER_ASAP7_75t_R FILLER_0_122_169 ();
 DECAPx6_ASAP7_75t_R FILLER_0_122_174 ();
 DECAPx2_ASAP7_75t_R FILLER_0_122_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_194 ();
 DECAPx6_ASAP7_75t_R FILLER_0_122_201 ();
 FILLER_ASAP7_75t_R FILLER_0_122_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_217 ();
 FILLER_ASAP7_75t_R FILLER_0_122_240 ();
 DECAPx2_ASAP7_75t_R FILLER_0_122_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_262 ();
 DECAPx1_ASAP7_75t_R FILLER_0_122_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_275 ();
 FILLER_ASAP7_75t_R FILLER_0_122_284 ();
 DECAPx4_ASAP7_75t_R FILLER_0_122_289 ();
 FILLER_ASAP7_75t_R FILLER_0_122_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_301 ();
 DECAPx2_ASAP7_75t_R FILLER_0_122_307 ();
 FILLER_ASAP7_75t_R FILLER_0_122_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_315 ();
 FILLER_ASAP7_75t_R FILLER_0_122_324 ();
 FILLER_ASAP7_75t_R FILLER_0_122_329 ();
 FILLER_ASAP7_75t_R FILLER_0_122_337 ();
 FILLER_ASAP7_75t_R FILLER_0_122_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_344 ();
 DECAPx1_ASAP7_75t_R FILLER_0_122_350 ();
 FILLER_ASAP7_75t_R FILLER_0_122_362 ();
 FILLER_ASAP7_75t_R FILLER_0_122_370 ();
 FILLER_ASAP7_75t_R FILLER_0_122_375 ();
 FILLER_ASAP7_75t_R FILLER_0_122_380 ();
 FILLER_ASAP7_75t_R FILLER_0_122_392 ();
 FILLER_ASAP7_75t_R FILLER_0_122_400 ();
 FILLER_ASAP7_75t_R FILLER_0_122_412 ();
 FILLER_ASAP7_75t_R FILLER_0_122_436 ();
 FILLER_ASAP7_75t_R FILLER_0_122_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_446 ();
 DECAPx2_ASAP7_75t_R FILLER_0_122_453 ();
 FILLER_ASAP7_75t_R FILLER_0_122_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_461 ();
 DECAPx4_ASAP7_75t_R FILLER_0_122_464 ();
 DECAPx2_ASAP7_75t_R FILLER_0_122_480 ();
 DECAPx2_ASAP7_75t_R FILLER_0_122_492 ();
 FILLER_ASAP7_75t_R FILLER_0_122_498 ();
 DECAPx2_ASAP7_75t_R FILLER_0_122_506 ();
 FILLER_ASAP7_75t_R FILLER_0_122_512 ();
 DECAPx2_ASAP7_75t_R FILLER_0_122_529 ();
 DECAPx2_ASAP7_75t_R FILLER_0_122_541 ();
 FILLER_ASAP7_75t_R FILLER_0_122_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_549 ();
 DECAPx2_ASAP7_75t_R FILLER_0_122_556 ();
 FILLER_ASAP7_75t_R FILLER_0_122_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_564 ();
 DECAPx1_ASAP7_75t_R FILLER_0_122_573 ();
 DECAPx1_ASAP7_75t_R FILLER_0_122_583 ();
 DECAPx2_ASAP7_75t_R FILLER_0_122_595 ();
 FILLER_ASAP7_75t_R FILLER_0_122_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_603 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_610 ();
 DECAPx2_ASAP7_75t_R FILLER_0_122_632 ();
 FILLER_ASAP7_75t_R FILLER_0_122_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_640 ();
 FILLER_ASAP7_75t_R FILLER_0_122_655 ();
 FILLER_ASAP7_75t_R FILLER_0_122_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_668 ();
 DECAPx2_ASAP7_75t_R FILLER_0_122_696 ();
 FILLER_ASAP7_75t_R FILLER_0_122_702 ();
 FILLER_ASAP7_75t_R FILLER_0_122_716 ();
 DECAPx6_ASAP7_75t_R FILLER_0_122_724 ();
 DECAPx1_ASAP7_75t_R FILLER_0_122_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_749 ();
 DECAPx4_ASAP7_75t_R FILLER_0_122_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_781 ();
 FILLER_ASAP7_75t_R FILLER_0_122_790 ();
 FILLER_ASAP7_75t_R FILLER_0_122_798 ();
 DECAPx1_ASAP7_75t_R FILLER_0_122_803 ();
 DECAPx2_ASAP7_75t_R FILLER_0_122_813 ();
 FILLER_ASAP7_75t_R FILLER_0_122_819 ();
 DECAPx4_ASAP7_75t_R FILLER_0_122_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_837 ();
 FILLER_ASAP7_75t_R FILLER_0_122_846 ();
 FILLER_ASAP7_75t_R FILLER_0_122_854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_886 ();
 DECAPx1_ASAP7_75t_R FILLER_0_122_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_912 ();
 FILLER_ASAP7_75t_R FILLER_0_122_919 ();
 FILLER_ASAP7_75t_R FILLER_0_122_931 ();
 FILLER_ASAP7_75t_R FILLER_0_122_943 ();
 FILLER_ASAP7_75t_R FILLER_0_122_955 ();
 FILLER_ASAP7_75t_R FILLER_0_122_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_962 ();
 FILLER_ASAP7_75t_R FILLER_0_122_967 ();
 DECAPx6_ASAP7_75t_R FILLER_0_122_977 ();
 DECAPx6_ASAP7_75t_R FILLER_0_122_999 ();
 FILLER_ASAP7_75t_R FILLER_0_122_1013 ();
 FILLER_ASAP7_75t_R FILLER_0_122_1018 ();
 DECAPx2_ASAP7_75t_R FILLER_0_122_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_1037 ();
 DECAPx6_ASAP7_75t_R FILLER_0_122_1049 ();
 FILLER_ASAP7_75t_R FILLER_0_122_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_1065 ();
 FILLER_ASAP7_75t_R FILLER_0_122_1072 ();
 FILLER_ASAP7_75t_R FILLER_0_122_1080 ();
 DECAPx6_ASAP7_75t_R FILLER_0_122_1088 ();
 DECAPx2_ASAP7_75t_R FILLER_0_122_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_1108 ();
 DECAPx6_ASAP7_75t_R FILLER_0_122_1117 ();
 DECAPx2_ASAP7_75t_R FILLER_0_122_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_1137 ();
 FILLER_ASAP7_75t_R FILLER_0_122_1162 ();
 FILLER_ASAP7_75t_R FILLER_0_122_1176 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_1178 ();
 FILLER_ASAP7_75t_R FILLER_0_122_1187 ();
 DECAPx1_ASAP7_75t_R FILLER_0_122_1195 ();
 DECAPx2_ASAP7_75t_R FILLER_0_122_1209 ();
 FILLER_ASAP7_75t_R FILLER_0_122_1222 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_1233 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_1255 ();
 FILLER_ASAP7_75t_R FILLER_0_122_1263 ();
 FILLER_ASAP7_75t_R FILLER_0_122_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_0_122_1280 ();
 FILLER_ASAP7_75t_R FILLER_0_122_1286 ();
 DECAPx6_ASAP7_75t_R FILLER_0_122_1298 ();
 DECAPx1_ASAP7_75t_R FILLER_0_122_1312 ();
 FILLER_ASAP7_75t_R FILLER_0_122_1319 ();
 FILLER_ASAP7_75t_R FILLER_0_122_1331 ();
 DECAPx1_ASAP7_75t_R FILLER_0_122_1336 ();
 FILLER_ASAP7_75t_R FILLER_0_122_1343 ();
 FILLER_ASAP7_75t_R FILLER_0_122_1350 ();
 FILLER_ASAP7_75t_R FILLER_0_122_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_122_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_123_2 ();
 FILLER_ASAP7_75t_R FILLER_0_123_26 ();
 FILLER_ASAP7_75t_R FILLER_0_123_34 ();
 FILLER_ASAP7_75t_R FILLER_0_123_42 ();
 FILLER_ASAP7_75t_R FILLER_0_123_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_69 ();
 FILLER_ASAP7_75t_R FILLER_0_123_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_93 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_122 ();
 FILLER_ASAP7_75t_R FILLER_0_123_133 ();
 FILLER_ASAP7_75t_R FILLER_0_123_140 ();
 FILLER_ASAP7_75t_R FILLER_0_123_147 ();
 FILLER_ASAP7_75t_R FILLER_0_123_155 ();
 FILLER_ASAP7_75t_R FILLER_0_123_160 ();
 FILLER_ASAP7_75t_R FILLER_0_123_168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_176 ();
 DECAPx6_ASAP7_75t_R FILLER_0_123_198 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_216 ();
 DECAPx2_ASAP7_75t_R FILLER_0_123_223 ();
 FILLER_ASAP7_75t_R FILLER_0_123_237 ();
 FILLER_ASAP7_75t_R FILLER_0_123_257 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_269 ();
 DECAPx6_ASAP7_75t_R FILLER_0_123_281 ();
 FILLER_ASAP7_75t_R FILLER_0_123_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_297 ();
 FILLER_ASAP7_75t_R FILLER_0_123_308 ();
 FILLER_ASAP7_75t_R FILLER_0_123_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_324 ();
 FILLER_ASAP7_75t_R FILLER_0_123_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_332 ();
 FILLER_ASAP7_75t_R FILLER_0_123_338 ();
 FILLER_ASAP7_75t_R FILLER_0_123_350 ();
 FILLER_ASAP7_75t_R FILLER_0_123_357 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_364 ();
 FILLER_ASAP7_75t_R FILLER_0_123_396 ();
 DECAPx6_ASAP7_75t_R FILLER_0_123_401 ();
 DECAPx4_ASAP7_75t_R FILLER_0_123_426 ();
 FILLER_ASAP7_75t_R FILLER_0_123_436 ();
 FILLER_ASAP7_75t_R FILLER_0_123_445 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_457 ();
 FILLER_ASAP7_75t_R FILLER_0_123_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_470 ();
 DECAPx2_ASAP7_75t_R FILLER_0_123_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_485 ();
 DECAPx2_ASAP7_75t_R FILLER_0_123_492 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_504 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_519 ();
 FILLER_ASAP7_75t_R FILLER_0_123_526 ();
 FILLER_ASAP7_75t_R FILLER_0_123_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_540 ();
 FILLER_ASAP7_75t_R FILLER_0_123_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_550 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_558 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_568 ();
 FILLER_ASAP7_75t_R FILLER_0_123_583 ();
 DECAPx6_ASAP7_75t_R FILLER_0_123_590 ();
 FILLER_ASAP7_75t_R FILLER_0_123_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_606 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_617 ();
 DECAPx2_ASAP7_75t_R FILLER_0_123_624 ();
 DECAPx2_ASAP7_75t_R FILLER_0_123_642 ();
 FILLER_ASAP7_75t_R FILLER_0_123_658 ();
 DECAPx6_ASAP7_75t_R FILLER_0_123_670 ();
 FILLER_ASAP7_75t_R FILLER_0_123_684 ();
 FILLER_ASAP7_75t_R FILLER_0_123_692 ();
 FILLER_ASAP7_75t_R FILLER_0_123_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_716 ();
 FILLER_ASAP7_75t_R FILLER_0_123_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_729 ();
 DECAPx6_ASAP7_75t_R FILLER_0_123_746 ();
 FILLER_ASAP7_75t_R FILLER_0_123_760 ();
 FILLER_ASAP7_75t_R FILLER_0_123_772 ();
 FILLER_ASAP7_75t_R FILLER_0_123_781 ();
 DECAPx6_ASAP7_75t_R FILLER_0_123_789 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_807 ();
 FILLER_ASAP7_75t_R FILLER_0_123_820 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_828 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_842 ();
 FILLER_ASAP7_75t_R FILLER_0_123_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_851 ();
 FILLER_ASAP7_75t_R FILLER_0_123_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_860 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_867 ();
 FILLER_ASAP7_75t_R FILLER_0_123_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_876 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_880 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_890 ();
 DECAPx2_ASAP7_75t_R FILLER_0_123_900 ();
 FILLER_ASAP7_75t_R FILLER_0_123_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_908 ();
 DECAPx4_ASAP7_75t_R FILLER_0_123_915 ();
 DECAPx4_ASAP7_75t_R FILLER_0_123_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_937 ();
 FILLER_ASAP7_75t_R FILLER_0_123_958 ();
 FILLER_ASAP7_75t_R FILLER_0_123_968 ();
 DECAPx4_ASAP7_75t_R FILLER_0_123_980 ();
 FILLER_ASAP7_75t_R FILLER_0_123_998 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_1007 ();
 FILLER_ASAP7_75t_R FILLER_0_123_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_1013 ();
 DECAPx2_ASAP7_75t_R FILLER_0_123_1025 ();
 FILLER_ASAP7_75t_R FILLER_0_123_1031 ();
 FILLER_ASAP7_75t_R FILLER_0_123_1039 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_1047 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_1059 ();
 FILLER_ASAP7_75t_R FILLER_0_123_1075 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_1083 ();
 FILLER_ASAP7_75t_R FILLER_0_123_1108 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_1117 ();
 DECAPx2_ASAP7_75t_R FILLER_0_123_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_1127 ();
 DECAPx4_ASAP7_75t_R FILLER_0_123_1134 ();
 FILLER_ASAP7_75t_R FILLER_0_123_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_1146 ();
 FILLER_ASAP7_75t_R FILLER_0_123_1157 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_1167 ();
 FILLER_ASAP7_75t_R FILLER_0_123_1181 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_1193 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_1200 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_1222 ();
 FILLER_ASAP7_75t_R FILLER_0_123_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_1243 ();
 DECAPx2_ASAP7_75t_R FILLER_0_123_1265 ();
 FILLER_ASAP7_75t_R FILLER_0_123_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_1301 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_1323 ();
 FILLER_ASAP7_75t_R FILLER_0_123_1327 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_1335 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_1339 ();
 FILLER_ASAP7_75t_R FILLER_0_123_1361 ();
 FILLER_ASAP7_75t_R FILLER_0_123_1369 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_124_2 ();
 FILLER_ASAP7_75t_R FILLER_0_124_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_11 ();
 FILLER_ASAP7_75t_R FILLER_0_124_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_19 ();
 FILLER_ASAP7_75t_R FILLER_0_124_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_27 ();
 FILLER_ASAP7_75t_R FILLER_0_124_34 ();
 FILLER_ASAP7_75t_R FILLER_0_124_41 ();
 FILLER_ASAP7_75t_R FILLER_0_124_53 ();
 FILLER_ASAP7_75t_R FILLER_0_124_61 ();
 DECAPx1_ASAP7_75t_R FILLER_0_124_69 ();
 FILLER_ASAP7_75t_R FILLER_0_124_76 ();
 DECAPx2_ASAP7_75t_R FILLER_0_124_84 ();
 FILLER_ASAP7_75t_R FILLER_0_124_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_92 ();
 DECAPx4_ASAP7_75t_R FILLER_0_124_96 ();
 FILLER_ASAP7_75t_R FILLER_0_124_106 ();
 DECAPx2_ASAP7_75t_R FILLER_0_124_118 ();
 DECAPx2_ASAP7_75t_R FILLER_0_124_136 ();
 FILLER_ASAP7_75t_R FILLER_0_124_142 ();
 DECAPx1_ASAP7_75t_R FILLER_0_124_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_151 ();
 FILLER_ASAP7_75t_R FILLER_0_124_158 ();
 FILLER_ASAP7_75t_R FILLER_0_124_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_175 ();
 DECAPx4_ASAP7_75t_R FILLER_0_124_203 ();
 FILLER_ASAP7_75t_R FILLER_0_124_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_223 ();
 FILLER_ASAP7_75t_R FILLER_0_124_227 ();
 FILLER_ASAP7_75t_R FILLER_0_124_232 ();
 DECAPx2_ASAP7_75t_R FILLER_0_124_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_252 ();
 FILLER_ASAP7_75t_R FILLER_0_124_271 ();
 DECAPx2_ASAP7_75t_R FILLER_0_124_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_287 ();
 FILLER_ASAP7_75t_R FILLER_0_124_293 ();
 DECAPx6_ASAP7_75t_R FILLER_0_124_310 ();
 FILLER_ASAP7_75t_R FILLER_0_124_330 ();
 FILLER_ASAP7_75t_R FILLER_0_124_337 ();
 FILLER_ASAP7_75t_R FILLER_0_124_349 ();
 FILLER_ASAP7_75t_R FILLER_0_124_355 ();
 DECAPx4_ASAP7_75t_R FILLER_0_124_368 ();
 FILLER_ASAP7_75t_R FILLER_0_124_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_386 ();
 DECAPx4_ASAP7_75t_R FILLER_0_124_408 ();
 FILLER_ASAP7_75t_R FILLER_0_124_418 ();
 DECAPx4_ASAP7_75t_R FILLER_0_124_430 ();
 FILLER_ASAP7_75t_R FILLER_0_124_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_442 ();
 FILLER_ASAP7_75t_R FILLER_0_124_449 ();
 DECAPx1_ASAP7_75t_R FILLER_0_124_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_461 ();
 DECAPx1_ASAP7_75t_R FILLER_0_124_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_468 ();
 FILLER_ASAP7_75t_R FILLER_0_124_476 ();
 DECAPx6_ASAP7_75t_R FILLER_0_124_484 ();
 FILLER_ASAP7_75t_R FILLER_0_124_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_500 ();
 FILLER_ASAP7_75t_R FILLER_0_124_507 ();
 DECAPx6_ASAP7_75t_R FILLER_0_124_517 ();
 FILLER_ASAP7_75t_R FILLER_0_124_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_533 ();
 DECAPx6_ASAP7_75t_R FILLER_0_124_544 ();
 FILLER_ASAP7_75t_R FILLER_0_124_568 ();
 DECAPx6_ASAP7_75t_R FILLER_0_124_575 ();
 FILLER_ASAP7_75t_R FILLER_0_124_589 ();
 DECAPx4_ASAP7_75t_R FILLER_0_124_597 ();
 FILLER_ASAP7_75t_R FILLER_0_124_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_615 ();
 FILLER_ASAP7_75t_R FILLER_0_124_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_624 ();
 FILLER_ASAP7_75t_R FILLER_0_124_631 ();
 DECAPx2_ASAP7_75t_R FILLER_0_124_645 ();
 FILLER_ASAP7_75t_R FILLER_0_124_661 ();
 FILLER_ASAP7_75t_R FILLER_0_124_669 ();
 FILLER_ASAP7_75t_R FILLER_0_124_677 ();
 DECAPx2_ASAP7_75t_R FILLER_0_124_691 ();
 FILLER_ASAP7_75t_R FILLER_0_124_697 ();
 FILLER_ASAP7_75t_R FILLER_0_124_705 ();
 DECAPx4_ASAP7_75t_R FILLER_0_124_713 ();
 FILLER_ASAP7_75t_R FILLER_0_124_723 ();
 FILLER_ASAP7_75t_R FILLER_0_124_736 ();
 FILLER_ASAP7_75t_R FILLER_0_124_746 ();
 DECAPx2_ASAP7_75t_R FILLER_0_124_754 ();
 FILLER_ASAP7_75t_R FILLER_0_124_760 ();
 FILLER_ASAP7_75t_R FILLER_0_124_770 ();
 DECAPx2_ASAP7_75t_R FILLER_0_124_776 ();
 FILLER_ASAP7_75t_R FILLER_0_124_782 ();
 DECAPx6_ASAP7_75t_R FILLER_0_124_790 ();
 DECAPx2_ASAP7_75t_R FILLER_0_124_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_810 ();
 DECAPx1_ASAP7_75t_R FILLER_0_124_817 ();
 FILLER_ASAP7_75t_R FILLER_0_124_827 ();
 DECAPx2_ASAP7_75t_R FILLER_0_124_835 ();
 DECAPx1_ASAP7_75t_R FILLER_0_124_851 ();
 FILLER_ASAP7_75t_R FILLER_0_124_860 ();
 FILLER_ASAP7_75t_R FILLER_0_124_874 ();
 FILLER_ASAP7_75t_R FILLER_0_124_882 ();
 FILLER_ASAP7_75t_R FILLER_0_124_891 ();
 DECAPx4_ASAP7_75t_R FILLER_0_124_901 ();
 FILLER_ASAP7_75t_R FILLER_0_124_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_913 ();
 FILLER_ASAP7_75t_R FILLER_0_124_917 ();
 DECAPx6_ASAP7_75t_R FILLER_0_124_925 ();
 DECAPx1_ASAP7_75t_R FILLER_0_124_939 ();
 DECAPx1_ASAP7_75t_R FILLER_0_124_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_957 ();
 FILLER_ASAP7_75t_R FILLER_0_124_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_970 ();
 DECAPx4_ASAP7_75t_R FILLER_0_124_979 ();
 FILLER_ASAP7_75t_R FILLER_0_124_1000 ();
 FILLER_ASAP7_75t_R FILLER_0_124_1010 ();
 FILLER_ASAP7_75t_R FILLER_0_124_1020 ();
 DECAPx2_ASAP7_75t_R FILLER_0_124_1028 ();
 FILLER_ASAP7_75t_R FILLER_0_124_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_1036 ();
 DECAPx1_ASAP7_75t_R FILLER_0_124_1040 ();
 DECAPx4_ASAP7_75t_R FILLER_0_124_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_1065 ();
 FILLER_ASAP7_75t_R FILLER_0_124_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_1080 ();
 FILLER_ASAP7_75t_R FILLER_0_124_1084 ();
 DECAPx2_ASAP7_75t_R FILLER_0_124_1098 ();
 FILLER_ASAP7_75t_R FILLER_0_124_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_1106 ();
 DECAPx2_ASAP7_75t_R FILLER_0_124_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_1137 ();
 FILLER_ASAP7_75t_R FILLER_0_124_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_1171 ();
 FILLER_ASAP7_75t_R FILLER_0_124_1182 ();
 FILLER_ASAP7_75t_R FILLER_0_124_1190 ();
 DECAPx2_ASAP7_75t_R FILLER_0_124_1198 ();
 DECAPx1_ASAP7_75t_R FILLER_0_124_1214 ();
 FILLER_ASAP7_75t_R FILLER_0_124_1228 ();
 FILLER_ASAP7_75t_R FILLER_0_124_1238 ();
 DECAPx2_ASAP7_75t_R FILLER_0_124_1245 ();
 DECAPx2_ASAP7_75t_R FILLER_0_124_1258 ();
 FILLER_ASAP7_75t_R FILLER_0_124_1270 ();
 DECAPx2_ASAP7_75t_R FILLER_0_124_1275 ();
 FILLER_ASAP7_75t_R FILLER_0_124_1281 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_1283 ();
 FILLER_ASAP7_75t_R FILLER_0_124_1294 ();
 DECAPx6_ASAP7_75t_R FILLER_0_124_1302 ();
 DECAPx2_ASAP7_75t_R FILLER_0_124_1316 ();
 FILLER_ASAP7_75t_R FILLER_0_124_1330 ();
 FILLER_ASAP7_75t_R FILLER_0_124_1338 ();
 FILLER_ASAP7_75t_R FILLER_0_124_1343 ();
 FILLER_ASAP7_75t_R FILLER_0_124_1351 ();
 FILLER_ASAP7_75t_R FILLER_0_124_1359 ();
 FILLER_ASAP7_75t_R FILLER_0_124_1366 ();
 FILLER_ASAP7_75t_R FILLER_0_124_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_124_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_125_2 ();
 FILLER_ASAP7_75t_R FILLER_0_125_25 ();
 FILLER_ASAP7_75t_R FILLER_0_125_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_125_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_125_59 ();
 FILLER_ASAP7_75t_R FILLER_0_125_70 ();
 FILLER_ASAP7_75t_R FILLER_0_125_78 ();
 DECAPx2_ASAP7_75t_R FILLER_0_125_83 ();
 FILLER_ASAP7_75t_R FILLER_0_125_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_125_91 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_112 ();
 DECAPx4_ASAP7_75t_R FILLER_0_125_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_125_144 ();
 DECAPx4_ASAP7_75t_R FILLER_0_125_155 ();
 FILLER_ASAP7_75t_R FILLER_0_125_165 ();
 DECAPx2_ASAP7_75t_R FILLER_0_125_173 ();
 FILLER_ASAP7_75t_R FILLER_0_125_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_125_181 ();
 FILLER_ASAP7_75t_R FILLER_0_125_187 ();
 DECAPx2_ASAP7_75t_R FILLER_0_125_209 ();
 FILLER_ASAP7_75t_R FILLER_0_125_215 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_125_247 ();
 FILLER_ASAP7_75t_R FILLER_0_125_259 ();
 FILLER_ASAP7_75t_R FILLER_0_125_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_125_271 ();
 DECAPx2_ASAP7_75t_R FILLER_0_125_282 ();
 FILLER_ASAP7_75t_R FILLER_0_125_288 ();
 FILLER_ASAP7_75t_R FILLER_0_125_298 ();
 FILLER_ASAP7_75t_R FILLER_0_125_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_125_312 ();
 DECAPx1_ASAP7_75t_R FILLER_0_125_337 ();
 DECAPx1_ASAP7_75t_R FILLER_0_125_351 ();
 DECAPx1_ASAP7_75t_R FILLER_0_125_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_125_369 ();
 FILLER_ASAP7_75t_R FILLER_0_125_378 ();
 FILLER_ASAP7_75t_R FILLER_0_125_383 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_393 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_415 ();
 DECAPx2_ASAP7_75t_R FILLER_0_125_437 ();
 FILLER_ASAP7_75t_R FILLER_0_125_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_125_445 ();
 DECAPx6_ASAP7_75t_R FILLER_0_125_452 ();
 DECAPx1_ASAP7_75t_R FILLER_0_125_466 ();
 FILLER_ASAP7_75t_R FILLER_0_125_480 ();
 DECAPx6_ASAP7_75t_R FILLER_0_125_487 ();
 FILLER_ASAP7_75t_R FILLER_0_125_501 ();
 FILLER_ASAP7_75t_R FILLER_0_125_509 ();
 FILLER_ASAP7_75t_R FILLER_0_125_517 ();
 DECAPx6_ASAP7_75t_R FILLER_0_125_522 ();
 DECAPx1_ASAP7_75t_R FILLER_0_125_536 ();
 FILLER_ASAP7_75t_R FILLER_0_125_550 ();
 DECAPx1_ASAP7_75t_R FILLER_0_125_558 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_125_562 ();
 DECAPx2_ASAP7_75t_R FILLER_0_125_568 ();
 FILLER_ASAP7_75t_R FILLER_0_125_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_581 ();
 FILLER_ASAP7_75t_R FILLER_0_125_609 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_617 ();
 FILLER_ASAP7_75t_R FILLER_0_125_639 ();
 FILLER_ASAP7_75t_R FILLER_0_125_647 ();
 FILLER_ASAP7_75t_R FILLER_0_125_659 ();
 FILLER_ASAP7_75t_R FILLER_0_125_669 ();
 FILLER_ASAP7_75t_R FILLER_0_125_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_125_678 ();
 DECAPx6_ASAP7_75t_R FILLER_0_125_685 ();
 DECAPx6_ASAP7_75t_R FILLER_0_125_705 ();
 FILLER_ASAP7_75t_R FILLER_0_125_719 ();
 DECAPx2_ASAP7_75t_R FILLER_0_125_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_125_739 ();
 FILLER_ASAP7_75t_R FILLER_0_125_746 ();
 FILLER_ASAP7_75t_R FILLER_0_125_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_125_756 ();
 DECAPx2_ASAP7_75t_R FILLER_0_125_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_125_766 ();
 DECAPx4_ASAP7_75t_R FILLER_0_125_773 ();
 DECAPx2_ASAP7_75t_R FILLER_0_125_794 ();
 FILLER_ASAP7_75t_R FILLER_0_125_800 ();
 FILLER_ASAP7_75t_R FILLER_0_125_808 ();
 DECAPx1_ASAP7_75t_R FILLER_0_125_816 ();
 DECAPx2_ASAP7_75t_R FILLER_0_125_831 ();
 FILLER_ASAP7_75t_R FILLER_0_125_837 ();
 DECAPx4_ASAP7_75t_R FILLER_0_125_845 ();
 DECAPx2_ASAP7_75t_R FILLER_0_125_875 ();
 FILLER_ASAP7_75t_R FILLER_0_125_881 ();
 FILLER_ASAP7_75t_R FILLER_0_125_889 ();
 DECAPx4_ASAP7_75t_R FILLER_0_125_897 ();
 FILLER_ASAP7_75t_R FILLER_0_125_907 ();
 DECAPx1_ASAP7_75t_R FILLER_0_125_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_125_916 ();
 FILLER_ASAP7_75t_R FILLER_0_125_923 ();
 DECAPx6_ASAP7_75t_R FILLER_0_125_927 ();
 DECAPx2_ASAP7_75t_R FILLER_0_125_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_125_947 ();
 DECAPx2_ASAP7_75t_R FILLER_0_125_953 ();
 DECAPx2_ASAP7_75t_R FILLER_0_125_967 ();
 FILLER_ASAP7_75t_R FILLER_0_125_973 ();
 FILLER_ASAP7_75t_R FILLER_0_125_985 ();
 FILLER_ASAP7_75t_R FILLER_0_125_995 ();
 DECAPx6_ASAP7_75t_R FILLER_0_125_1005 ();
 DECAPx1_ASAP7_75t_R FILLER_0_125_1019 ();
 FILLER_ASAP7_75t_R FILLER_0_125_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_125_1046 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_1053 ();
 DECAPx1_ASAP7_75t_R FILLER_0_125_1075 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_1091 ();
 DECAPx6_ASAP7_75t_R FILLER_0_125_1113 ();
 DECAPx2_ASAP7_75t_R FILLER_0_125_1127 ();
 DECAPx2_ASAP7_75t_R FILLER_0_125_1153 ();
 FILLER_ASAP7_75t_R FILLER_0_125_1169 ();
 DECAPx2_ASAP7_75t_R FILLER_0_125_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_125_1187 ();
 FILLER_ASAP7_75t_R FILLER_0_125_1193 ();
 DECAPx1_ASAP7_75t_R FILLER_0_125_1205 ();
 FILLER_ASAP7_75t_R FILLER_0_125_1219 ();
 FILLER_ASAP7_75t_R FILLER_0_125_1227 ();
 DECAPx1_ASAP7_75t_R FILLER_0_125_1239 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_125_1243 ();
 FILLER_ASAP7_75t_R FILLER_0_125_1254 ();
 FILLER_ASAP7_75t_R FILLER_0_125_1266 ();
 FILLER_ASAP7_75t_R FILLER_0_125_1276 ();
 DECAPx2_ASAP7_75t_R FILLER_0_125_1285 ();
 FILLER_ASAP7_75t_R FILLER_0_125_1291 ();
 FILLER_ASAP7_75t_R FILLER_0_125_1303 ();
 FILLER_ASAP7_75t_R FILLER_0_125_1311 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_125_1313 ();
 FILLER_ASAP7_75t_R FILLER_0_125_1320 ();
 DECAPx2_ASAP7_75t_R FILLER_0_125_1342 ();
 DECAPx1_ASAP7_75t_R FILLER_0_125_1370 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_125_1374 ();
 FILLER_ASAP7_75t_R FILLER_0_125_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_126_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_4 ();
 FILLER_ASAP7_75t_R FILLER_0_126_11 ();
 FILLER_ASAP7_75t_R FILLER_0_126_18 ();
 FILLER_ASAP7_75t_R FILLER_0_126_26 ();
 FILLER_ASAP7_75t_R FILLER_0_126_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_35 ();
 FILLER_ASAP7_75t_R FILLER_0_126_42 ();
 FILLER_ASAP7_75t_R FILLER_0_126_50 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_62 ();
 DECAPx4_ASAP7_75t_R FILLER_0_126_84 ();
 FILLER_ASAP7_75t_R FILLER_0_126_94 ();
 FILLER_ASAP7_75t_R FILLER_0_126_102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_114 ();
 DECAPx6_ASAP7_75t_R FILLER_0_126_136 ();
 FILLER_ASAP7_75t_R FILLER_0_126_150 ();
 FILLER_ASAP7_75t_R FILLER_0_126_162 ();
 FILLER_ASAP7_75t_R FILLER_0_126_167 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_175 ();
 DECAPx2_ASAP7_75t_R FILLER_0_126_197 ();
 FILLER_ASAP7_75t_R FILLER_0_126_203 ();
 FILLER_ASAP7_75t_R FILLER_0_126_211 ();
 DECAPx6_ASAP7_75t_R FILLER_0_126_219 ();
 FILLER_ASAP7_75t_R FILLER_0_126_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_235 ();
 FILLER_ASAP7_75t_R FILLER_0_126_247 ();
 FILLER_ASAP7_75t_R FILLER_0_126_259 ();
 FILLER_ASAP7_75t_R FILLER_0_126_271 ();
 DECAPx2_ASAP7_75t_R FILLER_0_126_279 ();
 FILLER_ASAP7_75t_R FILLER_0_126_285 ();
 FILLER_ASAP7_75t_R FILLER_0_126_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_295 ();
 DECAPx1_ASAP7_75t_R FILLER_0_126_304 ();
 DECAPx1_ASAP7_75t_R FILLER_0_126_319 ();
 FILLER_ASAP7_75t_R FILLER_0_126_329 ();
 FILLER_ASAP7_75t_R FILLER_0_126_341 ();
 DECAPx1_ASAP7_75t_R FILLER_0_126_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_353 ();
 FILLER_ASAP7_75t_R FILLER_0_126_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_366 ();
 DECAPx1_ASAP7_75t_R FILLER_0_126_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_376 ();
 FILLER_ASAP7_75t_R FILLER_0_126_383 ();
 FILLER_ASAP7_75t_R FILLER_0_126_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_393 ();
 FILLER_ASAP7_75t_R FILLER_0_126_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_404 ();
 FILLER_ASAP7_75t_R FILLER_0_126_411 ();
 FILLER_ASAP7_75t_R FILLER_0_126_416 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_424 ();
 FILLER_ASAP7_75t_R FILLER_0_126_446 ();
 DECAPx2_ASAP7_75t_R FILLER_0_126_454 ();
 FILLER_ASAP7_75t_R FILLER_0_126_460 ();
 DECAPx1_ASAP7_75t_R FILLER_0_126_464 ();
 FILLER_ASAP7_75t_R FILLER_0_126_478 ();
 FILLER_ASAP7_75t_R FILLER_0_126_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_488 ();
 DECAPx4_ASAP7_75t_R FILLER_0_126_495 ();
 DECAPx2_ASAP7_75t_R FILLER_0_126_511 ();
 FILLER_ASAP7_75t_R FILLER_0_126_523 ();
 FILLER_ASAP7_75t_R FILLER_0_126_531 ();
 FILLER_ASAP7_75t_R FILLER_0_126_553 ();
 FILLER_ASAP7_75t_R FILLER_0_126_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_563 ();
 FILLER_ASAP7_75t_R FILLER_0_126_572 ();
 DECAPx1_ASAP7_75t_R FILLER_0_126_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_584 ();
 FILLER_ASAP7_75t_R FILLER_0_126_591 ();
 DECAPx4_ASAP7_75t_R FILLER_0_126_599 ();
 FILLER_ASAP7_75t_R FILLER_0_126_609 ();
 FILLER_ASAP7_75t_R FILLER_0_126_617 ();
 DECAPx4_ASAP7_75t_R FILLER_0_126_625 ();
 FILLER_ASAP7_75t_R FILLER_0_126_641 ();
 FILLER_ASAP7_75t_R FILLER_0_126_653 ();
 FILLER_ASAP7_75t_R FILLER_0_126_661 ();
 DECAPx4_ASAP7_75t_R FILLER_0_126_668 ();
 FILLER_ASAP7_75t_R FILLER_0_126_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_680 ();
 FILLER_ASAP7_75t_R FILLER_0_126_693 ();
 DECAPx2_ASAP7_75t_R FILLER_0_126_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_711 ();
 DECAPx1_ASAP7_75t_R FILLER_0_126_722 ();
 DECAPx1_ASAP7_75t_R FILLER_0_126_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_736 ();
 FILLER_ASAP7_75t_R FILLER_0_126_743 ();
 FILLER_ASAP7_75t_R FILLER_0_126_751 ();
 DECAPx1_ASAP7_75t_R FILLER_0_126_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_763 ();
 FILLER_ASAP7_75t_R FILLER_0_126_770 ();
 DECAPx1_ASAP7_75t_R FILLER_0_126_778 ();
 DECAPx4_ASAP7_75t_R FILLER_0_126_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_798 ();
 DECAPx6_ASAP7_75t_R FILLER_0_126_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_819 ();
 FILLER_ASAP7_75t_R FILLER_0_126_826 ();
 DECAPx6_ASAP7_75t_R FILLER_0_126_834 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_848 ();
 FILLER_ASAP7_75t_R FILLER_0_126_855 ();
 FILLER_ASAP7_75t_R FILLER_0_126_867 ();
 FILLER_ASAP7_75t_R FILLER_0_126_875 ();
 DECAPx4_ASAP7_75t_R FILLER_0_126_883 ();
 FILLER_ASAP7_75t_R FILLER_0_126_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_895 ();
 FILLER_ASAP7_75t_R FILLER_0_126_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_904 ();
 DECAPx6_ASAP7_75t_R FILLER_0_126_911 ();
 FILLER_ASAP7_75t_R FILLER_0_126_935 ();
 FILLER_ASAP7_75t_R FILLER_0_126_945 ();
 DECAPx2_ASAP7_75t_R FILLER_0_126_950 ();
 FILLER_ASAP7_75t_R FILLER_0_126_956 ();
 DECAPx2_ASAP7_75t_R FILLER_0_126_968 ();
 FILLER_ASAP7_75t_R FILLER_0_126_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_976 ();
 DECAPx6_ASAP7_75t_R FILLER_0_126_987 ();
 DECAPx6_ASAP7_75t_R FILLER_0_126_1009 ();
 FILLER_ASAP7_75t_R FILLER_0_126_1023 ();
 DECAPx4_ASAP7_75t_R FILLER_0_126_1028 ();
 FILLER_ASAP7_75t_R FILLER_0_126_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_1040 ();
 DECAPx2_ASAP7_75t_R FILLER_0_126_1051 ();
 FILLER_ASAP7_75t_R FILLER_0_126_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_1059 ();
 DECAPx4_ASAP7_75t_R FILLER_0_126_1068 ();
 FILLER_ASAP7_75t_R FILLER_0_126_1084 ();
 FILLER_ASAP7_75t_R FILLER_0_126_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_1096 ();
 DECAPx1_ASAP7_75t_R FILLER_0_126_1105 ();
 FILLER_ASAP7_75t_R FILLER_0_126_1119 ();
 FILLER_ASAP7_75t_R FILLER_0_126_1131 ();
 FILLER_ASAP7_75t_R FILLER_0_126_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_1141 ();
 FILLER_ASAP7_75t_R FILLER_0_126_1154 ();
 FILLER_ASAP7_75t_R FILLER_0_126_1166 ();
 FILLER_ASAP7_75t_R FILLER_0_126_1178 ();
 FILLER_ASAP7_75t_R FILLER_0_126_1186 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_1188 ();
 FILLER_ASAP7_75t_R FILLER_0_126_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_1213 ();
 DECAPx1_ASAP7_75t_R FILLER_0_126_1224 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_1228 ();
 DECAPx1_ASAP7_75t_R FILLER_0_126_1237 ();
 DECAPx1_ASAP7_75t_R FILLER_0_126_1251 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_126_1255 ();
 FILLER_ASAP7_75t_R FILLER_0_126_1266 ();
 FILLER_ASAP7_75t_R FILLER_0_126_1274 ();
 FILLER_ASAP7_75t_R FILLER_0_126_1282 ();
 DECAPx1_ASAP7_75t_R FILLER_0_126_1290 ();
 DECAPx1_ASAP7_75t_R FILLER_0_126_1304 ();
 FILLER_ASAP7_75t_R FILLER_0_126_1318 ();
 DECAPx1_ASAP7_75t_R FILLER_0_126_1326 ();
 FILLER_ASAP7_75t_R FILLER_0_126_1333 ();
 FILLER_ASAP7_75t_R FILLER_0_126_1338 ();
 DECAPx2_ASAP7_75t_R FILLER_0_126_1362 ();
 FILLER_ASAP7_75t_R FILLER_0_126_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_126_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_127_2 ();
 FILLER_ASAP7_75t_R FILLER_0_127_9 ();
 FILLER_ASAP7_75t_R FILLER_0_127_33 ();
 FILLER_ASAP7_75t_R FILLER_0_127_40 ();
 DECAPx2_ASAP7_75t_R FILLER_0_127_45 ();
 FILLER_ASAP7_75t_R FILLER_0_127_57 ();
 DECAPx4_ASAP7_75t_R FILLER_0_127_62 ();
 FILLER_ASAP7_75t_R FILLER_0_127_72 ();
 DECAPx2_ASAP7_75t_R FILLER_0_127_84 ();
 FILLER_ASAP7_75t_R FILLER_0_127_100 ();
 FILLER_ASAP7_75t_R FILLER_0_127_105 ();
 DECAPx6_ASAP7_75t_R FILLER_0_127_113 ();
 DECAPx1_ASAP7_75t_R FILLER_0_127_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_131 ();
 DECAPx4_ASAP7_75t_R FILLER_0_127_156 ();
 DECAPx1_ASAP7_75t_R FILLER_0_127_172 ();
 DECAPx1_ASAP7_75t_R FILLER_0_127_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_183 ();
 FILLER_ASAP7_75t_R FILLER_0_127_194 ();
 FILLER_ASAP7_75t_R FILLER_0_127_208 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_235 ();
 FILLER_ASAP7_75t_R FILLER_0_127_247 ();
 DECAPx1_ASAP7_75t_R FILLER_0_127_255 ();
 FILLER_ASAP7_75t_R FILLER_0_127_269 ();
 DECAPx6_ASAP7_75t_R FILLER_0_127_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_291 ();
 DECAPx6_ASAP7_75t_R FILLER_0_127_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_312 ();
 FILLER_ASAP7_75t_R FILLER_0_127_323 ();
 FILLER_ASAP7_75t_R FILLER_0_127_330 ();
 DECAPx2_ASAP7_75t_R FILLER_0_127_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_348 ();
 FILLER_ASAP7_75t_R FILLER_0_127_359 ();
 DECAPx4_ASAP7_75t_R FILLER_0_127_366 ();
 FILLER_ASAP7_75t_R FILLER_0_127_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_384 ();
 FILLER_ASAP7_75t_R FILLER_0_127_395 ();
 DECAPx1_ASAP7_75t_R FILLER_0_127_400 ();
 FILLER_ASAP7_75t_R FILLER_0_127_407 ();
 FILLER_ASAP7_75t_R FILLER_0_127_415 ();
 FILLER_ASAP7_75t_R FILLER_0_127_425 ();
 FILLER_ASAP7_75t_R FILLER_0_127_432 ();
 DECAPx4_ASAP7_75t_R FILLER_0_127_437 ();
 FILLER_ASAP7_75t_R FILLER_0_127_447 ();
 DECAPx6_ASAP7_75t_R FILLER_0_127_457 ();
 FILLER_ASAP7_75t_R FILLER_0_127_471 ();
 DECAPx2_ASAP7_75t_R FILLER_0_127_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_482 ();
 DECAPx2_ASAP7_75t_R FILLER_0_127_489 ();
 FILLER_ASAP7_75t_R FILLER_0_127_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_497 ();
 DECAPx2_ASAP7_75t_R FILLER_0_127_506 ();
 DECAPx2_ASAP7_75t_R FILLER_0_127_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_522 ();
 FILLER_ASAP7_75t_R FILLER_0_127_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_531 ();
 DECAPx1_ASAP7_75t_R FILLER_0_127_538 ();
 DECAPx1_ASAP7_75t_R FILLER_0_127_548 ();
 DECAPx1_ASAP7_75t_R FILLER_0_127_558 ();
 FILLER_ASAP7_75t_R FILLER_0_127_565 ();
 DECAPx1_ASAP7_75t_R FILLER_0_127_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_578 ();
 FILLER_ASAP7_75t_R FILLER_0_127_586 ();
 DECAPx1_ASAP7_75t_R FILLER_0_127_599 ();
 DECAPx2_ASAP7_75t_R FILLER_0_127_613 ();
 FILLER_ASAP7_75t_R FILLER_0_127_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_621 ();
 DECAPx4_ASAP7_75t_R FILLER_0_127_628 ();
 FILLER_ASAP7_75t_R FILLER_0_127_644 ();
 FILLER_ASAP7_75t_R FILLER_0_127_656 ();
 DECAPx4_ASAP7_75t_R FILLER_0_127_664 ();
 FILLER_ASAP7_75t_R FILLER_0_127_677 ();
 DECAPx1_ASAP7_75t_R FILLER_0_127_691 ();
 DECAPx6_ASAP7_75t_R FILLER_0_127_701 ();
 DECAPx2_ASAP7_75t_R FILLER_0_127_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_721 ();
 FILLER_ASAP7_75t_R FILLER_0_127_732 ();
 FILLER_ASAP7_75t_R FILLER_0_127_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_739 ();
 FILLER_ASAP7_75t_R FILLER_0_127_746 ();
 DECAPx2_ASAP7_75t_R FILLER_0_127_754 ();
 FILLER_ASAP7_75t_R FILLER_0_127_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_762 ();
 DECAPx4_ASAP7_75t_R FILLER_0_127_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_779 ();
 FILLER_ASAP7_75t_R FILLER_0_127_786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_793 ();
 DECAPx4_ASAP7_75t_R FILLER_0_127_815 ();
 FILLER_ASAP7_75t_R FILLER_0_127_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_827 ();
 FILLER_ASAP7_75t_R FILLER_0_127_838 ();
 FILLER_ASAP7_75t_R FILLER_0_127_844 ();
 FILLER_ASAP7_75t_R FILLER_0_127_852 ();
 DECAPx2_ASAP7_75t_R FILLER_0_127_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_866 ();
 FILLER_ASAP7_75t_R FILLER_0_127_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_875 ();
 FILLER_ASAP7_75t_R FILLER_0_127_886 ();
 FILLER_ASAP7_75t_R FILLER_0_127_894 ();
 FILLER_ASAP7_75t_R FILLER_0_127_901 ();
 DECAPx1_ASAP7_75t_R FILLER_0_127_909 ();
 DECAPx2_ASAP7_75t_R FILLER_0_127_919 ();
 DECAPx4_ASAP7_75t_R FILLER_0_127_927 ();
 FILLER_ASAP7_75t_R FILLER_0_127_948 ();
 DECAPx1_ASAP7_75t_R FILLER_0_127_953 ();
 DECAPx1_ASAP7_75t_R FILLER_0_127_965 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_975 ();
 FILLER_ASAP7_75t_R FILLER_0_127_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_999 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_1011 ();
 DECAPx4_ASAP7_75t_R FILLER_0_127_1033 ();
 FILLER_ASAP7_75t_R FILLER_0_127_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_1045 ();
 FILLER_ASAP7_75t_R FILLER_0_127_1058 ();
 DECAPx1_ASAP7_75t_R FILLER_0_127_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_1067 ();
 DECAPx6_ASAP7_75t_R FILLER_0_127_1076 ();
 FILLER_ASAP7_75t_R FILLER_0_127_1090 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_1092 ();
 FILLER_ASAP7_75t_R FILLER_0_127_1103 ();
 FILLER_ASAP7_75t_R FILLER_0_127_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_1137 ();
 FILLER_ASAP7_75t_R FILLER_0_127_1159 ();
 DECAPx2_ASAP7_75t_R FILLER_0_127_1171 ();
 FILLER_ASAP7_75t_R FILLER_0_127_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_1179 ();
 DECAPx1_ASAP7_75t_R FILLER_0_127_1190 ();
 FILLER_ASAP7_75t_R FILLER_0_127_1199 ();
 DECAPx1_ASAP7_75t_R FILLER_0_127_1207 ();
 FILLER_ASAP7_75t_R FILLER_0_127_1219 ();
 DECAPx1_ASAP7_75t_R FILLER_0_127_1227 ();
 DECAPx4_ASAP7_75t_R FILLER_0_127_1241 ();
 FILLER_ASAP7_75t_R FILLER_0_127_1251 ();
 FILLER_ASAP7_75t_R FILLER_0_127_1259 ();
 FILLER_ASAP7_75t_R FILLER_0_127_1271 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_1273 ();
 DECAPx1_ASAP7_75t_R FILLER_0_127_1284 ();
 DECAPx2_ASAP7_75t_R FILLER_0_127_1308 ();
 FILLER_ASAP7_75t_R FILLER_0_127_1321 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_1323 ();
 DECAPx2_ASAP7_75t_R FILLER_0_127_1335 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_1341 ();
 DECAPx2_ASAP7_75t_R FILLER_0_127_1345 ();
 FILLER_ASAP7_75t_R FILLER_0_127_1356 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_127_1358 ();
 FILLER_ASAP7_75t_R FILLER_0_127_1364 ();
 DECAPx1_ASAP7_75t_R FILLER_0_127_1371 ();
 FILLER_ASAP7_75t_R FILLER_0_127_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_128_2 ();
 FILLER_ASAP7_75t_R FILLER_0_128_9 ();
 FILLER_ASAP7_75t_R FILLER_0_128_16 ();
 FILLER_ASAP7_75t_R FILLER_0_128_23 ();
 FILLER_ASAP7_75t_R FILLER_0_128_30 ();
 FILLER_ASAP7_75t_R FILLER_0_128_37 ();
 FILLER_ASAP7_75t_R FILLER_0_128_44 ();
 FILLER_ASAP7_75t_R FILLER_0_128_49 ();
 DECAPx4_ASAP7_75t_R FILLER_0_128_54 ();
 FILLER_ASAP7_75t_R FILLER_0_128_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_66 ();
 FILLER_ASAP7_75t_R FILLER_0_128_77 ();
 DECAPx6_ASAP7_75t_R FILLER_0_128_83 ();
 DECAPx1_ASAP7_75t_R FILLER_0_128_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_101 ();
 FILLER_ASAP7_75t_R FILLER_0_128_123 ();
 FILLER_ASAP7_75t_R FILLER_0_128_131 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_136 ();
 FILLER_ASAP7_75t_R FILLER_0_128_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_160 ();
 DECAPx1_ASAP7_75t_R FILLER_0_128_167 ();
 FILLER_ASAP7_75t_R FILLER_0_128_177 ();
 FILLER_ASAP7_75t_R FILLER_0_128_199 ();
 FILLER_ASAP7_75t_R FILLER_0_128_206 ();
 DECAPx2_ASAP7_75t_R FILLER_0_128_213 ();
 FILLER_ASAP7_75t_R FILLER_0_128_222 ();
 FILLER_ASAP7_75t_R FILLER_0_128_232 ();
 FILLER_ASAP7_75t_R FILLER_0_128_244 ();
 FILLER_ASAP7_75t_R FILLER_0_128_256 ();
 DECAPx4_ASAP7_75t_R FILLER_0_128_265 ();
 FILLER_ASAP7_75t_R FILLER_0_128_283 ();
 DECAPx4_ASAP7_75t_R FILLER_0_128_293 ();
 FILLER_ASAP7_75t_R FILLER_0_128_303 ();
 FILLER_ASAP7_75t_R FILLER_0_128_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_317 ();
 DECAPx2_ASAP7_75t_R FILLER_0_128_328 ();
 FILLER_ASAP7_75t_R FILLER_0_128_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_336 ();
 DECAPx1_ASAP7_75t_R FILLER_0_128_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_351 ();
 FILLER_ASAP7_75t_R FILLER_0_128_358 ();
 DECAPx1_ASAP7_75t_R FILLER_0_128_363 ();
 DECAPx4_ASAP7_75t_R FILLER_0_128_373 ();
 FILLER_ASAP7_75t_R FILLER_0_128_389 ();
 FILLER_ASAP7_75t_R FILLER_0_128_396 ();
 DECAPx1_ASAP7_75t_R FILLER_0_128_401 ();
 FILLER_ASAP7_75t_R FILLER_0_128_413 ();
 FILLER_ASAP7_75t_R FILLER_0_128_423 ();
 DECAPx2_ASAP7_75t_R FILLER_0_128_428 ();
 FILLER_ASAP7_75t_R FILLER_0_128_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_436 ();
 FILLER_ASAP7_75t_R FILLER_0_128_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_446 ();
 DECAPx2_ASAP7_75t_R FILLER_0_128_453 ();
 FILLER_ASAP7_75t_R FILLER_0_128_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_461 ();
 DECAPx2_ASAP7_75t_R FILLER_0_128_464 ();
 FILLER_ASAP7_75t_R FILLER_0_128_470 ();
 DECAPx4_ASAP7_75t_R FILLER_0_128_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_488 ();
 DECAPx4_ASAP7_75t_R FILLER_0_128_495 ();
 FILLER_ASAP7_75t_R FILLER_0_128_505 ();
 DECAPx2_ASAP7_75t_R FILLER_0_128_513 ();
 FILLER_ASAP7_75t_R FILLER_0_128_519 ();
 FILLER_ASAP7_75t_R FILLER_0_128_527 ();
 FILLER_ASAP7_75t_R FILLER_0_128_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_537 ();
 DECAPx2_ASAP7_75t_R FILLER_0_128_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_548 ();
 DECAPx4_ASAP7_75t_R FILLER_0_128_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_571 ();
 FILLER_ASAP7_75t_R FILLER_0_128_584 ();
 FILLER_ASAP7_75t_R FILLER_0_128_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_594 ();
 DECAPx2_ASAP7_75t_R FILLER_0_128_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_607 ();
 DECAPx4_ASAP7_75t_R FILLER_0_128_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_624 ();
 DECAPx1_ASAP7_75t_R FILLER_0_128_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_635 ();
 FILLER_ASAP7_75t_R FILLER_0_128_642 ();
 FILLER_ASAP7_75t_R FILLER_0_128_656 ();
 DECAPx1_ASAP7_75t_R FILLER_0_128_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_670 ();
 DECAPx1_ASAP7_75t_R FILLER_0_128_681 ();
 DECAPx6_ASAP7_75t_R FILLER_0_128_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_713 ();
 DECAPx1_ASAP7_75t_R FILLER_0_128_722 ();
 FILLER_ASAP7_75t_R FILLER_0_128_731 ();
 DECAPx6_ASAP7_75t_R FILLER_0_128_753 ();
 DECAPx1_ASAP7_75t_R FILLER_0_128_767 ();
 FILLER_ASAP7_75t_R FILLER_0_128_776 ();
 DECAPx4_ASAP7_75t_R FILLER_0_128_790 ();
 FILLER_ASAP7_75t_R FILLER_0_128_800 ();
 FILLER_ASAP7_75t_R FILLER_0_128_808 ();
 FILLER_ASAP7_75t_R FILLER_0_128_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_818 ();
 DECAPx2_ASAP7_75t_R FILLER_0_128_825 ();
 FILLER_ASAP7_75t_R FILLER_0_128_831 ();
 DECAPx2_ASAP7_75t_R FILLER_0_128_840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_854 ();
 DECAPx2_ASAP7_75t_R FILLER_0_128_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_889 ();
 FILLER_ASAP7_75t_R FILLER_0_128_896 ();
 FILLER_ASAP7_75t_R FILLER_0_128_904 ();
 FILLER_ASAP7_75t_R FILLER_0_128_912 ();
 FILLER_ASAP7_75t_R FILLER_0_128_920 ();
 FILLER_ASAP7_75t_R FILLER_0_128_928 ();
 DECAPx2_ASAP7_75t_R FILLER_0_128_934 ();
 FILLER_ASAP7_75t_R FILLER_0_128_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_942 ();
 FILLER_ASAP7_75t_R FILLER_0_128_947 ();
 FILLER_ASAP7_75t_R FILLER_0_128_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_959 ();
 DECAPx6_ASAP7_75t_R FILLER_0_128_963 ();
 DECAPx1_ASAP7_75t_R FILLER_0_128_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_981 ();
 FILLER_ASAP7_75t_R FILLER_0_128_990 ();
 DECAPx2_ASAP7_75t_R FILLER_0_128_995 ();
 FILLER_ASAP7_75t_R FILLER_0_128_1007 ();
 FILLER_ASAP7_75t_R FILLER_0_128_1017 ();
 DECAPx1_ASAP7_75t_R FILLER_0_128_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_1035 ();
 DECAPx4_ASAP7_75t_R FILLER_0_128_1048 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_1058 ();
 FILLER_ASAP7_75t_R FILLER_0_128_1067 ();
 FILLER_ASAP7_75t_R FILLER_0_128_1075 ();
 DECAPx6_ASAP7_75t_R FILLER_0_128_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_0_128_1103 ();
 DECAPx1_ASAP7_75t_R FILLER_0_128_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_1117 ();
 DECAPx4_ASAP7_75t_R FILLER_0_128_1138 ();
 FILLER_ASAP7_75t_R FILLER_0_128_1148 ();
 FILLER_ASAP7_75t_R FILLER_0_128_1160 ();
 FILLER_ASAP7_75t_R FILLER_0_128_1172 ();
 DECAPx4_ASAP7_75t_R FILLER_0_128_1184 ();
 FILLER_ASAP7_75t_R FILLER_0_128_1200 ();
 FILLER_ASAP7_75t_R FILLER_0_128_1208 ();
 FILLER_ASAP7_75t_R FILLER_0_128_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_1224 ();
 DECAPx2_ASAP7_75t_R FILLER_0_128_1246 ();
 DECAPx2_ASAP7_75t_R FILLER_0_128_1258 ();
 FILLER_ASAP7_75t_R FILLER_0_128_1270 ();
 DECAPx6_ASAP7_75t_R FILLER_0_128_1278 ();
 FILLER_ASAP7_75t_R FILLER_0_128_1302 ();
 DECAPx1_ASAP7_75t_R FILLER_0_128_1310 ();
 DECAPx6_ASAP7_75t_R FILLER_0_128_1324 ();
 DECAPx1_ASAP7_75t_R FILLER_0_128_1338 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_1342 ();
 FILLER_ASAP7_75t_R FILLER_0_128_1346 ();
 FILLER_ASAP7_75t_R FILLER_0_128_1369 ();
 DECAPx2_ASAP7_75t_R FILLER_0_128_1376 ();
 FILLER_ASAP7_75t_R FILLER_0_129_2 ();
 FILLER_ASAP7_75t_R FILLER_0_129_25 ();
 FILLER_ASAP7_75t_R FILLER_0_129_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_34 ();
 FILLER_ASAP7_75t_R FILLER_0_129_40 ();
 FILLER_ASAP7_75t_R FILLER_0_129_47 ();
 DECAPx6_ASAP7_75t_R FILLER_0_129_52 ();
 DECAPx1_ASAP7_75t_R FILLER_0_129_66 ();
 DECAPx6_ASAP7_75t_R FILLER_0_129_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_94 ();
 FILLER_ASAP7_75t_R FILLER_0_129_107 ();
 DECAPx4_ASAP7_75t_R FILLER_0_129_112 ();
 FILLER_ASAP7_75t_R FILLER_0_129_122 ();
 FILLER_ASAP7_75t_R FILLER_0_129_130 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_140 ();
 FILLER_ASAP7_75t_R FILLER_0_129_162 ();
 FILLER_ASAP7_75t_R FILLER_0_129_185 ();
 FILLER_ASAP7_75t_R FILLER_0_129_197 ();
 FILLER_ASAP7_75t_R FILLER_0_129_210 ();
 DECAPx1_ASAP7_75t_R FILLER_0_129_218 ();
 DECAPx2_ASAP7_75t_R FILLER_0_129_230 ();
 DECAPx1_ASAP7_75t_R FILLER_0_129_247 ();
 DECAPx2_ASAP7_75t_R FILLER_0_129_263 ();
 DECAPx1_ASAP7_75t_R FILLER_0_129_275 ();
 FILLER_ASAP7_75t_R FILLER_0_129_287 ();
 DECAPx4_ASAP7_75t_R FILLER_0_129_297 ();
 FILLER_ASAP7_75t_R FILLER_0_129_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_309 ();
 FILLER_ASAP7_75t_R FILLER_0_129_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_317 ();
 FILLER_ASAP7_75t_R FILLER_0_129_328 ();
 FILLER_ASAP7_75t_R FILLER_0_129_354 ();
 FILLER_ASAP7_75t_R FILLER_0_129_362 ();
 DECAPx6_ASAP7_75t_R FILLER_0_129_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_381 ();
 DECAPx2_ASAP7_75t_R FILLER_0_129_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_396 ();
 FILLER_ASAP7_75t_R FILLER_0_129_403 ();
 DECAPx4_ASAP7_75t_R FILLER_0_129_408 ();
 FILLER_ASAP7_75t_R FILLER_0_129_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_441 ();
 FILLER_ASAP7_75t_R FILLER_0_129_463 ();
 FILLER_ASAP7_75t_R FILLER_0_129_472 ();
 DECAPx2_ASAP7_75t_R FILLER_0_129_480 ();
 FILLER_ASAP7_75t_R FILLER_0_129_486 ();
 FILLER_ASAP7_75t_R FILLER_0_129_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_496 ();
 DECAPx1_ASAP7_75t_R FILLER_0_129_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_521 ();
 DECAPx4_ASAP7_75t_R FILLER_0_129_529 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_559 ();
 DECAPx6_ASAP7_75t_R FILLER_0_129_581 ();
 FILLER_ASAP7_75t_R FILLER_0_129_595 ();
 FILLER_ASAP7_75t_R FILLER_0_129_603 ();
 DECAPx4_ASAP7_75t_R FILLER_0_129_611 ();
 DECAPx2_ASAP7_75t_R FILLER_0_129_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_634 ();
 DECAPx4_ASAP7_75t_R FILLER_0_129_641 ();
 FILLER_ASAP7_75t_R FILLER_0_129_651 ();
 FILLER_ASAP7_75t_R FILLER_0_129_673 ();
 DECAPx2_ASAP7_75t_R FILLER_0_129_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_684 ();
 FILLER_ASAP7_75t_R FILLER_0_129_705 ();
 DECAPx6_ASAP7_75t_R FILLER_0_129_713 ();
 DECAPx2_ASAP7_75t_R FILLER_0_129_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_733 ();
 FILLER_ASAP7_75t_R FILLER_0_129_742 ();
 FILLER_ASAP7_75t_R FILLER_0_129_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_751 ();
 DECAPx2_ASAP7_75t_R FILLER_0_129_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_764 ();
 DECAPx4_ASAP7_75t_R FILLER_0_129_771 ();
 FILLER_ASAP7_75t_R FILLER_0_129_781 ();
 DECAPx2_ASAP7_75t_R FILLER_0_129_789 ();
 FILLER_ASAP7_75t_R FILLER_0_129_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_797 ();
 FILLER_ASAP7_75t_R FILLER_0_129_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_806 ();
 DECAPx2_ASAP7_75t_R FILLER_0_129_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_819 ();
 DECAPx2_ASAP7_75t_R FILLER_0_129_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_836 ();
 DECAPx2_ASAP7_75t_R FILLER_0_129_843 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_855 ();
 DECAPx6_ASAP7_75t_R FILLER_0_129_877 ();
 DECAPx1_ASAP7_75t_R FILLER_0_129_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_895 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_903 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_927 ();
 DECAPx4_ASAP7_75t_R FILLER_0_129_949 ();
 FILLER_ASAP7_75t_R FILLER_0_129_959 ();
 DECAPx1_ASAP7_75t_R FILLER_0_129_967 ();
 FILLER_ASAP7_75t_R FILLER_0_129_983 ();
 DECAPx1_ASAP7_75t_R FILLER_0_129_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_995 ();
 FILLER_ASAP7_75t_R FILLER_0_129_1006 ();
 DECAPx4_ASAP7_75t_R FILLER_0_129_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_1039 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_1046 ();
 DECAPx1_ASAP7_75t_R FILLER_0_129_1068 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_1084 ();
 DECAPx6_ASAP7_75t_R FILLER_0_129_1106 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_1120 ();
 FILLER_ASAP7_75t_R FILLER_0_129_1126 ();
 DECAPx6_ASAP7_75t_R FILLER_0_129_1135 ();
 DECAPx1_ASAP7_75t_R FILLER_0_129_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_1153 ();
 DECAPx2_ASAP7_75t_R FILLER_0_129_1160 ();
 FILLER_ASAP7_75t_R FILLER_0_129_1166 ();
 FILLER_ASAP7_75t_R FILLER_0_129_1173 ();
 DECAPx2_ASAP7_75t_R FILLER_0_129_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_1184 ();
 FILLER_ASAP7_75t_R FILLER_0_129_1195 ();
 DECAPx4_ASAP7_75t_R FILLER_0_129_1203 ();
 FILLER_ASAP7_75t_R FILLER_0_129_1213 ();
 DECAPx2_ASAP7_75t_R FILLER_0_129_1225 ();
 FILLER_ASAP7_75t_R FILLER_0_129_1231 ();
 DECAPx2_ASAP7_75t_R FILLER_0_129_1239 ();
 FILLER_ASAP7_75t_R FILLER_0_129_1245 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_1247 ();
 FILLER_ASAP7_75t_R FILLER_0_129_1254 ();
 DECAPx1_ASAP7_75t_R FILLER_0_129_1262 ();
 DECAPx6_ASAP7_75t_R FILLER_0_129_1272 ();
 FILLER_ASAP7_75t_R FILLER_0_129_1286 ();
 FILLER_ASAP7_75t_R FILLER_0_129_1308 ();
 FILLER_ASAP7_75t_R FILLER_0_129_1322 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_1324 ();
 FILLER_ASAP7_75t_R FILLER_0_129_1331 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_1333 ();
 FILLER_ASAP7_75t_R FILLER_0_129_1337 ();
 FILLER_ASAP7_75t_R FILLER_0_129_1342 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_1344 ();
 FILLER_ASAP7_75t_R FILLER_0_129_1350 ();
 FILLER_ASAP7_75t_R FILLER_0_129_1358 ();
 FILLER_ASAP7_75t_R FILLER_0_129_1366 ();
 FILLER_ASAP7_75t_R FILLER_0_129_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_129_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_130_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_130_10 ();
 FILLER_ASAP7_75t_R FILLER_0_130_22 ();
 FILLER_ASAP7_75t_R FILLER_0_130_46 ();
 DECAPx2_ASAP7_75t_R FILLER_0_130_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_60 ();
 DECAPx2_ASAP7_75t_R FILLER_0_130_67 ();
 FILLER_ASAP7_75t_R FILLER_0_130_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_75 ();
 DECAPx2_ASAP7_75t_R FILLER_0_130_88 ();
 DECAPx4_ASAP7_75t_R FILLER_0_130_102 ();
 FILLER_ASAP7_75t_R FILLER_0_130_112 ();
 DECAPx6_ASAP7_75t_R FILLER_0_130_120 ();
 DECAPx1_ASAP7_75t_R FILLER_0_130_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_138 ();
 FILLER_ASAP7_75t_R FILLER_0_130_147 ();
 DECAPx4_ASAP7_75t_R FILLER_0_130_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_165 ();
 DECAPx4_ASAP7_75t_R FILLER_0_130_169 ();
 FILLER_ASAP7_75t_R FILLER_0_130_179 ();
 FILLER_ASAP7_75t_R FILLER_0_130_191 ();
 FILLER_ASAP7_75t_R FILLER_0_130_197 ();
 DECAPx4_ASAP7_75t_R FILLER_0_130_207 ();
 FILLER_ASAP7_75t_R FILLER_0_130_223 ();
 DECAPx6_ASAP7_75t_R FILLER_0_130_231 ();
 FILLER_ASAP7_75t_R FILLER_0_130_245 ();
 DECAPx6_ASAP7_75t_R FILLER_0_130_255 ();
 FILLER_ASAP7_75t_R FILLER_0_130_269 ();
 FILLER_ASAP7_75t_R FILLER_0_130_277 ();
 DECAPx4_ASAP7_75t_R FILLER_0_130_287 ();
 FILLER_ASAP7_75t_R FILLER_0_130_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_299 ();
 FILLER_ASAP7_75t_R FILLER_0_130_304 ();
 FILLER_ASAP7_75t_R FILLER_0_130_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_318 ();
 DECAPx2_ASAP7_75t_R FILLER_0_130_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_335 ();
 FILLER_ASAP7_75t_R FILLER_0_130_344 ();
 FILLER_ASAP7_75t_R FILLER_0_130_349 ();
 FILLER_ASAP7_75t_R FILLER_0_130_357 ();
 FILLER_ASAP7_75t_R FILLER_0_130_365 ();
 DECAPx2_ASAP7_75t_R FILLER_0_130_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_382 ();
 DECAPx1_ASAP7_75t_R FILLER_0_130_393 ();
 FILLER_ASAP7_75t_R FILLER_0_130_405 ();
 FILLER_ASAP7_75t_R FILLER_0_130_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_415 ();
 DECAPx4_ASAP7_75t_R FILLER_0_130_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_429 ();
 FILLER_ASAP7_75t_R FILLER_0_130_438 ();
 DECAPx6_ASAP7_75t_R FILLER_0_130_445 ();
 FILLER_ASAP7_75t_R FILLER_0_130_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_461 ();
 DECAPx2_ASAP7_75t_R FILLER_0_130_464 ();
 FILLER_ASAP7_75t_R FILLER_0_130_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_472 ();
 DECAPx1_ASAP7_75t_R FILLER_0_130_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_487 ();
 FILLER_ASAP7_75t_R FILLER_0_130_494 ();
 DECAPx1_ASAP7_75t_R FILLER_0_130_502 ();
 DECAPx4_ASAP7_75t_R FILLER_0_130_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_519 ();
 DECAPx2_ASAP7_75t_R FILLER_0_130_526 ();
 FILLER_ASAP7_75t_R FILLER_0_130_538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_568 ();
 DECAPx2_ASAP7_75t_R FILLER_0_130_577 ();
 FILLER_ASAP7_75t_R FILLER_0_130_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_585 ();
 FILLER_ASAP7_75t_R FILLER_0_130_592 ();
 FILLER_ASAP7_75t_R FILLER_0_130_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_607 ();
 DECAPx2_ASAP7_75t_R FILLER_0_130_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_620 ();
 FILLER_ASAP7_75t_R FILLER_0_130_627 ();
 DECAPx6_ASAP7_75t_R FILLER_0_130_635 ();
 DECAPx1_ASAP7_75t_R FILLER_0_130_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_653 ();
 FILLER_ASAP7_75t_R FILLER_0_130_659 ();
 FILLER_ASAP7_75t_R FILLER_0_130_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_666 ();
 DECAPx1_ASAP7_75t_R FILLER_0_130_677 ();
 FILLER_ASAP7_75t_R FILLER_0_130_693 ();
 DECAPx1_ASAP7_75t_R FILLER_0_130_700 ();
 DECAPx6_ASAP7_75t_R FILLER_0_130_710 ();
 DECAPx2_ASAP7_75t_R FILLER_0_130_724 ();
 FILLER_ASAP7_75t_R FILLER_0_130_736 ();
 DECAPx2_ASAP7_75t_R FILLER_0_130_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_749 ();
 DECAPx2_ASAP7_75t_R FILLER_0_130_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_763 ();
 DECAPx2_ASAP7_75t_R FILLER_0_130_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_776 ();
 DECAPx4_ASAP7_75t_R FILLER_0_130_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_798 ();
 DECAPx1_ASAP7_75t_R FILLER_0_130_805 ();
 FILLER_ASAP7_75t_R FILLER_0_130_816 ();
 DECAPx2_ASAP7_75t_R FILLER_0_130_823 ();
 FILLER_ASAP7_75t_R FILLER_0_130_829 ();
 FILLER_ASAP7_75t_R FILLER_0_130_837 ();
 DECAPx2_ASAP7_75t_R FILLER_0_130_844 ();
 DECAPx6_ASAP7_75t_R FILLER_0_130_856 ();
 FILLER_ASAP7_75t_R FILLER_0_130_870 ();
 FILLER_ASAP7_75t_R FILLER_0_130_878 ();
 DECAPx6_ASAP7_75t_R FILLER_0_130_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_899 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_906 ();
 FILLER_ASAP7_75t_R FILLER_0_130_939 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_944 ();
 FILLER_ASAP7_75t_R FILLER_0_130_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_980 ();
 DECAPx4_ASAP7_75t_R FILLER_0_130_985 ();
 FILLER_ASAP7_75t_R FILLER_0_130_995 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_997 ();
 DECAPx1_ASAP7_75t_R FILLER_0_130_1006 ();
 DECAPx6_ASAP7_75t_R FILLER_0_130_1013 ();
 DECAPx1_ASAP7_75t_R FILLER_0_130_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_1031 ();
 FILLER_ASAP7_75t_R FILLER_0_130_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_1040 ();
 FILLER_ASAP7_75t_R FILLER_0_130_1048 ();
 DECAPx2_ASAP7_75t_R FILLER_0_130_1054 ();
 FILLER_ASAP7_75t_R FILLER_0_130_1066 ();
 FILLER_ASAP7_75t_R FILLER_0_130_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_1076 ();
 FILLER_ASAP7_75t_R FILLER_0_130_1084 ();
 FILLER_ASAP7_75t_R FILLER_0_130_1096 ();
 DECAPx4_ASAP7_75t_R FILLER_0_130_1108 ();
 FILLER_ASAP7_75t_R FILLER_0_130_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_1120 ();
 FILLER_ASAP7_75t_R FILLER_0_130_1127 ();
 FILLER_ASAP7_75t_R FILLER_0_130_1139 ();
 FILLER_ASAP7_75t_R FILLER_0_130_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_1153 ();
 FILLER_ASAP7_75t_R FILLER_0_130_1166 ();
 FILLER_ASAP7_75t_R FILLER_0_130_1178 ();
 DECAPx1_ASAP7_75t_R FILLER_0_130_1190 ();
 DECAPx4_ASAP7_75t_R FILLER_0_130_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_1214 ();
 DECAPx1_ASAP7_75t_R FILLER_0_130_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_1225 ();
 FILLER_ASAP7_75t_R FILLER_0_130_1236 ();
 FILLER_ASAP7_75t_R FILLER_0_130_1244 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_1246 ();
 FILLER_ASAP7_75t_R FILLER_0_130_1257 ();
 DECAPx1_ASAP7_75t_R FILLER_0_130_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_1273 ();
 DECAPx4_ASAP7_75t_R FILLER_0_130_1284 ();
 DECAPx4_ASAP7_75t_R FILLER_0_130_1304 ();
 FILLER_ASAP7_75t_R FILLER_0_130_1320 ();
 DECAPx2_ASAP7_75t_R FILLER_0_130_1328 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_1334 ();
 DECAPx2_ASAP7_75t_R FILLER_0_130_1341 ();
 FILLER_ASAP7_75t_R FILLER_0_130_1352 ();
 FILLER_ASAP7_75t_R FILLER_0_130_1359 ();
 FILLER_ASAP7_75t_R FILLER_0_130_1367 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_1369 ();
 FILLER_ASAP7_75t_R FILLER_0_130_1375 ();
 FILLER_ASAP7_75t_R FILLER_0_130_1380 ();
 DECAPx2_ASAP7_75t_R FILLER_0_131_2 ();
 FILLER_ASAP7_75t_R FILLER_0_131_13 ();
 DECAPx2_ASAP7_75t_R FILLER_0_131_20 ();
 FILLER_ASAP7_75t_R FILLER_0_131_32 ();
 FILLER_ASAP7_75t_R FILLER_0_131_55 ();
 FILLER_ASAP7_75t_R FILLER_0_131_60 ();
 DECAPx2_ASAP7_75t_R FILLER_0_131_65 ();
 FILLER_ASAP7_75t_R FILLER_0_131_71 ();
 FILLER_ASAP7_75t_R FILLER_0_131_79 ();
 DECAPx2_ASAP7_75t_R FILLER_0_131_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_131_93 ();
 DECAPx6_ASAP7_75t_R FILLER_0_131_100 ();
 DECAPx1_ASAP7_75t_R FILLER_0_131_114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_124 ();
 DECAPx2_ASAP7_75t_R FILLER_0_131_146 ();
 FILLER_ASAP7_75t_R FILLER_0_131_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_131_154 ();
 FILLER_ASAP7_75t_R FILLER_0_131_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_131_167 ();
 FILLER_ASAP7_75t_R FILLER_0_131_188 ();
 DECAPx1_ASAP7_75t_R FILLER_0_131_200 ();
 DECAPx4_ASAP7_75t_R FILLER_0_131_210 ();
 FILLER_ASAP7_75t_R FILLER_0_131_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_131_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_229 ();
 DECAPx1_ASAP7_75t_R FILLER_0_131_251 ();
 DECAPx4_ASAP7_75t_R FILLER_0_131_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_131_268 ();
 FILLER_ASAP7_75t_R FILLER_0_131_273 ();
 FILLER_ASAP7_75t_R FILLER_0_131_285 ();
 DECAPx6_ASAP7_75t_R FILLER_0_131_295 ();
 FILLER_ASAP7_75t_R FILLER_0_131_309 ();
 FILLER_ASAP7_75t_R FILLER_0_131_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_131_323 ();
 FILLER_ASAP7_75t_R FILLER_0_131_334 ();
 DECAPx1_ASAP7_75t_R FILLER_0_131_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_131_346 ();
 FILLER_ASAP7_75t_R FILLER_0_131_353 ();
 FILLER_ASAP7_75t_R FILLER_0_131_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_131_363 ();
 DECAPx4_ASAP7_75t_R FILLER_0_131_371 ();
 FILLER_ASAP7_75t_R FILLER_0_131_386 ();
 DECAPx4_ASAP7_75t_R FILLER_0_131_394 ();
 FILLER_ASAP7_75t_R FILLER_0_131_411 ();
 DECAPx4_ASAP7_75t_R FILLER_0_131_419 ();
 FILLER_ASAP7_75t_R FILLER_0_131_435 ();
 FILLER_ASAP7_75t_R FILLER_0_131_443 ();
 FILLER_ASAP7_75t_R FILLER_0_131_454 ();
 FILLER_ASAP7_75t_R FILLER_0_131_466 ();
 DECAPx4_ASAP7_75t_R FILLER_0_131_475 ();
 FILLER_ASAP7_75t_R FILLER_0_131_485 ();
 FILLER_ASAP7_75t_R FILLER_0_131_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_131_495 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_504 ();
 DECAPx4_ASAP7_75t_R FILLER_0_131_526 ();
 FILLER_ASAP7_75t_R FILLER_0_131_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_131_538 ();
 DECAPx2_ASAP7_75t_R FILLER_0_131_545 ();
 DECAPx4_ASAP7_75t_R FILLER_0_131_561 ();
 DECAPx2_ASAP7_75t_R FILLER_0_131_581 ();
 DECAPx1_ASAP7_75t_R FILLER_0_131_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_131_598 ();
 FILLER_ASAP7_75t_R FILLER_0_131_610 ();
 FILLER_ASAP7_75t_R FILLER_0_131_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_631 ();
 FILLER_ASAP7_75t_R FILLER_0_131_663 ();
 DECAPx1_ASAP7_75t_R FILLER_0_131_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_131_672 ();
 FILLER_ASAP7_75t_R FILLER_0_131_693 ();
 FILLER_ASAP7_75t_R FILLER_0_131_698 ();
 FILLER_ASAP7_75t_R FILLER_0_131_706 ();
 DECAPx4_ASAP7_75t_R FILLER_0_131_714 ();
 FILLER_ASAP7_75t_R FILLER_0_131_724 ();
 DECAPx1_ASAP7_75t_R FILLER_0_131_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_131_750 ();
 FILLER_ASAP7_75t_R FILLER_0_131_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_131_759 ();
 DECAPx2_ASAP7_75t_R FILLER_0_131_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_131_772 ();
 DECAPx6_ASAP7_75t_R FILLER_0_131_779 ();
 DECAPx2_ASAP7_75t_R FILLER_0_131_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_131_799 ();
 FILLER_ASAP7_75t_R FILLER_0_131_806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_131_813 ();
 FILLER_ASAP7_75t_R FILLER_0_131_832 ();
 DECAPx4_ASAP7_75t_R FILLER_0_131_840 ();
 FILLER_ASAP7_75t_R FILLER_0_131_850 ();
 FILLER_ASAP7_75t_R FILLER_0_131_858 ();
 FILLER_ASAP7_75t_R FILLER_0_131_872 ();
 FILLER_ASAP7_75t_R FILLER_0_131_880 ();
 DECAPx1_ASAP7_75t_R FILLER_0_131_888 ();
 FILLER_ASAP7_75t_R FILLER_0_131_898 ();
 DECAPx1_ASAP7_75t_R FILLER_0_131_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_131_924 ();
 FILLER_ASAP7_75t_R FILLER_0_131_927 ();
 FILLER_ASAP7_75t_R FILLER_0_131_932 ();
 FILLER_ASAP7_75t_R FILLER_0_131_942 ();
 FILLER_ASAP7_75t_R FILLER_0_131_947 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_131_949 ();
 FILLER_ASAP7_75t_R FILLER_0_131_971 ();
 FILLER_ASAP7_75t_R FILLER_0_131_985 ();
 FILLER_ASAP7_75t_R FILLER_0_131_997 ();
 DECAPx4_ASAP7_75t_R FILLER_0_131_1009 ();
 DECAPx4_ASAP7_75t_R FILLER_0_131_1029 ();
 FILLER_ASAP7_75t_R FILLER_0_131_1039 ();
 DECAPx2_ASAP7_75t_R FILLER_0_131_1047 ();
 FILLER_ASAP7_75t_R FILLER_0_131_1053 ();
 FILLER_ASAP7_75t_R FILLER_0_131_1063 ();
 FILLER_ASAP7_75t_R FILLER_0_131_1071 ();
 DECAPx1_ASAP7_75t_R FILLER_0_131_1076 ();
 DECAPx4_ASAP7_75t_R FILLER_0_131_1090 ();
 FILLER_ASAP7_75t_R FILLER_0_131_1100 ();
 DECAPx2_ASAP7_75t_R FILLER_0_131_1123 ();
 DECAPx2_ASAP7_75t_R FILLER_0_131_1139 ();
 FILLER_ASAP7_75t_R FILLER_0_131_1145 ();
 FILLER_ASAP7_75t_R FILLER_0_131_1151 ();
 DECAPx2_ASAP7_75t_R FILLER_0_131_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_1179 ();
 DECAPx1_ASAP7_75t_R FILLER_0_131_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_131_1205 ();
 FILLER_ASAP7_75t_R FILLER_0_131_1212 ();
 DECAPx6_ASAP7_75t_R FILLER_0_131_1220 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_131_1234 ();
 FILLER_ASAP7_75t_R FILLER_0_131_1245 ();
 FILLER_ASAP7_75t_R FILLER_0_131_1257 ();
 FILLER_ASAP7_75t_R FILLER_0_131_1269 ();
 DECAPx1_ASAP7_75t_R FILLER_0_131_1281 ();
 DECAPx1_ASAP7_75t_R FILLER_0_131_1291 ();
 DECAPx2_ASAP7_75t_R FILLER_0_131_1305 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_131_1311 ();
 FILLER_ASAP7_75t_R FILLER_0_131_1318 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_131_1320 ();
 FILLER_ASAP7_75t_R FILLER_0_131_1327 ();
 DECAPx1_ASAP7_75t_R FILLER_0_131_1335 ();
 FILLER_ASAP7_75t_R FILLER_0_131_1350 ();
 FILLER_ASAP7_75t_R FILLER_0_131_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_131_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_132_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_132_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_13 ();
 DECAPx1_ASAP7_75t_R FILLER_0_132_19 ();
 FILLER_ASAP7_75t_R FILLER_0_132_45 ();
 FILLER_ASAP7_75t_R FILLER_0_132_50 ();
 FILLER_ASAP7_75t_R FILLER_0_132_55 ();
 DECAPx2_ASAP7_75t_R FILLER_0_132_60 ();
 DECAPx1_ASAP7_75t_R FILLER_0_132_69 ();
 DECAPx2_ASAP7_75t_R FILLER_0_132_81 ();
 FILLER_ASAP7_75t_R FILLER_0_132_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_89 ();
 FILLER_ASAP7_75t_R FILLER_0_132_98 ();
 FILLER_ASAP7_75t_R FILLER_0_132_112 ();
 FILLER_ASAP7_75t_R FILLER_0_132_125 ();
 FILLER_ASAP7_75t_R FILLER_0_132_135 ();
 DECAPx2_ASAP7_75t_R FILLER_0_132_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_155 ();
 DECAPx4_ASAP7_75t_R FILLER_0_132_162 ();
 FILLER_ASAP7_75t_R FILLER_0_132_172 ();
 DECAPx4_ASAP7_75t_R FILLER_0_132_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_190 ();
 FILLER_ASAP7_75t_R FILLER_0_132_197 ();
 DECAPx2_ASAP7_75t_R FILLER_0_132_210 ();
 FILLER_ASAP7_75t_R FILLER_0_132_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_218 ();
 DECAPx2_ASAP7_75t_R FILLER_0_132_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_237 ();
 FILLER_ASAP7_75t_R FILLER_0_132_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_246 ();
 FILLER_ASAP7_75t_R FILLER_0_132_253 ();
 DECAPx4_ASAP7_75t_R FILLER_0_132_263 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_283 ();
 DECAPx2_ASAP7_75t_R FILLER_0_132_305 ();
 FILLER_ASAP7_75t_R FILLER_0_132_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_318 ();
 FILLER_ASAP7_75t_R FILLER_0_132_324 ();
 DECAPx2_ASAP7_75t_R FILLER_0_132_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_340 ();
 FILLER_ASAP7_75t_R FILLER_0_132_348 ();
 DECAPx4_ASAP7_75t_R FILLER_0_132_356 ();
 FILLER_ASAP7_75t_R FILLER_0_132_366 ();
 FILLER_ASAP7_75t_R FILLER_0_132_374 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_384 ();
 FILLER_ASAP7_75t_R FILLER_0_132_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_408 ();
 DECAPx2_ASAP7_75t_R FILLER_0_132_415 ();
 FILLER_ASAP7_75t_R FILLER_0_132_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_429 ();
 FILLER_ASAP7_75t_R FILLER_0_132_440 ();
 FILLER_ASAP7_75t_R FILLER_0_132_448 ();
 FILLER_ASAP7_75t_R FILLER_0_132_460 ();
 FILLER_ASAP7_75t_R FILLER_0_132_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_466 ();
 FILLER_ASAP7_75t_R FILLER_0_132_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_489 ();
 DECAPx2_ASAP7_75t_R FILLER_0_132_500 ();
 FILLER_ASAP7_75t_R FILLER_0_132_506 ();
 FILLER_ASAP7_75t_R FILLER_0_132_518 ();
 FILLER_ASAP7_75t_R FILLER_0_132_526 ();
 DECAPx1_ASAP7_75t_R FILLER_0_132_534 ();
 FILLER_ASAP7_75t_R FILLER_0_132_544 ();
 DECAPx2_ASAP7_75t_R FILLER_0_132_556 ();
 FILLER_ASAP7_75t_R FILLER_0_132_562 ();
 FILLER_ASAP7_75t_R FILLER_0_132_584 ();
 DECAPx4_ASAP7_75t_R FILLER_0_132_592 ();
 DECAPx4_ASAP7_75t_R FILLER_0_132_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_618 ();
 DECAPx1_ASAP7_75t_R FILLER_0_132_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_629 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_636 ();
 DECAPx2_ASAP7_75t_R FILLER_0_132_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_664 ();
 DECAPx1_ASAP7_75t_R FILLER_0_132_685 ();
 DECAPx4_ASAP7_75t_R FILLER_0_132_694 ();
 FILLER_ASAP7_75t_R FILLER_0_132_704 ();
 FILLER_ASAP7_75t_R FILLER_0_132_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_714 ();
 DECAPx2_ASAP7_75t_R FILLER_0_132_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_728 ();
 FILLER_ASAP7_75t_R FILLER_0_132_735 ();
 DECAPx2_ASAP7_75t_R FILLER_0_132_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_753 ();
 DECAPx1_ASAP7_75t_R FILLER_0_132_759 ();
 FILLER_ASAP7_75t_R FILLER_0_132_766 ();
 DECAPx1_ASAP7_75t_R FILLER_0_132_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_784 ();
 FILLER_ASAP7_75t_R FILLER_0_132_791 ();
 DECAPx2_ASAP7_75t_R FILLER_0_132_798 ();
 FILLER_ASAP7_75t_R FILLER_0_132_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_806 ();
 DECAPx1_ASAP7_75t_R FILLER_0_132_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_817 ();
 FILLER_ASAP7_75t_R FILLER_0_132_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_826 ();
 DECAPx1_ASAP7_75t_R FILLER_0_132_833 ();
 FILLER_ASAP7_75t_R FILLER_0_132_851 ();
 FILLER_ASAP7_75t_R FILLER_0_132_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_863 ();
 FILLER_ASAP7_75t_R FILLER_0_132_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_871 ();
 DECAPx2_ASAP7_75t_R FILLER_0_132_879 ();
 DECAPx2_ASAP7_75t_R FILLER_0_132_891 ();
 DECAPx2_ASAP7_75t_R FILLER_0_132_907 ();
 DECAPx6_ASAP7_75t_R FILLER_0_132_919 ();
 DECAPx1_ASAP7_75t_R FILLER_0_132_933 ();
 DECAPx2_ASAP7_75t_R FILLER_0_132_943 ();
 FILLER_ASAP7_75t_R FILLER_0_132_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_951 ();
 DECAPx4_ASAP7_75t_R FILLER_0_132_955 ();
 FILLER_ASAP7_75t_R FILLER_0_132_965 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_967 ();
 DECAPx4_ASAP7_75t_R FILLER_0_132_974 ();
 FILLER_ASAP7_75t_R FILLER_0_132_987 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_989 ();
 FILLER_ASAP7_75t_R FILLER_0_132_998 ();
 FILLER_ASAP7_75t_R FILLER_0_132_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_1010 ();
 DECAPx1_ASAP7_75t_R FILLER_0_132_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_1021 ();
 DECAPx4_ASAP7_75t_R FILLER_0_132_1030 ();
 FILLER_ASAP7_75t_R FILLER_0_132_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_1042 ();
 DECAPx4_ASAP7_75t_R FILLER_0_132_1054 ();
 FILLER_ASAP7_75t_R FILLER_0_132_1067 ();
 FILLER_ASAP7_75t_R FILLER_0_132_1079 ();
 FILLER_ASAP7_75t_R FILLER_0_132_1089 ();
 FILLER_ASAP7_75t_R FILLER_0_132_1099 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_1112 ();
 DECAPx2_ASAP7_75t_R FILLER_0_132_1134 ();
 FILLER_ASAP7_75t_R FILLER_0_132_1140 ();
 FILLER_ASAP7_75t_R FILLER_0_132_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_1150 ();
 DECAPx1_ASAP7_75t_R FILLER_0_132_1161 ();
 FILLER_ASAP7_75t_R FILLER_0_132_1175 ();
 FILLER_ASAP7_75t_R FILLER_0_132_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_1189 ();
 FILLER_ASAP7_75t_R FILLER_0_132_1196 ();
 DECAPx1_ASAP7_75t_R FILLER_0_132_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_1208 ();
 FILLER_ASAP7_75t_R FILLER_0_132_1215 ();
 DECAPx4_ASAP7_75t_R FILLER_0_132_1223 ();
 FILLER_ASAP7_75t_R FILLER_0_132_1233 ();
 DECAPx1_ASAP7_75t_R FILLER_0_132_1245 ();
 FILLER_ASAP7_75t_R FILLER_0_132_1259 ();
 DECAPx2_ASAP7_75t_R FILLER_0_132_1267 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_1273 ();
 FILLER_ASAP7_75t_R FILLER_0_132_1281 ();
 DECAPx2_ASAP7_75t_R FILLER_0_132_1289 ();
 FILLER_ASAP7_75t_R FILLER_0_132_1295 ();
 DECAPx4_ASAP7_75t_R FILLER_0_132_1304 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_1314 ();
 DECAPx4_ASAP7_75t_R FILLER_0_132_1323 ();
 DECAPx1_ASAP7_75t_R FILLER_0_132_1345 ();
 FILLER_ASAP7_75t_R FILLER_0_132_1371 ();
 DECAPx1_ASAP7_75t_R FILLER_0_132_1378 ();
 FILLER_ASAP7_75t_R FILLER_0_133_2 ();
 FILLER_ASAP7_75t_R FILLER_0_133_9 ();
 FILLER_ASAP7_75t_R FILLER_0_133_16 ();
 FILLER_ASAP7_75t_R FILLER_0_133_23 ();
 FILLER_ASAP7_75t_R FILLER_0_133_30 ();
 FILLER_ASAP7_75t_R FILLER_0_133_38 ();
 FILLER_ASAP7_75t_R FILLER_0_133_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_48 ();
 FILLER_ASAP7_75t_R FILLER_0_133_55 ();
 DECAPx4_ASAP7_75t_R FILLER_0_133_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_70 ();
 FILLER_ASAP7_75t_R FILLER_0_133_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_79 ();
 DECAPx4_ASAP7_75t_R FILLER_0_133_86 ();
 FILLER_ASAP7_75t_R FILLER_0_133_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_98 ();
 DECAPx2_ASAP7_75t_R FILLER_0_133_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_111 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_120 ();
 DECAPx4_ASAP7_75t_R FILLER_0_133_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_152 ();
 DECAPx4_ASAP7_75t_R FILLER_0_133_163 ();
 FILLER_ASAP7_75t_R FILLER_0_133_173 ();
 FILLER_ASAP7_75t_R FILLER_0_133_183 ();
 FILLER_ASAP7_75t_R FILLER_0_133_193 ();
 DECAPx6_ASAP7_75t_R FILLER_0_133_205 ();
 DECAPx2_ASAP7_75t_R FILLER_0_133_231 ();
 DECAPx4_ASAP7_75t_R FILLER_0_133_245 ();
 FILLER_ASAP7_75t_R FILLER_0_133_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_264 ();
 FILLER_ASAP7_75t_R FILLER_0_133_286 ();
 DECAPx6_ASAP7_75t_R FILLER_0_133_296 ();
 FILLER_ASAP7_75t_R FILLER_0_133_310 ();
 FILLER_ASAP7_75t_R FILLER_0_133_322 ();
 FILLER_ASAP7_75t_R FILLER_0_133_332 ();
 FILLER_ASAP7_75t_R FILLER_0_133_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_342 ();
 FILLER_ASAP7_75t_R FILLER_0_133_351 ();
 DECAPx2_ASAP7_75t_R FILLER_0_133_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_365 ();
 FILLER_ASAP7_75t_R FILLER_0_133_369 ();
 DECAPx4_ASAP7_75t_R FILLER_0_133_377 ();
 FILLER_ASAP7_75t_R FILLER_0_133_387 ();
 FILLER_ASAP7_75t_R FILLER_0_133_395 ();
 DECAPx2_ASAP7_75t_R FILLER_0_133_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_410 ();
 DECAPx2_ASAP7_75t_R FILLER_0_133_418 ();
 FILLER_ASAP7_75t_R FILLER_0_133_424 ();
 FILLER_ASAP7_75t_R FILLER_0_133_432 ();
 FILLER_ASAP7_75t_R FILLER_0_133_445 ();
 DECAPx6_ASAP7_75t_R FILLER_0_133_453 ();
 DECAPx1_ASAP7_75t_R FILLER_0_133_467 ();
 DECAPx2_ASAP7_75t_R FILLER_0_133_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_487 ();
 FILLER_ASAP7_75t_R FILLER_0_133_493 ();
 DECAPx2_ASAP7_75t_R FILLER_0_133_501 ();
 FILLER_ASAP7_75t_R FILLER_0_133_510 ();
 DECAPx6_ASAP7_75t_R FILLER_0_133_515 ();
 DECAPx2_ASAP7_75t_R FILLER_0_133_539 ();
 FILLER_ASAP7_75t_R FILLER_0_133_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_547 ();
 DECAPx2_ASAP7_75t_R FILLER_0_133_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_561 ();
 FILLER_ASAP7_75t_R FILLER_0_133_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_570 ();
 FILLER_ASAP7_75t_R FILLER_0_133_577 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_579 ();
 FILLER_ASAP7_75t_R FILLER_0_133_588 ();
 DECAPx1_ASAP7_75t_R FILLER_0_133_598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_605 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_627 ();
 DECAPx4_ASAP7_75t_R FILLER_0_133_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_659 ();
 DECAPx6_ASAP7_75t_R FILLER_0_133_670 ();
 DECAPx1_ASAP7_75t_R FILLER_0_133_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_688 ();
 FILLER_ASAP7_75t_R FILLER_0_133_692 ();
 FILLER_ASAP7_75t_R FILLER_0_133_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_707 ();
 DECAPx4_ASAP7_75t_R FILLER_0_133_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_724 ();
 FILLER_ASAP7_75t_R FILLER_0_133_731 ();
 FILLER_ASAP7_75t_R FILLER_0_133_739 ();
 FILLER_ASAP7_75t_R FILLER_0_133_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_749 ();
 DECAPx2_ASAP7_75t_R FILLER_0_133_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_766 ();
 DECAPx4_ASAP7_75t_R FILLER_0_133_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_780 ();
 FILLER_ASAP7_75t_R FILLER_0_133_789 ();
 DECAPx2_ASAP7_75t_R FILLER_0_133_796 ();
 FILLER_ASAP7_75t_R FILLER_0_133_809 ();
 FILLER_ASAP7_75t_R FILLER_0_133_816 ();
 FILLER_ASAP7_75t_R FILLER_0_133_823 ();
 DECAPx1_ASAP7_75t_R FILLER_0_133_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_835 ();
 FILLER_ASAP7_75t_R FILLER_0_133_842 ();
 DECAPx2_ASAP7_75t_R FILLER_0_133_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_855 ();
 DECAPx6_ASAP7_75t_R FILLER_0_133_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_876 ();
 FILLER_ASAP7_75t_R FILLER_0_133_882 ();
 DECAPx4_ASAP7_75t_R FILLER_0_133_892 ();
 FILLER_ASAP7_75t_R FILLER_0_133_902 ();
 DECAPx4_ASAP7_75t_R FILLER_0_133_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_924 ();
 DECAPx6_ASAP7_75t_R FILLER_0_133_927 ();
 FILLER_ASAP7_75t_R FILLER_0_133_941 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_943 ();
 DECAPx6_ASAP7_75t_R FILLER_0_133_954 ();
 FILLER_ASAP7_75t_R FILLER_0_133_968 ();
 DECAPx2_ASAP7_75t_R FILLER_0_133_978 ();
 DECAPx2_ASAP7_75t_R FILLER_0_133_992 ();
 FILLER_ASAP7_75t_R FILLER_0_133_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_1000 ();
 DECAPx6_ASAP7_75t_R FILLER_0_133_1007 ();
 FILLER_ASAP7_75t_R FILLER_0_133_1029 ();
 FILLER_ASAP7_75t_R FILLER_0_133_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_1043 ();
 DECAPx1_ASAP7_75t_R FILLER_0_133_1065 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_1069 ();
 FILLER_ASAP7_75t_R FILLER_0_133_1090 ();
 DECAPx2_ASAP7_75t_R FILLER_0_133_1098 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_1107 ();
 DECAPx4_ASAP7_75t_R FILLER_0_133_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_1139 ();
 DECAPx1_ASAP7_75t_R FILLER_0_133_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_1149 ();
 DECAPx4_ASAP7_75t_R FILLER_0_133_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_1170 ();
 FILLER_ASAP7_75t_R FILLER_0_133_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_1183 ();
 FILLER_ASAP7_75t_R FILLER_0_133_1192 ();
 FILLER_ASAP7_75t_R FILLER_0_133_1202 ();
 FILLER_ASAP7_75t_R FILLER_0_133_1210 ();
 FILLER_ASAP7_75t_R FILLER_0_133_1218 ();
 DECAPx2_ASAP7_75t_R FILLER_0_133_1226 ();
 FILLER_ASAP7_75t_R FILLER_0_133_1232 ();
 FILLER_ASAP7_75t_R FILLER_0_133_1240 ();
 DECAPx2_ASAP7_75t_R FILLER_0_133_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_1264 ();
 DECAPx4_ASAP7_75t_R FILLER_0_133_1286 ();
 FILLER_ASAP7_75t_R FILLER_0_133_1296 ();
 DECAPx2_ASAP7_75t_R FILLER_0_133_1306 ();
 FILLER_ASAP7_75t_R FILLER_0_133_1312 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_1314 ();
 FILLER_ASAP7_75t_R FILLER_0_133_1321 ();
 DECAPx4_ASAP7_75t_R FILLER_0_133_1331 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133_1341 ();
 FILLER_ASAP7_75t_R FILLER_0_133_1345 ();
 FILLER_ASAP7_75t_R FILLER_0_133_1352 ();
 FILLER_ASAP7_75t_R FILLER_0_133_1360 ();
 FILLER_ASAP7_75t_R FILLER_0_133_1368 ();
 DECAPx2_ASAP7_75t_R FILLER_0_133_1376 ();
 FILLER_ASAP7_75t_R FILLER_0_134_2 ();
 FILLER_ASAP7_75t_R FILLER_0_134_9 ();
 FILLER_ASAP7_75t_R FILLER_0_134_16 ();
 DECAPx2_ASAP7_75t_R FILLER_0_134_23 ();
 FILLER_ASAP7_75t_R FILLER_0_134_50 ();
 DECAPx2_ASAP7_75t_R FILLER_0_134_57 ();
 FILLER_ASAP7_75t_R FILLER_0_134_63 ();
 FILLER_ASAP7_75t_R FILLER_0_134_71 ();
 DECAPx6_ASAP7_75t_R FILLER_0_134_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_95 ();
 FILLER_ASAP7_75t_R FILLER_0_134_108 ();
 FILLER_ASAP7_75t_R FILLER_0_134_116 ();
 DECAPx2_ASAP7_75t_R FILLER_0_134_124 ();
 FILLER_ASAP7_75t_R FILLER_0_134_130 ();
 DECAPx1_ASAP7_75t_R FILLER_0_134_138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_134_150 ();
 DECAPx6_ASAP7_75t_R FILLER_0_134_166 ();
 DECAPx2_ASAP7_75t_R FILLER_0_134_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_186 ();
 DECAPx1_ASAP7_75t_R FILLER_0_134_193 ();
 DECAPx2_ASAP7_75t_R FILLER_0_134_203 ();
 DECAPx1_ASAP7_75t_R FILLER_0_134_231 ();
 DECAPx2_ASAP7_75t_R FILLER_0_134_241 ();
 FILLER_ASAP7_75t_R FILLER_0_134_257 ();
 DECAPx4_ASAP7_75t_R FILLER_0_134_269 ();
 FILLER_ASAP7_75t_R FILLER_0_134_279 ();
 FILLER_ASAP7_75t_R FILLER_0_134_291 ();
 FILLER_ASAP7_75t_R FILLER_0_134_298 ();
 FILLER_ASAP7_75t_R FILLER_0_134_305 ();
 FILLER_ASAP7_75t_R FILLER_0_134_310 ();
 DECAPx1_ASAP7_75t_R FILLER_0_134_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_326 ();
 FILLER_ASAP7_75t_R FILLER_0_134_337 ();
 DECAPx1_ASAP7_75t_R FILLER_0_134_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_351 ();
 FILLER_ASAP7_75t_R FILLER_0_134_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_360 ();
 FILLER_ASAP7_75t_R FILLER_0_134_367 ();
 DECAPx2_ASAP7_75t_R FILLER_0_134_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_381 ();
 FILLER_ASAP7_75t_R FILLER_0_134_388 ();
 FILLER_ASAP7_75t_R FILLER_0_134_396 ();
 DECAPx2_ASAP7_75t_R FILLER_0_134_418 ();
 FILLER_ASAP7_75t_R FILLER_0_134_424 ();
 FILLER_ASAP7_75t_R FILLER_0_134_432 ();
 DECAPx2_ASAP7_75t_R FILLER_0_134_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_446 ();
 DECAPx2_ASAP7_75t_R FILLER_0_134_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_461 ();
 FILLER_ASAP7_75t_R FILLER_0_134_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_466 ();
 DECAPx2_ASAP7_75t_R FILLER_0_134_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_476 ();
 DECAPx6_ASAP7_75t_R FILLER_0_134_487 ();
 FILLER_ASAP7_75t_R FILLER_0_134_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_523 ();
 FILLER_ASAP7_75t_R FILLER_0_134_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_532 ();
 FILLER_ASAP7_75t_R FILLER_0_134_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_541 ();
 DECAPx1_ASAP7_75t_R FILLER_0_134_548 ();
 DECAPx1_ASAP7_75t_R FILLER_0_134_558 ();
 FILLER_ASAP7_75t_R FILLER_0_134_568 ();
 DECAPx4_ASAP7_75t_R FILLER_0_134_576 ();
 FILLER_ASAP7_75t_R FILLER_0_134_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_588 ();
 DECAPx6_ASAP7_75t_R FILLER_0_134_600 ();
 DECAPx1_ASAP7_75t_R FILLER_0_134_614 ();
 DECAPx4_ASAP7_75t_R FILLER_0_134_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_650 ();
 FILLER_ASAP7_75t_R FILLER_0_134_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_661 ();
 DECAPx6_ASAP7_75t_R FILLER_0_134_665 ();
 DECAPx2_ASAP7_75t_R FILLER_0_134_679 ();
 DECAPx1_ASAP7_75t_R FILLER_0_134_693 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_707 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_736 ();
 DECAPx1_ASAP7_75t_R FILLER_0_134_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_762 ();
 DECAPx2_ASAP7_75t_R FILLER_0_134_770 ();
 FILLER_ASAP7_75t_R FILLER_0_134_781 ();
 DECAPx2_ASAP7_75t_R FILLER_0_134_793 ();
 DECAPx1_ASAP7_75t_R FILLER_0_134_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_813 ();
 FILLER_ASAP7_75t_R FILLER_0_134_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_826 ();
 FILLER_ASAP7_75t_R FILLER_0_134_837 ();
 FILLER_ASAP7_75t_R FILLER_0_134_844 ();
 DECAPx6_ASAP7_75t_R FILLER_0_134_851 ();
 DECAPx1_ASAP7_75t_R FILLER_0_134_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_869 ();
 FILLER_ASAP7_75t_R FILLER_0_134_878 ();
 FILLER_ASAP7_75t_R FILLER_0_134_886 ();
 FILLER_ASAP7_75t_R FILLER_0_134_894 ();
 DECAPx1_ASAP7_75t_R FILLER_0_134_902 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_916 ();
 DECAPx2_ASAP7_75t_R FILLER_0_134_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_944 ();
 DECAPx4_ASAP7_75t_R FILLER_0_134_956 ();
 FILLER_ASAP7_75t_R FILLER_0_134_966 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_968 ();
 DECAPx2_ASAP7_75t_R FILLER_0_134_975 ();
 FILLER_ASAP7_75t_R FILLER_0_134_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_983 ();
 FILLER_ASAP7_75t_R FILLER_0_134_992 ();
 DECAPx6_ASAP7_75t_R FILLER_0_134_1002 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_1024 ();
 FILLER_ASAP7_75t_R FILLER_0_134_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_1048 ();
 DECAPx4_ASAP7_75t_R FILLER_0_134_1061 ();
 FILLER_ASAP7_75t_R FILLER_0_134_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_1073 ();
 DECAPx1_ASAP7_75t_R FILLER_0_134_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_1090 ();
 FILLER_ASAP7_75t_R FILLER_0_134_1103 ();
 FILLER_ASAP7_75t_R FILLER_0_134_1117 ();
 FILLER_ASAP7_75t_R FILLER_0_134_1141 ();
 DECAPx6_ASAP7_75t_R FILLER_0_134_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_1163 ();
 FILLER_ASAP7_75t_R FILLER_0_134_1169 ();
 FILLER_ASAP7_75t_R FILLER_0_134_1177 ();
 FILLER_ASAP7_75t_R FILLER_0_134_1189 ();
 FILLER_ASAP7_75t_R FILLER_0_134_1195 ();
 FILLER_ASAP7_75t_R FILLER_0_134_1207 ();
 FILLER_ASAP7_75t_R FILLER_0_134_1215 ();
 FILLER_ASAP7_75t_R FILLER_0_134_1223 ();
 FILLER_ASAP7_75t_R FILLER_0_134_1230 ();
 DECAPx4_ASAP7_75t_R FILLER_0_134_1244 ();
 FILLER_ASAP7_75t_R FILLER_0_134_1264 ();
 DECAPx1_ASAP7_75t_R FILLER_0_134_1274 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_1278 ();
 DECAPx2_ASAP7_75t_R FILLER_0_134_1285 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_1291 ();
 FILLER_ASAP7_75t_R FILLER_0_134_1298 ();
 DECAPx4_ASAP7_75t_R FILLER_0_134_1306 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_1322 ();
 DECAPx1_ASAP7_75t_R FILLER_0_134_1344 ();
 FILLER_ASAP7_75t_R FILLER_0_134_1351 ();
 FILLER_ASAP7_75t_R FILLER_0_134_1374 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_1376 ();
 FILLER_ASAP7_75t_R FILLER_0_134_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_135_2 ();
 FILLER_ASAP7_75t_R FILLER_0_135_26 ();
 FILLER_ASAP7_75t_R FILLER_0_135_31 ();
 FILLER_ASAP7_75t_R FILLER_0_135_38 ();
 FILLER_ASAP7_75t_R FILLER_0_135_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_48 ();
 FILLER_ASAP7_75t_R FILLER_0_135_70 ();
 DECAPx1_ASAP7_75t_R FILLER_0_135_78 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_110 ();
 DECAPx6_ASAP7_75t_R FILLER_0_135_119 ();
 DECAPx4_ASAP7_75t_R FILLER_0_135_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_154 ();
 FILLER_ASAP7_75t_R FILLER_0_135_163 ();
 DECAPx2_ASAP7_75t_R FILLER_0_135_175 ();
 FILLER_ASAP7_75t_R FILLER_0_135_181 ();
 FILLER_ASAP7_75t_R FILLER_0_135_186 ();
 FILLER_ASAP7_75t_R FILLER_0_135_196 ();
 DECAPx6_ASAP7_75t_R FILLER_0_135_204 ();
 DECAPx2_ASAP7_75t_R FILLER_0_135_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_224 ();
 FILLER_ASAP7_75t_R FILLER_0_135_231 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_239 ();
 DECAPx1_ASAP7_75t_R FILLER_0_135_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_265 ();
 FILLER_ASAP7_75t_R FILLER_0_135_271 ();
 FILLER_ASAP7_75t_R FILLER_0_135_283 ();
 FILLER_ASAP7_75t_R FILLER_0_135_291 ();
 FILLER_ASAP7_75t_R FILLER_0_135_303 ();
 FILLER_ASAP7_75t_R FILLER_0_135_315 ();
 FILLER_ASAP7_75t_R FILLER_0_135_322 ();
 FILLER_ASAP7_75t_R FILLER_0_135_330 ();
 FILLER_ASAP7_75t_R FILLER_0_135_342 ();
 FILLER_ASAP7_75t_R FILLER_0_135_350 ();
 FILLER_ASAP7_75t_R FILLER_0_135_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_360 ();
 FILLER_ASAP7_75t_R FILLER_0_135_367 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_377 ();
 DECAPx2_ASAP7_75t_R FILLER_0_135_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_405 ();
 FILLER_ASAP7_75t_R FILLER_0_135_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_416 ();
 FILLER_ASAP7_75t_R FILLER_0_135_424 ();
 DECAPx2_ASAP7_75t_R FILLER_0_135_431 ();
 FILLER_ASAP7_75t_R FILLER_0_135_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_445 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_449 ();
 DECAPx2_ASAP7_75t_R FILLER_0_135_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_477 ();
 DECAPx6_ASAP7_75t_R FILLER_0_135_488 ();
 DECAPx1_ASAP7_75t_R FILLER_0_135_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_506 ();
 DECAPx6_ASAP7_75t_R FILLER_0_135_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_527 ();
 DECAPx2_ASAP7_75t_R FILLER_0_135_531 ();
 FILLER_ASAP7_75t_R FILLER_0_135_537 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_547 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_569 ();
 FILLER_ASAP7_75t_R FILLER_0_135_591 ();
 DECAPx6_ASAP7_75t_R FILLER_0_135_599 ();
 DECAPx2_ASAP7_75t_R FILLER_0_135_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_619 ();
 DECAPx1_ASAP7_75t_R FILLER_0_135_628 ();
 FILLER_ASAP7_75t_R FILLER_0_135_638 ();
 FILLER_ASAP7_75t_R FILLER_0_135_645 ();
 DECAPx2_ASAP7_75t_R FILLER_0_135_650 ();
 DECAPx6_ASAP7_75t_R FILLER_0_135_676 ();
 DECAPx1_ASAP7_75t_R FILLER_0_135_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_694 ();
 DECAPx1_ASAP7_75t_R FILLER_0_135_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_705 ();
 FILLER_ASAP7_75t_R FILLER_0_135_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_714 ();
 DECAPx1_ASAP7_75t_R FILLER_0_135_721 ();
 DECAPx1_ASAP7_75t_R FILLER_0_135_731 ();
 FILLER_ASAP7_75t_R FILLER_0_135_741 ();
 DECAPx2_ASAP7_75t_R FILLER_0_135_749 ();
 FILLER_ASAP7_75t_R FILLER_0_135_755 ();
 FILLER_ASAP7_75t_R FILLER_0_135_763 ();
 FILLER_ASAP7_75t_R FILLER_0_135_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_774 ();
 FILLER_ASAP7_75t_R FILLER_0_135_785 ();
 DECAPx2_ASAP7_75t_R FILLER_0_135_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_798 ();
 DECAPx2_ASAP7_75t_R FILLER_0_135_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_815 ();
 FILLER_ASAP7_75t_R FILLER_0_135_826 ();
 FILLER_ASAP7_75t_R FILLER_0_135_838 ();
 FILLER_ASAP7_75t_R FILLER_0_135_846 ();
 FILLER_ASAP7_75t_R FILLER_0_135_854 ();
 FILLER_ASAP7_75t_R FILLER_0_135_862 ();
 DECAPx1_ASAP7_75t_R FILLER_0_135_870 ();
 DECAPx2_ASAP7_75t_R FILLER_0_135_884 ();
 DECAPx2_ASAP7_75t_R FILLER_0_135_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_902 ();
 FILLER_ASAP7_75t_R FILLER_0_135_923 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_927 ();
 DECAPx6_ASAP7_75t_R FILLER_0_135_949 ();
 DECAPx2_ASAP7_75t_R FILLER_0_135_963 ();
 FILLER_ASAP7_75t_R FILLER_0_135_973 ();
 FILLER_ASAP7_75t_R FILLER_0_135_981 ();
 DECAPx2_ASAP7_75t_R FILLER_0_135_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_995 ();
 FILLER_ASAP7_75t_R FILLER_0_135_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_1008 ();
 FILLER_ASAP7_75t_R FILLER_0_135_1017 ();
 FILLER_ASAP7_75t_R FILLER_0_135_1027 ();
 DECAPx1_ASAP7_75t_R FILLER_0_135_1032 ();
 FILLER_ASAP7_75t_R FILLER_0_135_1048 ();
 DECAPx1_ASAP7_75t_R FILLER_0_135_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_1066 ();
 DECAPx2_ASAP7_75t_R FILLER_0_135_1079 ();
 FILLER_ASAP7_75t_R FILLER_0_135_1085 ();
 FILLER_ASAP7_75t_R FILLER_0_135_1090 ();
 DECAPx1_ASAP7_75t_R FILLER_0_135_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_1104 ();
 DECAPx4_ASAP7_75t_R FILLER_0_135_1111 ();
 DECAPx1_ASAP7_75t_R FILLER_0_135_1124 ();
 FILLER_ASAP7_75t_R FILLER_0_135_1138 ();
 FILLER_ASAP7_75t_R FILLER_0_135_1158 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_1160 ();
 DECAPx2_ASAP7_75t_R FILLER_0_135_1171 ();
 FILLER_ASAP7_75t_R FILLER_0_135_1187 ();
 FILLER_ASAP7_75t_R FILLER_0_135_1199 ();
 FILLER_ASAP7_75t_R FILLER_0_135_1207 ();
 FILLER_ASAP7_75t_R FILLER_0_135_1215 ();
 FILLER_ASAP7_75t_R FILLER_0_135_1223 ();
 DECAPx2_ASAP7_75t_R FILLER_0_135_1231 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_1237 ();
 DECAPx4_ASAP7_75t_R FILLER_0_135_1241 ();
 FILLER_ASAP7_75t_R FILLER_0_135_1263 ();
 FILLER_ASAP7_75t_R FILLER_0_135_1271 ();
 FILLER_ASAP7_75t_R FILLER_0_135_1281 ();
 DECAPx2_ASAP7_75t_R FILLER_0_135_1289 ();
 DECAPx2_ASAP7_75t_R FILLER_0_135_1306 ();
 FILLER_ASAP7_75t_R FILLER_0_135_1312 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_1314 ();
 DECAPx4_ASAP7_75t_R FILLER_0_135_1321 ();
 FILLER_ASAP7_75t_R FILLER_0_135_1343 ();
 FILLER_ASAP7_75t_R FILLER_0_135_1350 ();
 FILLER_ASAP7_75t_R FILLER_0_135_1357 ();
 DECAPx2_ASAP7_75t_R FILLER_0_135_1364 ();
 FILLER_ASAP7_75t_R FILLER_0_135_1375 ();
 FILLER_ASAP7_75t_R FILLER_0_135_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_136_2 ();
 FILLER_ASAP7_75t_R FILLER_0_136_7 ();
 FILLER_ASAP7_75t_R FILLER_0_136_14 ();
 FILLER_ASAP7_75t_R FILLER_0_136_21 ();
 FILLER_ASAP7_75t_R FILLER_0_136_28 ();
 FILLER_ASAP7_75t_R FILLER_0_136_35 ();
 DECAPx1_ASAP7_75t_R FILLER_0_136_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_44 ();
 FILLER_ASAP7_75t_R FILLER_0_136_53 ();
 FILLER_ASAP7_75t_R FILLER_0_136_58 ();
 FILLER_ASAP7_75t_R FILLER_0_136_72 ();
 DECAPx6_ASAP7_75t_R FILLER_0_136_82 ();
 DECAPx1_ASAP7_75t_R FILLER_0_136_96 ();
 DECAPx4_ASAP7_75t_R FILLER_0_136_106 ();
 FILLER_ASAP7_75t_R FILLER_0_136_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_118 ();
 DECAPx2_ASAP7_75t_R FILLER_0_136_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_137 ();
 FILLER_ASAP7_75t_R FILLER_0_136_146 ();
 FILLER_ASAP7_75t_R FILLER_0_136_154 ();
 FILLER_ASAP7_75t_R FILLER_0_136_162 ();
 DECAPx4_ASAP7_75t_R FILLER_0_136_170 ();
 DECAPx2_ASAP7_75t_R FILLER_0_136_192 ();
 FILLER_ASAP7_75t_R FILLER_0_136_198 ();
 DECAPx2_ASAP7_75t_R FILLER_0_136_206 ();
 DECAPx4_ASAP7_75t_R FILLER_0_136_220 ();
 FILLER_ASAP7_75t_R FILLER_0_136_236 ();
 FILLER_ASAP7_75t_R FILLER_0_136_244 ();
 DECAPx6_ASAP7_75t_R FILLER_0_136_257 ();
 FILLER_ASAP7_75t_R FILLER_0_136_282 ();
 DECAPx4_ASAP7_75t_R FILLER_0_136_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_304 ();
 FILLER_ASAP7_75t_R FILLER_0_136_315 ();
 DECAPx1_ASAP7_75t_R FILLER_0_136_322 ();
 FILLER_ASAP7_75t_R FILLER_0_136_334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_342 ();
 FILLER_ASAP7_75t_R FILLER_0_136_364 ();
 DECAPx4_ASAP7_75t_R FILLER_0_136_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_382 ();
 FILLER_ASAP7_75t_R FILLER_0_136_389 ();
 DECAPx4_ASAP7_75t_R FILLER_0_136_397 ();
 FILLER_ASAP7_75t_R FILLER_0_136_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_415 ();
 FILLER_ASAP7_75t_R FILLER_0_136_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_425 ();
 DECAPx2_ASAP7_75t_R FILLER_0_136_432 ();
 FILLER_ASAP7_75t_R FILLER_0_136_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_440 ();
 FILLER_ASAP7_75t_R FILLER_0_136_447 ();
 FILLER_ASAP7_75t_R FILLER_0_136_452 ();
 FILLER_ASAP7_75t_R FILLER_0_136_460 ();
 FILLER_ASAP7_75t_R FILLER_0_136_464 ();
 DECAPx1_ASAP7_75t_R FILLER_0_136_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_476 ();
 FILLER_ASAP7_75t_R FILLER_0_136_488 ();
 DECAPx6_ASAP7_75t_R FILLER_0_136_496 ();
 DECAPx4_ASAP7_75t_R FILLER_0_136_516 ();
 FILLER_ASAP7_75t_R FILLER_0_136_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_528 ();
 FILLER_ASAP7_75t_R FILLER_0_136_533 ();
 FILLER_ASAP7_75t_R FILLER_0_136_541 ();
 DECAPx1_ASAP7_75t_R FILLER_0_136_549 ();
 DECAPx2_ASAP7_75t_R FILLER_0_136_559 ();
 FILLER_ASAP7_75t_R FILLER_0_136_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_567 ();
 DECAPx2_ASAP7_75t_R FILLER_0_136_574 ();
 FILLER_ASAP7_75t_R FILLER_0_136_580 ();
 DECAPx2_ASAP7_75t_R FILLER_0_136_603 ();
 FILLER_ASAP7_75t_R FILLER_0_136_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_611 ();
 FILLER_ASAP7_75t_R FILLER_0_136_617 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_640 ();
 DECAPx6_ASAP7_75t_R FILLER_0_136_662 ();
 FILLER_ASAP7_75t_R FILLER_0_136_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_678 ();
 DECAPx1_ASAP7_75t_R FILLER_0_136_689 ();
 FILLER_ASAP7_75t_R FILLER_0_136_703 ();
 FILLER_ASAP7_75t_R FILLER_0_136_713 ();
 DECAPx1_ASAP7_75t_R FILLER_0_136_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_725 ();
 DECAPx1_ASAP7_75t_R FILLER_0_136_736 ();
 DECAPx2_ASAP7_75t_R FILLER_0_136_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_753 ();
 FILLER_ASAP7_75t_R FILLER_0_136_765 ();
 FILLER_ASAP7_75t_R FILLER_0_136_772 ();
 FILLER_ASAP7_75t_R FILLER_0_136_781 ();
 DECAPx2_ASAP7_75t_R FILLER_0_136_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_807 ();
 DECAPx2_ASAP7_75t_R FILLER_0_136_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_820 ();
 FILLER_ASAP7_75t_R FILLER_0_136_829 ();
 FILLER_ASAP7_75t_R FILLER_0_136_837 ();
 FILLER_ASAP7_75t_R FILLER_0_136_845 ();
 FILLER_ASAP7_75t_R FILLER_0_136_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_855 ();
 DECAPx1_ASAP7_75t_R FILLER_0_136_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_866 ();
 FILLER_ASAP7_75t_R FILLER_0_136_873 ();
 FILLER_ASAP7_75t_R FILLER_0_136_882 ();
 DECAPx1_ASAP7_75t_R FILLER_0_136_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_898 ();
 DECAPx1_ASAP7_75t_R FILLER_0_136_905 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_915 ();
 FILLER_ASAP7_75t_R FILLER_0_136_937 ();
 FILLER_ASAP7_75t_R FILLER_0_136_945 ();
 DECAPx2_ASAP7_75t_R FILLER_0_136_957 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_963 ();
 DECAPx1_ASAP7_75t_R FILLER_0_136_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_976 ();
 DECAPx6_ASAP7_75t_R FILLER_0_136_983 ();
 FILLER_ASAP7_75t_R FILLER_0_136_1007 ();
 FILLER_ASAP7_75t_R FILLER_0_136_1019 ();
 FILLER_ASAP7_75t_R FILLER_0_136_1029 ();
 DECAPx6_ASAP7_75t_R FILLER_0_136_1037 ();
 DECAPx6_ASAP7_75t_R FILLER_0_136_1062 ();
 DECAPx1_ASAP7_75t_R FILLER_0_136_1076 ();
 FILLER_ASAP7_75t_R FILLER_0_136_1088 ();
 DECAPx1_ASAP7_75t_R FILLER_0_136_1100 ();
 DECAPx6_ASAP7_75t_R FILLER_0_136_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_1129 ();
 DECAPx1_ASAP7_75t_R FILLER_0_136_1136 ();
 DECAPx1_ASAP7_75t_R FILLER_0_136_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_1154 ();
 FILLER_ASAP7_75t_R FILLER_0_136_1160 ();
 DECAPx1_ASAP7_75t_R FILLER_0_136_1172 ();
 FILLER_ASAP7_75t_R FILLER_0_136_1182 ();
 FILLER_ASAP7_75t_R FILLER_0_136_1198 ();
 FILLER_ASAP7_75t_R FILLER_0_136_1206 ();
 FILLER_ASAP7_75t_R FILLER_0_136_1215 ();
 FILLER_ASAP7_75t_R FILLER_0_136_1223 ();
 DECAPx2_ASAP7_75t_R FILLER_0_136_1230 ();
 DECAPx4_ASAP7_75t_R FILLER_0_136_1242 ();
 DECAPx4_ASAP7_75t_R FILLER_0_136_1264 ();
 FILLER_ASAP7_75t_R FILLER_0_136_1274 ();
 FILLER_ASAP7_75t_R FILLER_0_136_1282 ();
 DECAPx4_ASAP7_75t_R FILLER_0_136_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_1300 ();
 FILLER_ASAP7_75t_R FILLER_0_136_1307 ();
 DECAPx2_ASAP7_75t_R FILLER_0_136_1315 ();
 FILLER_ASAP7_75t_R FILLER_0_136_1321 ();
 FILLER_ASAP7_75t_R FILLER_0_136_1329 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_1331 ();
 FILLER_ASAP7_75t_R FILLER_0_136_1335 ();
 FILLER_ASAP7_75t_R FILLER_0_136_1342 ();
 FILLER_ASAP7_75t_R FILLER_0_136_1365 ();
 FILLER_ASAP7_75t_R FILLER_0_136_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_136_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_137_2 ();
 FILLER_ASAP7_75t_R FILLER_0_137_26 ();
 FILLER_ASAP7_75t_R FILLER_0_137_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_36 ();
 DECAPx1_ASAP7_75t_R FILLER_0_137_43 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_74 ();
 FILLER_ASAP7_75t_R FILLER_0_137_78 ();
 FILLER_ASAP7_75t_R FILLER_0_137_86 ();
 FILLER_ASAP7_75t_R FILLER_0_137_100 ();
 DECAPx2_ASAP7_75t_R FILLER_0_137_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_114 ();
 DECAPx2_ASAP7_75t_R FILLER_0_137_126 ();
 FILLER_ASAP7_75t_R FILLER_0_137_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_134 ();
 DECAPx4_ASAP7_75t_R FILLER_0_137_141 ();
 FILLER_ASAP7_75t_R FILLER_0_137_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_153 ();
 DECAPx6_ASAP7_75t_R FILLER_0_137_164 ();
 DECAPx1_ASAP7_75t_R FILLER_0_137_178 ();
 FILLER_ASAP7_75t_R FILLER_0_137_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_196 ();
 FILLER_ASAP7_75t_R FILLER_0_137_207 ();
 FILLER_ASAP7_75t_R FILLER_0_137_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_222 ();
 FILLER_ASAP7_75t_R FILLER_0_137_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_237 ();
 FILLER_ASAP7_75t_R FILLER_0_137_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_246 ();
 FILLER_ASAP7_75t_R FILLER_0_137_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_255 ();
 FILLER_ASAP7_75t_R FILLER_0_137_268 ();
 DECAPx1_ASAP7_75t_R FILLER_0_137_276 ();
 DECAPx2_ASAP7_75t_R FILLER_0_137_285 ();
 FILLER_ASAP7_75t_R FILLER_0_137_291 ();
 DECAPx2_ASAP7_75t_R FILLER_0_137_303 ();
 FILLER_ASAP7_75t_R FILLER_0_137_319 ();
 DECAPx2_ASAP7_75t_R FILLER_0_137_329 ();
 DECAPx4_ASAP7_75t_R FILLER_0_137_343 ();
 FILLER_ASAP7_75t_R FILLER_0_137_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_355 ();
 DECAPx2_ASAP7_75t_R FILLER_0_137_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_368 ();
 DECAPx4_ASAP7_75t_R FILLER_0_137_375 ();
 FILLER_ASAP7_75t_R FILLER_0_137_393 ();
 DECAPx2_ASAP7_75t_R FILLER_0_137_401 ();
 FILLER_ASAP7_75t_R FILLER_0_137_407 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_415 ();
 DECAPx2_ASAP7_75t_R FILLER_0_137_437 ();
 FILLER_ASAP7_75t_R FILLER_0_137_443 ();
 FILLER_ASAP7_75t_R FILLER_0_137_451 ();
 DECAPx6_ASAP7_75t_R FILLER_0_137_459 ();
 FILLER_ASAP7_75t_R FILLER_0_137_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_475 ();
 FILLER_ASAP7_75t_R FILLER_0_137_482 ();
 FILLER_ASAP7_75t_R FILLER_0_137_487 ();
 DECAPx2_ASAP7_75t_R FILLER_0_137_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_501 ();
 FILLER_ASAP7_75t_R FILLER_0_137_513 ();
 DECAPx1_ASAP7_75t_R FILLER_0_137_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_525 ();
 DECAPx6_ASAP7_75t_R FILLER_0_137_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_550 ();
 FILLER_ASAP7_75t_R FILLER_0_137_557 ();
 FILLER_ASAP7_75t_R FILLER_0_137_565 ();
 DECAPx2_ASAP7_75t_R FILLER_0_137_570 ();
 FILLER_ASAP7_75t_R FILLER_0_137_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_578 ();
 FILLER_ASAP7_75t_R FILLER_0_137_582 ();
 DECAPx4_ASAP7_75t_R FILLER_0_137_592 ();
 FILLER_ASAP7_75t_R FILLER_0_137_602 ();
 DECAPx1_ASAP7_75t_R FILLER_0_137_615 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_630 ();
 FILLER_ASAP7_75t_R FILLER_0_137_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_654 ();
 FILLER_ASAP7_75t_R FILLER_0_137_675 ();
 FILLER_ASAP7_75t_R FILLER_0_137_680 ();
 FILLER_ASAP7_75t_R FILLER_0_137_692 ();
 FILLER_ASAP7_75t_R FILLER_0_137_704 ();
 DECAPx1_ASAP7_75t_R FILLER_0_137_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_718 ();
 FILLER_ASAP7_75t_R FILLER_0_137_725 ();
 FILLER_ASAP7_75t_R FILLER_0_137_733 ();
 FILLER_ASAP7_75t_R FILLER_0_137_741 ();
 FILLER_ASAP7_75t_R FILLER_0_137_749 ();
 DECAPx2_ASAP7_75t_R FILLER_0_137_757 ();
 FILLER_ASAP7_75t_R FILLER_0_137_763 ();
 FILLER_ASAP7_75t_R FILLER_0_137_775 ();
 FILLER_ASAP7_75t_R FILLER_0_137_787 ();
 FILLER_ASAP7_75t_R FILLER_0_137_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_801 ();
 DECAPx2_ASAP7_75t_R FILLER_0_137_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_818 ();
 FILLER_ASAP7_75t_R FILLER_0_137_826 ();
 FILLER_ASAP7_75t_R FILLER_0_137_834 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_836 ();
 FILLER_ASAP7_75t_R FILLER_0_137_843 ();
 FILLER_ASAP7_75t_R FILLER_0_137_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_853 ();
 FILLER_ASAP7_75t_R FILLER_0_137_860 ();
 FILLER_ASAP7_75t_R FILLER_0_137_868 ();
 DECAPx1_ASAP7_75t_R FILLER_0_137_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_880 ();
 FILLER_ASAP7_75t_R FILLER_0_137_886 ();
 FILLER_ASAP7_75t_R FILLER_0_137_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_896 ();
 FILLER_ASAP7_75t_R FILLER_0_137_903 ();
 FILLER_ASAP7_75t_R FILLER_0_137_911 ();
 DECAPx2_ASAP7_75t_R FILLER_0_137_916 ();
 FILLER_ASAP7_75t_R FILLER_0_137_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_924 ();
 FILLER_ASAP7_75t_R FILLER_0_137_927 ();
 FILLER_ASAP7_75t_R FILLER_0_137_949 ();
 FILLER_ASAP7_75t_R FILLER_0_137_959 ();
 DECAPx2_ASAP7_75t_R FILLER_0_137_969 ();
 FILLER_ASAP7_75t_R FILLER_0_137_983 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_995 ();
 DECAPx1_ASAP7_75t_R FILLER_0_137_1017 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_1029 ();
 DECAPx6_ASAP7_75t_R FILLER_0_137_1051 ();
 DECAPx1_ASAP7_75t_R FILLER_0_137_1065 ();
 FILLER_ASAP7_75t_R FILLER_0_137_1079 ();
 FILLER_ASAP7_75t_R FILLER_0_137_1092 ();
 FILLER_ASAP7_75t_R FILLER_0_137_1102 ();
 FILLER_ASAP7_75t_R FILLER_0_137_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_1114 ();
 DECAPx4_ASAP7_75t_R FILLER_0_137_1118 ();
 FILLER_ASAP7_75t_R FILLER_0_137_1128 ();
 DECAPx1_ASAP7_75t_R FILLER_0_137_1140 ();
 DECAPx1_ASAP7_75t_R FILLER_0_137_1150 ();
 FILLER_ASAP7_75t_R FILLER_0_137_1160 ();
 FILLER_ASAP7_75t_R FILLER_0_137_1172 ();
 FILLER_ASAP7_75t_R FILLER_0_137_1180 ();
 FILLER_ASAP7_75t_R FILLER_0_137_1198 ();
 FILLER_ASAP7_75t_R FILLER_0_137_1210 ();
 DECAPx2_ASAP7_75t_R FILLER_0_137_1218 ();
 DECAPx1_ASAP7_75t_R FILLER_0_137_1232 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_1236 ();
 DECAPx2_ASAP7_75t_R FILLER_0_137_1247 ();
 FILLER_ASAP7_75t_R FILLER_0_137_1253 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_1255 ();
 FILLER_ASAP7_75t_R FILLER_0_137_1262 ();
 DECAPx2_ASAP7_75t_R FILLER_0_137_1269 ();
 FILLER_ASAP7_75t_R FILLER_0_137_1275 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_1277 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_1283 ();
 FILLER_ASAP7_75t_R FILLER_0_137_1305 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_1307 ();
 DECAPx2_ASAP7_75t_R FILLER_0_137_1314 ();
 FILLER_ASAP7_75t_R FILLER_0_137_1336 ();
 FILLER_ASAP7_75t_R FILLER_0_137_1349 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_1351 ();
 FILLER_ASAP7_75t_R FILLER_0_137_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_137_1365 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137_1367 ();
 FILLER_ASAP7_75t_R FILLER_0_137_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_137_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_138_2 ();
 FILLER_ASAP7_75t_R FILLER_0_138_9 ();
 FILLER_ASAP7_75t_R FILLER_0_138_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_18 ();
 FILLER_ASAP7_75t_R FILLER_0_138_25 ();
 FILLER_ASAP7_75t_R FILLER_0_138_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_138_56 ();
 DECAPx2_ASAP7_75t_R FILLER_0_138_66 ();
 FILLER_ASAP7_75t_R FILLER_0_138_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_74 ();
 FILLER_ASAP7_75t_R FILLER_0_138_80 ();
 FILLER_ASAP7_75t_R FILLER_0_138_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_96 ();
 DECAPx6_ASAP7_75t_R FILLER_0_138_105 ();
 FILLER_ASAP7_75t_R FILLER_0_138_119 ();
 DECAPx6_ASAP7_75t_R FILLER_0_138_133 ();
 FILLER_ASAP7_75t_R FILLER_0_138_153 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_165 ();
 DECAPx2_ASAP7_75t_R FILLER_0_138_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_193 ();
 FILLER_ASAP7_75t_R FILLER_0_138_204 ();
 FILLER_ASAP7_75t_R FILLER_0_138_209 ();
 DECAPx4_ASAP7_75t_R FILLER_0_138_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_227 ();
 DECAPx2_ASAP7_75t_R FILLER_0_138_233 ();
 FILLER_ASAP7_75t_R FILLER_0_138_247 ();
 DECAPx1_ASAP7_75t_R FILLER_0_138_252 ();
 FILLER_ASAP7_75t_R FILLER_0_138_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_270 ();
 FILLER_ASAP7_75t_R FILLER_0_138_295 ();
 DECAPx2_ASAP7_75t_R FILLER_0_138_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_313 ();
 FILLER_ASAP7_75t_R FILLER_0_138_324 ();
 FILLER_ASAP7_75t_R FILLER_0_138_333 ();
 FILLER_ASAP7_75t_R FILLER_0_138_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_343 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_364 ();
 DECAPx4_ASAP7_75t_R FILLER_0_138_386 ();
 DECAPx6_ASAP7_75t_R FILLER_0_138_402 ();
 DECAPx1_ASAP7_75t_R FILLER_0_138_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_420 ();
 DECAPx4_ASAP7_75t_R FILLER_0_138_427 ();
 FILLER_ASAP7_75t_R FILLER_0_138_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_445 ();
 DECAPx4_ASAP7_75t_R FILLER_0_138_452 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_464 ();
 DECAPx2_ASAP7_75t_R FILLER_0_138_486 ();
 FILLER_ASAP7_75t_R FILLER_0_138_492 ();
 DECAPx1_ASAP7_75t_R FILLER_0_138_500 ();
 FILLER_ASAP7_75t_R FILLER_0_138_507 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_515 ();
 DECAPx6_ASAP7_75t_R FILLER_0_138_537 ();
 DECAPx1_ASAP7_75t_R FILLER_0_138_551 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_588 ();
 DECAPx4_ASAP7_75t_R FILLER_0_138_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_624 ();
 DECAPx4_ASAP7_75t_R FILLER_0_138_646 ();
 FILLER_ASAP7_75t_R FILLER_0_138_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_658 ();
 FILLER_ASAP7_75t_R FILLER_0_138_664 ();
 DECAPx2_ASAP7_75t_R FILLER_0_138_676 ();
 FILLER_ASAP7_75t_R FILLER_0_138_688 ();
 DECAPx2_ASAP7_75t_R FILLER_0_138_700 ();
 FILLER_ASAP7_75t_R FILLER_0_138_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_708 ();
 FILLER_ASAP7_75t_R FILLER_0_138_719 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_727 ();
 DECAPx4_ASAP7_75t_R FILLER_0_138_749 ();
 FILLER_ASAP7_75t_R FILLER_0_138_759 ();
 DECAPx1_ASAP7_75t_R FILLER_0_138_767 ();
 FILLER_ASAP7_75t_R FILLER_0_138_776 ();
 FILLER_ASAP7_75t_R FILLER_0_138_796 ();
 DECAPx1_ASAP7_75t_R FILLER_0_138_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_820 ();
 FILLER_ASAP7_75t_R FILLER_0_138_826 ();
 FILLER_ASAP7_75t_R FILLER_0_138_833 ();
 DECAPx2_ASAP7_75t_R FILLER_0_138_840 ();
 FILLER_ASAP7_75t_R FILLER_0_138_852 ();
 FILLER_ASAP7_75t_R FILLER_0_138_858 ();
 FILLER_ASAP7_75t_R FILLER_0_138_870 ();
 FILLER_ASAP7_75t_R FILLER_0_138_878 ();
 FILLER_ASAP7_75t_R FILLER_0_138_886 ();
 FILLER_ASAP7_75t_R FILLER_0_138_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_895 ();
 FILLER_ASAP7_75t_R FILLER_0_138_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_904 ();
 DECAPx4_ASAP7_75t_R FILLER_0_138_913 ();
 DECAPx1_ASAP7_75t_R FILLER_0_138_944 ();
 FILLER_ASAP7_75t_R FILLER_0_138_953 ();
 DECAPx1_ASAP7_75t_R FILLER_0_138_958 ();
 DECAPx6_ASAP7_75t_R FILLER_0_138_970 ();
 DECAPx2_ASAP7_75t_R FILLER_0_138_992 ();
 FILLER_ASAP7_75t_R FILLER_0_138_998 ();
 DECAPx6_ASAP7_75t_R FILLER_0_138_1007 ();
 DECAPx2_ASAP7_75t_R FILLER_0_138_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_1037 ();
 DECAPx1_ASAP7_75t_R FILLER_0_138_1044 ();
 DECAPx6_ASAP7_75t_R FILLER_0_138_1054 ();
 DECAPx2_ASAP7_75t_R FILLER_0_138_1068 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_1074 ();
 FILLER_ASAP7_75t_R FILLER_0_138_1078 ();
 DECAPx2_ASAP7_75t_R FILLER_0_138_1086 ();
 DECAPx2_ASAP7_75t_R FILLER_0_138_1098 ();
 DECAPx2_ASAP7_75t_R FILLER_0_138_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_1113 ();
 DECAPx2_ASAP7_75t_R FILLER_0_138_1120 ();
 FILLER_ASAP7_75t_R FILLER_0_138_1148 ();
 FILLER_ASAP7_75t_R FILLER_0_138_1160 ();
 FILLER_ASAP7_75t_R FILLER_0_138_1172 ();
 FILLER_ASAP7_75t_R FILLER_0_138_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_138_1205 ();
 DECAPx2_ASAP7_75t_R FILLER_0_138_1213 ();
 FILLER_ASAP7_75t_R FILLER_0_138_1219 ();
 FILLER_ASAP7_75t_R FILLER_0_138_1228 ();
 FILLER_ASAP7_75t_R FILLER_0_138_1235 ();
 DECAPx4_ASAP7_75t_R FILLER_0_138_1242 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_1252 ();
 FILLER_ASAP7_75t_R FILLER_0_138_1259 ();
 DECAPx2_ASAP7_75t_R FILLER_0_138_1267 ();
 FILLER_ASAP7_75t_R FILLER_0_138_1273 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_1275 ();
 DECAPx2_ASAP7_75t_R FILLER_0_138_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_1292 ();
 FILLER_ASAP7_75t_R FILLER_0_138_1301 ();
 DECAPx2_ASAP7_75t_R FILLER_0_138_1308 ();
 FILLER_ASAP7_75t_R FILLER_0_138_1314 ();
 DECAPx4_ASAP7_75t_R FILLER_0_138_1326 ();
 FILLER_ASAP7_75t_R FILLER_0_138_1342 ();
 FILLER_ASAP7_75t_R FILLER_0_138_1350 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_1352 ();
 FILLER_ASAP7_75t_R FILLER_0_138_1356 ();
 FILLER_ASAP7_75t_R FILLER_0_138_1363 ();
 DECAPx1_ASAP7_75t_R FILLER_0_138_1371 ();
 FILLER_ASAP7_75t_R FILLER_0_138_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_139_2 ();
 FILLER_ASAP7_75t_R FILLER_0_139_9 ();
 FILLER_ASAP7_75t_R FILLER_0_139_33 ();
 FILLER_ASAP7_75t_R FILLER_0_139_40 ();
 FILLER_ASAP7_75t_R FILLER_0_139_46 ();
 DECAPx6_ASAP7_75t_R FILLER_0_139_51 ();
 FILLER_ASAP7_75t_R FILLER_0_139_65 ();
 DECAPx1_ASAP7_75t_R FILLER_0_139_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_76 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_85 ();
 FILLER_ASAP7_75t_R FILLER_0_139_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_93 ();
 FILLER_ASAP7_75t_R FILLER_0_139_104 ();
 DECAPx6_ASAP7_75t_R FILLER_0_139_117 ();
 FILLER_ASAP7_75t_R FILLER_0_139_143 ();
 FILLER_ASAP7_75t_R FILLER_0_139_153 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_171 ();
 FILLER_ASAP7_75t_R FILLER_0_139_178 ();
 FILLER_ASAP7_75t_R FILLER_0_139_190 ();
 DECAPx4_ASAP7_75t_R FILLER_0_139_212 ();
 FILLER_ASAP7_75t_R FILLER_0_139_222 ();
 FILLER_ASAP7_75t_R FILLER_0_139_236 ();
 DECAPx6_ASAP7_75t_R FILLER_0_139_246 ();
 DECAPx6_ASAP7_75t_R FILLER_0_139_263 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_283 ();
 FILLER_ASAP7_75t_R FILLER_0_139_290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_304 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_317 ();
 FILLER_ASAP7_75t_R FILLER_0_139_328 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_336 ();
 FILLER_ASAP7_75t_R FILLER_0_139_342 ();
 FILLER_ASAP7_75t_R FILLER_0_139_350 ();
 FILLER_ASAP7_75t_R FILLER_0_139_357 ();
 FILLER_ASAP7_75t_R FILLER_0_139_369 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_377 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_389 ();
 FILLER_ASAP7_75t_R FILLER_0_139_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_397 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_404 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_416 ();
 FILLER_ASAP7_75t_R FILLER_0_139_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_424 ();
 FILLER_ASAP7_75t_R FILLER_0_139_431 ();
 DECAPx6_ASAP7_75t_R FILLER_0_139_441 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_455 ();
 FILLER_ASAP7_75t_R FILLER_0_139_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_139_514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_139_528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_544 ();
 DECAPx1_ASAP7_75t_R FILLER_0_139_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_555 ();
 DECAPx4_ASAP7_75t_R FILLER_0_139_568 ();
 FILLER_ASAP7_75t_R FILLER_0_139_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_580 ();
 FILLER_ASAP7_75t_R FILLER_0_139_593 ();
 FILLER_ASAP7_75t_R FILLER_0_139_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_609 ();
 DECAPx6_ASAP7_75t_R FILLER_0_139_622 ();
 FILLER_ASAP7_75t_R FILLER_0_139_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_638 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_650 ();
 FILLER_ASAP7_75t_R FILLER_0_139_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_658 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_665 ();
 FILLER_ASAP7_75t_R FILLER_0_139_681 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_688 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_710 ();
 FILLER_ASAP7_75t_R FILLER_0_139_719 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_727 ();
 FILLER_ASAP7_75t_R FILLER_0_139_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_735 ();
 FILLER_ASAP7_75t_R FILLER_0_139_743 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_757 ();
 FILLER_ASAP7_75t_R FILLER_0_139_765 ();
 FILLER_ASAP7_75t_R FILLER_0_139_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_776 ();
 FILLER_ASAP7_75t_R FILLER_0_139_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_789 ();
 FILLER_ASAP7_75t_R FILLER_0_139_800 ();
 FILLER_ASAP7_75t_R FILLER_0_139_812 ();
 FILLER_ASAP7_75t_R FILLER_0_139_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_826 ();
 FILLER_ASAP7_75t_R FILLER_0_139_833 ();
 FILLER_ASAP7_75t_R FILLER_0_139_840 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_852 ();
 FILLER_ASAP7_75t_R FILLER_0_139_858 ();
 FILLER_ASAP7_75t_R FILLER_0_139_870 ();
 DECAPx1_ASAP7_75t_R FILLER_0_139_877 ();
 FILLER_ASAP7_75t_R FILLER_0_139_891 ();
 FILLER_ASAP7_75t_R FILLER_0_139_896 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_910 ();
 FILLER_ASAP7_75t_R FILLER_0_139_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_919 ();
 FILLER_ASAP7_75t_R FILLER_0_139_923 ();
 FILLER_ASAP7_75t_R FILLER_0_139_927 ();
 DECAPx1_ASAP7_75t_R FILLER_0_139_937 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_947 ();
 FILLER_ASAP7_75t_R FILLER_0_139_953 ();
 FILLER_ASAP7_75t_R FILLER_0_139_963 ();
 FILLER_ASAP7_75t_R FILLER_0_139_973 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_991 ();
 FILLER_ASAP7_75t_R FILLER_0_139_999 ();
 DECAPx4_ASAP7_75t_R FILLER_0_139_1008 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_1020 ();
 DECAPx1_ASAP7_75t_R FILLER_0_139_1032 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1042 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_1055 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_1079 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1092 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_1100 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1106 ();
 DECAPx6_ASAP7_75t_R FILLER_0_139_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_1125 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1131 ();
 DECAPx1_ASAP7_75t_R FILLER_0_139_1136 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1145 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1157 ();
 DECAPx1_ASAP7_75t_R FILLER_0_139_1164 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1182 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1194 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1206 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1211 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1219 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1231 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1239 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1247 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1255 ();
 DECAPx4_ASAP7_75t_R FILLER_0_139_1260 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_1272 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1283 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1295 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1303 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_1305 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1313 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_1315 ();
 DECAPx4_ASAP7_75t_R FILLER_0_139_1326 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1342 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_1344 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1350 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_139_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_140_2 ();
 FILLER_ASAP7_75t_R FILLER_0_140_7 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_12 ();
 FILLER_ASAP7_75t_R FILLER_0_140_18 ();
 FILLER_ASAP7_75t_R FILLER_0_140_26 ();
 FILLER_ASAP7_75t_R FILLER_0_140_34 ();
 FILLER_ASAP7_75t_R FILLER_0_140_42 ();
 FILLER_ASAP7_75t_R FILLER_0_140_47 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_55 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_71 ();
 FILLER_ASAP7_75t_R FILLER_0_140_77 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_89 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_111 ();
 FILLER_ASAP7_75t_R FILLER_0_140_117 ();
 DECAPx6_ASAP7_75t_R FILLER_0_140_122 ();
 FILLER_ASAP7_75t_R FILLER_0_140_136 ();
 FILLER_ASAP7_75t_R FILLER_0_140_144 ();
 FILLER_ASAP7_75t_R FILLER_0_140_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_154 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_165 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_197 ();
 FILLER_ASAP7_75t_R FILLER_0_140_206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_214 ();
 DECAPx1_ASAP7_75t_R FILLER_0_140_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_240 ();
 DECAPx4_ASAP7_75t_R FILLER_0_140_249 ();
 FILLER_ASAP7_75t_R FILLER_0_140_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_261 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_268 ();
 FILLER_ASAP7_75t_R FILLER_0_140_285 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_301 ();
 FILLER_ASAP7_75t_R FILLER_0_140_324 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_344 ();
 DECAPx4_ASAP7_75t_R FILLER_0_140_351 ();
 FILLER_ASAP7_75t_R FILLER_0_140_367 ();
 FILLER_ASAP7_75t_R FILLER_0_140_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_379 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_386 ();
 FILLER_ASAP7_75t_R FILLER_0_140_392 ();
 FILLER_ASAP7_75t_R FILLER_0_140_400 ();
 FILLER_ASAP7_75t_R FILLER_0_140_408 ();
 DECAPx1_ASAP7_75t_R FILLER_0_140_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_421 ();
 FILLER_ASAP7_75t_R FILLER_0_140_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_430 ();
 FILLER_ASAP7_75t_R FILLER_0_140_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_439 ();
 DECAPx6_ASAP7_75t_R FILLER_0_140_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_461 ();
 DECAPx4_ASAP7_75t_R FILLER_0_140_464 ();
 DECAPx6_ASAP7_75t_R FILLER_0_140_480 ();
 FILLER_ASAP7_75t_R FILLER_0_140_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_496 ();
 FILLER_ASAP7_75t_R FILLER_0_140_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_511 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_524 ();
 FILLER_ASAP7_75t_R FILLER_0_140_530 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_538 ();
 FILLER_ASAP7_75t_R FILLER_0_140_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_546 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_561 ();
 FILLER_ASAP7_75t_R FILLER_0_140_574 ();
 FILLER_ASAP7_75t_R FILLER_0_140_588 ();
 FILLER_ASAP7_75t_R FILLER_0_140_602 ();
 FILLER_ASAP7_75t_R FILLER_0_140_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_618 ();
 DECAPx1_ASAP7_75t_R FILLER_0_140_631 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_647 ();
 FILLER_ASAP7_75t_R FILLER_0_140_653 ();
 FILLER_ASAP7_75t_R FILLER_0_140_675 ();
 FILLER_ASAP7_75t_R FILLER_0_140_687 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_700 ();
 FILLER_ASAP7_75t_R FILLER_0_140_707 ();
 DECAPx1_ASAP7_75t_R FILLER_0_140_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_717 ();
 FILLER_ASAP7_75t_R FILLER_0_140_724 ();
 DECAPx1_ASAP7_75t_R FILLER_0_140_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_733 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_740 ();
 FILLER_ASAP7_75t_R FILLER_0_140_746 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_755 ();
 DECAPx1_ASAP7_75t_R FILLER_0_140_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_781 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_793 ();
 FILLER_ASAP7_75t_R FILLER_0_140_800 ();
 FILLER_ASAP7_75t_R FILLER_0_140_812 ();
 FILLER_ASAP7_75t_R FILLER_0_140_820 ();
 FILLER_ASAP7_75t_R FILLER_0_140_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_834 ();
 FILLER_ASAP7_75t_R FILLER_0_140_845 ();
 FILLER_ASAP7_75t_R FILLER_0_140_857 ();
 FILLER_ASAP7_75t_R FILLER_0_140_869 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_885 ();
 FILLER_ASAP7_75t_R FILLER_0_140_896 ();
 FILLER_ASAP7_75t_R FILLER_0_140_906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_916 ();
 DECAPx1_ASAP7_75t_R FILLER_0_140_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_942 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_961 ();
 DECAPx1_ASAP7_75t_R FILLER_0_140_970 ();
 FILLER_ASAP7_75t_R FILLER_0_140_980 ();
 FILLER_ASAP7_75t_R FILLER_0_140_990 ();
 DECAPx1_ASAP7_75t_R FILLER_0_140_999 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_1011 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_1033 ();
 FILLER_ASAP7_75t_R FILLER_0_140_1045 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_1053 ();
 FILLER_ASAP7_75t_R FILLER_0_140_1067 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_1080 ();
 FILLER_ASAP7_75t_R FILLER_0_140_1096 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_1104 ();
 FILLER_ASAP7_75t_R FILLER_0_140_1116 ();
 FILLER_ASAP7_75t_R FILLER_0_140_1129 ();
 DECAPx4_ASAP7_75t_R FILLER_0_140_1139 ();
 FILLER_ASAP7_75t_R FILLER_0_140_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_1151 ();
 FILLER_ASAP7_75t_R FILLER_0_140_1162 ();
 FILLER_ASAP7_75t_R FILLER_0_140_1174 ();
 FILLER_ASAP7_75t_R FILLER_0_140_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_140_1198 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_1210 ();
 FILLER_ASAP7_75t_R FILLER_0_140_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_1224 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_1246 ();
 FILLER_ASAP7_75t_R FILLER_0_140_1257 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_1265 ();
 FILLER_ASAP7_75t_R FILLER_0_140_1281 ();
 FILLER_ASAP7_75t_R FILLER_0_140_1293 ();
 DECAPx1_ASAP7_75t_R FILLER_0_140_1301 ();
 DECAPx1_ASAP7_75t_R FILLER_0_140_1315 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_1319 ();
 FILLER_ASAP7_75t_R FILLER_0_140_1326 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_1328 ();
 FILLER_ASAP7_75t_R FILLER_0_140_1335 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_1337 ();
 FILLER_ASAP7_75t_R FILLER_0_140_1344 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_1346 ();
 FILLER_ASAP7_75t_R FILLER_0_140_1350 ();
 FILLER_ASAP7_75t_R FILLER_0_140_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_140_1364 ();
 FILLER_ASAP7_75t_R FILLER_0_140_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_1374 ();
 FILLER_ASAP7_75t_R FILLER_0_140_1380 ();
 DECAPx6_ASAP7_75t_R FILLER_0_141_2 ();
 FILLER_ASAP7_75t_R FILLER_0_141_21 ();
 DECAPx1_ASAP7_75t_R FILLER_0_141_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_48 ();
 FILLER_ASAP7_75t_R FILLER_0_141_55 ();
 DECAPx6_ASAP7_75t_R FILLER_0_141_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_79 ();
 DECAPx1_ASAP7_75t_R FILLER_0_141_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_94 ();
 DECAPx1_ASAP7_75t_R FILLER_0_141_105 ();
 FILLER_ASAP7_75t_R FILLER_0_141_112 ();
 FILLER_ASAP7_75t_R FILLER_0_141_122 ();
 FILLER_ASAP7_75t_R FILLER_0_141_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_143 ();
 DECAPx6_ASAP7_75t_R FILLER_0_141_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_179 ();
 DECAPx4_ASAP7_75t_R FILLER_0_141_191 ();
 DECAPx1_ASAP7_75t_R FILLER_0_141_211 ();
 DECAPx6_ASAP7_75t_R FILLER_0_141_226 ();
 DECAPx2_ASAP7_75t_R FILLER_0_141_240 ();
 DECAPx2_ASAP7_75t_R FILLER_0_141_249 ();
 FILLER_ASAP7_75t_R FILLER_0_141_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_257 ();
 DECAPx6_ASAP7_75t_R FILLER_0_141_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_278 ();
 FILLER_ASAP7_75t_R FILLER_0_141_289 ();
 FILLER_ASAP7_75t_R FILLER_0_141_301 ();
 FILLER_ASAP7_75t_R FILLER_0_141_308 ();
 FILLER_ASAP7_75t_R FILLER_0_141_320 ();
 FILLER_ASAP7_75t_R FILLER_0_141_332 ();
 FILLER_ASAP7_75t_R FILLER_0_141_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_342 ();
 DECAPx1_ASAP7_75t_R FILLER_0_141_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_353 ();
 FILLER_ASAP7_75t_R FILLER_0_141_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_366 ();
 FILLER_ASAP7_75t_R FILLER_0_141_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_375 ();
 DECAPx1_ASAP7_75t_R FILLER_0_141_396 ();
 DECAPx1_ASAP7_75t_R FILLER_0_141_407 ();
 DECAPx1_ASAP7_75t_R FILLER_0_141_417 ();
 FILLER_ASAP7_75t_R FILLER_0_141_441 ();
 FILLER_ASAP7_75t_R FILLER_0_141_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_451 ();
 DECAPx4_ASAP7_75t_R FILLER_0_141_458 ();
 FILLER_ASAP7_75t_R FILLER_0_141_468 ();
 DECAPx1_ASAP7_75t_R FILLER_0_141_491 ();
 DECAPx2_ASAP7_75t_R FILLER_0_141_507 ();
 DECAPx2_ASAP7_75t_R FILLER_0_141_525 ();
 DECAPx2_ASAP7_75t_R FILLER_0_141_539 ();
 DECAPx2_ASAP7_75t_R FILLER_0_141_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_572 ();
 DECAPx4_ASAP7_75t_R FILLER_0_141_585 ();
 FILLER_ASAP7_75t_R FILLER_0_141_595 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_608 ();
 DECAPx2_ASAP7_75t_R FILLER_0_141_630 ();
 FILLER_ASAP7_75t_R FILLER_0_141_636 ();
 DECAPx2_ASAP7_75t_R FILLER_0_141_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_656 ();
 DECAPx2_ASAP7_75t_R FILLER_0_141_664 ();
 FILLER_ASAP7_75t_R FILLER_0_141_670 ();
 FILLER_ASAP7_75t_R FILLER_0_141_682 ();
 FILLER_ASAP7_75t_R FILLER_0_141_694 ();
 DECAPx2_ASAP7_75t_R FILLER_0_141_701 ();
 FILLER_ASAP7_75t_R FILLER_0_141_715 ();
 DECAPx4_ASAP7_75t_R FILLER_0_141_723 ();
 FILLER_ASAP7_75t_R FILLER_0_141_733 ();
 FILLER_ASAP7_75t_R FILLER_0_141_755 ();
 FILLER_ASAP7_75t_R FILLER_0_141_769 ();
 DECAPx1_ASAP7_75t_R FILLER_0_141_777 ();
 FILLER_ASAP7_75t_R FILLER_0_141_788 ();
 DECAPx1_ASAP7_75t_R FILLER_0_141_798 ();
 FILLER_ASAP7_75t_R FILLER_0_141_808 ();
 FILLER_ASAP7_75t_R FILLER_0_141_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_815 ();
 FILLER_ASAP7_75t_R FILLER_0_141_826 ();
 FILLER_ASAP7_75t_R FILLER_0_141_838 ();
 FILLER_ASAP7_75t_R FILLER_0_141_848 ();
 DECAPx2_ASAP7_75t_R FILLER_0_141_855 ();
 FILLER_ASAP7_75t_R FILLER_0_141_861 ();
 FILLER_ASAP7_75t_R FILLER_0_141_873 ();
 FILLER_ASAP7_75t_R FILLER_0_141_885 ();
 DECAPx1_ASAP7_75t_R FILLER_0_141_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_897 ();
 DECAPx6_ASAP7_75t_R FILLER_0_141_906 ();
 DECAPx1_ASAP7_75t_R FILLER_0_141_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_924 ();
 DECAPx6_ASAP7_75t_R FILLER_0_141_927 ();
 FILLER_ASAP7_75t_R FILLER_0_141_941 ();
 FILLER_ASAP7_75t_R FILLER_0_141_953 ();
 DECAPx6_ASAP7_75t_R FILLER_0_141_961 ();
 DECAPx4_ASAP7_75t_R FILLER_0_141_980 ();
 FILLER_ASAP7_75t_R FILLER_0_141_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_992 ();
 FILLER_ASAP7_75t_R FILLER_0_141_1001 ();
 FILLER_ASAP7_75t_R FILLER_0_141_1011 ();
 FILLER_ASAP7_75t_R FILLER_0_141_1016 ();
 DECAPx6_ASAP7_75t_R FILLER_0_141_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_1043 ();
 DECAPx6_ASAP7_75t_R FILLER_0_141_1050 ();
 DECAPx1_ASAP7_75t_R FILLER_0_141_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_1079 ();
 DECAPx2_ASAP7_75t_R FILLER_0_141_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_1094 ();
 DECAPx2_ASAP7_75t_R FILLER_0_141_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_1113 ();
 DECAPx2_ASAP7_75t_R FILLER_0_141_1122 ();
 DECAPx4_ASAP7_75t_R FILLER_0_141_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_1145 ();
 FILLER_ASAP7_75t_R FILLER_0_141_1151 ();
 FILLER_ASAP7_75t_R FILLER_0_141_1159 ();
 FILLER_ASAP7_75t_R FILLER_0_141_1169 ();
 DECAPx2_ASAP7_75t_R FILLER_0_141_1181 ();
 FILLER_ASAP7_75t_R FILLER_0_141_1187 ();
 FILLER_ASAP7_75t_R FILLER_0_141_1200 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_1202 ();
 FILLER_ASAP7_75t_R FILLER_0_141_1210 ();
 FILLER_ASAP7_75t_R FILLER_0_141_1218 ();
 DECAPx4_ASAP7_75t_R FILLER_0_141_1226 ();
 FILLER_ASAP7_75t_R FILLER_0_141_1236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_1248 ();
 DECAPx2_ASAP7_75t_R FILLER_0_141_1270 ();
 DECAPx2_ASAP7_75t_R FILLER_0_141_1286 ();
 FILLER_ASAP7_75t_R FILLER_0_141_1292 ();
 FILLER_ASAP7_75t_R FILLER_0_141_1300 ();
 DECAPx2_ASAP7_75t_R FILLER_0_141_1308 ();
 FILLER_ASAP7_75t_R FILLER_0_141_1314 ();
 FILLER_ASAP7_75t_R FILLER_0_141_1328 ();
 FILLER_ASAP7_75t_R FILLER_0_141_1336 ();
 FILLER_ASAP7_75t_R FILLER_0_141_1341 ();
 DECAPx1_ASAP7_75t_R FILLER_0_141_1349 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_1353 ();
 DECAPx2_ASAP7_75t_R FILLER_0_141_1376 ();
 DECAPx4_ASAP7_75t_R FILLER_0_142_2 ();
 FILLER_ASAP7_75t_R FILLER_0_142_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_14 ();
 FILLER_ASAP7_75t_R FILLER_0_142_18 ();
 FILLER_ASAP7_75t_R FILLER_0_142_26 ();
 FILLER_ASAP7_75t_R FILLER_0_142_34 ();
 DECAPx4_ASAP7_75t_R FILLER_0_142_42 ();
 FILLER_ASAP7_75t_R FILLER_0_142_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_54 ();
 DECAPx6_ASAP7_75t_R FILLER_0_142_63 ();
 DECAPx2_ASAP7_75t_R FILLER_0_142_77 ();
 FILLER_ASAP7_75t_R FILLER_0_142_94 ();
 DECAPx2_ASAP7_75t_R FILLER_0_142_104 ();
 FILLER_ASAP7_75t_R FILLER_0_142_110 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_123 ();
 DECAPx2_ASAP7_75t_R FILLER_0_142_145 ();
 FILLER_ASAP7_75t_R FILLER_0_142_151 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_165 ();
 DECAPx4_ASAP7_75t_R FILLER_0_142_187 ();
 DECAPx1_ASAP7_75t_R FILLER_0_142_201 ();
 DECAPx1_ASAP7_75t_R FILLER_0_142_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_215 ();
 DECAPx6_ASAP7_75t_R FILLER_0_142_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_236 ();
 DECAPx4_ASAP7_75t_R FILLER_0_142_248 ();
 FILLER_ASAP7_75t_R FILLER_0_142_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_260 ();
 DECAPx2_ASAP7_75t_R FILLER_0_142_267 ();
 FILLER_ASAP7_75t_R FILLER_0_142_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_275 ();
 DECAPx6_ASAP7_75t_R FILLER_0_142_286 ();
 DECAPx1_ASAP7_75t_R FILLER_0_142_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_304 ();
 FILLER_ASAP7_75t_R FILLER_0_142_316 ();
 FILLER_ASAP7_75t_R FILLER_0_142_322 ();
 FILLER_ASAP7_75t_R FILLER_0_142_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_336 ();
 FILLER_ASAP7_75t_R FILLER_0_142_343 ();
 FILLER_ASAP7_75t_R FILLER_0_142_352 ();
 FILLER_ASAP7_75t_R FILLER_0_142_360 ();
 FILLER_ASAP7_75t_R FILLER_0_142_369 ();
 DECAPx1_ASAP7_75t_R FILLER_0_142_377 ();
 DECAPx6_ASAP7_75t_R FILLER_0_142_388 ();
 DECAPx1_ASAP7_75t_R FILLER_0_142_402 ();
 FILLER_ASAP7_75t_R FILLER_0_142_412 ();
 FILLER_ASAP7_75t_R FILLER_0_142_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_421 ();
 FILLER_ASAP7_75t_R FILLER_0_142_442 ();
 FILLER_ASAP7_75t_R FILLER_0_142_450 ();
 DECAPx1_ASAP7_75t_R FILLER_0_142_458 ();
 DECAPx1_ASAP7_75t_R FILLER_0_142_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_468 ();
 FILLER_ASAP7_75t_R FILLER_0_142_474 ();
 FILLER_ASAP7_75t_R FILLER_0_142_479 ();
 FILLER_ASAP7_75t_R FILLER_0_142_486 ();
 DECAPx1_ASAP7_75t_R FILLER_0_142_494 ();
 DECAPx4_ASAP7_75t_R FILLER_0_142_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_520 ();
 DECAPx1_ASAP7_75t_R FILLER_0_142_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_533 ();
 FILLER_ASAP7_75t_R FILLER_0_142_545 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_550 ();
 DECAPx1_ASAP7_75t_R FILLER_0_142_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_632 ();
 FILLER_ASAP7_75t_R FILLER_0_142_645 ();
 DECAPx1_ASAP7_75t_R FILLER_0_142_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_663 ();
 FILLER_ASAP7_75t_R FILLER_0_142_668 ();
 FILLER_ASAP7_75t_R FILLER_0_142_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_682 ();
 DECAPx2_ASAP7_75t_R FILLER_0_142_693 ();
 FILLER_ASAP7_75t_R FILLER_0_142_709 ();
 FILLER_ASAP7_75t_R FILLER_0_142_719 ();
 DECAPx2_ASAP7_75t_R FILLER_0_142_726 ();
 DECAPx2_ASAP7_75t_R FILLER_0_142_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_744 ();
 FILLER_ASAP7_75t_R FILLER_0_142_755 ();
 FILLER_ASAP7_75t_R FILLER_0_142_765 ();
 DECAPx2_ASAP7_75t_R FILLER_0_142_777 ();
 FILLER_ASAP7_75t_R FILLER_0_142_783 ();
 FILLER_ASAP7_75t_R FILLER_0_142_795 ();
 FILLER_ASAP7_75t_R FILLER_0_142_807 ();
 FILLER_ASAP7_75t_R FILLER_0_142_819 ();
 FILLER_ASAP7_75t_R FILLER_0_142_829 ();
 FILLER_ASAP7_75t_R FILLER_0_142_838 ();
 FILLER_ASAP7_75t_R FILLER_0_142_847 ();
 FILLER_ASAP7_75t_R FILLER_0_142_855 ();
 DECAPx1_ASAP7_75t_R FILLER_0_142_862 ();
 FILLER_ASAP7_75t_R FILLER_0_142_876 ();
 FILLER_ASAP7_75t_R FILLER_0_142_884 ();
 FILLER_ASAP7_75t_R FILLER_0_142_891 ();
 FILLER_ASAP7_75t_R FILLER_0_142_898 ();
 DECAPx6_ASAP7_75t_R FILLER_0_142_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_919 ();
 DECAPx1_ASAP7_75t_R FILLER_0_142_930 ();
 FILLER_ASAP7_75t_R FILLER_0_142_955 ();
 DECAPx6_ASAP7_75t_R FILLER_0_142_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_974 ();
 FILLER_ASAP7_75t_R FILLER_0_142_986 ();
 DECAPx1_ASAP7_75t_R FILLER_0_142_999 ();
 DECAPx2_ASAP7_75t_R FILLER_0_142_1011 ();
 FILLER_ASAP7_75t_R FILLER_0_142_1017 ();
 DECAPx4_ASAP7_75t_R FILLER_0_142_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_1041 ();
 DECAPx6_ASAP7_75t_R FILLER_0_142_1050 ();
 DECAPx2_ASAP7_75t_R FILLER_0_142_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_1070 ();
 FILLER_ASAP7_75t_R FILLER_0_142_1076 ();
 DECAPx6_ASAP7_75t_R FILLER_0_142_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_1102 ();
 FILLER_ASAP7_75t_R FILLER_0_142_1115 ();
 DECAPx2_ASAP7_75t_R FILLER_0_142_1123 ();
 FILLER_ASAP7_75t_R FILLER_0_142_1129 ();
 DECAPx4_ASAP7_75t_R FILLER_0_142_1139 ();
 FILLER_ASAP7_75t_R FILLER_0_142_1154 ();
 FILLER_ASAP7_75t_R FILLER_0_142_1162 ();
 DECAPx2_ASAP7_75t_R FILLER_0_142_1170 ();
 DECAPx1_ASAP7_75t_R FILLER_0_142_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_142_1201 ();
 FILLER_ASAP7_75t_R FILLER_0_142_1209 ();
 DECAPx2_ASAP7_75t_R FILLER_0_142_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_1223 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_1235 ();
 DECAPx1_ASAP7_75t_R FILLER_0_142_1257 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_1261 ();
 FILLER_ASAP7_75t_R FILLER_0_142_1272 ();
 FILLER_ASAP7_75t_R FILLER_0_142_1279 ();
 FILLER_ASAP7_75t_R FILLER_0_142_1286 ();
 DECAPx2_ASAP7_75t_R FILLER_0_142_1293 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_1299 ();
 DECAPx1_ASAP7_75t_R FILLER_0_142_1306 ();
 FILLER_ASAP7_75t_R FILLER_0_142_1320 ();
 DECAPx1_ASAP7_75t_R FILLER_0_142_1329 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_1333 ();
 DECAPx1_ASAP7_75t_R FILLER_0_142_1354 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_1358 ();
 FILLER_ASAP7_75t_R FILLER_0_142_1364 ();
 FILLER_ASAP7_75t_R FILLER_0_142_1371 ();
 DECAPx1_ASAP7_75t_R FILLER_0_142_1378 ();
 DECAPx2_ASAP7_75t_R FILLER_0_143_2 ();
 FILLER_ASAP7_75t_R FILLER_0_143_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143_10 ();
 DECAPx1_ASAP7_75t_R FILLER_0_143_16 ();
 FILLER_ASAP7_75t_R FILLER_0_143_41 ();
 DECAPx6_ASAP7_75t_R FILLER_0_143_48 ();
 FILLER_ASAP7_75t_R FILLER_0_143_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_70 ();
 DECAPx1_ASAP7_75t_R FILLER_0_143_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143_96 ();
 FILLER_ASAP7_75t_R FILLER_0_143_103 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_111 ();
 FILLER_ASAP7_75t_R FILLER_0_143_133 ();
 DECAPx6_ASAP7_75t_R FILLER_0_143_142 ();
 FILLER_ASAP7_75t_R FILLER_0_143_156 ();
 DECAPx1_ASAP7_75t_R FILLER_0_143_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143_168 ();
 FILLER_ASAP7_75t_R FILLER_0_143_177 ();
 DECAPx1_ASAP7_75t_R FILLER_0_143_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143_194 ();
 FILLER_ASAP7_75t_R FILLER_0_143_201 ();
 DECAPx2_ASAP7_75t_R FILLER_0_143_209 ();
 FILLER_ASAP7_75t_R FILLER_0_143_215 ();
 DECAPx6_ASAP7_75t_R FILLER_0_143_225 ();
 FILLER_ASAP7_75t_R FILLER_0_143_239 ();
 FILLER_ASAP7_75t_R FILLER_0_143_252 ();
 FILLER_ASAP7_75t_R FILLER_0_143_257 ();
 DECAPx4_ASAP7_75t_R FILLER_0_143_267 ();
 FILLER_ASAP7_75t_R FILLER_0_143_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143_279 ();
 DECAPx1_ASAP7_75t_R FILLER_0_143_286 ();
 DECAPx4_ASAP7_75t_R FILLER_0_143_300 ();
 FILLER_ASAP7_75t_R FILLER_0_143_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143_312 ();
 FILLER_ASAP7_75t_R FILLER_0_143_327 ();
 DECAPx2_ASAP7_75t_R FILLER_0_143_349 ();
 FILLER_ASAP7_75t_R FILLER_0_143_360 ();
 FILLER_ASAP7_75t_R FILLER_0_143_367 ();
 FILLER_ASAP7_75t_R FILLER_0_143_379 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_387 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_409 ();
 FILLER_ASAP7_75t_R FILLER_0_143_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143_433 ();
 FILLER_ASAP7_75t_R FILLER_0_143_440 ();
 FILLER_ASAP7_75t_R FILLER_0_143_448 ();
 DECAPx1_ASAP7_75t_R FILLER_0_143_458 ();
 DECAPx6_ASAP7_75t_R FILLER_0_143_468 ();
 DECAPx1_ASAP7_75t_R FILLER_0_143_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143_486 ();
 DECAPx4_ASAP7_75t_R FILLER_0_143_508 ();
 FILLER_ASAP7_75t_R FILLER_0_143_518 ();
 FILLER_ASAP7_75t_R FILLER_0_143_541 ();
 DECAPx2_ASAP7_75t_R FILLER_0_143_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143_552 ();
 DECAPx6_ASAP7_75t_R FILLER_0_143_574 ();
 DECAPx2_ASAP7_75t_R FILLER_0_143_588 ();
 FILLER_ASAP7_75t_R FILLER_0_143_615 ();
 DECAPx2_ASAP7_75t_R FILLER_0_143_629 ();
 FILLER_ASAP7_75t_R FILLER_0_143_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143_637 ();
 FILLER_ASAP7_75t_R FILLER_0_143_650 ();
 DECAPx1_ASAP7_75t_R FILLER_0_143_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143_667 ();
 FILLER_ASAP7_75t_R FILLER_0_143_675 ();
 DECAPx1_ASAP7_75t_R FILLER_0_143_687 ();
 FILLER_ASAP7_75t_R FILLER_0_143_696 ();
 FILLER_ASAP7_75t_R FILLER_0_143_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143_710 ();
 FILLER_ASAP7_75t_R FILLER_0_143_721 ();
 FILLER_ASAP7_75t_R FILLER_0_143_728 ();
 FILLER_ASAP7_75t_R FILLER_0_143_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143_742 ();
 DECAPx4_ASAP7_75t_R FILLER_0_143_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143_763 ();
 DECAPx1_ASAP7_75t_R FILLER_0_143_774 ();
 FILLER_ASAP7_75t_R FILLER_0_143_783 ();
 FILLER_ASAP7_75t_R FILLER_0_143_795 ();
 FILLER_ASAP7_75t_R FILLER_0_143_807 ();
 FILLER_ASAP7_75t_R FILLER_0_143_819 ();
 FILLER_ASAP7_75t_R FILLER_0_143_831 ();
 FILLER_ASAP7_75t_R FILLER_0_143_838 ();
 FILLER_ASAP7_75t_R FILLER_0_143_852 ();
 DECAPx2_ASAP7_75t_R FILLER_0_143_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143_870 ();
 FILLER_ASAP7_75t_R FILLER_0_143_885 ();
 FILLER_ASAP7_75t_R FILLER_0_143_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143_899 ();
 DECAPx4_ASAP7_75t_R FILLER_0_143_906 ();
 FILLER_ASAP7_75t_R FILLER_0_143_916 ();
 FILLER_ASAP7_75t_R FILLER_0_143_923 ();
 FILLER_ASAP7_75t_R FILLER_0_143_927 ();
 FILLER_ASAP7_75t_R FILLER_0_143_947 ();
 DECAPx1_ASAP7_75t_R FILLER_0_143_955 ();
 DECAPx6_ASAP7_75t_R FILLER_0_143_969 ();
 DECAPx1_ASAP7_75t_R FILLER_0_143_983 ();
 DECAPx2_ASAP7_75t_R FILLER_0_143_995 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1001 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_1011 ();
 DECAPx2_ASAP7_75t_R FILLER_0_143_1033 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1039 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1047 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1057 ();
 DECAPx4_ASAP7_75t_R FILLER_0_143_1064 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_1082 ();
 DECAPx1_ASAP7_75t_R FILLER_0_143_1104 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1120 ();
 DECAPx4_ASAP7_75t_R FILLER_0_143_1132 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1147 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1154 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1161 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143_1175 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1188 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1200 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1209 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1222 ();
 DECAPx1_ASAP7_75t_R FILLER_0_143_1230 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1240 ();
 DECAPx6_ASAP7_75t_R FILLER_0_143_1248 ();
 DECAPx2_ASAP7_75t_R FILLER_0_143_1262 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143_1268 ();
 DECAPx2_ASAP7_75t_R FILLER_0_143_1275 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143_1281 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1294 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1307 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1314 ();
 DECAPx2_ASAP7_75t_R FILLER_0_143_1322 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1331 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1345 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1353 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143_1355 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1361 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1368 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_143_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_144_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_144_9 ();
 FILLER_ASAP7_75t_R FILLER_0_144_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_17 ();
 FILLER_ASAP7_75t_R FILLER_0_144_21 ();
 FILLER_ASAP7_75t_R FILLER_0_144_45 ();
 FILLER_ASAP7_75t_R FILLER_0_144_55 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_65 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_87 ();
 FILLER_ASAP7_75t_R FILLER_0_144_121 ();
 FILLER_ASAP7_75t_R FILLER_0_144_134 ();
 DECAPx4_ASAP7_75t_R FILLER_0_144_142 ();
 FILLER_ASAP7_75t_R FILLER_0_144_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_154 ();
 DECAPx2_ASAP7_75t_R FILLER_0_144_163 ();
 DECAPx6_ASAP7_75t_R FILLER_0_144_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_191 ();
 DECAPx2_ASAP7_75t_R FILLER_0_144_198 ();
 FILLER_ASAP7_75t_R FILLER_0_144_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_241 ();
 DECAPx1_ASAP7_75t_R FILLER_0_144_248 ();
 DECAPx6_ASAP7_75t_R FILLER_0_144_260 ();
 DECAPx2_ASAP7_75t_R FILLER_0_144_274 ();
 DECAPx4_ASAP7_75t_R FILLER_0_144_290 ();
 FILLER_ASAP7_75t_R FILLER_0_144_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_302 ();
 DECAPx1_ASAP7_75t_R FILLER_0_144_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_313 ();
 FILLER_ASAP7_75t_R FILLER_0_144_320 ();
 DECAPx1_ASAP7_75t_R FILLER_0_144_332 ();
 FILLER_ASAP7_75t_R FILLER_0_144_339 ();
 FILLER_ASAP7_75t_R FILLER_0_144_347 ();
 DECAPx2_ASAP7_75t_R FILLER_0_144_357 ();
 FILLER_ASAP7_75t_R FILLER_0_144_368 ();
 FILLER_ASAP7_75t_R FILLER_0_144_380 ();
 DECAPx6_ASAP7_75t_R FILLER_0_144_386 ();
 DECAPx1_ASAP7_75t_R FILLER_0_144_400 ();
 FILLER_ASAP7_75t_R FILLER_0_144_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_416 ();
 FILLER_ASAP7_75t_R FILLER_0_144_423 ();
 FILLER_ASAP7_75t_R FILLER_0_144_431 ();
 FILLER_ASAP7_75t_R FILLER_0_144_440 ();
 FILLER_ASAP7_75t_R FILLER_0_144_447 ();
 DECAPx1_ASAP7_75t_R FILLER_0_144_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_461 ();
 DECAPx1_ASAP7_75t_R FILLER_0_144_464 ();
 DECAPx6_ASAP7_75t_R FILLER_0_144_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_144_514 ();
 FILLER_ASAP7_75t_R FILLER_0_144_520 ();
 DECAPx4_ASAP7_75t_R FILLER_0_144_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_535 ();
 DECAPx2_ASAP7_75t_R FILLER_0_144_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_554 ();
 DECAPx6_ASAP7_75t_R FILLER_0_144_558 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_572 ();
 DECAPx6_ASAP7_75t_R FILLER_0_144_579 ();
 FILLER_ASAP7_75t_R FILLER_0_144_593 ();
 DECAPx2_ASAP7_75t_R FILLER_0_144_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_612 ();
 FILLER_ASAP7_75t_R FILLER_0_144_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_618 ();
 DECAPx2_ASAP7_75t_R FILLER_0_144_625 ();
 FILLER_ASAP7_75t_R FILLER_0_144_631 ();
 DECAPx4_ASAP7_75t_R FILLER_0_144_645 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_655 ();
 FILLER_ASAP7_75t_R FILLER_0_144_661 ();
 FILLER_ASAP7_75t_R FILLER_0_144_669 ();
 FILLER_ASAP7_75t_R FILLER_0_144_681 ();
 DECAPx1_ASAP7_75t_R FILLER_0_144_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_692 ();
 FILLER_ASAP7_75t_R FILLER_0_144_703 ();
 DECAPx1_ASAP7_75t_R FILLER_0_144_711 ();
 DECAPx2_ASAP7_75t_R FILLER_0_144_725 ();
 FILLER_ASAP7_75t_R FILLER_0_144_731 ();
 FILLER_ASAP7_75t_R FILLER_0_144_743 ();
 DECAPx6_ASAP7_75t_R FILLER_0_144_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_769 ();
 FILLER_ASAP7_75t_R FILLER_0_144_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_778 ();
 FILLER_ASAP7_75t_R FILLER_0_144_789 ();
 FILLER_ASAP7_75t_R FILLER_0_144_801 ();
 DECAPx1_ASAP7_75t_R FILLER_0_144_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_813 ();
 FILLER_ASAP7_75t_R FILLER_0_144_824 ();
 DECAPx1_ASAP7_75t_R FILLER_0_144_836 ();
 DECAPx2_ASAP7_75t_R FILLER_0_144_852 ();
 FILLER_ASAP7_75t_R FILLER_0_144_864 ();
 DECAPx2_ASAP7_75t_R FILLER_0_144_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_877 ();
 FILLER_ASAP7_75t_R FILLER_0_144_898 ();
 DECAPx2_ASAP7_75t_R FILLER_0_144_911 ();
 FILLER_ASAP7_75t_R FILLER_0_144_917 ();
 FILLER_ASAP7_75t_R FILLER_0_144_922 ();
 FILLER_ASAP7_75t_R FILLER_0_144_934 ();
 DECAPx1_ASAP7_75t_R FILLER_0_144_939 ();
 FILLER_ASAP7_75t_R FILLER_0_144_949 ();
 FILLER_ASAP7_75t_R FILLER_0_144_956 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_969 ();
 DECAPx6_ASAP7_75t_R FILLER_0_144_991 ();
 DECAPx6_ASAP7_75t_R FILLER_0_144_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_1027 ();
 DECAPx4_ASAP7_75t_R FILLER_0_144_1049 ();
 FILLER_ASAP7_75t_R FILLER_0_144_1059 ();
 FILLER_ASAP7_75t_R FILLER_0_144_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_1071 ();
 FILLER_ASAP7_75t_R FILLER_0_144_1082 ();
 DECAPx6_ASAP7_75t_R FILLER_0_144_1095 ();
 DECAPx1_ASAP7_75t_R FILLER_0_144_1109 ();
 DECAPx6_ASAP7_75t_R FILLER_0_144_1118 ();
 FILLER_ASAP7_75t_R FILLER_0_144_1132 ();
 FILLER_ASAP7_75t_R FILLER_0_144_1155 ();
 DECAPx1_ASAP7_75t_R FILLER_0_144_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_1167 ();
 FILLER_ASAP7_75t_R FILLER_0_144_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_144_1198 ();
 DECAPx6_ASAP7_75t_R FILLER_0_144_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_1221 ();
 DECAPx2_ASAP7_75t_R FILLER_0_144_1228 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_1234 ();
 DECAPx2_ASAP7_75t_R FILLER_0_144_1241 ();
 FILLER_ASAP7_75t_R FILLER_0_144_1251 ();
 FILLER_ASAP7_75t_R FILLER_0_144_1265 ();
 DECAPx2_ASAP7_75t_R FILLER_0_144_1273 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_1279 ();
 FILLER_ASAP7_75t_R FILLER_0_144_1292 ();
 FILLER_ASAP7_75t_R FILLER_0_144_1304 ();
 FILLER_ASAP7_75t_R FILLER_0_144_1312 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_1314 ();
 FILLER_ASAP7_75t_R FILLER_0_144_1327 ();
 FILLER_ASAP7_75t_R FILLER_0_144_1341 ();
 FILLER_ASAP7_75t_R FILLER_0_144_1351 ();
 FILLER_ASAP7_75t_R FILLER_0_144_1356 ();
 FILLER_ASAP7_75t_R FILLER_0_144_1363 ();
 FILLER_ASAP7_75t_R FILLER_0_144_1370 ();
 DECAPx1_ASAP7_75t_R FILLER_0_144_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_145_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_4 ();
 FILLER_ASAP7_75t_R FILLER_0_145_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_12 ();
 DECAPx2_ASAP7_75t_R FILLER_0_145_17 ();
 FILLER_ASAP7_75t_R FILLER_0_145_23 ();
 DECAPx4_ASAP7_75t_R FILLER_0_145_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_38 ();
 DECAPx2_ASAP7_75t_R FILLER_0_145_42 ();
 FILLER_ASAP7_75t_R FILLER_0_145_48 ();
 FILLER_ASAP7_75t_R FILLER_0_145_56 ();
 DECAPx1_ASAP7_75t_R FILLER_0_145_64 ();
 DECAPx1_ASAP7_75t_R FILLER_0_145_80 ();
 DECAPx1_ASAP7_75t_R FILLER_0_145_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_94 ();
 FILLER_ASAP7_75t_R FILLER_0_145_105 ();
 FILLER_ASAP7_75t_R FILLER_0_145_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_119 ();
 DECAPx1_ASAP7_75t_R FILLER_0_145_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_130 ();
 DECAPx6_ASAP7_75t_R FILLER_0_145_137 ();
 FILLER_ASAP7_75t_R FILLER_0_145_157 ();
 FILLER_ASAP7_75t_R FILLER_0_145_165 ();
 DECAPx2_ASAP7_75t_R FILLER_0_145_170 ();
 FILLER_ASAP7_75t_R FILLER_0_145_176 ();
 FILLER_ASAP7_75t_R FILLER_0_145_190 ();
 FILLER_ASAP7_75t_R FILLER_0_145_202 ();
 DECAPx1_ASAP7_75t_R FILLER_0_145_212 ();
 DECAPx2_ASAP7_75t_R FILLER_0_145_224 ();
 FILLER_ASAP7_75t_R FILLER_0_145_230 ();
 DECAPx1_ASAP7_75t_R FILLER_0_145_238 ();
 DECAPx6_ASAP7_75t_R FILLER_0_145_250 ();
 DECAPx2_ASAP7_75t_R FILLER_0_145_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_270 ();
 FILLER_ASAP7_75t_R FILLER_0_145_295 ();
 FILLER_ASAP7_75t_R FILLER_0_145_300 ();
 DECAPx2_ASAP7_75t_R FILLER_0_145_308 ();
 FILLER_ASAP7_75t_R FILLER_0_145_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_316 ();
 DECAPx2_ASAP7_75t_R FILLER_0_145_329 ();
 FILLER_ASAP7_75t_R FILLER_0_145_335 ();
 FILLER_ASAP7_75t_R FILLER_0_145_342 ();
 FILLER_ASAP7_75t_R FILLER_0_145_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_356 ();
 FILLER_ASAP7_75t_R FILLER_0_145_367 ();
 FILLER_ASAP7_75t_R FILLER_0_145_375 ();
 FILLER_ASAP7_75t_R FILLER_0_145_383 ();
 DECAPx4_ASAP7_75t_R FILLER_0_145_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_402 ();
 FILLER_ASAP7_75t_R FILLER_0_145_409 ();
 DECAPx1_ASAP7_75t_R FILLER_0_145_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_421 ();
 FILLER_ASAP7_75t_R FILLER_0_145_428 ();
 DECAPx4_ASAP7_75t_R FILLER_0_145_438 ();
 FILLER_ASAP7_75t_R FILLER_0_145_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_450 ();
 FILLER_ASAP7_75t_R FILLER_0_145_459 ();
 FILLER_ASAP7_75t_R FILLER_0_145_467 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_501 ();
 DECAPx2_ASAP7_75t_R FILLER_0_145_524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_552 ();
 DECAPx6_ASAP7_75t_R FILLER_0_145_595 ();
 DECAPx2_ASAP7_75t_R FILLER_0_145_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_615 ();
 FILLER_ASAP7_75t_R FILLER_0_145_628 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_641 ();
 DECAPx6_ASAP7_75t_R FILLER_0_145_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_687 ();
 FILLER_ASAP7_75t_R FILLER_0_145_693 ();
 FILLER_ASAP7_75t_R FILLER_0_145_705 ();
 FILLER_ASAP7_75t_R FILLER_0_145_717 ();
 DECAPx6_ASAP7_75t_R FILLER_0_145_724 ();
 DECAPx2_ASAP7_75t_R FILLER_0_145_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_744 ();
 DECAPx2_ASAP7_75t_R FILLER_0_145_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_761 ();
 DECAPx2_ASAP7_75t_R FILLER_0_145_772 ();
 FILLER_ASAP7_75t_R FILLER_0_145_788 ();
 DECAPx2_ASAP7_75t_R FILLER_0_145_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_806 ();
 FILLER_ASAP7_75t_R FILLER_0_145_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_816 ();
 FILLER_ASAP7_75t_R FILLER_0_145_827 ();
 FILLER_ASAP7_75t_R FILLER_0_145_837 ();
 FILLER_ASAP7_75t_R FILLER_0_145_844 ();
 FILLER_ASAP7_75t_R FILLER_0_145_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_853 ();
 FILLER_ASAP7_75t_R FILLER_0_145_860 ();
 FILLER_ASAP7_75t_R FILLER_0_145_868 ();
 DECAPx2_ASAP7_75t_R FILLER_0_145_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_882 ();
 DECAPx4_ASAP7_75t_R FILLER_0_145_890 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_900 ();
 DECAPx6_ASAP7_75t_R FILLER_0_145_907 ();
 DECAPx1_ASAP7_75t_R FILLER_0_145_921 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_927 ();
 DECAPx2_ASAP7_75t_R FILLER_0_145_949 ();
 FILLER_ASAP7_75t_R FILLER_0_145_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_978 ();
 DECAPx1_ASAP7_75t_R FILLER_0_145_1001 ();
 FILLER_ASAP7_75t_R FILLER_0_145_1013 ();
 FILLER_ASAP7_75t_R FILLER_0_145_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_1022 ();
 FILLER_ASAP7_75t_R FILLER_0_145_1035 ();
 DECAPx6_ASAP7_75t_R FILLER_0_145_1040 ();
 DECAPx1_ASAP7_75t_R FILLER_0_145_1054 ();
 DECAPx2_ASAP7_75t_R FILLER_0_145_1068 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_0_145_1079 ();
 FILLER_ASAP7_75t_R FILLER_0_145_1085 ();
 FILLER_ASAP7_75t_R FILLER_0_145_1095 ();
 DECAPx1_ASAP7_75t_R FILLER_0_145_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_1112 ();
 DECAPx4_ASAP7_75t_R FILLER_0_145_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_1128 ();
 FILLER_ASAP7_75t_R FILLER_0_145_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_1152 ();
 FILLER_ASAP7_75t_R FILLER_0_145_1158 ();
 DECAPx1_ASAP7_75t_R FILLER_0_145_1170 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_1174 ();
 FILLER_ASAP7_75t_R FILLER_0_145_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_1189 ();
 DECAPx1_ASAP7_75t_R FILLER_0_145_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_1212 ();
 FILLER_ASAP7_75t_R FILLER_0_145_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_1224 ();
 DECAPx6_ASAP7_75t_R FILLER_0_145_1246 ();
 FILLER_ASAP7_75t_R FILLER_0_145_1260 ();
 FILLER_ASAP7_75t_R FILLER_0_145_1269 ();
 DECAPx6_ASAP7_75t_R FILLER_0_145_1277 ();
 DECAPx1_ASAP7_75t_R FILLER_0_145_1291 ();
 DECAPx6_ASAP7_75t_R FILLER_0_145_1301 ();
 FILLER_ASAP7_75t_R FILLER_0_145_1315 ();
 FILLER_ASAP7_75t_R FILLER_0_145_1327 ();
 DECAPx2_ASAP7_75t_R FILLER_0_145_1334 ();
 FILLER_ASAP7_75t_R FILLER_0_145_1346 ();
 FILLER_ASAP7_75t_R FILLER_0_145_1351 ();
 FILLER_ASAP7_75t_R FILLER_0_145_1359 ();
 FILLER_ASAP7_75t_R FILLER_0_145_1367 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_1369 ();
 DECAPx2_ASAP7_75t_R FILLER_0_145_1376 ();
 FILLER_ASAP7_75t_R FILLER_0_146_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_146_9 ();
 FILLER_ASAP7_75t_R FILLER_0_146_15 ();
 FILLER_ASAP7_75t_R FILLER_0_146_22 ();
 DECAPx1_ASAP7_75t_R FILLER_0_146_30 ();
 DECAPx4_ASAP7_75t_R FILLER_0_146_40 ();
 FILLER_ASAP7_75t_R FILLER_0_146_56 ();
 FILLER_ASAP7_75t_R FILLER_0_146_64 ();
 DECAPx2_ASAP7_75t_R FILLER_0_146_78 ();
 FILLER_ASAP7_75t_R FILLER_0_146_95 ();
 DECAPx1_ASAP7_75t_R FILLER_0_146_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_111 ();
 FILLER_ASAP7_75t_R FILLER_0_146_122 ();
 DECAPx2_ASAP7_75t_R FILLER_0_146_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_136 ();
 FILLER_ASAP7_75t_R FILLER_0_146_149 ();
 FILLER_ASAP7_75t_R FILLER_0_146_163 ();
 DECAPx2_ASAP7_75t_R FILLER_0_146_173 ();
 DECAPx2_ASAP7_75t_R FILLER_0_146_191 ();
 DECAPx4_ASAP7_75t_R FILLER_0_146_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_213 ();
 DECAPx4_ASAP7_75t_R FILLER_0_146_221 ();
 FILLER_ASAP7_75t_R FILLER_0_146_231 ();
 FILLER_ASAP7_75t_R FILLER_0_146_241 ();
 DECAPx6_ASAP7_75t_R FILLER_0_146_251 ();
 DECAPx1_ASAP7_75t_R FILLER_0_146_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_269 ();
 FILLER_ASAP7_75t_R FILLER_0_146_276 ();
 DECAPx1_ASAP7_75t_R FILLER_0_146_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_289 ();
 FILLER_ASAP7_75t_R FILLER_0_146_296 ();
 DECAPx2_ASAP7_75t_R FILLER_0_146_305 ();
 FILLER_ASAP7_75t_R FILLER_0_146_311 ();
 DECAPx4_ASAP7_75t_R FILLER_0_146_319 ();
 FILLER_ASAP7_75t_R FILLER_0_146_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_341 ();
 FILLER_ASAP7_75t_R FILLER_0_146_347 ();
 DECAPx2_ASAP7_75t_R FILLER_0_146_355 ();
 FILLER_ASAP7_75t_R FILLER_0_146_371 ();
 DECAPx1_ASAP7_75t_R FILLER_0_146_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_385 ();
 DECAPx6_ASAP7_75t_R FILLER_0_146_392 ();
 FILLER_ASAP7_75t_R FILLER_0_146_412 ();
 DECAPx2_ASAP7_75t_R FILLER_0_146_422 ();
 DECAPx1_ASAP7_75t_R FILLER_0_146_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_438 ();
 DECAPx1_ASAP7_75t_R FILLER_0_146_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_449 ();
 DECAPx1_ASAP7_75t_R FILLER_0_146_458 ();
 DECAPx2_ASAP7_75t_R FILLER_0_146_464 ();
 DECAPx6_ASAP7_75t_R FILLER_0_146_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_490 ();
 FILLER_ASAP7_75t_R FILLER_0_146_512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_522 ();
 DECAPx2_ASAP7_75t_R FILLER_0_146_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_550 ();
 DECAPx1_ASAP7_75t_R FILLER_0_146_572 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_579 ();
 DECAPx6_ASAP7_75t_R FILLER_0_146_601 ();
 FILLER_ASAP7_75t_R FILLER_0_146_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_617 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_624 ();
 DECAPx1_ASAP7_75t_R FILLER_0_146_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_650 ();
 DECAPx6_ASAP7_75t_R FILLER_0_146_657 ();
 DECAPx1_ASAP7_75t_R FILLER_0_146_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_685 ();
 FILLER_ASAP7_75t_R FILLER_0_146_696 ();
 FILLER_ASAP7_75t_R FILLER_0_146_708 ();
 FILLER_ASAP7_75t_R FILLER_0_146_715 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_723 ();
 DECAPx4_ASAP7_75t_R FILLER_0_146_745 ();
 FILLER_ASAP7_75t_R FILLER_0_146_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_757 ();
 FILLER_ASAP7_75t_R FILLER_0_146_766 ();
 DECAPx1_ASAP7_75t_R FILLER_0_146_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_777 ();
 DECAPx2_ASAP7_75t_R FILLER_0_146_788 ();
 FILLER_ASAP7_75t_R FILLER_0_146_806 ();
 FILLER_ASAP7_75t_R FILLER_0_146_814 ();
 FILLER_ASAP7_75t_R FILLER_0_146_824 ();
 FILLER_ASAP7_75t_R FILLER_0_146_832 ();
 FILLER_ASAP7_75t_R FILLER_0_146_840 ();
 FILLER_ASAP7_75t_R FILLER_0_146_848 ();
 FILLER_ASAP7_75t_R FILLER_0_146_856 ();
 FILLER_ASAP7_75t_R FILLER_0_146_864 ();
 FILLER_ASAP7_75t_R FILLER_0_146_876 ();
 DECAPx4_ASAP7_75t_R FILLER_0_146_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_894 ();
 DECAPx6_ASAP7_75t_R FILLER_0_146_901 ();
 DECAPx1_ASAP7_75t_R FILLER_0_146_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_919 ();
 DECAPx1_ASAP7_75t_R FILLER_0_146_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_936 ();
 FILLER_ASAP7_75t_R FILLER_0_146_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_951 ();
 FILLER_ASAP7_75t_R FILLER_0_146_958 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_960 ();
 DECAPx2_ASAP7_75t_R FILLER_0_146_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_973 ();
 DECAPx1_ASAP7_75t_R FILLER_0_146_977 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_981 ();
 FILLER_ASAP7_75t_R FILLER_0_146_1003 ();
 FILLER_ASAP7_75t_R FILLER_0_146_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_1010 ();
 DECAPx2_ASAP7_75t_R FILLER_0_146_1019 ();
 DECAPx1_ASAP7_75t_R FILLER_0_146_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_1035 ();
 DECAPx2_ASAP7_75t_R FILLER_0_146_1056 ();
 DECAPx1_ASAP7_75t_R FILLER_0_146_1070 ();
 FILLER_ASAP7_75t_R FILLER_0_146_1080 ();
 DECAPx1_ASAP7_75t_R FILLER_0_146_1088 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_1092 ();
 FILLER_ASAP7_75t_R FILLER_0_146_1096 ();
 FILLER_ASAP7_75t_R FILLER_0_146_1106 ();
 FILLER_ASAP7_75t_R FILLER_0_146_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_1113 ();
 FILLER_ASAP7_75t_R FILLER_0_146_1117 ();
 FILLER_ASAP7_75t_R FILLER_0_146_1122 ();
 FILLER_ASAP7_75t_R FILLER_0_146_1132 ();
 DECAPx1_ASAP7_75t_R FILLER_0_146_1137 ();
 FILLER_ASAP7_75t_R FILLER_0_146_1146 ();
 DECAPx1_ASAP7_75t_R FILLER_0_146_1154 ();
 FILLER_ASAP7_75t_R FILLER_0_146_1168 ();
 FILLER_ASAP7_75t_R FILLER_0_146_1180 ();
 FILLER_ASAP7_75t_R FILLER_0_146_1187 ();
 FILLER_ASAP7_75t_R FILLER_0_146_1197 ();
 DECAPx2_ASAP7_75t_R FILLER_0_146_1206 ();
 DECAPx1_ASAP7_75t_R FILLER_0_146_1226 ();
 FILLER_ASAP7_75t_R FILLER_0_146_1236 ();
 FILLER_ASAP7_75t_R FILLER_0_146_1244 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_1246 ();
 DECAPx1_ASAP7_75t_R FILLER_0_146_1253 ();
 DECAPx2_ASAP7_75t_R FILLER_0_146_1267 ();
 FILLER_ASAP7_75t_R FILLER_0_146_1279 ();
 DECAPx6_ASAP7_75t_R FILLER_0_146_1286 ();
 DECAPx1_ASAP7_75t_R FILLER_0_146_1300 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_1304 ();
 FILLER_ASAP7_75t_R FILLER_0_146_1310 ();
 FILLER_ASAP7_75t_R FILLER_0_146_1340 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_1342 ();
 FILLER_ASAP7_75t_R FILLER_0_146_1349 ();
 FILLER_ASAP7_75t_R FILLER_0_146_1372 ();
 FILLER_ASAP7_75t_R FILLER_0_146_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_147_2 ();
 FILLER_ASAP7_75t_R FILLER_0_147_9 ();
 FILLER_ASAP7_75t_R FILLER_0_147_16 ();
 FILLER_ASAP7_75t_R FILLER_0_147_21 ();
 DECAPx4_ASAP7_75t_R FILLER_0_147_44 ();
 DECAPx2_ASAP7_75t_R FILLER_0_147_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_72 ();
 DECAPx1_ASAP7_75t_R FILLER_0_147_85 ();
 DECAPx2_ASAP7_75t_R FILLER_0_147_100 ();
 FILLER_ASAP7_75t_R FILLER_0_147_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_108 ();
 DECAPx1_ASAP7_75t_R FILLER_0_147_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_119 ();
 DECAPx2_ASAP7_75t_R FILLER_0_147_128 ();
 DECAPx2_ASAP7_75t_R FILLER_0_147_146 ();
 FILLER_ASAP7_75t_R FILLER_0_147_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_154 ();
 FILLER_ASAP7_75t_R FILLER_0_147_161 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_166 ();
 DECAPx2_ASAP7_75t_R FILLER_0_147_188 ();
 FILLER_ASAP7_75t_R FILLER_0_147_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_196 ();
 DECAPx2_ASAP7_75t_R FILLER_0_147_205 ();
 DECAPx2_ASAP7_75t_R FILLER_0_147_222 ();
 FILLER_ASAP7_75t_R FILLER_0_147_228 ();
 FILLER_ASAP7_75t_R FILLER_0_147_240 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_250 ();
 FILLER_ASAP7_75t_R FILLER_0_147_275 ();
 FILLER_ASAP7_75t_R FILLER_0_147_283 ();
 DECAPx1_ASAP7_75t_R FILLER_0_147_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_292 ();
 DECAPx1_ASAP7_75t_R FILLER_0_147_303 ();
 FILLER_ASAP7_75t_R FILLER_0_147_313 ();
 DECAPx4_ASAP7_75t_R FILLER_0_147_321 ();
 DECAPx1_ASAP7_75t_R FILLER_0_147_334 ();
 FILLER_ASAP7_75t_R FILLER_0_147_346 ();
 DECAPx2_ASAP7_75t_R FILLER_0_147_358 ();
 FILLER_ASAP7_75t_R FILLER_0_147_364 ();
 FILLER_ASAP7_75t_R FILLER_0_147_376 ();
 FILLER_ASAP7_75t_R FILLER_0_147_384 ();
 FILLER_ASAP7_75t_R FILLER_0_147_391 ();
 DECAPx1_ASAP7_75t_R FILLER_0_147_396 ();
 FILLER_ASAP7_75t_R FILLER_0_147_406 ();
 DECAPx4_ASAP7_75t_R FILLER_0_147_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_426 ();
 DECAPx4_ASAP7_75t_R FILLER_0_147_434 ();
 FILLER_ASAP7_75t_R FILLER_0_147_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_446 ();
 FILLER_ASAP7_75t_R FILLER_0_147_453 ();
 DECAPx2_ASAP7_75t_R FILLER_0_147_462 ();
 DECAPx6_ASAP7_75t_R FILLER_0_147_471 ();
 DECAPx2_ASAP7_75t_R FILLER_0_147_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_491 ();
 FILLER_ASAP7_75t_R FILLER_0_147_495 ();
 DECAPx2_ASAP7_75t_R FILLER_0_147_505 ();
 FILLER_ASAP7_75t_R FILLER_0_147_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_513 ();
 FILLER_ASAP7_75t_R FILLER_0_147_522 ();
 FILLER_ASAP7_75t_R FILLER_0_147_532 ();
 DECAPx1_ASAP7_75t_R FILLER_0_147_540 ();
 FILLER_ASAP7_75t_R FILLER_0_147_565 ();
 DECAPx1_ASAP7_75t_R FILLER_0_147_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_583 ();
 DECAPx6_ASAP7_75t_R FILLER_0_147_595 ();
 FILLER_ASAP7_75t_R FILLER_0_147_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_623 ();
 DECAPx4_ASAP7_75t_R FILLER_0_147_631 ();
 FILLER_ASAP7_75t_R FILLER_0_147_641 ();
 FILLER_ASAP7_75t_R FILLER_0_147_664 ();
 FILLER_ASAP7_75t_R FILLER_0_147_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_678 ();
 FILLER_ASAP7_75t_R FILLER_0_147_684 ();
 DECAPx2_ASAP7_75t_R FILLER_0_147_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_702 ();
 FILLER_ASAP7_75t_R FILLER_0_147_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_710 ();
 DECAPx4_ASAP7_75t_R FILLER_0_147_723 ();
 FILLER_ASAP7_75t_R FILLER_0_147_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_735 ();
 DECAPx1_ASAP7_75t_R FILLER_0_147_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_745 ();
 FILLER_ASAP7_75t_R FILLER_0_147_753 ();
 FILLER_ASAP7_75t_R FILLER_0_147_758 ();
 DECAPx1_ASAP7_75t_R FILLER_0_147_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_770 ();
 FILLER_ASAP7_75t_R FILLER_0_147_781 ();
 FILLER_ASAP7_75t_R FILLER_0_147_793 ();
 FILLER_ASAP7_75t_R FILLER_0_147_813 ();
 FILLER_ASAP7_75t_R FILLER_0_147_821 ();
 DECAPx1_ASAP7_75t_R FILLER_0_147_829 ();
 DECAPx1_ASAP7_75t_R FILLER_0_147_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_843 ();
 FILLER_ASAP7_75t_R FILLER_0_147_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_856 ();
 FILLER_ASAP7_75t_R FILLER_0_147_863 ();
 FILLER_ASAP7_75t_R FILLER_0_147_871 ();
 DECAPx2_ASAP7_75t_R FILLER_0_147_878 ();
 DECAPx2_ASAP7_75t_R FILLER_0_147_890 ();
 FILLER_ASAP7_75t_R FILLER_0_147_902 ();
 DECAPx6_ASAP7_75t_R FILLER_0_147_911 ();
 FILLER_ASAP7_75t_R FILLER_0_147_927 ();
 FILLER_ASAP7_75t_R FILLER_0_147_941 ();
 DECAPx1_ASAP7_75t_R FILLER_0_147_955 ();
 DECAPx4_ASAP7_75t_R FILLER_0_147_966 ();
 FILLER_ASAP7_75t_R FILLER_0_147_988 ();
 DECAPx6_ASAP7_75t_R FILLER_0_147_996 ();
 DECAPx1_ASAP7_75t_R FILLER_0_147_1010 ();
 FILLER_ASAP7_75t_R FILLER_0_147_1020 ();
 FILLER_ASAP7_75t_R FILLER_0_147_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_1032 ();
 FILLER_ASAP7_75t_R FILLER_0_147_1053 ();
 FILLER_ASAP7_75t_R FILLER_0_147_1063 ();
 DECAPx2_ASAP7_75t_R FILLER_0_147_1073 ();
 FILLER_ASAP7_75t_R FILLER_0_147_1079 ();
 DECAPx2_ASAP7_75t_R FILLER_0_147_1089 ();
 DECAPx4_ASAP7_75t_R FILLER_0_147_1106 ();
 FILLER_ASAP7_75t_R FILLER_0_147_1127 ();
 DECAPx1_ASAP7_75t_R FILLER_0_147_1135 ();
 DECAPx2_ASAP7_75t_R FILLER_0_147_1142 ();
 FILLER_ASAP7_75t_R FILLER_0_147_1148 ();
 FILLER_ASAP7_75t_R FILLER_0_147_1155 ();
 FILLER_ASAP7_75t_R FILLER_0_147_1167 ();
 FILLER_ASAP7_75t_R FILLER_0_147_1179 ();
 FILLER_ASAP7_75t_R FILLER_0_147_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_147_1195 ();
 FILLER_ASAP7_75t_R FILLER_0_147_1203 ();
 FILLER_ASAP7_75t_R FILLER_0_147_1211 ();
 DECAPx6_ASAP7_75t_R FILLER_0_147_1218 ();
 DECAPx1_ASAP7_75t_R FILLER_0_147_1232 ();
 FILLER_ASAP7_75t_R FILLER_0_147_1242 ();
 FILLER_ASAP7_75t_R FILLER_0_147_1249 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_1251 ();
 DECAPx2_ASAP7_75t_R FILLER_0_147_1258 ();
 FILLER_ASAP7_75t_R FILLER_0_147_1264 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_1266 ();
 FILLER_ASAP7_75t_R FILLER_0_147_1274 ();
 DECAPx2_ASAP7_75t_R FILLER_0_147_1282 ();
 DECAPx2_ASAP7_75t_R FILLER_0_147_1300 ();
 FILLER_ASAP7_75t_R FILLER_0_147_1306 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_1308 ();
 FILLER_ASAP7_75t_R FILLER_0_147_1315 ();
 FILLER_ASAP7_75t_R FILLER_0_147_1322 ();
 FILLER_ASAP7_75t_R FILLER_0_147_1362 ();
 DECAPx2_ASAP7_75t_R FILLER_0_147_1369 ();
 FILLER_ASAP7_75t_R FILLER_0_147_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_148_2 ();
 FILLER_ASAP7_75t_R FILLER_0_148_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_28 ();
 FILLER_ASAP7_75t_R FILLER_0_148_34 ();
 DECAPx6_ASAP7_75t_R FILLER_0_148_39 ();
 DECAPx4_ASAP7_75t_R FILLER_0_148_59 ();
 DECAPx6_ASAP7_75t_R FILLER_0_148_77 ();
 FILLER_ASAP7_75t_R FILLER_0_148_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_93 ();
 DECAPx2_ASAP7_75t_R FILLER_0_148_102 ();
 FILLER_ASAP7_75t_R FILLER_0_148_114 ();
 DECAPx2_ASAP7_75t_R FILLER_0_148_122 ();
 FILLER_ASAP7_75t_R FILLER_0_148_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_130 ();
 DECAPx4_ASAP7_75t_R FILLER_0_148_143 ();
 FILLER_ASAP7_75t_R FILLER_0_148_153 ();
 DECAPx2_ASAP7_75t_R FILLER_0_148_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_169 ();
 DECAPx6_ASAP7_75t_R FILLER_0_148_181 ();
 DECAPx2_ASAP7_75t_R FILLER_0_148_195 ();
 DECAPx6_ASAP7_75t_R FILLER_0_148_207 ();
 DECAPx2_ASAP7_75t_R FILLER_0_148_221 ();
 FILLER_ASAP7_75t_R FILLER_0_148_232 ();
 FILLER_ASAP7_75t_R FILLER_0_148_244 ();
 DECAPx6_ASAP7_75t_R FILLER_0_148_254 ();
 FILLER_ASAP7_75t_R FILLER_0_148_274 ();
 FILLER_ASAP7_75t_R FILLER_0_148_282 ();
 FILLER_ASAP7_75t_R FILLER_0_148_290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_298 ();
 DECAPx6_ASAP7_75t_R FILLER_0_148_320 ();
 DECAPx1_ASAP7_75t_R FILLER_0_148_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_338 ();
 DECAPx1_ASAP7_75t_R FILLER_0_148_344 ();
 FILLER_ASAP7_75t_R FILLER_0_148_354 ();
 FILLER_ASAP7_75t_R FILLER_0_148_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_365 ();
 FILLER_ASAP7_75t_R FILLER_0_148_371 ();
 DECAPx1_ASAP7_75t_R FILLER_0_148_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_383 ();
 DECAPx4_ASAP7_75t_R FILLER_0_148_387 ();
 FILLER_ASAP7_75t_R FILLER_0_148_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_405 ();
 DECAPx4_ASAP7_75t_R FILLER_0_148_412 ();
 FILLER_ASAP7_75t_R FILLER_0_148_422 ();
 DECAPx4_ASAP7_75t_R FILLER_0_148_432 ();
 FILLER_ASAP7_75t_R FILLER_0_148_442 ();
 FILLER_ASAP7_75t_R FILLER_0_148_450 ();
 FILLER_ASAP7_75t_R FILLER_0_148_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_461 ();
 FILLER_ASAP7_75t_R FILLER_0_148_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_466 ();
 DECAPx6_ASAP7_75t_R FILLER_0_148_473 ();
 DECAPx2_ASAP7_75t_R FILLER_0_148_487 ();
 DECAPx2_ASAP7_75t_R FILLER_0_148_503 ();
 FILLER_ASAP7_75t_R FILLER_0_148_509 ();
 DECAPx1_ASAP7_75t_R FILLER_0_148_517 ();
 FILLER_ASAP7_75t_R FILLER_0_148_533 ();
 FILLER_ASAP7_75t_R FILLER_0_148_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_545 ();
 FILLER_ASAP7_75t_R FILLER_0_148_557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_148_562 ();
 FILLER_ASAP7_75t_R FILLER_0_148_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_570 ();
 FILLER_ASAP7_75t_R FILLER_0_148_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_585 ();
 FILLER_ASAP7_75t_R FILLER_0_148_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_148_607 ();
 FILLER_ASAP7_75t_R FILLER_0_148_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_615 ();
 FILLER_ASAP7_75t_R FILLER_0_148_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_639 ();
 FILLER_ASAP7_75t_R FILLER_0_148_643 ();
 DECAPx4_ASAP7_75t_R FILLER_0_148_653 ();
 FILLER_ASAP7_75t_R FILLER_0_148_663 ();
 DECAPx4_ASAP7_75t_R FILLER_0_148_675 ();
 FILLER_ASAP7_75t_R FILLER_0_148_685 ();
 DECAPx1_ASAP7_75t_R FILLER_0_148_697 ();
 DECAPx1_ASAP7_75t_R FILLER_0_148_711 ();
 FILLER_ASAP7_75t_R FILLER_0_148_721 ();
 DECAPx2_ASAP7_75t_R FILLER_0_148_729 ();
 FILLER_ASAP7_75t_R FILLER_0_148_735 ();
 DECAPx1_ASAP7_75t_R FILLER_0_148_749 ();
 DECAPx6_ASAP7_75t_R FILLER_0_148_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_773 ();
 FILLER_ASAP7_75t_R FILLER_0_148_781 ();
 FILLER_ASAP7_75t_R FILLER_0_148_793 ();
 DECAPx1_ASAP7_75t_R FILLER_0_148_805 ();
 FILLER_ASAP7_75t_R FILLER_0_148_815 ();
 DECAPx6_ASAP7_75t_R FILLER_0_148_822 ();
 FILLER_ASAP7_75t_R FILLER_0_148_836 ();
 DECAPx6_ASAP7_75t_R FILLER_0_148_844 ();
 DECAPx1_ASAP7_75t_R FILLER_0_148_858 ();
 FILLER_ASAP7_75t_R FILLER_0_148_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_870 ();
 FILLER_ASAP7_75t_R FILLER_0_148_879 ();
 FILLER_ASAP7_75t_R FILLER_0_148_887 ();
 FILLER_ASAP7_75t_R FILLER_0_148_895 ();
 FILLER_ASAP7_75t_R FILLER_0_148_907 ();
 DECAPx6_ASAP7_75t_R FILLER_0_148_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_926 ();
 DECAPx1_ASAP7_75t_R FILLER_0_148_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_943 ();
 DECAPx1_ASAP7_75t_R FILLER_0_148_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_959 ();
 FILLER_ASAP7_75t_R FILLER_0_148_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_973 ();
 FILLER_ASAP7_75t_R FILLER_0_148_982 ();
 DECAPx4_ASAP7_75t_R FILLER_0_148_987 ();
 FILLER_ASAP7_75t_R FILLER_0_148_997 ();
 DECAPx4_ASAP7_75t_R FILLER_0_148_1004 ();
 FILLER_ASAP7_75t_R FILLER_0_148_1014 ();
 FILLER_ASAP7_75t_R FILLER_0_148_1019 ();
 DECAPx2_ASAP7_75t_R FILLER_0_148_1027 ();
 FILLER_ASAP7_75t_R FILLER_0_148_1033 ();
 FILLER_ASAP7_75t_R FILLER_0_148_1045 ();
 FILLER_ASAP7_75t_R FILLER_0_148_1053 ();
 FILLER_ASAP7_75t_R FILLER_0_148_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_1065 ();
 DECAPx4_ASAP7_75t_R FILLER_0_148_1072 ();
 FILLER_ASAP7_75t_R FILLER_0_148_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_0_148_1096 ();
 DECAPx4_ASAP7_75t_R FILLER_0_148_1110 ();
 DECAPx1_ASAP7_75t_R FILLER_0_148_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_1127 ();
 DECAPx2_ASAP7_75t_R FILLER_0_148_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_1146 ();
 FILLER_ASAP7_75t_R FILLER_0_148_1168 ();
 FILLER_ASAP7_75t_R FILLER_0_148_1178 ();
 FILLER_ASAP7_75t_R FILLER_0_148_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_148_1194 ();
 DECAPx6_ASAP7_75t_R FILLER_0_148_1202 ();
 FILLER_ASAP7_75t_R FILLER_0_148_1216 ();
 FILLER_ASAP7_75t_R FILLER_0_148_1226 ();
 DECAPx1_ASAP7_75t_R FILLER_0_148_1234 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_1238 ();
 DECAPx2_ASAP7_75t_R FILLER_0_148_1245 ();
 FILLER_ASAP7_75t_R FILLER_0_148_1257 ();
 DECAPx2_ASAP7_75t_R FILLER_0_148_1265 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_1271 ();
 DECAPx1_ASAP7_75t_R FILLER_0_148_1279 ();
 FILLER_ASAP7_75t_R FILLER_0_148_1289 ();
 DECAPx4_ASAP7_75t_R FILLER_0_148_1298 ();
 FILLER_ASAP7_75t_R FILLER_0_148_1308 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_1310 ();
 DECAPx1_ASAP7_75t_R FILLER_0_148_1321 ();
 FILLER_ASAP7_75t_R FILLER_0_148_1333 ();
 FILLER_ASAP7_75t_R FILLER_0_148_1338 ();
 FILLER_ASAP7_75t_R FILLER_0_148_1351 ();
 FILLER_ASAP7_75t_R FILLER_0_148_1363 ();
 FILLER_ASAP7_75t_R FILLER_0_148_1371 ();
 FILLER_ASAP7_75t_R FILLER_0_148_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_149_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_4 ();
 DECAPx1_ASAP7_75t_R FILLER_0_149_11 ();
 FILLER_ASAP7_75t_R FILLER_0_149_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_149_49 ();
 DECAPx2_ASAP7_75t_R FILLER_0_149_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_69 ();
 FILLER_ASAP7_75t_R FILLER_0_149_74 ();
 DECAPx1_ASAP7_75t_R FILLER_0_149_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_86 ();
 FILLER_ASAP7_75t_R FILLER_0_149_93 ();
 DECAPx4_ASAP7_75t_R FILLER_0_149_103 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_149_138 ();
 FILLER_ASAP7_75t_R FILLER_0_149_163 ();
 FILLER_ASAP7_75t_R FILLER_0_149_171 ();
 DECAPx6_ASAP7_75t_R FILLER_0_149_176 ();
 DECAPx2_ASAP7_75t_R FILLER_0_149_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_196 ();
 DECAPx6_ASAP7_75t_R FILLER_0_149_209 ();
 FILLER_ASAP7_75t_R FILLER_0_149_223 ();
 DECAPx4_ASAP7_75t_R FILLER_0_149_231 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_271 ();
 DECAPx2_ASAP7_75t_R FILLER_0_149_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_285 ();
 FILLER_ASAP7_75t_R FILLER_0_149_293 ();
 DECAPx1_ASAP7_75t_R FILLER_0_149_301 ();
 FILLER_ASAP7_75t_R FILLER_0_149_311 ();
 DECAPx6_ASAP7_75t_R FILLER_0_149_319 ();
 DECAPx1_ASAP7_75t_R FILLER_0_149_343 ();
 DECAPx1_ASAP7_75t_R FILLER_0_149_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_361 ();
 DECAPx1_ASAP7_75t_R FILLER_0_149_368 ();
 DECAPx2_ASAP7_75t_R FILLER_0_149_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_384 ();
 FILLER_ASAP7_75t_R FILLER_0_149_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_395 ();
 DECAPx1_ASAP7_75t_R FILLER_0_149_399 ();
 DECAPx2_ASAP7_75t_R FILLER_0_149_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_415 ();
 FILLER_ASAP7_75t_R FILLER_0_149_422 ();
 DECAPx1_ASAP7_75t_R FILLER_0_149_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_434 ();
 DECAPx4_ASAP7_75t_R FILLER_0_149_441 ();
 FILLER_ASAP7_75t_R FILLER_0_149_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_453 ();
 FILLER_ASAP7_75t_R FILLER_0_149_457 ();
 FILLER_ASAP7_75t_R FILLER_0_149_465 ();
 DECAPx6_ASAP7_75t_R FILLER_0_149_473 ();
 FILLER_ASAP7_75t_R FILLER_0_149_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_489 ();
 DECAPx2_ASAP7_75t_R FILLER_0_149_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_517 ();
 DECAPx4_ASAP7_75t_R FILLER_0_149_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_535 ();
 DECAPx1_ASAP7_75t_R FILLER_0_149_542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_549 ();
 FILLER_ASAP7_75t_R FILLER_0_149_571 ();
 FILLER_ASAP7_75t_R FILLER_0_149_585 ();
 FILLER_ASAP7_75t_R FILLER_0_149_599 ();
 FILLER_ASAP7_75t_R FILLER_0_149_607 ();
 FILLER_ASAP7_75t_R FILLER_0_149_612 ();
 DECAPx4_ASAP7_75t_R FILLER_0_149_626 ();
 FILLER_ASAP7_75t_R FILLER_0_149_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_638 ();
 DECAPx6_ASAP7_75t_R FILLER_0_149_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_665 ();
 DECAPx2_ASAP7_75t_R FILLER_0_149_676 ();
 FILLER_ASAP7_75t_R FILLER_0_149_687 ();
 FILLER_ASAP7_75t_R FILLER_0_149_699 ();
 DECAPx1_ASAP7_75t_R FILLER_0_149_706 ();
 FILLER_ASAP7_75t_R FILLER_0_149_716 ();
 DECAPx4_ASAP7_75t_R FILLER_0_149_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_734 ();
 DECAPx2_ASAP7_75t_R FILLER_0_149_747 ();
 FILLER_ASAP7_75t_R FILLER_0_149_760 ();
 DECAPx1_ASAP7_75t_R FILLER_0_149_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_772 ();
 FILLER_ASAP7_75t_R FILLER_0_149_781 ();
 DECAPx1_ASAP7_75t_R FILLER_0_149_793 ();
 FILLER_ASAP7_75t_R FILLER_0_149_807 ();
 FILLER_ASAP7_75t_R FILLER_0_149_817 ();
 DECAPx6_ASAP7_75t_R FILLER_0_149_824 ();
 DECAPx6_ASAP7_75t_R FILLER_0_149_846 ();
 DECAPx2_ASAP7_75t_R FILLER_0_149_860 ();
 DECAPx4_ASAP7_75t_R FILLER_0_149_872 ();
 FILLER_ASAP7_75t_R FILLER_0_149_882 ();
 FILLER_ASAP7_75t_R FILLER_0_149_890 ();
 FILLER_ASAP7_75t_R FILLER_0_149_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_900 ();
 FILLER_ASAP7_75t_R FILLER_0_149_907 ();
 DECAPx4_ASAP7_75t_R FILLER_0_149_915 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_927 ();
 FILLER_ASAP7_75t_R FILLER_0_149_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_951 ();
 DECAPx1_ASAP7_75t_R FILLER_0_149_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_966 ();
 DECAPx6_ASAP7_75t_R FILLER_0_149_974 ();
 FILLER_ASAP7_75t_R FILLER_0_149_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_990 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_999 ();
 DECAPx4_ASAP7_75t_R FILLER_0_149_1021 ();
 FILLER_ASAP7_75t_R FILLER_0_149_1031 ();
 FILLER_ASAP7_75t_R FILLER_0_149_1039 ();
 FILLER_ASAP7_75t_R FILLER_0_149_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_1064 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_1086 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_1108 ();
 DECAPx6_ASAP7_75t_R FILLER_0_149_1130 ();
 DECAPx1_ASAP7_75t_R FILLER_0_149_1144 ();
 FILLER_ASAP7_75t_R FILLER_0_149_1151 ();
 FILLER_ASAP7_75t_R FILLER_0_149_1179 ();
 FILLER_ASAP7_75t_R FILLER_0_149_1187 ();
 DECAPx6_ASAP7_75t_R FILLER_0_149_1194 ();
 FILLER_ASAP7_75t_R FILLER_0_149_1220 ();
 FILLER_ASAP7_75t_R FILLER_0_149_1232 ();
 FILLER_ASAP7_75t_R FILLER_0_149_1244 ();
 FILLER_ASAP7_75t_R FILLER_0_149_1252 ();
 FILLER_ASAP7_75t_R FILLER_0_149_1260 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_1262 ();
 DECAPx1_ASAP7_75t_R FILLER_0_149_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_1273 ();
 FILLER_ASAP7_75t_R FILLER_0_149_1280 ();
 FILLER_ASAP7_75t_R FILLER_0_149_1294 ();
 DECAPx1_ASAP7_75t_R FILLER_0_149_1304 ();
 DECAPx1_ASAP7_75t_R FILLER_0_149_1318 ();
 DECAPx2_ASAP7_75t_R FILLER_0_149_1328 ();
 DECAPx1_ASAP7_75t_R FILLER_0_149_1345 ();
 DECAPx1_ASAP7_75t_R FILLER_0_149_1370 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_1374 ();
 FILLER_ASAP7_75t_R FILLER_0_149_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_150_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_150_25 ();
 DECAPx6_ASAP7_75t_R FILLER_0_150_34 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_48 ();
 FILLER_ASAP7_75t_R FILLER_0_150_65 ();
 FILLER_ASAP7_75t_R FILLER_0_150_73 ();
 FILLER_ASAP7_75t_R FILLER_0_150_83 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_91 ();
 FILLER_ASAP7_75t_R FILLER_0_150_97 ();
 FILLER_ASAP7_75t_R FILLER_0_150_110 ();
 DECAPx6_ASAP7_75t_R FILLER_0_150_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_134 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_149 ();
 FILLER_ASAP7_75t_R FILLER_0_150_154 ();
 DECAPx4_ASAP7_75t_R FILLER_0_150_162 ();
 FILLER_ASAP7_75t_R FILLER_0_150_172 ();
 FILLER_ASAP7_75t_R FILLER_0_150_182 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_198 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_210 ();
 FILLER_ASAP7_75t_R FILLER_0_150_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_218 ();
 FILLER_ASAP7_75t_R FILLER_0_150_225 ();
 FILLER_ASAP7_75t_R FILLER_0_150_235 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_245 ();
 DECAPx1_ASAP7_75t_R FILLER_0_150_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_271 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_278 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_290 ();
 FILLER_ASAP7_75t_R FILLER_0_150_296 ();
 FILLER_ASAP7_75t_R FILLER_0_150_304 ();
 FILLER_ASAP7_75t_R FILLER_0_150_312 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_320 ();
 FILLER_ASAP7_75t_R FILLER_0_150_336 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_348 ();
 FILLER_ASAP7_75t_R FILLER_0_150_354 ();
 FILLER_ASAP7_75t_R FILLER_0_150_364 ();
 FILLER_ASAP7_75t_R FILLER_0_150_369 ();
 FILLER_ASAP7_75t_R FILLER_0_150_377 ();
 DECAPx6_ASAP7_75t_R FILLER_0_150_384 ();
 FILLER_ASAP7_75t_R FILLER_0_150_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_408 ();
 FILLER_ASAP7_75t_R FILLER_0_150_417 ();
 FILLER_ASAP7_75t_R FILLER_0_150_425 ();
 FILLER_ASAP7_75t_R FILLER_0_150_433 ();
 DECAPx6_ASAP7_75t_R FILLER_0_150_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_486 ();
 FILLER_ASAP7_75t_R FILLER_0_150_499 ();
 DECAPx1_ASAP7_75t_R FILLER_0_150_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_508 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_523 ();
 FILLER_ASAP7_75t_R FILLER_0_150_529 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_541 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_569 ();
 DECAPx6_ASAP7_75t_R FILLER_0_150_582 ();
 DECAPx1_ASAP7_75t_R FILLER_0_150_596 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_608 ();
 FILLER_ASAP7_75t_R FILLER_0_150_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_616 ();
 DECAPx4_ASAP7_75t_R FILLER_0_150_629 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_651 ();
 FILLER_ASAP7_75t_R FILLER_0_150_665 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_670 ();
 FILLER_ASAP7_75t_R FILLER_0_150_676 ();
 FILLER_ASAP7_75t_R FILLER_0_150_688 ();
 FILLER_ASAP7_75t_R FILLER_0_150_700 ();
 FILLER_ASAP7_75t_R FILLER_0_150_710 ();
 DECAPx6_ASAP7_75t_R FILLER_0_150_718 ();
 FILLER_ASAP7_75t_R FILLER_0_150_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_734 ();
 FILLER_ASAP7_75t_R FILLER_0_150_741 ();
 FILLER_ASAP7_75t_R FILLER_0_150_749 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_757 ();
 FILLER_ASAP7_75t_R FILLER_0_150_763 ();
 FILLER_ASAP7_75t_R FILLER_0_150_772 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_787 ();
 FILLER_ASAP7_75t_R FILLER_0_150_795 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_810 ();
 FILLER_ASAP7_75t_R FILLER_0_150_823 ();
 DECAPx1_ASAP7_75t_R FILLER_0_150_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_832 ();
 FILLER_ASAP7_75t_R FILLER_0_150_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_841 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_848 ();
 FILLER_ASAP7_75t_R FILLER_0_150_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_856 ();
 FILLER_ASAP7_75t_R FILLER_0_150_863 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_894 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_916 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_922 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_935 ();
 DECAPx6_ASAP7_75t_R FILLER_0_150_957 ();
 FILLER_ASAP7_75t_R FILLER_0_150_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_1015 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_1037 ();
 FILLER_ASAP7_75t_R FILLER_0_150_1046 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_1053 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_1075 ();
 FILLER_ASAP7_75t_R FILLER_0_150_1081 ();
 DECAPx4_ASAP7_75t_R FILLER_0_150_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_1104 ();
 DECAPx6_ASAP7_75t_R FILLER_0_150_1113 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_1127 ();
 DECAPx4_ASAP7_75t_R FILLER_0_150_1143 ();
 FILLER_ASAP7_75t_R FILLER_0_150_1158 ();
 FILLER_ASAP7_75t_R FILLER_0_150_1170 ();
 FILLER_ASAP7_75t_R FILLER_0_150_1182 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_1190 ();
 FILLER_ASAP7_75t_R FILLER_0_150_1196 ();
 DECAPx6_ASAP7_75t_R FILLER_0_150_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_1218 ();
 DECAPx4_ASAP7_75t_R FILLER_0_150_1225 ();
 FILLER_ASAP7_75t_R FILLER_0_150_1235 ();
 DECAPx4_ASAP7_75t_R FILLER_0_150_1241 ();
 FILLER_ASAP7_75t_R FILLER_0_150_1251 ();
 DECAPx6_ASAP7_75t_R FILLER_0_150_1259 ();
 FILLER_ASAP7_75t_R FILLER_0_150_1273 ();
 DECAPx4_ASAP7_75t_R FILLER_0_150_1281 ();
 FILLER_ASAP7_75t_R FILLER_0_150_1291 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_1293 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_1304 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_1310 ();
 DECAPx2_ASAP7_75t_R FILLER_0_150_1321 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_1327 ();
 DECAPx1_ASAP7_75t_R FILLER_0_150_1339 ();
 FILLER_ASAP7_75t_R FILLER_0_150_1351 ();
 FILLER_ASAP7_75t_R FILLER_0_150_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_150_1365 ();
 FILLER_ASAP7_75t_R FILLER_0_150_1372 ();
 FILLER_ASAP7_75t_R FILLER_0_150_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_151_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_4 ();
 FILLER_ASAP7_75t_R FILLER_0_151_8 ();
 FILLER_ASAP7_75t_R FILLER_0_151_15 ();
 FILLER_ASAP7_75t_R FILLER_0_151_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_22 ();
 DECAPx2_ASAP7_75t_R FILLER_0_151_29 ();
 FILLER_ASAP7_75t_R FILLER_0_151_35 ();
 DECAPx2_ASAP7_75t_R FILLER_0_151_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_49 ();
 DECAPx2_ASAP7_75t_R FILLER_0_151_62 ();
 FILLER_ASAP7_75t_R FILLER_0_151_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_70 ();
 DECAPx1_ASAP7_75t_R FILLER_0_151_81 ();
 DECAPx6_ASAP7_75t_R FILLER_0_151_93 ();
 DECAPx1_ASAP7_75t_R FILLER_0_151_107 ();
 DECAPx2_ASAP7_75t_R FILLER_0_151_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_123 ();
 FILLER_ASAP7_75t_R FILLER_0_151_132 ();
 FILLER_ASAP7_75t_R FILLER_0_151_142 ();
 DECAPx2_ASAP7_75t_R FILLER_0_151_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_156 ();
 DECAPx2_ASAP7_75t_R FILLER_0_151_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_169 ();
 FILLER_ASAP7_75t_R FILLER_0_151_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_184 ();
 DECAPx4_ASAP7_75t_R FILLER_0_151_191 ();
 FILLER_ASAP7_75t_R FILLER_0_151_207 ();
 DECAPx6_ASAP7_75t_R FILLER_0_151_217 ();
 FILLER_ASAP7_75t_R FILLER_0_151_231 ();
 DECAPx6_ASAP7_75t_R FILLER_0_151_239 ();
 FILLER_ASAP7_75t_R FILLER_0_151_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_255 ();
 DECAPx4_ASAP7_75t_R FILLER_0_151_259 ();
 FILLER_ASAP7_75t_R FILLER_0_151_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_271 ();
 DECAPx2_ASAP7_75t_R FILLER_0_151_278 ();
 FILLER_ASAP7_75t_R FILLER_0_151_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_286 ();
 DECAPx4_ASAP7_75t_R FILLER_0_151_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_305 ();
 DECAPx6_ASAP7_75t_R FILLER_0_151_314 ();
 FILLER_ASAP7_75t_R FILLER_0_151_328 ();
 FILLER_ASAP7_75t_R FILLER_0_151_340 ();
 FILLER_ASAP7_75t_R FILLER_0_151_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_374 ();
 DECAPx6_ASAP7_75t_R FILLER_0_151_396 ();
 FILLER_ASAP7_75t_R FILLER_0_151_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_412 ();
 DECAPx6_ASAP7_75t_R FILLER_0_151_423 ();
 FILLER_ASAP7_75t_R FILLER_0_151_437 ();
 FILLER_ASAP7_75t_R FILLER_0_151_442 ();
 DECAPx6_ASAP7_75t_R FILLER_0_151_452 ();
 FILLER_ASAP7_75t_R FILLER_0_151_466 ();
 FILLER_ASAP7_75t_R FILLER_0_151_474 ();
 FILLER_ASAP7_75t_R FILLER_0_151_482 ();
 DECAPx2_ASAP7_75t_R FILLER_0_151_490 ();
 FILLER_ASAP7_75t_R FILLER_0_151_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_498 ();
 DECAPx2_ASAP7_75t_R FILLER_0_151_520 ();
 FILLER_ASAP7_75t_R FILLER_0_151_538 ();
 DECAPx2_ASAP7_75t_R FILLER_0_151_561 ();
 FILLER_ASAP7_75t_R FILLER_0_151_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_569 ();
 DECAPx4_ASAP7_75t_R FILLER_0_151_592 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_610 ();
 DECAPx4_ASAP7_75t_R FILLER_0_151_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_642 ();
 FILLER_ASAP7_75t_R FILLER_0_151_655 ();
 DECAPx2_ASAP7_75t_R FILLER_0_151_660 ();
 FILLER_ASAP7_75t_R FILLER_0_151_672 ();
 DECAPx1_ASAP7_75t_R FILLER_0_151_686 ();
 FILLER_ASAP7_75t_R FILLER_0_151_702 ();
 FILLER_ASAP7_75t_R FILLER_0_151_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_712 ();
 FILLER_ASAP7_75t_R FILLER_0_151_725 ();
 FILLER_ASAP7_75t_R FILLER_0_151_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_734 ();
 FILLER_ASAP7_75t_R FILLER_0_151_745 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_754 ();
 FILLER_ASAP7_75t_R FILLER_0_151_776 ();
 FILLER_ASAP7_75t_R FILLER_0_151_789 ();
 FILLER_ASAP7_75t_R FILLER_0_151_797 ();
 FILLER_ASAP7_75t_R FILLER_0_151_805 ();
 FILLER_ASAP7_75t_R FILLER_0_151_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_815 ();
 DECAPx1_ASAP7_75t_R FILLER_0_151_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_826 ();
 FILLER_ASAP7_75t_R FILLER_0_151_830 ();
 FILLER_ASAP7_75t_R FILLER_0_151_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_845 ();
 DECAPx1_ASAP7_75t_R FILLER_0_151_853 ();
 DECAPx1_ASAP7_75t_R FILLER_0_151_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_873 ();
 FILLER_ASAP7_75t_R FILLER_0_151_880 ();
 DECAPx2_ASAP7_75t_R FILLER_0_151_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_894 ();
 FILLER_ASAP7_75t_R FILLER_0_151_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_903 ();
 FILLER_ASAP7_75t_R FILLER_0_151_910 ();
 FILLER_ASAP7_75t_R FILLER_0_151_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_924 ();
 DECAPx1_ASAP7_75t_R FILLER_0_151_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_931 ();
 FILLER_ASAP7_75t_R FILLER_0_151_938 ();
 DECAPx1_ASAP7_75t_R FILLER_0_151_946 ();
 FILLER_ASAP7_75t_R FILLER_0_151_958 ();
 DECAPx2_ASAP7_75t_R FILLER_0_151_968 ();
 DECAPx2_ASAP7_75t_R FILLER_0_151_982 ();
 FILLER_ASAP7_75t_R FILLER_0_151_988 ();
 FILLER_ASAP7_75t_R FILLER_0_151_993 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1003 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_1008 ();
 DECAPx2_ASAP7_75t_R FILLER_0_151_1030 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1036 ();
 DECAPx4_ASAP7_75t_R FILLER_0_151_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_1054 ();
 DECAPx4_ASAP7_75t_R FILLER_0_151_1061 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1081 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1094 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1104 ();
 DECAPx2_ASAP7_75t_R FILLER_0_151_1112 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_1118 ();
 DECAPx2_ASAP7_75t_R FILLER_0_151_1129 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_1137 ();
 DECAPx2_ASAP7_75t_R FILLER_0_151_1148 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1154 ();
 DECAPx2_ASAP7_75t_R FILLER_0_151_1166 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1172 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1180 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1188 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1196 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1204 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1212 ();
 DECAPx2_ASAP7_75t_R FILLER_0_151_1220 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1233 ();
 DECAPx4_ASAP7_75t_R FILLER_0_151_1242 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_1252 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1259 ();
 DECAPx2_ASAP7_75t_R FILLER_0_151_1271 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_1277 ();
 DECAPx2_ASAP7_75t_R FILLER_0_151_1288 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1299 ();
 DECAPx2_ASAP7_75t_R FILLER_0_151_1311 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1325 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1333 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1341 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_1343 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1347 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1354 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1360 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1367 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1374 ();
 FILLER_ASAP7_75t_R FILLER_0_151_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_152_2 ();
 FILLER_ASAP7_75t_R FILLER_0_152_9 ();
 FILLER_ASAP7_75t_R FILLER_0_152_16 ();
 FILLER_ASAP7_75t_R FILLER_0_152_23 ();
 FILLER_ASAP7_75t_R FILLER_0_152_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_152_61 ();
 DECAPx1_ASAP7_75t_R FILLER_0_152_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_77 ();
 DECAPx1_ASAP7_75t_R FILLER_0_152_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_90 ();
 DECAPx4_ASAP7_75t_R FILLER_0_152_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_112 ();
 FILLER_ASAP7_75t_R FILLER_0_152_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_122 ();
 FILLER_ASAP7_75t_R FILLER_0_152_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_133 ();
 FILLER_ASAP7_75t_R FILLER_0_152_142 ();
 FILLER_ASAP7_75t_R FILLER_0_152_155 ();
 DECAPx2_ASAP7_75t_R FILLER_0_152_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_169 ();
 DECAPx6_ASAP7_75t_R FILLER_0_152_182 ();
 FILLER_ASAP7_75t_R FILLER_0_152_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_198 ();
 DECAPx6_ASAP7_75t_R FILLER_0_152_205 ();
 FILLER_ASAP7_75t_R FILLER_0_152_219 ();
 DECAPx1_ASAP7_75t_R FILLER_0_152_231 ();
 FILLER_ASAP7_75t_R FILLER_0_152_257 ();
 FILLER_ASAP7_75t_R FILLER_0_152_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_272 ();
 FILLER_ASAP7_75t_R FILLER_0_152_276 ();
 FILLER_ASAP7_75t_R FILLER_0_152_284 ();
 DECAPx10_ASAP7_75t_R FILLER_0_152_292 ();
 FILLER_ASAP7_75t_R FILLER_0_152_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_316 ();
 DECAPx2_ASAP7_75t_R FILLER_0_152_322 ();
 FILLER_ASAP7_75t_R FILLER_0_152_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_330 ();
 FILLER_ASAP7_75t_R FILLER_0_152_336 ();
 FILLER_ASAP7_75t_R FILLER_0_152_348 ();
 DECAPx6_ASAP7_75t_R FILLER_0_152_356 ();
 FILLER_ASAP7_75t_R FILLER_0_152_370 ();
 DECAPx1_ASAP7_75t_R FILLER_0_152_380 ();
 FILLER_ASAP7_75t_R FILLER_0_152_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_396 ();
 FILLER_ASAP7_75t_R FILLER_0_152_405 ();
 FILLER_ASAP7_75t_R FILLER_0_152_414 ();
 FILLER_ASAP7_75t_R FILLER_0_152_422 ();
 DECAPx1_ASAP7_75t_R FILLER_0_152_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_436 ();
 FILLER_ASAP7_75t_R FILLER_0_152_442 ();
 DECAPx4_ASAP7_75t_R FILLER_0_152_450 ();
 FILLER_ASAP7_75t_R FILLER_0_152_460 ();
 FILLER_ASAP7_75t_R FILLER_0_152_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_152_473 ();
 FILLER_ASAP7_75t_R FILLER_0_152_495 ();
 FILLER_ASAP7_75t_R FILLER_0_152_505 ();
 DECAPx2_ASAP7_75t_R FILLER_0_152_519 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_525 ();
 FILLER_ASAP7_75t_R FILLER_0_152_538 ();
 DECAPx1_ASAP7_75t_R FILLER_0_152_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_550 ();
 DECAPx2_ASAP7_75t_R FILLER_0_152_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_578 ();
 FILLER_ASAP7_75t_R FILLER_0_152_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_587 ();
 FILLER_ASAP7_75t_R FILLER_0_152_591 ();
 FILLER_ASAP7_75t_R FILLER_0_152_615 ();
 FILLER_ASAP7_75t_R FILLER_0_152_638 ();
 FILLER_ASAP7_75t_R FILLER_0_152_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_653 ();
 FILLER_ASAP7_75t_R FILLER_0_152_675 ();
 FILLER_ASAP7_75t_R FILLER_0_152_687 ();
 FILLER_ASAP7_75t_R FILLER_0_152_697 ();
 DECAPx1_ASAP7_75t_R FILLER_0_152_705 ();
 DECAPx1_ASAP7_75t_R FILLER_0_152_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_720 ();
 FILLER_ASAP7_75t_R FILLER_0_152_739 ();
 FILLER_ASAP7_75t_R FILLER_0_152_747 ();
 DECAPx4_ASAP7_75t_R FILLER_0_152_754 ();
 FILLER_ASAP7_75t_R FILLER_0_152_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_766 ();
 FILLER_ASAP7_75t_R FILLER_0_152_774 ();
 DECAPx6_ASAP7_75t_R FILLER_0_152_783 ();
 DECAPx1_ASAP7_75t_R FILLER_0_152_797 ();
 DECAPx4_ASAP7_75t_R FILLER_0_152_807 ();
 FILLER_ASAP7_75t_R FILLER_0_152_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_819 ();
 DECAPx2_ASAP7_75t_R FILLER_0_152_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_832 ();
 FILLER_ASAP7_75t_R FILLER_0_152_843 ();
 DECAPx4_ASAP7_75t_R FILLER_0_152_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_861 ();
 DECAPx1_ASAP7_75t_R FILLER_0_152_868 ();
 DECAPx1_ASAP7_75t_R FILLER_0_152_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_882 ();
 DECAPx1_ASAP7_75t_R FILLER_0_152_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_897 ();
 DECAPx1_ASAP7_75t_R FILLER_0_152_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_908 ();
 DECAPx2_ASAP7_75t_R FILLER_0_152_915 ();
 FILLER_ASAP7_75t_R FILLER_0_152_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_923 ();
 FILLER_ASAP7_75t_R FILLER_0_152_936 ();
 DECAPx6_ASAP7_75t_R FILLER_0_152_946 ();
 DECAPx1_ASAP7_75t_R FILLER_0_152_960 ();
 DECAPx4_ASAP7_75t_R FILLER_0_152_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_980 ();
 DECAPx6_ASAP7_75t_R FILLER_0_152_987 ();
 DECAPx2_ASAP7_75t_R FILLER_0_152_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_1007 ();
 FILLER_ASAP7_75t_R FILLER_0_152_1014 ();
 FILLER_ASAP7_75t_R FILLER_0_152_1037 ();
 DECAPx6_ASAP7_75t_R FILLER_0_152_1049 ();
 FILLER_ASAP7_75t_R FILLER_0_152_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_0_152_1086 ();
 FILLER_ASAP7_75t_R FILLER_0_152_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_1094 ();
 FILLER_ASAP7_75t_R FILLER_0_152_1103 ();
 DECAPx1_ASAP7_75t_R FILLER_0_152_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_1115 ();
 DECAPx2_ASAP7_75t_R FILLER_0_152_1124 ();
 FILLER_ASAP7_75t_R FILLER_0_152_1130 ();
 DECAPx6_ASAP7_75t_R FILLER_0_152_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_1154 ();
 DECAPx1_ASAP7_75t_R FILLER_0_152_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_1169 ();
 FILLER_ASAP7_75t_R FILLER_0_152_1180 ();
 DECAPx1_ASAP7_75t_R FILLER_0_152_1188 ();
 FILLER_ASAP7_75t_R FILLER_0_152_1199 ();
 DECAPx4_ASAP7_75t_R FILLER_0_152_1207 ();
 FILLER_ASAP7_75t_R FILLER_0_152_1223 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_1225 ();
 FILLER_ASAP7_75t_R FILLER_0_152_1232 ();
 DECAPx6_ASAP7_75t_R FILLER_0_152_1241 ();
 FILLER_ASAP7_75t_R FILLER_0_152_1255 ();
 DECAPx1_ASAP7_75t_R FILLER_0_152_1265 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_1269 ();
 DECAPx4_ASAP7_75t_R FILLER_0_152_1278 ();
 FILLER_ASAP7_75t_R FILLER_0_152_1288 ();
 DECAPx1_ASAP7_75t_R FILLER_0_152_1298 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_1302 ();
 FILLER_ASAP7_75t_R FILLER_0_152_1310 ();
 DECAPx2_ASAP7_75t_R FILLER_0_152_1318 ();
 FILLER_ASAP7_75t_R FILLER_0_152_1329 ();
 FILLER_ASAP7_75t_R FILLER_0_152_1343 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152_1345 ();
 FILLER_ASAP7_75t_R FILLER_0_152_1349 ();
 FILLER_ASAP7_75t_R FILLER_0_152_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_152_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_153_2 ();
 FILLER_ASAP7_75t_R FILLER_0_153_9 ();
 FILLER_ASAP7_75t_R FILLER_0_153_16 ();
 DECAPx1_ASAP7_75t_R FILLER_0_153_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_153_27 ();
 FILLER_ASAP7_75t_R FILLER_0_153_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_153_52 ();
 DECAPx1_ASAP7_75t_R FILLER_0_153_59 ();
 DECAPx10_ASAP7_75t_R FILLER_0_153_69 ();
 DECAPx10_ASAP7_75t_R FILLER_0_153_91 ();
 DECAPx6_ASAP7_75t_R FILLER_0_153_113 ();
 DECAPx2_ASAP7_75t_R FILLER_0_153_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_153_133 ();
 DECAPx6_ASAP7_75t_R FILLER_0_153_142 ();
 DECAPx10_ASAP7_75t_R FILLER_0_153_164 ();
 DECAPx2_ASAP7_75t_R FILLER_0_153_186 ();
 FILLER_ASAP7_75t_R FILLER_0_153_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_153_194 ();
 FILLER_ASAP7_75t_R FILLER_0_153_207 ();
 DECAPx4_ASAP7_75t_R FILLER_0_153_219 ();
 DECAPx1_ASAP7_75t_R FILLER_0_153_233 ();
 DECAPx2_ASAP7_75t_R FILLER_0_153_240 ();
 FILLER_ASAP7_75t_R FILLER_0_153_254 ();
 FILLER_ASAP7_75t_R FILLER_0_153_274 ();
 FILLER_ASAP7_75t_R FILLER_0_153_284 ();
 DECAPx6_ASAP7_75t_R FILLER_0_153_292 ();
 DECAPx4_ASAP7_75t_R FILLER_0_153_312 ();
 FILLER_ASAP7_75t_R FILLER_0_153_322 ();
 DECAPx2_ASAP7_75t_R FILLER_0_153_330 ();
 FILLER_ASAP7_75t_R FILLER_0_153_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_153_338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_153_344 ();
 FILLER_ASAP7_75t_R FILLER_0_153_366 ();
 FILLER_ASAP7_75t_R FILLER_0_153_375 ();
 DECAPx4_ASAP7_75t_R FILLER_0_153_387 ();
 FILLER_ASAP7_75t_R FILLER_0_153_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_153_399 ();
 FILLER_ASAP7_75t_R FILLER_0_153_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_153_408 ();
 FILLER_ASAP7_75t_R FILLER_0_153_415 ();
 DECAPx1_ASAP7_75t_R FILLER_0_153_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_153_429 ();
 DECAPx2_ASAP7_75t_R FILLER_0_153_436 ();
 FILLER_ASAP7_75t_R FILLER_0_153_442 ();
 FILLER_ASAP7_75t_R FILLER_0_153_450 ();
 DECAPx2_ASAP7_75t_R FILLER_0_153_455 ();
 FILLER_ASAP7_75t_R FILLER_0_153_461 ();
 FILLER_ASAP7_75t_R FILLER_0_153_471 ();
 DECAPx6_ASAP7_75t_R FILLER_0_153_476 ();
 DECAPx1_ASAP7_75t_R FILLER_0_153_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_153_494 ();
 FILLER_ASAP7_75t_R FILLER_0_153_501 ();
 DECAPx2_ASAP7_75t_R FILLER_0_153_508 ();
 DECAPx2_ASAP7_75t_R FILLER_0_153_526 ();
 DECAPx1_ASAP7_75t_R FILLER_0_153_544 ();
 DECAPx4_ASAP7_75t_R FILLER_0_153_554 ();
 FILLER_ASAP7_75t_R FILLER_0_153_564 ();
 FILLER_ASAP7_75t_R FILLER_0_153_569 ();
 DECAPx6_ASAP7_75t_R FILLER_0_153_592 ();
 FILLER_ASAP7_75t_R FILLER_0_153_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_153_608 ();
 FILLER_ASAP7_75t_R FILLER_0_153_612 ();
 FILLER_ASAP7_75t_R FILLER_0_153_619 ();
 DECAPx6_ASAP7_75t_R FILLER_0_153_624 ();
 FILLER_ASAP7_75t_R FILLER_0_153_644 ();
 FILLER_ASAP7_75t_R FILLER_0_153_667 ();
 FILLER_ASAP7_75t_R FILLER_0_153_675 ();
 DECAPx2_ASAP7_75t_R FILLER_0_153_687 ();
 FILLER_ASAP7_75t_R FILLER_0_153_693 ();
 FILLER_ASAP7_75t_R FILLER_0_153_701 ();
 FILLER_ASAP7_75t_R FILLER_0_153_709 ();
 FILLER_ASAP7_75t_R FILLER_0_153_716 ();
 FILLER_ASAP7_75t_R FILLER_0_153_724 ();
 FILLER_ASAP7_75t_R FILLER_0_153_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_153_731 ();
 FILLER_ASAP7_75t_R FILLER_0_153_738 ();
 FILLER_ASAP7_75t_R FILLER_0_153_746 ();
 DECAPx4_ASAP7_75t_R FILLER_0_153_753 ();
 FILLER_ASAP7_75t_R FILLER_0_153_763 ();
 DECAPx6_ASAP7_75t_R FILLER_0_153_771 ();
 FILLER_ASAP7_75t_R FILLER_0_153_788 ();
 FILLER_ASAP7_75t_R FILLER_0_153_800 ();
 DECAPx6_ASAP7_75t_R FILLER_0_153_812 ();
 FILLER_ASAP7_75t_R FILLER_0_153_826 ();
 DECAPx10_ASAP7_75t_R FILLER_0_153_834 ();
 DECAPx10_ASAP7_75t_R FILLER_0_153_856 ();
 DECAPx2_ASAP7_75t_R FILLER_0_153_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_153_890 ();
 DECAPx6_ASAP7_75t_R FILLER_0_153_897 ();
 FILLER_ASAP7_75t_R FILLER_0_153_911 ();
 FILLER_ASAP7_75t_R FILLER_0_153_923 ();
 DECAPx4_ASAP7_75t_R FILLER_0_153_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_153_937 ();
 DECAPx2_ASAP7_75t_R FILLER_0_153_944 ();
 FILLER_ASAP7_75t_R FILLER_0_153_958 ();
 FILLER_ASAP7_75t_R FILLER_0_153_966 ();
 FILLER_ASAP7_75t_R FILLER_0_153_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_153_976 ();
 DECAPx1_ASAP7_75t_R FILLER_0_153_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_153_988 ();
 DECAPx2_ASAP7_75t_R FILLER_0_153_997 ();
 FILLER_ASAP7_75t_R FILLER_0_153_1003 ();
 DECAPx1_ASAP7_75t_R FILLER_0_153_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_153_1017 ();
 DECAPx4_ASAP7_75t_R FILLER_0_153_1021 ();
 FILLER_ASAP7_75t_R FILLER_0_153_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_153_1033 ();
 FILLER_ASAP7_75t_R FILLER_0_153_1044 ();
 FILLER_ASAP7_75t_R FILLER_0_153_1064 ();
 FILLER_ASAP7_75t_R FILLER_0_153_1074 ();
 DECAPx4_ASAP7_75t_R FILLER_0_153_1082 ();
 FILLER_ASAP7_75t_R FILLER_0_153_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_153_1094 ();
 DECAPx4_ASAP7_75t_R FILLER_0_153_1105 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_153_1115 ();
 DECAPx10_ASAP7_75t_R FILLER_0_153_1122 ();
 DECAPx6_ASAP7_75t_R FILLER_0_153_1144 ();
 FILLER_ASAP7_75t_R FILLER_0_153_1158 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_153_1160 ();
 FILLER_ASAP7_75t_R FILLER_0_153_1171 ();
 DECAPx2_ASAP7_75t_R FILLER_0_153_1178 ();
 FILLER_ASAP7_75t_R FILLER_0_153_1190 ();
 FILLER_ASAP7_75t_R FILLER_0_153_1198 ();
 FILLER_ASAP7_75t_R FILLER_0_153_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_153_1208 ();
 FILLER_ASAP7_75t_R FILLER_0_153_1216 ();
 DECAPx1_ASAP7_75t_R FILLER_0_153_1225 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_153_1229 ();
 DECAPx4_ASAP7_75t_R FILLER_0_153_1237 ();
 FILLER_ASAP7_75t_R FILLER_0_153_1247 ();
 FILLER_ASAP7_75t_R FILLER_0_153_1254 ();
 DECAPx2_ASAP7_75t_R FILLER_0_153_1264 ();
 FILLER_ASAP7_75t_R FILLER_0_153_1270 ();
 DECAPx1_ASAP7_75t_R FILLER_0_153_1283 ();
 FILLER_ASAP7_75t_R FILLER_0_153_1294 ();
 DECAPx2_ASAP7_75t_R FILLER_0_153_1302 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_153_1308 ();
 FILLER_ASAP7_75t_R FILLER_0_153_1314 ();
 FILLER_ASAP7_75t_R FILLER_0_153_1338 ();
 FILLER_ASAP7_75t_R FILLER_0_153_1361 ();
 FILLER_ASAP7_75t_R FILLER_0_153_1366 ();
 FILLER_ASAP7_75t_R FILLER_0_153_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_153_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_154_2 ();
 FILLER_ASAP7_75t_R FILLER_0_154_9 ();
 FILLER_ASAP7_75t_R FILLER_0_154_16 ();
 DECAPx1_ASAP7_75t_R FILLER_0_154_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_27 ();
 FILLER_ASAP7_75t_R FILLER_0_154_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_52 ();
 FILLER_ASAP7_75t_R FILLER_0_154_65 ();
 DECAPx10_ASAP7_75t_R FILLER_0_154_73 ();
 FILLER_ASAP7_75t_R FILLER_0_154_101 ();
 FILLER_ASAP7_75t_R FILLER_0_154_109 ();
 DECAPx4_ASAP7_75t_R FILLER_0_154_123 ();
 FILLER_ASAP7_75t_R FILLER_0_154_133 ();
 DECAPx10_ASAP7_75t_R FILLER_0_154_145 ();
 DECAPx4_ASAP7_75t_R FILLER_0_154_167 ();
 FILLER_ASAP7_75t_R FILLER_0_154_177 ();
 DECAPx4_ASAP7_75t_R FILLER_0_154_182 ();
 FILLER_ASAP7_75t_R FILLER_0_154_204 ();
 DECAPx2_ASAP7_75t_R FILLER_0_154_212 ();
 FILLER_ASAP7_75t_R FILLER_0_154_230 ();
 DECAPx6_ASAP7_75t_R FILLER_0_154_242 ();
 FILLER_ASAP7_75t_R FILLER_0_154_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_258 ();
 FILLER_ASAP7_75t_R FILLER_0_154_265 ();
 DECAPx6_ASAP7_75t_R FILLER_0_154_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_287 ();
 FILLER_ASAP7_75t_R FILLER_0_154_295 ();
 DECAPx6_ASAP7_75t_R FILLER_0_154_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_317 ();
 FILLER_ASAP7_75t_R FILLER_0_154_324 ();
 DECAPx2_ASAP7_75t_R FILLER_0_154_329 ();
 DECAPx1_ASAP7_75t_R FILLER_0_154_341 ();
 DECAPx6_ASAP7_75t_R FILLER_0_154_355 ();
 DECAPx2_ASAP7_75t_R FILLER_0_154_369 ();
 DECAPx2_ASAP7_75t_R FILLER_0_154_381 ();
 DECAPx6_ASAP7_75t_R FILLER_0_154_393 ();
 FILLER_ASAP7_75t_R FILLER_0_154_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_409 ();
 DECAPx1_ASAP7_75t_R FILLER_0_154_416 ();
 FILLER_ASAP7_75t_R FILLER_0_154_426 ();
 FILLER_ASAP7_75t_R FILLER_0_154_434 ();
 DECAPx2_ASAP7_75t_R FILLER_0_154_442 ();
 FILLER_ASAP7_75t_R FILLER_0_154_448 ();
 DECAPx1_ASAP7_75t_R FILLER_0_154_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_461 ();
 FILLER_ASAP7_75t_R FILLER_0_154_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_154_474 ();
 DECAPx2_ASAP7_75t_R FILLER_0_154_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_154_506 ();
 DECAPx6_ASAP7_75t_R FILLER_0_154_528 ();
 DECAPx10_ASAP7_75t_R FILLER_0_154_545 ();
 DECAPx1_ASAP7_75t_R FILLER_0_154_567 ();
 FILLER_ASAP7_75t_R FILLER_0_154_574 ();
 DECAPx4_ASAP7_75t_R FILLER_0_154_581 ();
 DECAPx10_ASAP7_75t_R FILLER_0_154_601 ();
 DECAPx10_ASAP7_75t_R FILLER_0_154_623 ();
 FILLER_ASAP7_75t_R FILLER_0_154_645 ();
 FILLER_ASAP7_75t_R FILLER_0_154_668 ();
 FILLER_ASAP7_75t_R FILLER_0_154_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_675 ();
 FILLER_ASAP7_75t_R FILLER_0_154_688 ();
 FILLER_ASAP7_75t_R FILLER_0_154_696 ();
 FILLER_ASAP7_75t_R FILLER_0_154_703 ();
 DECAPx2_ASAP7_75t_R FILLER_0_154_711 ();
 FILLER_ASAP7_75t_R FILLER_0_154_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_719 ();
 FILLER_ASAP7_75t_R FILLER_0_154_726 ();
 DECAPx2_ASAP7_75t_R FILLER_0_154_734 ();
 FILLER_ASAP7_75t_R FILLER_0_154_740 ();
 DECAPx2_ASAP7_75t_R FILLER_0_154_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_756 ();
 FILLER_ASAP7_75t_R FILLER_0_154_764 ();
 DECAPx4_ASAP7_75t_R FILLER_0_154_773 ();
 FILLER_ASAP7_75t_R FILLER_0_154_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_785 ();
 DECAPx2_ASAP7_75t_R FILLER_0_154_792 ();
 FILLER_ASAP7_75t_R FILLER_0_154_798 ();
 DECAPx6_ASAP7_75t_R FILLER_0_154_810 ();
 FILLER_ASAP7_75t_R FILLER_0_154_830 ();
 FILLER_ASAP7_75t_R FILLER_0_154_839 ();
 DECAPx1_ASAP7_75t_R FILLER_0_154_847 ();
 FILLER_ASAP7_75t_R FILLER_0_154_858 ();
 FILLER_ASAP7_75t_R FILLER_0_154_866 ();
 DECAPx4_ASAP7_75t_R FILLER_0_154_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_884 ();
 FILLER_ASAP7_75t_R FILLER_0_154_905 ();
 DECAPx1_ASAP7_75t_R FILLER_0_154_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_917 ();
 FILLER_ASAP7_75t_R FILLER_0_154_928 ();
 FILLER_ASAP7_75t_R FILLER_0_154_940 ();
 DECAPx2_ASAP7_75t_R FILLER_0_154_952 ();
 FILLER_ASAP7_75t_R FILLER_0_154_958 ();
 DECAPx2_ASAP7_75t_R FILLER_0_154_966 ();
 DECAPx1_ASAP7_75t_R FILLER_0_154_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_987 ();
 DECAPx6_ASAP7_75t_R FILLER_0_154_994 ();
 FILLER_ASAP7_75t_R FILLER_0_154_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_1010 ();
 FILLER_ASAP7_75t_R FILLER_0_154_1017 ();
 FILLER_ASAP7_75t_R FILLER_0_154_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_1032 ();
 FILLER_ASAP7_75t_R FILLER_0_154_1041 ();
 DECAPx2_ASAP7_75t_R FILLER_0_154_1049 ();
 FILLER_ASAP7_75t_R FILLER_0_154_1055 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_1057 ();
 DECAPx1_ASAP7_75t_R FILLER_0_154_1066 ();
 DECAPx6_ASAP7_75t_R FILLER_0_154_1081 ();
 FILLER_ASAP7_75t_R FILLER_0_154_1095 ();
 FILLER_ASAP7_75t_R FILLER_0_154_1108 ();
 DECAPx4_ASAP7_75t_R FILLER_0_154_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_1131 ();
 FILLER_ASAP7_75t_R FILLER_0_154_1142 ();
 DECAPx2_ASAP7_75t_R FILLER_0_154_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_1156 ();
 DECAPx1_ASAP7_75t_R FILLER_0_154_1177 ();
 FILLER_ASAP7_75t_R FILLER_0_154_1191 ();
 FILLER_ASAP7_75t_R FILLER_0_154_1199 ();
 DECAPx1_ASAP7_75t_R FILLER_0_154_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_1211 ();
 DECAPx4_ASAP7_75t_R FILLER_0_154_1223 ();
 FILLER_ASAP7_75t_R FILLER_0_154_1233 ();
 FILLER_ASAP7_75t_R FILLER_0_154_1241 ();
 DECAPx2_ASAP7_75t_R FILLER_0_154_1249 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_1255 ();
 DECAPx1_ASAP7_75t_R FILLER_0_154_1262 ();
 FILLER_ASAP7_75t_R FILLER_0_154_1273 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_1275 ();
 FILLER_ASAP7_75t_R FILLER_0_154_1282 ();
 DECAPx2_ASAP7_75t_R FILLER_0_154_1289 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_1295 ();
 FILLER_ASAP7_75t_R FILLER_0_154_1302 ();
 FILLER_ASAP7_75t_R FILLER_0_154_1310 ();
 FILLER_ASAP7_75t_R FILLER_0_154_1317 ();
 FILLER_ASAP7_75t_R FILLER_0_154_1325 ();
 FILLER_ASAP7_75t_R FILLER_0_154_1338 ();
 FILLER_ASAP7_75t_R FILLER_0_154_1343 ();
 FILLER_ASAP7_75t_R FILLER_0_154_1351 ();
 FILLER_ASAP7_75t_R FILLER_0_154_1356 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154_1358 ();
 FILLER_ASAP7_75t_R FILLER_0_154_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_155_2 ();
 FILLER_ASAP7_75t_R FILLER_0_155_9 ();
 FILLER_ASAP7_75t_R FILLER_0_155_16 ();
 FILLER_ASAP7_75t_R FILLER_0_155_21 ();
 FILLER_ASAP7_75t_R FILLER_0_155_28 ();
 DECAPx1_ASAP7_75t_R FILLER_0_155_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_37 ();
 FILLER_ASAP7_75t_R FILLER_0_155_41 ();
 FILLER_ASAP7_75t_R FILLER_0_155_46 ();
 DECAPx2_ASAP7_75t_R FILLER_0_155_51 ();
 FILLER_ASAP7_75t_R FILLER_0_155_69 ();
 DECAPx2_ASAP7_75t_R FILLER_0_155_79 ();
 FILLER_ASAP7_75t_R FILLER_0_155_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_87 ();
 FILLER_ASAP7_75t_R FILLER_0_155_99 ();
 FILLER_ASAP7_75t_R FILLER_0_155_109 ();
 DECAPx4_ASAP7_75t_R FILLER_0_155_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_129 ();
 FILLER_ASAP7_75t_R FILLER_0_155_136 ();
 DECAPx1_ASAP7_75t_R FILLER_0_155_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_148 ();
 FILLER_ASAP7_75t_R FILLER_0_155_154 ();
 DECAPx1_ASAP7_75t_R FILLER_0_155_166 ();
 FILLER_ASAP7_75t_R FILLER_0_155_180 ();
 DECAPx6_ASAP7_75t_R FILLER_0_155_190 ();
 FILLER_ASAP7_75t_R FILLER_0_155_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_206 ();
 DECAPx4_ASAP7_75t_R FILLER_0_155_218 ();
 FILLER_ASAP7_75t_R FILLER_0_155_228 ();
 DECAPx6_ASAP7_75t_R FILLER_0_155_242 ();
 DECAPx1_ASAP7_75t_R FILLER_0_155_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_260 ();
 DECAPx2_ASAP7_75t_R FILLER_0_155_269 ();
 FILLER_ASAP7_75t_R FILLER_0_155_275 ();
 DECAPx2_ASAP7_75t_R FILLER_0_155_283 ();
 FILLER_ASAP7_75t_R FILLER_0_155_289 ();
 FILLER_ASAP7_75t_R FILLER_0_155_297 ();
 FILLER_ASAP7_75t_R FILLER_0_155_307 ();
 DECAPx2_ASAP7_75t_R FILLER_0_155_312 ();
 FILLER_ASAP7_75t_R FILLER_0_155_326 ();
 FILLER_ASAP7_75t_R FILLER_0_155_335 ();
 DECAPx2_ASAP7_75t_R FILLER_0_155_343 ();
 FILLER_ASAP7_75t_R FILLER_0_155_349 ();
 DECAPx1_ASAP7_75t_R FILLER_0_155_361 ();
 DECAPx2_ASAP7_75t_R FILLER_0_155_375 ();
 FILLER_ASAP7_75t_R FILLER_0_155_381 ();
 FILLER_ASAP7_75t_R FILLER_0_155_389 ();
 FILLER_ASAP7_75t_R FILLER_0_155_399 ();
 DECAPx1_ASAP7_75t_R FILLER_0_155_407 ();
 FILLER_ASAP7_75t_R FILLER_0_155_416 ();
 DECAPx6_ASAP7_75t_R FILLER_0_155_421 ();
 DECAPx2_ASAP7_75t_R FILLER_0_155_442 ();
 DECAPx1_ASAP7_75t_R FILLER_0_155_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_460 ();
 DECAPx10_ASAP7_75t_R FILLER_0_155_467 ();
 DECAPx4_ASAP7_75t_R FILLER_0_155_489 ();
 FILLER_ASAP7_75t_R FILLER_0_155_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_501 ();
 FILLER_ASAP7_75t_R FILLER_0_155_505 ();
 DECAPx10_ASAP7_75t_R FILLER_0_155_513 ();
 DECAPx4_ASAP7_75t_R FILLER_0_155_535 ();
 FILLER_ASAP7_75t_R FILLER_0_155_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_155_556 ();
 DECAPx2_ASAP7_75t_R FILLER_0_155_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_572 ();
 DECAPx10_ASAP7_75t_R FILLER_0_155_576 ();
 DECAPx1_ASAP7_75t_R FILLER_0_155_598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_155_622 ();
 DECAPx6_ASAP7_75t_R FILLER_0_155_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_658 ();
 FILLER_ASAP7_75t_R FILLER_0_155_662 ();
 FILLER_ASAP7_75t_R FILLER_0_155_694 ();
 FILLER_ASAP7_75t_R FILLER_0_155_702 ();
 FILLER_ASAP7_75t_R FILLER_0_155_710 ();
 DECAPx1_ASAP7_75t_R FILLER_0_155_718 ();
 DECAPx2_ASAP7_75t_R FILLER_0_155_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_734 ();
 DECAPx2_ASAP7_75t_R FILLER_0_155_740 ();
 FILLER_ASAP7_75t_R FILLER_0_155_746 ();
 FILLER_ASAP7_75t_R FILLER_0_155_760 ();
 DECAPx6_ASAP7_75t_R FILLER_0_155_769 ();
 FILLER_ASAP7_75t_R FILLER_0_155_791 ();
 DECAPx2_ASAP7_75t_R FILLER_0_155_805 ();
 FILLER_ASAP7_75t_R FILLER_0_155_811 ();
 DECAPx2_ASAP7_75t_R FILLER_0_155_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_825 ();
 FILLER_ASAP7_75t_R FILLER_0_155_832 ();
 DECAPx1_ASAP7_75t_R FILLER_0_155_845 ();
 FILLER_ASAP7_75t_R FILLER_0_155_855 ();
 FILLER_ASAP7_75t_R FILLER_0_155_863 ();
 FILLER_ASAP7_75t_R FILLER_0_155_873 ();
 DECAPx6_ASAP7_75t_R FILLER_0_155_881 ();
 DECAPx1_ASAP7_75t_R FILLER_0_155_895 ();
 DECAPx4_ASAP7_75t_R FILLER_0_155_905 ();
 DECAPx1_ASAP7_75t_R FILLER_0_155_921 ();
 DECAPx2_ASAP7_75t_R FILLER_0_155_927 ();
 FILLER_ASAP7_75t_R FILLER_0_155_939 ();
 DECAPx4_ASAP7_75t_R FILLER_0_155_944 ();
 FILLER_ASAP7_75t_R FILLER_0_155_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_956 ();
 FILLER_ASAP7_75t_R FILLER_0_155_969 ();
 FILLER_ASAP7_75t_R FILLER_0_155_982 ();
 DECAPx2_ASAP7_75t_R FILLER_0_155_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_1002 ();
 DECAPx1_ASAP7_75t_R FILLER_0_155_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_1029 ();
 DECAPx2_ASAP7_75t_R FILLER_0_155_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_1047 ();
 FILLER_ASAP7_75t_R FILLER_0_155_1059 ();
 FILLER_ASAP7_75t_R FILLER_0_155_1064 ();
 DECAPx1_ASAP7_75t_R FILLER_0_155_1069 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_1073 ();
 DECAPx10_ASAP7_75t_R FILLER_0_155_1082 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_1104 ();
 FILLER_ASAP7_75t_R FILLER_0_155_1111 ();
 DECAPx10_ASAP7_75t_R FILLER_0_155_1119 ();
 DECAPx10_ASAP7_75t_R FILLER_0_155_1141 ();
 FILLER_ASAP7_75t_R FILLER_0_155_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_1165 ();
 DECAPx6_ASAP7_75t_R FILLER_0_155_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_1185 ();
 FILLER_ASAP7_75t_R FILLER_0_155_1204 ();
 FILLER_ASAP7_75t_R FILLER_0_155_1212 ();
 DECAPx6_ASAP7_75t_R FILLER_0_155_1220 ();
 FILLER_ASAP7_75t_R FILLER_0_155_1234 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_1236 ();
 DECAPx4_ASAP7_75t_R FILLER_0_155_1243 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_1253 ();
 DECAPx6_ASAP7_75t_R FILLER_0_155_1265 ();
 DECAPx1_ASAP7_75t_R FILLER_0_155_1279 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_1283 ();
 DECAPx1_ASAP7_75t_R FILLER_0_155_1294 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_1298 ();
 FILLER_ASAP7_75t_R FILLER_0_155_1304 ();
 FILLER_ASAP7_75t_R FILLER_0_155_1314 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_1316 ();
 FILLER_ASAP7_75t_R FILLER_0_155_1320 ();
 FILLER_ASAP7_75t_R FILLER_0_155_1328 ();
 FILLER_ASAP7_75t_R FILLER_0_155_1335 ();
 FILLER_ASAP7_75t_R FILLER_0_155_1342 ();
 FILLER_ASAP7_75t_R FILLER_0_155_1350 ();
 FILLER_ASAP7_75t_R FILLER_0_155_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_155_1365 ();
 FILLER_ASAP7_75t_R FILLER_0_155_1372 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155_1374 ();
 FILLER_ASAP7_75t_R FILLER_0_155_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_156_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_4 ();
 FILLER_ASAP7_75t_R FILLER_0_156_11 ();
 FILLER_ASAP7_75t_R FILLER_0_156_16 ();
 FILLER_ASAP7_75t_R FILLER_0_156_23 ();
 FILLER_ASAP7_75t_R FILLER_0_156_30 ();
 FILLER_ASAP7_75t_R FILLER_0_156_35 ();
 DECAPx4_ASAP7_75t_R FILLER_0_156_40 ();
 DECAPx2_ASAP7_75t_R FILLER_0_156_62 ();
 FILLER_ASAP7_75t_R FILLER_0_156_68 ();
 FILLER_ASAP7_75t_R FILLER_0_156_81 ();
 DECAPx2_ASAP7_75t_R FILLER_0_156_93 ();
 FILLER_ASAP7_75t_R FILLER_0_156_99 ();
 FILLER_ASAP7_75t_R FILLER_0_156_107 ();
 DECAPx6_ASAP7_75t_R FILLER_0_156_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_131 ();
 FILLER_ASAP7_75t_R FILLER_0_156_142 ();
 FILLER_ASAP7_75t_R FILLER_0_156_154 ();
 FILLER_ASAP7_75t_R FILLER_0_156_166 ();
 FILLER_ASAP7_75t_R FILLER_0_156_178 ();
 DECAPx6_ASAP7_75t_R FILLER_0_156_188 ();
 DECAPx1_ASAP7_75t_R FILLER_0_156_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_206 ();
 FILLER_ASAP7_75t_R FILLER_0_156_215 ();
 DECAPx4_ASAP7_75t_R FILLER_0_156_224 ();
 FILLER_ASAP7_75t_R FILLER_0_156_240 ();
 DECAPx6_ASAP7_75t_R FILLER_0_156_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_259 ();
 DECAPx2_ASAP7_75t_R FILLER_0_156_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_276 ();
 FILLER_ASAP7_75t_R FILLER_0_156_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_287 ();
 DECAPx1_ASAP7_75t_R FILLER_0_156_294 ();
 FILLER_ASAP7_75t_R FILLER_0_156_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_308 ();
 DECAPx1_ASAP7_75t_R FILLER_0_156_317 ();
 FILLER_ASAP7_75t_R FILLER_0_156_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_329 ();
 DECAPx6_ASAP7_75t_R FILLER_0_156_336 ();
 FILLER_ASAP7_75t_R FILLER_0_156_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_362 ();
 FILLER_ASAP7_75t_R FILLER_0_156_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_375 ();
 DECAPx2_ASAP7_75t_R FILLER_0_156_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_388 ();
 FILLER_ASAP7_75t_R FILLER_0_156_395 ();
 FILLER_ASAP7_75t_R FILLER_0_156_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_405 ();
 DECAPx2_ASAP7_75t_R FILLER_0_156_412 ();
 FILLER_ASAP7_75t_R FILLER_0_156_424 ();
 FILLER_ASAP7_75t_R FILLER_0_156_432 ();
 DECAPx4_ASAP7_75t_R FILLER_0_156_440 ();
 FILLER_ASAP7_75t_R FILLER_0_156_450 ();
 FILLER_ASAP7_75t_R FILLER_0_156_460 ();
 DECAPx10_ASAP7_75t_R FILLER_0_156_464 ();
 FILLER_ASAP7_75t_R FILLER_0_156_486 ();
 FILLER_ASAP7_75t_R FILLER_0_156_495 ();
 FILLER_ASAP7_75t_R FILLER_0_156_500 ();
 FILLER_ASAP7_75t_R FILLER_0_156_510 ();
 FILLER_ASAP7_75t_R FILLER_0_156_518 ();
 FILLER_ASAP7_75t_R FILLER_0_156_526 ();
 FILLER_ASAP7_75t_R FILLER_0_156_550 ();
 FILLER_ASAP7_75t_R FILLER_0_156_559 ();
 FILLER_ASAP7_75t_R FILLER_0_156_568 ();
 FILLER_ASAP7_75t_R FILLER_0_156_576 ();
 FILLER_ASAP7_75t_R FILLER_0_156_581 ();
 DECAPx6_ASAP7_75t_R FILLER_0_156_589 ();
 FILLER_ASAP7_75t_R FILLER_0_156_609 ();
 DECAPx2_ASAP7_75t_R FILLER_0_156_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_620 ();
 DECAPx6_ASAP7_75t_R FILLER_0_156_628 ();
 DECAPx1_ASAP7_75t_R FILLER_0_156_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_646 ();
 DECAPx4_ASAP7_75t_R FILLER_0_156_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_678 ();
 DECAPx2_ASAP7_75t_R FILLER_0_156_697 ();
 FILLER_ASAP7_75t_R FILLER_0_156_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_705 ();
 DECAPx2_ASAP7_75t_R FILLER_0_156_712 ();
 FILLER_ASAP7_75t_R FILLER_0_156_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_720 ();
 DECAPx4_ASAP7_75t_R FILLER_0_156_727 ();
 FILLER_ASAP7_75t_R FILLER_0_156_743 ();
 DECAPx10_ASAP7_75t_R FILLER_0_156_751 ();
 DECAPx2_ASAP7_75t_R FILLER_0_156_773 ();
 FILLER_ASAP7_75t_R FILLER_0_156_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_781 ();
 FILLER_ASAP7_75t_R FILLER_0_156_788 ();
 FILLER_ASAP7_75t_R FILLER_0_156_802 ();
 DECAPx10_ASAP7_75t_R FILLER_0_156_811 ();
 FILLER_ASAP7_75t_R FILLER_0_156_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_835 ();
 DECAPx4_ASAP7_75t_R FILLER_0_156_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_853 ();
 DECAPx2_ASAP7_75t_R FILLER_0_156_865 ();
 FILLER_ASAP7_75t_R FILLER_0_156_877 ();
 DECAPx2_ASAP7_75t_R FILLER_0_156_886 ();
 FILLER_ASAP7_75t_R FILLER_0_156_892 ();
 FILLER_ASAP7_75t_R FILLER_0_156_900 ();
 DECAPx10_ASAP7_75t_R FILLER_0_156_908 ();
 DECAPx1_ASAP7_75t_R FILLER_0_156_930 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_934 ();
 DECAPx10_ASAP7_75t_R FILLER_0_156_938 ();
 DECAPx2_ASAP7_75t_R FILLER_0_156_960 ();
 FILLER_ASAP7_75t_R FILLER_0_156_978 ();
 DECAPx4_ASAP7_75t_R FILLER_0_156_986 ();
 FILLER_ASAP7_75t_R FILLER_0_156_996 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_998 ();
 FILLER_ASAP7_75t_R FILLER_0_156_1002 ();
 FILLER_ASAP7_75t_R FILLER_0_156_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_1014 ();
 FILLER_ASAP7_75t_R FILLER_0_156_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_1023 ();
 FILLER_ASAP7_75t_R FILLER_0_156_1035 ();
 DECAPx10_ASAP7_75t_R FILLER_0_156_1043 ();
 DECAPx10_ASAP7_75t_R FILLER_0_156_1065 ();
 DECAPx2_ASAP7_75t_R FILLER_0_156_1087 ();
 FILLER_ASAP7_75t_R FILLER_0_156_1093 ();
 DECAPx1_ASAP7_75t_R FILLER_0_156_1107 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_1111 ();
 FILLER_ASAP7_75t_R FILLER_0_156_1124 ();
 FILLER_ASAP7_75t_R FILLER_0_156_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_156_1146 ();
 FILLER_ASAP7_75t_R FILLER_0_156_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_1170 ();
 DECAPx2_ASAP7_75t_R FILLER_0_156_1179 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_1185 ();
 FILLER_ASAP7_75t_R FILLER_0_156_1196 ();
 DECAPx6_ASAP7_75t_R FILLER_0_156_1206 ();
 FILLER_ASAP7_75t_R FILLER_0_156_1220 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_1222 ();
 DECAPx6_ASAP7_75t_R FILLER_0_156_1229 ();
 DECAPx2_ASAP7_75t_R FILLER_0_156_1243 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_1249 ();
 FILLER_ASAP7_75t_R FILLER_0_156_1256 ();
 FILLER_ASAP7_75t_R FILLER_0_156_1274 ();
 DECAPx4_ASAP7_75t_R FILLER_0_156_1282 ();
 FILLER_ASAP7_75t_R FILLER_0_156_1292 ();
 FILLER_ASAP7_75t_R FILLER_0_156_1304 ();
 FILLER_ASAP7_75t_R FILLER_0_156_1312 ();
 DECAPx2_ASAP7_75t_R FILLER_0_156_1324 ();
 FILLER_ASAP7_75t_R FILLER_0_156_1336 ();
 FILLER_ASAP7_75t_R FILLER_0_156_1341 ();
 FILLER_ASAP7_75t_R FILLER_0_156_1348 ();
 FILLER_ASAP7_75t_R FILLER_0_156_1355 ();
 DECAPx1_ASAP7_75t_R FILLER_0_156_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156_1367 ();
 FILLER_ASAP7_75t_R FILLER_0_156_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_156_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_157_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_4 ();
 FILLER_ASAP7_75t_R FILLER_0_157_8 ();
 DECAPx1_ASAP7_75t_R FILLER_0_157_16 ();
 FILLER_ASAP7_75t_R FILLER_0_157_42 ();
 DECAPx6_ASAP7_75t_R FILLER_0_157_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_61 ();
 DECAPx2_ASAP7_75t_R FILLER_0_157_74 ();
 DECAPx4_ASAP7_75t_R FILLER_0_157_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_111 ();
 DECAPx10_ASAP7_75t_R FILLER_0_157_118 ();
 DECAPx2_ASAP7_75t_R FILLER_0_157_140 ();
 FILLER_ASAP7_75t_R FILLER_0_157_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_148 ();
 DECAPx4_ASAP7_75t_R FILLER_0_157_160 ();
 FILLER_ASAP7_75t_R FILLER_0_157_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_172 ();
 FILLER_ASAP7_75t_R FILLER_0_157_181 ();
 DECAPx6_ASAP7_75t_R FILLER_0_157_191 ();
 DECAPx2_ASAP7_75t_R FILLER_0_157_205 ();
 FILLER_ASAP7_75t_R FILLER_0_157_214 ();
 DECAPx4_ASAP7_75t_R FILLER_0_157_224 ();
 DECAPx6_ASAP7_75t_R FILLER_0_157_245 ();
 DECAPx1_ASAP7_75t_R FILLER_0_157_259 ();
 DECAPx4_ASAP7_75t_R FILLER_0_157_269 ();
 DECAPx4_ASAP7_75t_R FILLER_0_157_285 ();
 FILLER_ASAP7_75t_R FILLER_0_157_295 ();
 FILLER_ASAP7_75t_R FILLER_0_157_303 ();
 DECAPx10_ASAP7_75t_R FILLER_0_157_311 ();
 DECAPx4_ASAP7_75t_R FILLER_0_157_333 ();
 FILLER_ASAP7_75t_R FILLER_0_157_353 ();
 FILLER_ASAP7_75t_R FILLER_0_157_365 ();
 DECAPx4_ASAP7_75t_R FILLER_0_157_377 ();
 DECAPx4_ASAP7_75t_R FILLER_0_157_393 ();
 FILLER_ASAP7_75t_R FILLER_0_157_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_405 ();
 DECAPx10_ASAP7_75t_R FILLER_0_157_412 ();
 DECAPx4_ASAP7_75t_R FILLER_0_157_440 ();
 DECAPx10_ASAP7_75t_R FILLER_0_157_456 ();
 DECAPx6_ASAP7_75t_R FILLER_0_157_478 ();
 FILLER_ASAP7_75t_R FILLER_0_157_492 ();
 FILLER_ASAP7_75t_R FILLER_0_157_500 ();
 DECAPx2_ASAP7_75t_R FILLER_0_157_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_516 ();
 DECAPx6_ASAP7_75t_R FILLER_0_157_525 ();
 DECAPx2_ASAP7_75t_R FILLER_0_157_539 ();
 DECAPx1_ASAP7_75t_R FILLER_0_157_551 ();
 FILLER_ASAP7_75t_R FILLER_0_157_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_563 ();
 FILLER_ASAP7_75t_R FILLER_0_157_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_574 ();
 DECAPx4_ASAP7_75t_R FILLER_0_157_583 ();
 FILLER_ASAP7_75t_R FILLER_0_157_593 ();
 FILLER_ASAP7_75t_R FILLER_0_157_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_609 ();
 FILLER_ASAP7_75t_R FILLER_0_157_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_619 ();
 FILLER_ASAP7_75t_R FILLER_0_157_627 ();
 FILLER_ASAP7_75t_R FILLER_0_157_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_637 ();
 DECAPx10_ASAP7_75t_R FILLER_0_157_641 ();
 FILLER_ASAP7_75t_R FILLER_0_157_666 ();
 DECAPx1_ASAP7_75t_R FILLER_0_157_680 ();
 FILLER_ASAP7_75t_R FILLER_0_157_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_704 ();
 FILLER_ASAP7_75t_R FILLER_0_157_711 ();
 DECAPx6_ASAP7_75t_R FILLER_0_157_719 ();
 DECAPx10_ASAP7_75t_R FILLER_0_157_739 ();
 DECAPx2_ASAP7_75t_R FILLER_0_157_761 ();
 DECAPx2_ASAP7_75t_R FILLER_0_157_775 ();
 FILLER_ASAP7_75t_R FILLER_0_157_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_783 ();
 DECAPx1_ASAP7_75t_R FILLER_0_157_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_795 ();
 DECAPx10_ASAP7_75t_R FILLER_0_157_802 ();
 DECAPx4_ASAP7_75t_R FILLER_0_157_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_834 ();
 DECAPx6_ASAP7_75t_R FILLER_0_157_841 ();
 FILLER_ASAP7_75t_R FILLER_0_157_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_857 ();
 DECAPx1_ASAP7_75t_R FILLER_0_157_864 ();
 DECAPx1_ASAP7_75t_R FILLER_0_157_876 ();
 DECAPx2_ASAP7_75t_R FILLER_0_157_887 ();
 FILLER_ASAP7_75t_R FILLER_0_157_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_902 ();
 FILLER_ASAP7_75t_R FILLER_0_157_923 ();
 DECAPx10_ASAP7_75t_R FILLER_0_157_927 ();
 FILLER_ASAP7_75t_R FILLER_0_157_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_951 ();
 DECAPx6_ASAP7_75t_R FILLER_0_157_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_976 ();
 DECAPx6_ASAP7_75t_R FILLER_0_157_989 ();
 FILLER_ASAP7_75t_R FILLER_0_157_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_1005 ();
 DECAPx10_ASAP7_75t_R FILLER_0_157_1014 ();
 DECAPx4_ASAP7_75t_R FILLER_0_157_1036 ();
 DECAPx1_ASAP7_75t_R FILLER_0_157_1050 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_1054 ();
 FILLER_ASAP7_75t_R FILLER_0_157_1063 ();
 DECAPx2_ASAP7_75t_R FILLER_0_157_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_1077 ();
 FILLER_ASAP7_75t_R FILLER_0_157_1090 ();
 DECAPx4_ASAP7_75t_R FILLER_0_157_1104 ();
 DECAPx2_ASAP7_75t_R FILLER_0_157_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_1132 ();
 FILLER_ASAP7_75t_R FILLER_0_157_1136 ();
 FILLER_ASAP7_75t_R FILLER_0_157_1146 ();
 DECAPx6_ASAP7_75t_R FILLER_0_157_1153 ();
 DECAPx1_ASAP7_75t_R FILLER_0_157_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_1171 ();
 FILLER_ASAP7_75t_R FILLER_0_157_1178 ();
 DECAPx6_ASAP7_75t_R FILLER_0_157_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_1204 ();
 DECAPx4_ASAP7_75t_R FILLER_0_157_1217 ();
 FILLER_ASAP7_75t_R FILLER_0_157_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_0_157_1246 ();
 DECAPx4_ASAP7_75t_R FILLER_0_157_1268 ();
 FILLER_ASAP7_75t_R FILLER_0_157_1278 ();
 FILLER_ASAP7_75t_R FILLER_0_157_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_1292 ();
 FILLER_ASAP7_75t_R FILLER_0_157_1296 ();
 FILLER_ASAP7_75t_R FILLER_0_157_1318 ();
 FILLER_ASAP7_75t_R FILLER_0_157_1326 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_1328 ();
 FILLER_ASAP7_75t_R FILLER_0_157_1335 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_1337 ();
 FILLER_ASAP7_75t_R FILLER_0_157_1360 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157_1362 ();
 FILLER_ASAP7_75t_R FILLER_0_157_1368 ();
 FILLER_ASAP7_75t_R FILLER_0_157_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_157_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_158_2 ();
 FILLER_ASAP7_75t_R FILLER_0_158_25 ();
 FILLER_ASAP7_75t_R FILLER_0_158_32 ();
 FILLER_ASAP7_75t_R FILLER_0_158_39 ();
 FILLER_ASAP7_75t_R FILLER_0_158_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_48 ();
 FILLER_ASAP7_75t_R FILLER_0_158_61 ();
 DECAPx4_ASAP7_75t_R FILLER_0_158_69 ();
 FILLER_ASAP7_75t_R FILLER_0_158_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_81 ();
 DECAPx2_ASAP7_75t_R FILLER_0_158_85 ();
 FILLER_ASAP7_75t_R FILLER_0_158_91 ();
 FILLER_ASAP7_75t_R FILLER_0_158_99 ();
 DECAPx1_ASAP7_75t_R FILLER_0_158_107 ();
 DECAPx4_ASAP7_75t_R FILLER_0_158_119 ();
 FILLER_ASAP7_75t_R FILLER_0_158_129 ();
 FILLER_ASAP7_75t_R FILLER_0_158_142 ();
 DECAPx6_ASAP7_75t_R FILLER_0_158_156 ();
 FILLER_ASAP7_75t_R FILLER_0_158_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_172 ();
 DECAPx2_ASAP7_75t_R FILLER_0_158_181 ();
 FILLER_ASAP7_75t_R FILLER_0_158_187 ();
 FILLER_ASAP7_75t_R FILLER_0_158_210 ();
 DECAPx6_ASAP7_75t_R FILLER_0_158_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_234 ();
 DECAPx4_ASAP7_75t_R FILLER_0_158_243 ();
 FILLER_ASAP7_75t_R FILLER_0_158_253 ();
 DECAPx2_ASAP7_75t_R FILLER_0_158_260 ();
 FILLER_ASAP7_75t_R FILLER_0_158_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_268 ();
 DECAPx1_ASAP7_75t_R FILLER_0_158_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_279 ();
 DECAPx1_ASAP7_75t_R FILLER_0_158_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_290 ();
 DECAPx4_ASAP7_75t_R FILLER_0_158_301 ();
 FILLER_ASAP7_75t_R FILLER_0_158_317 ();
 DECAPx4_ASAP7_75t_R FILLER_0_158_329 ();
 FILLER_ASAP7_75t_R FILLER_0_158_339 ();
 FILLER_ASAP7_75t_R FILLER_0_158_347 ();
 DECAPx1_ASAP7_75t_R FILLER_0_158_354 ();
 FILLER_ASAP7_75t_R FILLER_0_158_368 ();
 DECAPx2_ASAP7_75t_R FILLER_0_158_376 ();
 FILLER_ASAP7_75t_R FILLER_0_158_382 ();
 DECAPx4_ASAP7_75t_R FILLER_0_158_394 ();
 FILLER_ASAP7_75t_R FILLER_0_158_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_406 ();
 FILLER_ASAP7_75t_R FILLER_0_158_415 ();
 DECAPx2_ASAP7_75t_R FILLER_0_158_423 ();
 FILLER_ASAP7_75t_R FILLER_0_158_429 ();
 FILLER_ASAP7_75t_R FILLER_0_158_437 ();
 DECAPx6_ASAP7_75t_R FILLER_0_158_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_158_464 ();
 DECAPx2_ASAP7_75t_R FILLER_0_158_486 ();
 FILLER_ASAP7_75t_R FILLER_0_158_492 ();
 FILLER_ASAP7_75t_R FILLER_0_158_500 ();
 DECAPx2_ASAP7_75t_R FILLER_0_158_508 ();
 FILLER_ASAP7_75t_R FILLER_0_158_514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_158_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_528 ();
 FILLER_ASAP7_75t_R FILLER_0_158_535 ();
 DECAPx10_ASAP7_75t_R FILLER_0_158_543 ();
 DECAPx2_ASAP7_75t_R FILLER_0_158_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_571 ();
 FILLER_ASAP7_75t_R FILLER_0_158_578 ();
 FILLER_ASAP7_75t_R FILLER_0_158_586 ();
 DECAPx1_ASAP7_75t_R FILLER_0_158_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_600 ();
 DECAPx4_ASAP7_75t_R FILLER_0_158_607 ();
 FILLER_ASAP7_75t_R FILLER_0_158_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_625 ();
 FILLER_ASAP7_75t_R FILLER_0_158_634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_158_642 ();
 DECAPx1_ASAP7_75t_R FILLER_0_158_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_668 ();
 FILLER_ASAP7_75t_R FILLER_0_158_707 ();
 DECAPx2_ASAP7_75t_R FILLER_0_158_720 ();
 FILLER_ASAP7_75t_R FILLER_0_158_731 ();
 FILLER_ASAP7_75t_R FILLER_0_158_739 ();
 DECAPx2_ASAP7_75t_R FILLER_0_158_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_759 ();
 FILLER_ASAP7_75t_R FILLER_0_158_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_772 ();
 FILLER_ASAP7_75t_R FILLER_0_158_783 ();
 FILLER_ASAP7_75t_R FILLER_0_158_795 ();
 DECAPx2_ASAP7_75t_R FILLER_0_158_803 ();
 FILLER_ASAP7_75t_R FILLER_0_158_809 ();
 DECAPx1_ASAP7_75t_R FILLER_0_158_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_827 ();
 DECAPx6_ASAP7_75t_R FILLER_0_158_834 ();
 DECAPx1_ASAP7_75t_R FILLER_0_158_854 ();
 DECAPx4_ASAP7_75t_R FILLER_0_158_864 ();
 FILLER_ASAP7_75t_R FILLER_0_158_874 ();
 DECAPx4_ASAP7_75t_R FILLER_0_158_887 ();
 FILLER_ASAP7_75t_R FILLER_0_158_897 ();
 DECAPx4_ASAP7_75t_R FILLER_0_158_905 ();
 DECAPx6_ASAP7_75t_R FILLER_0_158_921 ();
 FILLER_ASAP7_75t_R FILLER_0_158_935 ();
 FILLER_ASAP7_75t_R FILLER_0_158_947 ();
 FILLER_ASAP7_75t_R FILLER_0_158_959 ();
 DECAPx2_ASAP7_75t_R FILLER_0_158_966 ();
 FILLER_ASAP7_75t_R FILLER_0_158_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_974 ();
 FILLER_ASAP7_75t_R FILLER_0_158_987 ();
 DECAPx2_ASAP7_75t_R FILLER_0_158_995 ();
 FILLER_ASAP7_75t_R FILLER_0_158_1001 ();
 FILLER_ASAP7_75t_R FILLER_0_158_1011 ();
 DECAPx2_ASAP7_75t_R FILLER_0_158_1024 ();
 FILLER_ASAP7_75t_R FILLER_0_158_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_1032 ();
 DECAPx4_ASAP7_75t_R FILLER_0_158_1043 ();
 FILLER_ASAP7_75t_R FILLER_0_158_1059 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_1061 ();
 DECAPx1_ASAP7_75t_R FILLER_0_158_1070 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_1074 ();
 DECAPx1_ASAP7_75t_R FILLER_0_158_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_0_158_1097 ();
 DECAPx2_ASAP7_75t_R FILLER_0_158_1119 ();
 FILLER_ASAP7_75t_R FILLER_0_158_1125 ();
 FILLER_ASAP7_75t_R FILLER_0_158_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_1137 ();
 FILLER_ASAP7_75t_R FILLER_0_158_1146 ();
 DECAPx6_ASAP7_75t_R FILLER_0_158_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_1168 ();
 DECAPx1_ASAP7_75t_R FILLER_0_158_1175 ();
 FILLER_ASAP7_75t_R FILLER_0_158_1185 ();
 FILLER_ASAP7_75t_R FILLER_0_158_1193 ();
 FILLER_ASAP7_75t_R FILLER_0_158_1215 ();
 DECAPx1_ASAP7_75t_R FILLER_0_158_1225 ();
 DECAPx2_ASAP7_75t_R FILLER_0_158_1235 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_1241 ();
 DECAPx6_ASAP7_75t_R FILLER_0_158_1248 ();
 DECAPx1_ASAP7_75t_R FILLER_0_158_1262 ();
 FILLER_ASAP7_75t_R FILLER_0_158_1272 ();
 DECAPx2_ASAP7_75t_R FILLER_0_158_1280 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_1286 ();
 FILLER_ASAP7_75t_R FILLER_0_158_1294 ();
 DECAPx1_ASAP7_75t_R FILLER_0_158_1306 ();
 FILLER_ASAP7_75t_R FILLER_0_158_1316 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_1318 ();
 FILLER_ASAP7_75t_R FILLER_0_158_1324 ();
 DECAPx1_ASAP7_75t_R FILLER_0_158_1337 ();
 FILLER_ASAP7_75t_R FILLER_0_158_1346 ();
 DECAPx1_ASAP7_75t_R FILLER_0_158_1354 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158_1358 ();
 FILLER_ASAP7_75t_R FILLER_0_158_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_159_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_4 ();
 FILLER_ASAP7_75t_R FILLER_0_159_8 ();
 FILLER_ASAP7_75t_R FILLER_0_159_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_17 ();
 FILLER_ASAP7_75t_R FILLER_0_159_21 ();
 DECAPx1_ASAP7_75t_R FILLER_0_159_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_32 ();
 FILLER_ASAP7_75t_R FILLER_0_159_55 ();
 FILLER_ASAP7_75t_R FILLER_0_159_63 ();
 DECAPx6_ASAP7_75t_R FILLER_0_159_68 ();
 DECAPx1_ASAP7_75t_R FILLER_0_159_82 ();
 FILLER_ASAP7_75t_R FILLER_0_159_92 ();
 DECAPx2_ASAP7_75t_R FILLER_0_159_102 ();
 FILLER_ASAP7_75t_R FILLER_0_159_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_110 ();
 FILLER_ASAP7_75t_R FILLER_0_159_117 ();
 FILLER_ASAP7_75t_R FILLER_0_159_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_127 ();
 DECAPx4_ASAP7_75t_R FILLER_0_159_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_149 ();
 FILLER_ASAP7_75t_R FILLER_0_159_160 ();
 DECAPx2_ASAP7_75t_R FILLER_0_159_167 ();
 DECAPx4_ASAP7_75t_R FILLER_0_159_181 ();
 DECAPx6_ASAP7_75t_R FILLER_0_159_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_208 ();
 FILLER_ASAP7_75t_R FILLER_0_159_219 ();
 DECAPx1_ASAP7_75t_R FILLER_0_159_227 ();
 FILLER_ASAP7_75t_R FILLER_0_159_237 ();
 DECAPx6_ASAP7_75t_R FILLER_0_159_247 ();
 FILLER_ASAP7_75t_R FILLER_0_159_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_263 ();
 DECAPx1_ASAP7_75t_R FILLER_0_159_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_274 ();
 FILLER_ASAP7_75t_R FILLER_0_159_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_285 ();
 DECAPx1_ASAP7_75t_R FILLER_0_159_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_296 ();
 DECAPx2_ASAP7_75t_R FILLER_0_159_303 ();
 FILLER_ASAP7_75t_R FILLER_0_159_309 ();
 DECAPx2_ASAP7_75t_R FILLER_0_159_317 ();
 FILLER_ASAP7_75t_R FILLER_0_159_323 ();
 DECAPx2_ASAP7_75t_R FILLER_0_159_331 ();
 DECAPx1_ASAP7_75t_R FILLER_0_159_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_349 ();
 DECAPx4_ASAP7_75t_R FILLER_0_159_356 ();
 DECAPx2_ASAP7_75t_R FILLER_0_159_376 ();
 FILLER_ASAP7_75t_R FILLER_0_159_382 ();
 FILLER_ASAP7_75t_R FILLER_0_159_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_396 ();
 FILLER_ASAP7_75t_R FILLER_0_159_403 ();
 DECAPx2_ASAP7_75t_R FILLER_0_159_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_417 ();
 FILLER_ASAP7_75t_R FILLER_0_159_424 ();
 DECAPx1_ASAP7_75t_R FILLER_0_159_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_436 ();
 DECAPx2_ASAP7_75t_R FILLER_0_159_443 ();
 DECAPx2_ASAP7_75t_R FILLER_0_159_455 ();
 FILLER_ASAP7_75t_R FILLER_0_159_461 ();
 DECAPx2_ASAP7_75t_R FILLER_0_159_485 ();
 FILLER_ASAP7_75t_R FILLER_0_159_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_493 ();
 FILLER_ASAP7_75t_R FILLER_0_159_500 ();
 DECAPx4_ASAP7_75t_R FILLER_0_159_508 ();
 DECAPx4_ASAP7_75t_R FILLER_0_159_525 ();
 FILLER_ASAP7_75t_R FILLER_0_159_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_537 ();
 FILLER_ASAP7_75t_R FILLER_0_159_544 ();
 DECAPx2_ASAP7_75t_R FILLER_0_159_552 ();
 DECAPx6_ASAP7_75t_R FILLER_0_159_568 ();
 DECAPx1_ASAP7_75t_R FILLER_0_159_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_586 ();
 DECAPx6_ASAP7_75t_R FILLER_0_159_593 ();
 DECAPx1_ASAP7_75t_R FILLER_0_159_607 ();
 FILLER_ASAP7_75t_R FILLER_0_159_617 ();
 FILLER_ASAP7_75t_R FILLER_0_159_625 ();
 DECAPx6_ASAP7_75t_R FILLER_0_159_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_647 ();
 FILLER_ASAP7_75t_R FILLER_0_159_670 ();
 FILLER_ASAP7_75t_R FILLER_0_159_677 ();
 FILLER_ASAP7_75t_R FILLER_0_159_689 ();
 DECAPx2_ASAP7_75t_R FILLER_0_159_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_713 ();
 DECAPx2_ASAP7_75t_R FILLER_0_159_720 ();
 FILLER_ASAP7_75t_R FILLER_0_159_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_734 ();
 DECAPx4_ASAP7_75t_R FILLER_0_159_745 ();
 FILLER_ASAP7_75t_R FILLER_0_159_755 ();
 FILLER_ASAP7_75t_R FILLER_0_159_763 ();
 DECAPx2_ASAP7_75t_R FILLER_0_159_771 ();
 FILLER_ASAP7_75t_R FILLER_0_159_783 ();
 FILLER_ASAP7_75t_R FILLER_0_159_791 ();
 FILLER_ASAP7_75t_R FILLER_0_159_803 ();
 FILLER_ASAP7_75t_R FILLER_0_159_817 ();
 FILLER_ASAP7_75t_R FILLER_0_159_825 ();
 DECAPx6_ASAP7_75t_R FILLER_0_159_838 ();
 DECAPx1_ASAP7_75t_R FILLER_0_159_852 ();
 FILLER_ASAP7_75t_R FILLER_0_159_862 ();
 DECAPx6_ASAP7_75t_R FILLER_0_159_874 ();
 FILLER_ASAP7_75t_R FILLER_0_159_888 ();
 DECAPx10_ASAP7_75t_R FILLER_0_159_896 ();
 FILLER_ASAP7_75t_R FILLER_0_159_918 ();
 FILLER_ASAP7_75t_R FILLER_0_159_923 ();
 FILLER_ASAP7_75t_R FILLER_0_159_927 ();
 FILLER_ASAP7_75t_R FILLER_0_159_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_941 ();
 DECAPx1_ASAP7_75t_R FILLER_0_159_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_952 ();
 DECAPx4_ASAP7_75t_R FILLER_0_159_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_966 ();
 FILLER_ASAP7_75t_R FILLER_0_159_972 ();
 FILLER_ASAP7_75t_R FILLER_0_159_986 ();
 DECAPx1_ASAP7_75t_R FILLER_0_159_1000 ();
 DECAPx1_ASAP7_75t_R FILLER_0_159_1010 ();
 DECAPx4_ASAP7_75t_R FILLER_0_159_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_1032 ();
 FILLER_ASAP7_75t_R FILLER_0_159_1041 ();
 FILLER_ASAP7_75t_R FILLER_0_159_1053 ();
 DECAPx2_ASAP7_75t_R FILLER_0_159_1061 ();
 FILLER_ASAP7_75t_R FILLER_0_159_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_1069 ();
 FILLER_ASAP7_75t_R FILLER_0_159_1078 ();
 DECAPx10_ASAP7_75t_R FILLER_0_159_1086 ();
 DECAPx2_ASAP7_75t_R FILLER_0_159_1108 ();
 FILLER_ASAP7_75t_R FILLER_0_159_1126 ();
 DECAPx4_ASAP7_75t_R FILLER_0_159_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_1144 ();
 DECAPx6_ASAP7_75t_R FILLER_0_159_1151 ();
 DECAPx1_ASAP7_75t_R FILLER_0_159_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_1169 ();
 DECAPx1_ASAP7_75t_R FILLER_0_159_1176 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_1180 ();
 FILLER_ASAP7_75t_R FILLER_0_159_1187 ();
 FILLER_ASAP7_75t_R FILLER_0_159_1196 ();
 FILLER_ASAP7_75t_R FILLER_0_159_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_1210 ();
 FILLER_ASAP7_75t_R FILLER_0_159_1217 ();
 DECAPx1_ASAP7_75t_R FILLER_0_159_1230 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_1234 ();
 FILLER_ASAP7_75t_R FILLER_0_159_1241 ();
 DECAPx2_ASAP7_75t_R FILLER_0_159_1249 ();
 FILLER_ASAP7_75t_R FILLER_0_159_1255 ();
 FILLER_ASAP7_75t_R FILLER_0_159_1263 ();
 FILLER_ASAP7_75t_R FILLER_0_159_1271 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_1273 ();
 FILLER_ASAP7_75t_R FILLER_0_159_1280 ();
 DECAPx2_ASAP7_75t_R FILLER_0_159_1288 ();
 FILLER_ASAP7_75t_R FILLER_0_159_1294 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_1296 ();
 FILLER_ASAP7_75t_R FILLER_0_159_1317 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159_1319 ();
 FILLER_ASAP7_75t_R FILLER_0_159_1323 ();
 DECAPx2_ASAP7_75t_R FILLER_0_159_1331 ();
 FILLER_ASAP7_75t_R FILLER_0_159_1358 ();
 FILLER_ASAP7_75t_R FILLER_0_159_1366 ();
 FILLER_ASAP7_75t_R FILLER_0_159_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_159_1380 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_13 ();
 FILLER_ASAP7_75t_R FILLER_0_160_41 ();
 FILLER_ASAP7_75t_R FILLER_0_160_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_55 ();
 FILLER_ASAP7_75t_R FILLER_0_160_69 ();
 FILLER_ASAP7_75t_R FILLER_0_160_74 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_88 ();
 FILLER_ASAP7_75t_R FILLER_0_160_100 ();
 DECAPx4_ASAP7_75t_R FILLER_0_160_107 ();
 FILLER_ASAP7_75t_R FILLER_0_160_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_119 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_138 ();
 DECAPx4_ASAP7_75t_R FILLER_0_160_143 ();
 FILLER_ASAP7_75t_R FILLER_0_160_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_167 ();
 FILLER_ASAP7_75t_R FILLER_0_160_174 ();
 FILLER_ASAP7_75t_R FILLER_0_160_184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_160_192 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_222 ();
 FILLER_ASAP7_75t_R FILLER_0_160_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_230 ();
 FILLER_ASAP7_75t_R FILLER_0_160_234 ();
 FILLER_ASAP7_75t_R FILLER_0_160_244 ();
 DECAPx4_ASAP7_75t_R FILLER_0_160_252 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_268 ();
 FILLER_ASAP7_75t_R FILLER_0_160_274 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_282 ();
 FILLER_ASAP7_75t_R FILLER_0_160_295 ();
 FILLER_ASAP7_75t_R FILLER_0_160_303 ();
 DECAPx1_ASAP7_75t_R FILLER_0_160_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_314 ();
 DECAPx6_ASAP7_75t_R FILLER_0_160_321 ();
 DECAPx1_ASAP7_75t_R FILLER_0_160_335 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_345 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_359 ();
 FILLER_ASAP7_75t_R FILLER_0_160_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_367 ();
 DECAPx4_ASAP7_75t_R FILLER_0_160_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_384 ();
 FILLER_ASAP7_75t_R FILLER_0_160_391 ();
 FILLER_ASAP7_75t_R FILLER_0_160_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_401 ();
 FILLER_ASAP7_75t_R FILLER_0_160_408 ();
 FILLER_ASAP7_75t_R FILLER_0_160_416 ();
 FILLER_ASAP7_75t_R FILLER_0_160_424 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_434 ();
 DECAPx6_ASAP7_75t_R FILLER_0_160_448 ();
 FILLER_ASAP7_75t_R FILLER_0_160_464 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_469 ();
 FILLER_ASAP7_75t_R FILLER_0_160_475 ();
 FILLER_ASAP7_75t_R FILLER_0_160_482 ();
 FILLER_ASAP7_75t_R FILLER_0_160_502 ();
 DECAPx1_ASAP7_75t_R FILLER_0_160_511 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_521 ();
 FILLER_ASAP7_75t_R FILLER_0_160_527 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_535 ();
 DECAPx4_ASAP7_75t_R FILLER_0_160_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_571 ();
 DECAPx6_ASAP7_75t_R FILLER_0_160_575 ();
 FILLER_ASAP7_75t_R FILLER_0_160_589 ();
 DECAPx10_ASAP7_75t_R FILLER_0_160_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_616 ();
 DECAPx4_ASAP7_75t_R FILLER_0_160_625 ();
 FILLER_ASAP7_75t_R FILLER_0_160_642 ();
 FILLER_ASAP7_75t_R FILLER_0_160_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_649 ();
 FILLER_ASAP7_75t_R FILLER_0_160_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_655 ();
 FILLER_ASAP7_75t_R FILLER_0_160_662 ();
 FILLER_ASAP7_75t_R FILLER_0_160_667 ();
 DECAPx1_ASAP7_75t_R FILLER_0_160_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_683 ();
 FILLER_ASAP7_75t_R FILLER_0_160_692 ();
 DECAPx4_ASAP7_75t_R FILLER_0_160_699 ();
 FILLER_ASAP7_75t_R FILLER_0_160_709 ();
 DECAPx1_ASAP7_75t_R FILLER_0_160_717 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_727 ();
 FILLER_ASAP7_75t_R FILLER_0_160_739 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_753 ();
 FILLER_ASAP7_75t_R FILLER_0_160_762 ();
 DECAPx6_ASAP7_75t_R FILLER_0_160_770 ();
 DECAPx1_ASAP7_75t_R FILLER_0_160_784 ();
 FILLER_ASAP7_75t_R FILLER_0_160_794 ();
 FILLER_ASAP7_75t_R FILLER_0_160_806 ();
 FILLER_ASAP7_75t_R FILLER_0_160_814 ();
 FILLER_ASAP7_75t_R FILLER_0_160_822 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_830 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_848 ();
 FILLER_ASAP7_75t_R FILLER_0_160_855 ();
 FILLER_ASAP7_75t_R FILLER_0_160_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_865 ();
 DECAPx4_ASAP7_75t_R FILLER_0_160_873 ();
 FILLER_ASAP7_75t_R FILLER_0_160_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_885 ();
 FILLER_ASAP7_75t_R FILLER_0_160_892 ();
 DECAPx4_ASAP7_75t_R FILLER_0_160_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_910 ();
 DECAPx1_ASAP7_75t_R FILLER_0_160_921 ();
 FILLER_ASAP7_75t_R FILLER_0_160_930 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_948 ();
 FILLER_ASAP7_75t_R FILLER_0_160_957 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_970 ();
 FILLER_ASAP7_75t_R FILLER_0_160_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_978 ();
 DECAPx1_ASAP7_75t_R FILLER_0_160_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_993 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_999 ();
 FILLER_ASAP7_75t_R FILLER_0_160_1005 ();
 DECAPx1_ASAP7_75t_R FILLER_0_160_1013 ();
 FILLER_ASAP7_75t_R FILLER_0_160_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_1025 ();
 FILLER_ASAP7_75t_R FILLER_0_160_1032 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_1044 ();
 FILLER_ASAP7_75t_R FILLER_0_160_1050 ();
 FILLER_ASAP7_75t_R FILLER_0_160_1058 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_1072 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_1083 ();
 FILLER_ASAP7_75t_R FILLER_0_160_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_1091 ();
 FILLER_ASAP7_75t_R FILLER_0_160_1104 ();
 FILLER_ASAP7_75t_R FILLER_0_160_1118 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_1126 ();
 FILLER_ASAP7_75t_R FILLER_0_160_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_0_160_1140 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_1162 ();
 FILLER_ASAP7_75t_R FILLER_0_160_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_1170 ();
 DECAPx6_ASAP7_75t_R FILLER_0_160_1177 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_1197 ();
 FILLER_ASAP7_75t_R FILLER_0_160_1204 ();
 DECAPx1_ASAP7_75t_R FILLER_0_160_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_1216 ();
 FILLER_ASAP7_75t_R FILLER_0_160_1223 ();
 DECAPx4_ASAP7_75t_R FILLER_0_160_1231 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_1247 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_1253 ();
 DECAPx1_ASAP7_75t_R FILLER_0_160_1260 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_1270 ();
 FILLER_ASAP7_75t_R FILLER_0_160_1276 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_1278 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_1288 ();
 FILLER_ASAP7_75t_R FILLER_0_160_1295 ();
 FILLER_ASAP7_75t_R FILLER_0_160_1303 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_1305 ();
 FILLER_ASAP7_75t_R FILLER_0_160_1309 ();
 FILLER_ASAP7_75t_R FILLER_0_160_1316 ();
 DECAPx1_ASAP7_75t_R FILLER_0_160_1324 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160_1328 ();
 FILLER_ASAP7_75t_R FILLER_0_160_1335 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_1342 ();
 FILLER_ASAP7_75t_R FILLER_0_160_1354 ();
 FILLER_ASAP7_75t_R FILLER_0_160_1361 ();
 FILLER_ASAP7_75t_R FILLER_0_160_1369 ();
 DECAPx2_ASAP7_75t_R FILLER_0_160_1376 ();
 FILLER_ASAP7_75t_R FILLER_0_161_2 ();
 FILLER_ASAP7_75t_R FILLER_0_161_9 ();
 FILLER_ASAP7_75t_R FILLER_0_161_16 ();
 FILLER_ASAP7_75t_R FILLER_0_161_28 ();
 FILLER_ASAP7_75t_R FILLER_0_161_35 ();
 DECAPx2_ASAP7_75t_R FILLER_0_161_59 ();
 FILLER_ASAP7_75t_R FILLER_0_161_73 ();
 FILLER_ASAP7_75t_R FILLER_0_161_81 ();
 DECAPx1_ASAP7_75t_R FILLER_0_161_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161_90 ();
 FILLER_ASAP7_75t_R FILLER_0_161_101 ();
 FILLER_ASAP7_75t_R FILLER_0_161_109 ();
 FILLER_ASAP7_75t_R FILLER_0_161_121 ();
 DECAPx2_ASAP7_75t_R FILLER_0_161_128 ();
 FILLER_ASAP7_75t_R FILLER_0_161_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161_136 ();
 DECAPx4_ASAP7_75t_R FILLER_0_161_147 ();
 DECAPx2_ASAP7_75t_R FILLER_0_161_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161_173 ();
 DECAPx2_ASAP7_75t_R FILLER_0_161_180 ();
 FILLER_ASAP7_75t_R FILLER_0_161_186 ();
 DECAPx4_ASAP7_75t_R FILLER_0_161_196 ();
 FILLER_ASAP7_75t_R FILLER_0_161_206 ();
 FILLER_ASAP7_75t_R FILLER_0_161_211 ();
 DECAPx2_ASAP7_75t_R FILLER_0_161_224 ();
 FILLER_ASAP7_75t_R FILLER_0_161_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161_232 ();
 DECAPx1_ASAP7_75t_R FILLER_0_161_243 ();
 DECAPx2_ASAP7_75t_R FILLER_0_161_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161_263 ();
 DECAPx6_ASAP7_75t_R FILLER_0_161_271 ();
 FILLER_ASAP7_75t_R FILLER_0_161_285 ();
 FILLER_ASAP7_75t_R FILLER_0_161_293 ();
 DECAPx6_ASAP7_75t_R FILLER_0_161_301 ();
 FILLER_ASAP7_75t_R FILLER_0_161_315 ();
 DECAPx6_ASAP7_75t_R FILLER_0_161_323 ();
 DECAPx1_ASAP7_75t_R FILLER_0_161_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161_341 ();
 FILLER_ASAP7_75t_R FILLER_0_161_348 ();
 DECAPx4_ASAP7_75t_R FILLER_0_161_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161_366 ();
 DECAPx4_ASAP7_75t_R FILLER_0_161_373 ();
 FILLER_ASAP7_75t_R FILLER_0_161_383 ();
 DECAPx4_ASAP7_75t_R FILLER_0_161_407 ();
 DECAPx1_ASAP7_75t_R FILLER_0_161_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161_431 ();
 FILLER_ASAP7_75t_R FILLER_0_161_438 ();
 DECAPx10_ASAP7_75t_R FILLER_0_161_446 ();
 DECAPx6_ASAP7_75t_R FILLER_0_161_468 ();
 FILLER_ASAP7_75t_R FILLER_0_161_482 ();
 FILLER_ASAP7_75t_R FILLER_0_161_498 ();
 DECAPx2_ASAP7_75t_R FILLER_0_161_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161_512 ();
 DECAPx2_ASAP7_75t_R FILLER_0_161_519 ();
 FILLER_ASAP7_75t_R FILLER_0_161_525 ();
 DECAPx1_ASAP7_75t_R FILLER_0_161_533 ();
 DECAPx1_ASAP7_75t_R FILLER_0_161_543 ();
 DECAPx1_ASAP7_75t_R FILLER_0_161_553 ();
 FILLER_ASAP7_75t_R FILLER_0_161_564 ();
 FILLER_ASAP7_75t_R FILLER_0_161_573 ();
 DECAPx1_ASAP7_75t_R FILLER_0_161_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161_585 ();
 DECAPx2_ASAP7_75t_R FILLER_0_161_594 ();
 FILLER_ASAP7_75t_R FILLER_0_161_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161_602 ();
 FILLER_ASAP7_75t_R FILLER_0_161_611 ();
 FILLER_ASAP7_75t_R FILLER_0_161_619 ();
 FILLER_ASAP7_75t_R FILLER_0_161_627 ();
 FILLER_ASAP7_75t_R FILLER_0_161_649 ();
 FILLER_ASAP7_75t_R FILLER_0_161_654 ();
 FILLER_ASAP7_75t_R FILLER_0_161_662 ();
 FILLER_ASAP7_75t_R FILLER_0_161_670 ();
 DECAPx6_ASAP7_75t_R FILLER_0_161_675 ();
 FILLER_ASAP7_75t_R FILLER_0_161_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161_691 ();
 DECAPx1_ASAP7_75t_R FILLER_0_161_698 ();
 DECAPx2_ASAP7_75t_R FILLER_0_161_712 ();
 FILLER_ASAP7_75t_R FILLER_0_161_718 ();
 FILLER_ASAP7_75t_R FILLER_0_161_726 ();
 DECAPx10_ASAP7_75t_R FILLER_0_161_733 ();
 FILLER_ASAP7_75t_R FILLER_0_161_755 ();
 DECAPx1_ASAP7_75t_R FILLER_0_161_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161_764 ();
 DECAPx2_ASAP7_75t_R FILLER_0_161_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161_777 ();
 FILLER_ASAP7_75t_R FILLER_0_161_784 ();
 DECAPx6_ASAP7_75t_R FILLER_0_161_796 ();
 FILLER_ASAP7_75t_R FILLER_0_161_810 ();
 DECAPx1_ASAP7_75t_R FILLER_0_161_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161_822 ();
 FILLER_ASAP7_75t_R FILLER_0_161_833 ();
 DECAPx10_ASAP7_75t_R FILLER_0_161_838 ();
 DECAPx6_ASAP7_75t_R FILLER_0_161_860 ();
 DECAPx2_ASAP7_75t_R FILLER_0_161_874 ();
 DECAPx4_ASAP7_75t_R FILLER_0_161_891 ();
 FILLER_ASAP7_75t_R FILLER_0_161_901 ();
 FILLER_ASAP7_75t_R FILLER_0_161_923 ();
 DECAPx2_ASAP7_75t_R FILLER_0_161_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161_933 ();
 DECAPx6_ASAP7_75t_R FILLER_0_161_942 ();
 DECAPx1_ASAP7_75t_R FILLER_0_161_956 ();
 DECAPx2_ASAP7_75t_R FILLER_0_161_966 ();
 FILLER_ASAP7_75t_R FILLER_0_161_972 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161_974 ();
 FILLER_ASAP7_75t_R FILLER_0_161_981 ();
 FILLER_ASAP7_75t_R FILLER_0_161_989 ();
 DECAPx1_ASAP7_75t_R FILLER_0_161_1002 ();
 DECAPx10_ASAP7_75t_R FILLER_0_161_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161_1039 ();
 DECAPx4_ASAP7_75t_R FILLER_0_161_1046 ();
 DECAPx1_ASAP7_75t_R FILLER_0_161_1068 ();
 DECAPx1_ASAP7_75t_R FILLER_0_161_1080 ();
 DECAPx4_ASAP7_75t_R FILLER_0_161_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161_1105 ();
 FILLER_ASAP7_75t_R FILLER_0_161_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161_1120 ();
 DECAPx2_ASAP7_75t_R FILLER_0_161_1127 ();
 FILLER_ASAP7_75t_R FILLER_0_161_1141 ();
 DECAPx6_ASAP7_75t_R FILLER_0_161_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161_1169 ();
 FILLER_ASAP7_75t_R FILLER_0_161_1176 ();
 DECAPx6_ASAP7_75t_R FILLER_0_161_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161_1198 ();
 DECAPx10_ASAP7_75t_R FILLER_0_161_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161_1231 ();
 FILLER_ASAP7_75t_R FILLER_0_161_1238 ();
 FILLER_ASAP7_75t_R FILLER_0_161_1246 ();
 DECAPx4_ASAP7_75t_R FILLER_0_161_1253 ();
 FILLER_ASAP7_75t_R FILLER_0_161_1270 ();
 FILLER_ASAP7_75t_R FILLER_0_161_1278 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161_1280 ();
 FILLER_ASAP7_75t_R FILLER_0_161_1293 ();
 DECAPx2_ASAP7_75t_R FILLER_0_161_1303 ();
 DECAPx1_ASAP7_75t_R FILLER_0_161_1315 ();
 FILLER_ASAP7_75t_R FILLER_0_161_1322 ();
 FILLER_ASAP7_75t_R FILLER_0_161_1329 ();
 FILLER_ASAP7_75t_R FILLER_0_161_1353 ();
 DECAPx2_ASAP7_75t_R FILLER_0_161_1376 ();
 DECAPx1_ASAP7_75t_R FILLER_0_162_2 ();
 FILLER_ASAP7_75t_R FILLER_0_162_11 ();
 FILLER_ASAP7_75t_R FILLER_0_162_19 ();
 FILLER_ASAP7_75t_R FILLER_0_162_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_28 ();
 FILLER_ASAP7_75t_R FILLER_0_162_35 ();
 FILLER_ASAP7_75t_R FILLER_0_162_42 ();
 FILLER_ASAP7_75t_R FILLER_0_162_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_49 ();
 FILLER_ASAP7_75t_R FILLER_0_162_55 ();
 FILLER_ASAP7_75t_R FILLER_0_162_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_62 ();
 FILLER_ASAP7_75t_R FILLER_0_162_69 ();
 FILLER_ASAP7_75t_R FILLER_0_162_79 ();
 FILLER_ASAP7_75t_R FILLER_0_162_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_88 ();
 FILLER_ASAP7_75t_R FILLER_0_162_97 ();
 FILLER_ASAP7_75t_R FILLER_0_162_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_111 ();
 FILLER_ASAP7_75t_R FILLER_0_162_122 ();
 FILLER_ASAP7_75t_R FILLER_0_162_134 ();
 FILLER_ASAP7_75t_R FILLER_0_162_146 ();
 DECAPx1_ASAP7_75t_R FILLER_0_162_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_158 ();
 DECAPx6_ASAP7_75t_R FILLER_0_162_169 ();
 FILLER_ASAP7_75t_R FILLER_0_162_195 ();
 DECAPx10_ASAP7_75t_R FILLER_0_162_218 ();
 DECAPx4_ASAP7_75t_R FILLER_0_162_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_270 ();
 FILLER_ASAP7_75t_R FILLER_0_162_295 ();
 FILLER_ASAP7_75t_R FILLER_0_162_304 ();
 DECAPx1_ASAP7_75t_R FILLER_0_162_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_316 ();
 DECAPx2_ASAP7_75t_R FILLER_0_162_325 ();
 FILLER_ASAP7_75t_R FILLER_0_162_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_333 ();
 FILLER_ASAP7_75t_R FILLER_0_162_340 ();
 DECAPx10_ASAP7_75t_R FILLER_0_162_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_370 ();
 FILLER_ASAP7_75t_R FILLER_0_162_391 ();
 DECAPx6_ASAP7_75t_R FILLER_0_162_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_413 ();
 DECAPx4_ASAP7_75t_R FILLER_0_162_417 ();
 FILLER_ASAP7_75t_R FILLER_0_162_433 ();
 DECAPx6_ASAP7_75t_R FILLER_0_162_441 ();
 DECAPx2_ASAP7_75t_R FILLER_0_162_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_461 ();
 DECAPx4_ASAP7_75t_R FILLER_0_162_464 ();
 FILLER_ASAP7_75t_R FILLER_0_162_482 ();
 FILLER_ASAP7_75t_R FILLER_0_162_487 ();
 DECAPx2_ASAP7_75t_R FILLER_0_162_495 ();
 FILLER_ASAP7_75t_R FILLER_0_162_501 ();
 FILLER_ASAP7_75t_R FILLER_0_162_514 ();
 FILLER_ASAP7_75t_R FILLER_0_162_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_524 ();
 FILLER_ASAP7_75t_R FILLER_0_162_530 ();
 FILLER_ASAP7_75t_R FILLER_0_162_540 ();
 FILLER_ASAP7_75t_R FILLER_0_162_548 ();
 FILLER_ASAP7_75t_R FILLER_0_162_553 ();
 DECAPx1_ASAP7_75t_R FILLER_0_162_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_565 ();
 FILLER_ASAP7_75t_R FILLER_0_162_572 ();
 DECAPx1_ASAP7_75t_R FILLER_0_162_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_584 ();
 DECAPx2_ASAP7_75t_R FILLER_0_162_591 ();
 FILLER_ASAP7_75t_R FILLER_0_162_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_605 ();
 FILLER_ASAP7_75t_R FILLER_0_162_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_616 ();
 FILLER_ASAP7_75t_R FILLER_0_162_623 ();
 DECAPx2_ASAP7_75t_R FILLER_0_162_628 ();
 DECAPx1_ASAP7_75t_R FILLER_0_162_637 ();
 DECAPx10_ASAP7_75t_R FILLER_0_162_647 ();
 DECAPx6_ASAP7_75t_R FILLER_0_162_669 ();
 DECAPx1_ASAP7_75t_R FILLER_0_162_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_687 ();
 FILLER_ASAP7_75t_R FILLER_0_162_708 ();
 FILLER_ASAP7_75t_R FILLER_0_162_720 ();
 DECAPx1_ASAP7_75t_R FILLER_0_162_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_162_738 ();
 FILLER_ASAP7_75t_R FILLER_0_162_744 ();
 DECAPx1_ASAP7_75t_R FILLER_0_162_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_753 ();
 DECAPx6_ASAP7_75t_R FILLER_0_162_760 ();
 DECAPx1_ASAP7_75t_R FILLER_0_162_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_778 ();
 FILLER_ASAP7_75t_R FILLER_0_162_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_801 ();
 FILLER_ASAP7_75t_R FILLER_0_162_808 ();
 DECAPx4_ASAP7_75t_R FILLER_0_162_821 ();
 DECAPx4_ASAP7_75t_R FILLER_0_162_841 ();
 FILLER_ASAP7_75t_R FILLER_0_162_851 ();
 DECAPx6_ASAP7_75t_R FILLER_0_162_861 ();
 FILLER_ASAP7_75t_R FILLER_0_162_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_877 ();
 FILLER_ASAP7_75t_R FILLER_0_162_884 ();
 DECAPx2_ASAP7_75t_R FILLER_0_162_892 ();
 FILLER_ASAP7_75t_R FILLER_0_162_898 ();
 DECAPx6_ASAP7_75t_R FILLER_0_162_906 ();
 FILLER_ASAP7_75t_R FILLER_0_162_920 ();
 FILLER_ASAP7_75t_R FILLER_0_162_930 ();
 DECAPx1_ASAP7_75t_R FILLER_0_162_938 ();
 DECAPx1_ASAP7_75t_R FILLER_0_162_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_950 ();
 FILLER_ASAP7_75t_R FILLER_0_162_961 ();
 DECAPx2_ASAP7_75t_R FILLER_0_162_971 ();
 DECAPx2_ASAP7_75t_R FILLER_0_162_985 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_991 ();
 DECAPx10_ASAP7_75t_R FILLER_0_162_1003 ();
 DECAPx6_ASAP7_75t_R FILLER_0_162_1025 ();
 FILLER_ASAP7_75t_R FILLER_0_162_1039 ();
 FILLER_ASAP7_75t_R FILLER_0_162_1053 ();
 FILLER_ASAP7_75t_R FILLER_0_162_1061 ();
 FILLER_ASAP7_75t_R FILLER_0_162_1069 ();
 FILLER_ASAP7_75t_R FILLER_0_162_1079 ();
 FILLER_ASAP7_75t_R FILLER_0_162_1092 ();
 DECAPx6_ASAP7_75t_R FILLER_0_162_1100 ();
 DECAPx1_ASAP7_75t_R FILLER_0_162_1114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_162_1124 ();
 FILLER_ASAP7_75t_R FILLER_0_162_1146 ();
 DECAPx1_ASAP7_75t_R FILLER_0_162_1169 ();
 DECAPx1_ASAP7_75t_R FILLER_0_162_1184 ();
 FILLER_ASAP7_75t_R FILLER_0_162_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_1196 ();
 FILLER_ASAP7_75t_R FILLER_0_162_1217 ();
 DECAPx4_ASAP7_75t_R FILLER_0_162_1226 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_1236 ();
 DECAPx1_ASAP7_75t_R FILLER_0_162_1243 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_1247 ();
 DECAPx6_ASAP7_75t_R FILLER_0_162_1254 ();
 DECAPx2_ASAP7_75t_R FILLER_0_162_1268 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_1274 ();
 DECAPx2_ASAP7_75t_R FILLER_0_162_1280 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_1286 ();
 FILLER_ASAP7_75t_R FILLER_0_162_1293 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_1295 ();
 FILLER_ASAP7_75t_R FILLER_0_162_1299 ();
 FILLER_ASAP7_75t_R FILLER_0_162_1307 ();
 FILLER_ASAP7_75t_R FILLER_0_162_1317 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_1319 ();
 FILLER_ASAP7_75t_R FILLER_0_162_1323 ();
 FILLER_ASAP7_75t_R FILLER_0_162_1331 ();
 DECAPx1_ASAP7_75t_R FILLER_0_162_1339 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_1343 ();
 FILLER_ASAP7_75t_R FILLER_0_162_1349 ();
 FILLER_ASAP7_75t_R FILLER_0_162_1356 ();
 FILLER_ASAP7_75t_R FILLER_0_162_1363 ();
 FILLER_ASAP7_75t_R FILLER_0_162_1370 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162_1372 ();
 DECAPx1_ASAP7_75t_R FILLER_0_162_1378 ();
 FILLER_ASAP7_75t_R FILLER_0_163_2 ();
 FILLER_ASAP7_75t_R FILLER_0_163_9 ();
 FILLER_ASAP7_75t_R FILLER_0_163_32 ();
 FILLER_ASAP7_75t_R FILLER_0_163_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_57 ();
 FILLER_ASAP7_75t_R FILLER_0_163_61 ();
 FILLER_ASAP7_75t_R FILLER_0_163_69 ();
 FILLER_ASAP7_75t_R FILLER_0_163_81 ();
 DECAPx1_ASAP7_75t_R FILLER_0_163_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_92 ();
 DECAPx4_ASAP7_75t_R FILLER_0_163_103 ();
 FILLER_ASAP7_75t_R FILLER_0_163_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_115 ();
 DECAPx1_ASAP7_75t_R FILLER_0_163_124 ();
 FILLER_ASAP7_75t_R FILLER_0_163_138 ();
 DECAPx1_ASAP7_75t_R FILLER_0_163_150 ();
 DECAPx6_ASAP7_75t_R FILLER_0_163_174 ();
 FILLER_ASAP7_75t_R FILLER_0_163_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_190 ();
 FILLER_ASAP7_75t_R FILLER_0_163_194 ();
 DECAPx1_ASAP7_75t_R FILLER_0_163_202 ();
 FILLER_ASAP7_75t_R FILLER_0_163_218 ();
 DECAPx6_ASAP7_75t_R FILLER_0_163_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_240 ();
 FILLER_ASAP7_75t_R FILLER_0_163_249 ();
 FILLER_ASAP7_75t_R FILLER_0_163_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_256 ();
 FILLER_ASAP7_75t_R FILLER_0_163_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_263 ();
 DECAPx6_ASAP7_75t_R FILLER_0_163_270 ();
 DECAPx2_ASAP7_75t_R FILLER_0_163_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_290 ();
 FILLER_ASAP7_75t_R FILLER_0_163_297 ();
 FILLER_ASAP7_75t_R FILLER_0_163_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_309 ();
 FILLER_ASAP7_75t_R FILLER_0_163_316 ();
 DECAPx1_ASAP7_75t_R FILLER_0_163_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_330 ();
 FILLER_ASAP7_75t_R FILLER_0_163_337 ();
 DECAPx2_ASAP7_75t_R FILLER_0_163_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_352 ();
 DECAPx1_ASAP7_75t_R FILLER_0_163_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_363 ();
 DECAPx4_ASAP7_75t_R FILLER_0_163_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_384 ();
 FILLER_ASAP7_75t_R FILLER_0_163_391 ();
 FILLER_ASAP7_75t_R FILLER_0_163_401 ();
 DECAPx1_ASAP7_75t_R FILLER_0_163_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_410 ();
 DECAPx6_ASAP7_75t_R FILLER_0_163_417 ();
 DECAPx2_ASAP7_75t_R FILLER_0_163_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_437 ();
 DECAPx10_ASAP7_75t_R FILLER_0_163_444 ();
 DECAPx1_ASAP7_75t_R FILLER_0_163_476 ();
 FILLER_ASAP7_75t_R FILLER_0_163_483 ();
 FILLER_ASAP7_75t_R FILLER_0_163_491 ();
 FILLER_ASAP7_75t_R FILLER_0_163_499 ();
 FILLER_ASAP7_75t_R FILLER_0_163_507 ();
 FILLER_ASAP7_75t_R FILLER_0_163_515 ();
 DECAPx6_ASAP7_75t_R FILLER_0_163_522 ();
 DECAPx2_ASAP7_75t_R FILLER_0_163_536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_163_548 ();
 DECAPx6_ASAP7_75t_R FILLER_0_163_570 ();
 DECAPx4_ASAP7_75t_R FILLER_0_163_592 ();
 FILLER_ASAP7_75t_R FILLER_0_163_602 ();
 DECAPx2_ASAP7_75t_R FILLER_0_163_610 ();
 FILLER_ASAP7_75t_R FILLER_0_163_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_163_626 ();
 DECAPx6_ASAP7_75t_R FILLER_0_163_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_662 ();
 DECAPx6_ASAP7_75t_R FILLER_0_163_666 ();
 DECAPx1_ASAP7_75t_R FILLER_0_163_680 ();
 FILLER_ASAP7_75t_R FILLER_0_163_690 ();
 FILLER_ASAP7_75t_R FILLER_0_163_698 ();
 FILLER_ASAP7_75t_R FILLER_0_163_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_709 ();
 DECAPx1_ASAP7_75t_R FILLER_0_163_716 ();
 DECAPx1_ASAP7_75t_R FILLER_0_163_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_730 ();
 FILLER_ASAP7_75t_R FILLER_0_163_737 ();
 FILLER_ASAP7_75t_R FILLER_0_163_745 ();
 FILLER_ASAP7_75t_R FILLER_0_163_753 ();
 FILLER_ASAP7_75t_R FILLER_0_163_761 ();
 DECAPx1_ASAP7_75t_R FILLER_0_163_769 ();
 FILLER_ASAP7_75t_R FILLER_0_163_779 ();
 DECAPx2_ASAP7_75t_R FILLER_0_163_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_793 ();
 FILLER_ASAP7_75t_R FILLER_0_163_800 ();
 FILLER_ASAP7_75t_R FILLER_0_163_810 ();
 FILLER_ASAP7_75t_R FILLER_0_163_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_821 ();
 DECAPx2_ASAP7_75t_R FILLER_0_163_827 ();
 FILLER_ASAP7_75t_R FILLER_0_163_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_835 ();
 DECAPx1_ASAP7_75t_R FILLER_0_163_844 ();
 FILLER_ASAP7_75t_R FILLER_0_163_859 ();
 FILLER_ASAP7_75t_R FILLER_0_163_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_870 ();
 FILLER_ASAP7_75t_R FILLER_0_163_877 ();
 FILLER_ASAP7_75t_R FILLER_0_163_885 ();
 FILLER_ASAP7_75t_R FILLER_0_163_893 ();
 FILLER_ASAP7_75t_R FILLER_0_163_901 ();
 FILLER_ASAP7_75t_R FILLER_0_163_923 ();
 DECAPx2_ASAP7_75t_R FILLER_0_163_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_933 ();
 FILLER_ASAP7_75t_R FILLER_0_163_954 ();
 FILLER_ASAP7_75t_R FILLER_0_163_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_966 ();
 DECAPx1_ASAP7_75t_R FILLER_0_163_973 ();
 DECAPx10_ASAP7_75t_R FILLER_0_163_985 ();
 DECAPx10_ASAP7_75t_R FILLER_0_163_1007 ();
 DECAPx2_ASAP7_75t_R FILLER_0_163_1029 ();
 FILLER_ASAP7_75t_R FILLER_0_163_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_1037 ();
 FILLER_ASAP7_75t_R FILLER_0_163_1049 ();
 FILLER_ASAP7_75t_R FILLER_0_163_1063 ();
 FILLER_ASAP7_75t_R FILLER_0_163_1073 ();
 DECAPx2_ASAP7_75t_R FILLER_0_163_1081 ();
 FILLER_ASAP7_75t_R FILLER_0_163_1087 ();
 DECAPx2_ASAP7_75t_R FILLER_0_163_1101 ();
 FILLER_ASAP7_75t_R FILLER_0_163_1112 ();
 FILLER_ASAP7_75t_R FILLER_0_163_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_1128 ();
 DECAPx2_ASAP7_75t_R FILLER_0_163_1137 ();
 FILLER_ASAP7_75t_R FILLER_0_163_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_1145 ();
 DECAPx2_ASAP7_75t_R FILLER_0_163_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_1173 ();
 FILLER_ASAP7_75t_R FILLER_0_163_1180 ();
 FILLER_ASAP7_75t_R FILLER_0_163_1188 ();
 FILLER_ASAP7_75t_R FILLER_0_163_1200 ();
 FILLER_ASAP7_75t_R FILLER_0_163_1208 ();
 FILLER_ASAP7_75t_R FILLER_0_163_1220 ();
 FILLER_ASAP7_75t_R FILLER_0_163_1228 ();
 DECAPx6_ASAP7_75t_R FILLER_0_163_1236 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_1250 ();
 DECAPx4_ASAP7_75t_R FILLER_0_163_1257 ();
 DECAPx2_ASAP7_75t_R FILLER_0_163_1273 ();
 FILLER_ASAP7_75t_R FILLER_0_163_1279 ();
 FILLER_ASAP7_75t_R FILLER_0_163_1287 ();
 DECAPx4_ASAP7_75t_R FILLER_0_163_1295 ();
 FILLER_ASAP7_75t_R FILLER_0_163_1305 ();
 FILLER_ASAP7_75t_R FILLER_0_163_1313 ();
 DECAPx2_ASAP7_75t_R FILLER_0_163_1321 ();
 FILLER_ASAP7_75t_R FILLER_0_163_1333 ();
 FILLER_ASAP7_75t_R FILLER_0_163_1341 ();
 DECAPx1_ASAP7_75t_R FILLER_0_163_1348 ();
 FILLER_ASAP7_75t_R FILLER_0_163_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_163_1364 ();
 FILLER_ASAP7_75t_R FILLER_0_163_1372 ();
 FILLER_ASAP7_75t_R FILLER_0_163_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_164_2 ();
 FILLER_ASAP7_75t_R FILLER_0_164_9 ();
 FILLER_ASAP7_75t_R FILLER_0_164_16 ();
 FILLER_ASAP7_75t_R FILLER_0_164_23 ();
 FILLER_ASAP7_75t_R FILLER_0_164_31 ();
 FILLER_ASAP7_75t_R FILLER_0_164_39 ();
 FILLER_ASAP7_75t_R FILLER_0_164_47 ();
 FILLER_ASAP7_75t_R FILLER_0_164_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_56 ();
 FILLER_ASAP7_75t_R FILLER_0_164_77 ();
 FILLER_ASAP7_75t_R FILLER_0_164_84 ();
 DECAPx2_ASAP7_75t_R FILLER_0_164_91 ();
 FILLER_ASAP7_75t_R FILLER_0_164_97 ();
 DECAPx4_ASAP7_75t_R FILLER_0_164_107 ();
 FILLER_ASAP7_75t_R FILLER_0_164_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_131 ();
 FILLER_ASAP7_75t_R FILLER_0_164_143 ();
 DECAPx2_ASAP7_75t_R FILLER_0_164_151 ();
 DECAPx6_ASAP7_75t_R FILLER_0_164_165 ();
 DECAPx6_ASAP7_75t_R FILLER_0_164_200 ();
 FILLER_ASAP7_75t_R FILLER_0_164_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_216 ();
 FILLER_ASAP7_75t_R FILLER_0_164_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_240 ();
 DECAPx6_ASAP7_75t_R FILLER_0_164_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_263 ();
 FILLER_ASAP7_75t_R FILLER_0_164_284 ();
 DECAPx6_ASAP7_75t_R FILLER_0_164_294 ();
 FILLER_ASAP7_75t_R FILLER_0_164_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_310 ();
 DECAPx4_ASAP7_75t_R FILLER_0_164_317 ();
 FILLER_ASAP7_75t_R FILLER_0_164_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_329 ();
 DECAPx2_ASAP7_75t_R FILLER_0_164_336 ();
 FILLER_ASAP7_75t_R FILLER_0_164_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_344 ();
 FILLER_ASAP7_75t_R FILLER_0_164_351 ();
 DECAPx1_ASAP7_75t_R FILLER_0_164_360 ();
 DECAPx2_ASAP7_75t_R FILLER_0_164_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_376 ();
 FILLER_ASAP7_75t_R FILLER_0_164_397 ();
 DECAPx1_ASAP7_75t_R FILLER_0_164_405 ();
 DECAPx2_ASAP7_75t_R FILLER_0_164_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_421 ();
 FILLER_ASAP7_75t_R FILLER_0_164_428 ();
 DECAPx4_ASAP7_75t_R FILLER_0_164_450 ();
 FILLER_ASAP7_75t_R FILLER_0_164_460 ();
 DECAPx6_ASAP7_75t_R FILLER_0_164_464 ();
 FILLER_ASAP7_75t_R FILLER_0_164_484 ();
 FILLER_ASAP7_75t_R FILLER_0_164_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_494 ();
 FILLER_ASAP7_75t_R FILLER_0_164_515 ();
 DECAPx4_ASAP7_75t_R FILLER_0_164_525 ();
 FILLER_ASAP7_75t_R FILLER_0_164_535 ();
 DECAPx2_ASAP7_75t_R FILLER_0_164_540 ();
 FILLER_ASAP7_75t_R FILLER_0_164_553 ();
 FILLER_ASAP7_75t_R FILLER_0_164_561 ();
 FILLER_ASAP7_75t_R FILLER_0_164_569 ();
 DECAPx10_ASAP7_75t_R FILLER_0_164_574 ();
 FILLER_ASAP7_75t_R FILLER_0_164_596 ();
 FILLER_ASAP7_75t_R FILLER_0_164_604 ();
 DECAPx6_ASAP7_75t_R FILLER_0_164_612 ();
 DECAPx1_ASAP7_75t_R FILLER_0_164_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_630 ();
 FILLER_ASAP7_75t_R FILLER_0_164_637 ();
 DECAPx4_ASAP7_75t_R FILLER_0_164_645 ();
 DECAPx10_ASAP7_75t_R FILLER_0_164_661 ();
 DECAPx1_ASAP7_75t_R FILLER_0_164_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_687 ();
 FILLER_ASAP7_75t_R FILLER_0_164_693 ();
 FILLER_ASAP7_75t_R FILLER_0_164_701 ();
 FILLER_ASAP7_75t_R FILLER_0_164_709 ();
 FILLER_ASAP7_75t_R FILLER_0_164_717 ();
 FILLER_ASAP7_75t_R FILLER_0_164_725 ();
 DECAPx1_ASAP7_75t_R FILLER_0_164_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_737 ();
 DECAPx10_ASAP7_75t_R FILLER_0_164_749 ();
 DECAPx4_ASAP7_75t_R FILLER_0_164_771 ();
 FILLER_ASAP7_75t_R FILLER_0_164_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_783 ();
 DECAPx2_ASAP7_75t_R FILLER_0_164_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_793 ();
 DECAPx4_ASAP7_75t_R FILLER_0_164_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_810 ();
 FILLER_ASAP7_75t_R FILLER_0_164_835 ();
 FILLER_ASAP7_75t_R FILLER_0_164_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_845 ();
 DECAPx2_ASAP7_75t_R FILLER_0_164_852 ();
 FILLER_ASAP7_75t_R FILLER_0_164_864 ();
 DECAPx1_ASAP7_75t_R FILLER_0_164_872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_164_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_904 ();
 DECAPx6_ASAP7_75t_R FILLER_0_164_908 ();
 FILLER_ASAP7_75t_R FILLER_0_164_922 ();
 FILLER_ASAP7_75t_R FILLER_0_164_930 ();
 DECAPx2_ASAP7_75t_R FILLER_0_164_938 ();
 FILLER_ASAP7_75t_R FILLER_0_164_944 ();
 FILLER_ASAP7_75t_R FILLER_0_164_956 ();
 FILLER_ASAP7_75t_R FILLER_0_164_966 ();
 FILLER_ASAP7_75t_R FILLER_0_164_976 ();
 FILLER_ASAP7_75t_R FILLER_0_164_984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_164_992 ();
 DECAPx2_ASAP7_75t_R FILLER_0_164_1014 ();
 DECAPx6_ASAP7_75t_R FILLER_0_164_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_1055 ();
 DECAPx6_ASAP7_75t_R FILLER_0_164_1068 ();
 DECAPx1_ASAP7_75t_R FILLER_0_164_1082 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_1086 ();
 FILLER_ASAP7_75t_R FILLER_0_164_1090 ();
 FILLER_ASAP7_75t_R FILLER_0_164_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_1102 ();
 FILLER_ASAP7_75t_R FILLER_0_164_1115 ();
 FILLER_ASAP7_75t_R FILLER_0_164_1129 ();
 DECAPx4_ASAP7_75t_R FILLER_0_164_1137 ();
 FILLER_ASAP7_75t_R FILLER_0_164_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_1149 ();
 FILLER_ASAP7_75t_R FILLER_0_164_1153 ();
 DECAPx2_ASAP7_75t_R FILLER_0_164_1158 ();
 FILLER_ASAP7_75t_R FILLER_0_164_1164 ();
 DECAPx2_ASAP7_75t_R FILLER_0_164_1176 ();
 FILLER_ASAP7_75t_R FILLER_0_164_1182 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_1184 ();
 DECAPx1_ASAP7_75t_R FILLER_0_164_1191 ();
 DECAPx2_ASAP7_75t_R FILLER_0_164_1201 ();
 FILLER_ASAP7_75t_R FILLER_0_164_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_1209 ();
 DECAPx2_ASAP7_75t_R FILLER_0_164_1216 ();
 FILLER_ASAP7_75t_R FILLER_0_164_1228 ();
 DECAPx6_ASAP7_75t_R FILLER_0_164_1233 ();
 DECAPx1_ASAP7_75t_R FILLER_0_164_1247 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_1251 ();
 DECAPx1_ASAP7_75t_R FILLER_0_164_1258 ();
 FILLER_ASAP7_75t_R FILLER_0_164_1268 ();
 FILLER_ASAP7_75t_R FILLER_0_164_1277 ();
 FILLER_ASAP7_75t_R FILLER_0_164_1285 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_1287 ();
 FILLER_ASAP7_75t_R FILLER_0_164_1294 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_1296 ();
 FILLER_ASAP7_75t_R FILLER_0_164_1307 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_1309 ();
 FILLER_ASAP7_75t_R FILLER_0_164_1313 ();
 FILLER_ASAP7_75t_R FILLER_0_164_1320 ();
 FILLER_ASAP7_75t_R FILLER_0_164_1327 ();
 FILLER_ASAP7_75t_R FILLER_0_164_1335 ();
 DECAPx1_ASAP7_75t_R FILLER_0_164_1343 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164_1347 ();
 DECAPx2_ASAP7_75t_R FILLER_0_164_1354 ();
 FILLER_ASAP7_75t_R FILLER_0_164_1365 ();
 FILLER_ASAP7_75t_R FILLER_0_164_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_164_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_165_2 ();
 FILLER_ASAP7_75t_R FILLER_0_165_9 ();
 FILLER_ASAP7_75t_R FILLER_0_165_16 ();
 FILLER_ASAP7_75t_R FILLER_0_165_24 ();
 FILLER_ASAP7_75t_R FILLER_0_165_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_33 ();
 FILLER_ASAP7_75t_R FILLER_0_165_37 ();
 FILLER_ASAP7_75t_R FILLER_0_165_44 ();
 FILLER_ASAP7_75t_R FILLER_0_165_51 ();
 FILLER_ASAP7_75t_R FILLER_0_165_58 ();
 FILLER_ASAP7_75t_R FILLER_0_165_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_67 ();
 FILLER_ASAP7_75t_R FILLER_0_165_80 ();
 FILLER_ASAP7_75t_R FILLER_0_165_87 ();
 FILLER_ASAP7_75t_R FILLER_0_165_92 ();
 FILLER_ASAP7_75t_R FILLER_0_165_104 ();
 FILLER_ASAP7_75t_R FILLER_0_165_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_129 ();
 FILLER_ASAP7_75t_R FILLER_0_165_136 ();
 DECAPx2_ASAP7_75t_R FILLER_0_165_146 ();
 FILLER_ASAP7_75t_R FILLER_0_165_155 ();
 DECAPx2_ASAP7_75t_R FILLER_0_165_163 ();
 FILLER_ASAP7_75t_R FILLER_0_165_169 ();
 FILLER_ASAP7_75t_R FILLER_0_165_177 ();
 FILLER_ASAP7_75t_R FILLER_0_165_185 ();
 DECAPx10_ASAP7_75t_R FILLER_0_165_190 ();
 DECAPx1_ASAP7_75t_R FILLER_0_165_212 ();
 FILLER_ASAP7_75t_R FILLER_0_165_219 ();
 FILLER_ASAP7_75t_R FILLER_0_165_231 ();
 FILLER_ASAP7_75t_R FILLER_0_165_239 ();
 DECAPx4_ASAP7_75t_R FILLER_0_165_247 ();
 FILLER_ASAP7_75t_R FILLER_0_165_257 ();
 FILLER_ASAP7_75t_R FILLER_0_165_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_271 ();
 FILLER_ASAP7_75t_R FILLER_0_165_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_280 ();
 FILLER_ASAP7_75t_R FILLER_0_165_287 ();
 FILLER_ASAP7_75t_R FILLER_0_165_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_311 ();
 DECAPx2_ASAP7_75t_R FILLER_0_165_318 ();
 FILLER_ASAP7_75t_R FILLER_0_165_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_326 ();
 FILLER_ASAP7_75t_R FILLER_0_165_333 ();
 DECAPx6_ASAP7_75t_R FILLER_0_165_341 ();
 DECAPx1_ASAP7_75t_R FILLER_0_165_355 ();
 FILLER_ASAP7_75t_R FILLER_0_165_362 ();
 DECAPx10_ASAP7_75t_R FILLER_0_165_370 ();
 DECAPx1_ASAP7_75t_R FILLER_0_165_398 ();
 FILLER_ASAP7_75t_R FILLER_0_165_408 ();
 DECAPx2_ASAP7_75t_R FILLER_0_165_418 ();
 FILLER_ASAP7_75t_R FILLER_0_165_424 ();
 FILLER_ASAP7_75t_R FILLER_0_165_432 ();
 FILLER_ASAP7_75t_R FILLER_0_165_440 ();
 FILLER_ASAP7_75t_R FILLER_0_165_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_450 ();
 DECAPx1_ASAP7_75t_R FILLER_0_165_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_461 ();
 FILLER_ASAP7_75t_R FILLER_0_165_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_470 ();
 DECAPx4_ASAP7_75t_R FILLER_0_165_474 ();
 FILLER_ASAP7_75t_R FILLER_0_165_484 ();
 FILLER_ASAP7_75t_R FILLER_0_165_492 ();
 FILLER_ASAP7_75t_R FILLER_0_165_500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_165_508 ();
 DECAPx1_ASAP7_75t_R FILLER_0_165_530 ();
 DECAPx2_ASAP7_75t_R FILLER_0_165_540 ();
 FILLER_ASAP7_75t_R FILLER_0_165_552 ();
 DECAPx4_ASAP7_75t_R FILLER_0_165_560 ();
 FILLER_ASAP7_75t_R FILLER_0_165_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_572 ();
 FILLER_ASAP7_75t_R FILLER_0_165_581 ();
 DECAPx2_ASAP7_75t_R FILLER_0_165_603 ();
 DECAPx6_ASAP7_75t_R FILLER_0_165_616 ();
 FILLER_ASAP7_75t_R FILLER_0_165_636 ();
 DECAPx1_ASAP7_75t_R FILLER_0_165_645 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_649 ();
 DECAPx10_ASAP7_75t_R FILLER_0_165_656 ();
 DECAPx2_ASAP7_75t_R FILLER_0_165_678 ();
 FILLER_ASAP7_75t_R FILLER_0_165_694 ();
 FILLER_ASAP7_75t_R FILLER_0_165_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_165_724 ();
 DECAPx10_ASAP7_75t_R FILLER_0_165_746 ();
 FILLER_ASAP7_75t_R FILLER_0_165_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_770 ();
 FILLER_ASAP7_75t_R FILLER_0_165_782 ();
 DECAPx6_ASAP7_75t_R FILLER_0_165_787 ();
 DECAPx1_ASAP7_75t_R FILLER_0_165_801 ();
 FILLER_ASAP7_75t_R FILLER_0_165_811 ();
 DECAPx10_ASAP7_75t_R FILLER_0_165_818 ();
 DECAPx6_ASAP7_75t_R FILLER_0_165_840 ();
 FILLER_ASAP7_75t_R FILLER_0_165_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_856 ();
 DECAPx2_ASAP7_75t_R FILLER_0_165_861 ();
 DECAPx10_ASAP7_75t_R FILLER_0_165_873 ();
 DECAPx1_ASAP7_75t_R FILLER_0_165_895 ();
 DECAPx2_ASAP7_75t_R FILLER_0_165_905 ();
 FILLER_ASAP7_75t_R FILLER_0_165_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_913 ();
 FILLER_ASAP7_75t_R FILLER_0_165_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_924 ();
 DECAPx6_ASAP7_75t_R FILLER_0_165_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_941 ();
 DECAPx2_ASAP7_75t_R FILLER_0_165_948 ();
 FILLER_ASAP7_75t_R FILLER_0_165_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_956 ();
 FILLER_ASAP7_75t_R FILLER_0_165_962 ();
 DECAPx2_ASAP7_75t_R FILLER_0_165_970 ();
 FILLER_ASAP7_75t_R FILLER_0_165_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_978 ();
 DECAPx4_ASAP7_75t_R FILLER_0_165_987 ();
 FILLER_ASAP7_75t_R FILLER_0_165_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_999 ();
 FILLER_ASAP7_75t_R FILLER_0_165_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_1010 ();
 FILLER_ASAP7_75t_R FILLER_0_165_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_1021 ();
 DECAPx10_ASAP7_75t_R FILLER_0_165_1025 ();
 DECAPx2_ASAP7_75t_R FILLER_0_165_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_1053 ();
 DECAPx6_ASAP7_75t_R FILLER_0_165_1058 ();
 FILLER_ASAP7_75t_R FILLER_0_165_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_1074 ();
 DECAPx1_ASAP7_75t_R FILLER_0_165_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_1089 ();
 FILLER_ASAP7_75t_R FILLER_0_165_1093 ();
 DECAPx6_ASAP7_75t_R FILLER_0_165_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_1115 ();
 DECAPx2_ASAP7_75t_R FILLER_0_165_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_1134 ();
 DECAPx2_ASAP7_75t_R FILLER_0_165_1140 ();
 FILLER_ASAP7_75t_R FILLER_0_165_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_1148 ();
 FILLER_ASAP7_75t_R FILLER_0_165_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_1157 ();
 FILLER_ASAP7_75t_R FILLER_0_165_1163 ();
 DECAPx10_ASAP7_75t_R FILLER_0_165_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_165_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_1210 ();
 FILLER_ASAP7_75t_R FILLER_0_165_1222 ();
 FILLER_ASAP7_75t_R FILLER_0_165_1231 ();
 FILLER_ASAP7_75t_R FILLER_0_165_1236 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_1238 ();
 FILLER_ASAP7_75t_R FILLER_0_165_1250 ();
 DECAPx6_ASAP7_75t_R FILLER_0_165_1262 ();
 DECAPx2_ASAP7_75t_R FILLER_0_165_1282 ();
 FILLER_ASAP7_75t_R FILLER_0_165_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_165_1294 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165_1316 ();
 FILLER_ASAP7_75t_R FILLER_0_165_1322 ();
 FILLER_ASAP7_75t_R FILLER_0_165_1329 ();
 FILLER_ASAP7_75t_R FILLER_0_165_1336 ();
 FILLER_ASAP7_75t_R FILLER_0_165_1359 ();
 FILLER_ASAP7_75t_R FILLER_0_165_1366 ();
 FILLER_ASAP7_75t_R FILLER_0_165_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_165_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_166_2 ();
 FILLER_ASAP7_75t_R FILLER_0_166_10 ();
 FILLER_ASAP7_75t_R FILLER_0_166_17 ();
 FILLER_ASAP7_75t_R FILLER_0_166_25 ();
 FILLER_ASAP7_75t_R FILLER_0_166_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_35 ();
 FILLER_ASAP7_75t_R FILLER_0_166_41 ();
 FILLER_ASAP7_75t_R FILLER_0_166_48 ();
 FILLER_ASAP7_75t_R FILLER_0_166_53 ();
 FILLER_ASAP7_75t_R FILLER_0_166_76 ();
 FILLER_ASAP7_75t_R FILLER_0_166_90 ();
 FILLER_ASAP7_75t_R FILLER_0_166_97 ();
 DECAPx2_ASAP7_75t_R FILLER_0_166_104 ();
 FILLER_ASAP7_75t_R FILLER_0_166_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_118 ();
 FILLER_ASAP7_75t_R FILLER_0_166_129 ();
 FILLER_ASAP7_75t_R FILLER_0_166_142 ();
 FILLER_ASAP7_75t_R FILLER_0_166_147 ();
 FILLER_ASAP7_75t_R FILLER_0_166_157 ();
 FILLER_ASAP7_75t_R FILLER_0_166_162 ();
 FILLER_ASAP7_75t_R FILLER_0_166_172 ();
 DECAPx4_ASAP7_75t_R FILLER_0_166_182 ();
 DECAPx4_ASAP7_75t_R FILLER_0_166_198 ();
 DECAPx10_ASAP7_75t_R FILLER_0_166_220 ();
 DECAPx10_ASAP7_75t_R FILLER_0_166_242 ();
 FILLER_ASAP7_75t_R FILLER_0_166_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_266 ();
 FILLER_ASAP7_75t_R FILLER_0_166_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_272 ();
 FILLER_ASAP7_75t_R FILLER_0_166_280 ();
 DECAPx2_ASAP7_75t_R FILLER_0_166_288 ();
 FILLER_ASAP7_75t_R FILLER_0_166_294 ();
 FILLER_ASAP7_75t_R FILLER_0_166_302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_166_310 ();
 FILLER_ASAP7_75t_R FILLER_0_166_338 ();
 DECAPx4_ASAP7_75t_R FILLER_0_166_346 ();
 DECAPx2_ASAP7_75t_R FILLER_0_166_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_368 ();
 FILLER_ASAP7_75t_R FILLER_0_166_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_374 ();
 DECAPx1_ASAP7_75t_R FILLER_0_166_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_389 ();
 FILLER_ASAP7_75t_R FILLER_0_166_393 ();
 DECAPx1_ASAP7_75t_R FILLER_0_166_400 ();
 DECAPx6_ASAP7_75t_R FILLER_0_166_411 ();
 DECAPx4_ASAP7_75t_R FILLER_0_166_449 ();
 FILLER_ASAP7_75t_R FILLER_0_166_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_461 ();
 DECAPx2_ASAP7_75t_R FILLER_0_166_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_470 ();
 DECAPx4_ASAP7_75t_R FILLER_0_166_478 ();
 FILLER_ASAP7_75t_R FILLER_0_166_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_490 ();
 FILLER_ASAP7_75t_R FILLER_0_166_498 ();
 FILLER_ASAP7_75t_R FILLER_0_166_503 ();
 FILLER_ASAP7_75t_R FILLER_0_166_511 ();
 DECAPx2_ASAP7_75t_R FILLER_0_166_519 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_525 ();
 FILLER_ASAP7_75t_R FILLER_0_166_534 ();
 FILLER_ASAP7_75t_R FILLER_0_166_544 ();
 FILLER_ASAP7_75t_R FILLER_0_166_553 ();
 DECAPx2_ASAP7_75t_R FILLER_0_166_561 ();
 FILLER_ASAP7_75t_R FILLER_0_166_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_569 ();
 DECAPx2_ASAP7_75t_R FILLER_0_166_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_582 ();
 FILLER_ASAP7_75t_R FILLER_0_166_605 ();
 DECAPx2_ASAP7_75t_R FILLER_0_166_617 ();
 FILLER_ASAP7_75t_R FILLER_0_166_623 ();
 FILLER_ASAP7_75t_R FILLER_0_166_631 ();
 FILLER_ASAP7_75t_R FILLER_0_166_640 ();
 DECAPx2_ASAP7_75t_R FILLER_0_166_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_656 ();
 FILLER_ASAP7_75t_R FILLER_0_166_678 ();
 DECAPx2_ASAP7_75t_R FILLER_0_166_686 ();
 FILLER_ASAP7_75t_R FILLER_0_166_692 ();
 DECAPx2_ASAP7_75t_R FILLER_0_166_699 ();
 FILLER_ASAP7_75t_R FILLER_0_166_705 ();
 DECAPx2_ASAP7_75t_R FILLER_0_166_713 ();
 FILLER_ASAP7_75t_R FILLER_0_166_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_721 ();
 FILLER_ASAP7_75t_R FILLER_0_166_738 ();
 FILLER_ASAP7_75t_R FILLER_0_166_746 ();
 FILLER_ASAP7_75t_R FILLER_0_166_754 ();
 DECAPx4_ASAP7_75t_R FILLER_0_166_762 ();
 FILLER_ASAP7_75t_R FILLER_0_166_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_780 ();
 DECAPx6_ASAP7_75t_R FILLER_0_166_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_801 ();
 FILLER_ASAP7_75t_R FILLER_0_166_808 ();
 FILLER_ASAP7_75t_R FILLER_0_166_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_820 ();
 FILLER_ASAP7_75t_R FILLER_0_166_829 ();
 DECAPx6_ASAP7_75t_R FILLER_0_166_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_851 ();
 FILLER_ASAP7_75t_R FILLER_0_166_858 ();
 FILLER_ASAP7_75t_R FILLER_0_166_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_868 ();
 DECAPx1_ASAP7_75t_R FILLER_0_166_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_880 ();
 DECAPx10_ASAP7_75t_R FILLER_0_166_884 ();
 DECAPx2_ASAP7_75t_R FILLER_0_166_906 ();
 FILLER_ASAP7_75t_R FILLER_0_166_912 ();
 DECAPx1_ASAP7_75t_R FILLER_0_166_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_939 ();
 DECAPx10_ASAP7_75t_R FILLER_0_166_948 ();
 DECAPx1_ASAP7_75t_R FILLER_0_166_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_974 ();
 FILLER_ASAP7_75t_R FILLER_0_166_986 ();
 FILLER_ASAP7_75t_R FILLER_0_166_1000 ();
 FILLER_ASAP7_75t_R FILLER_0_166_1008 ();
 FILLER_ASAP7_75t_R FILLER_0_166_1018 ();
 FILLER_ASAP7_75t_R FILLER_0_166_1031 ();
 FILLER_ASAP7_75t_R FILLER_0_166_1039 ();
 DECAPx4_ASAP7_75t_R FILLER_0_166_1047 ();
 FILLER_ASAP7_75t_R FILLER_0_166_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_1059 ();
 DECAPx2_ASAP7_75t_R FILLER_0_166_1068 ();
 FILLER_ASAP7_75t_R FILLER_0_166_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_0_166_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_0_166_1102 ();
 DECAPx6_ASAP7_75t_R FILLER_0_166_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_1138 ();
 FILLER_ASAP7_75t_R FILLER_0_166_1147 ();
 FILLER_ASAP7_75t_R FILLER_0_166_1157 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_1159 ();
 FILLER_ASAP7_75t_R FILLER_0_166_1181 ();
 DECAPx10_ASAP7_75t_R FILLER_0_166_1186 ();
 DECAPx4_ASAP7_75t_R FILLER_0_166_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_0_166_1225 ();
 DECAPx10_ASAP7_75t_R FILLER_0_166_1247 ();
 DECAPx10_ASAP7_75t_R FILLER_0_166_1269 ();
 DECAPx6_ASAP7_75t_R FILLER_0_166_1291 ();
 DECAPx1_ASAP7_75t_R FILLER_0_166_1305 ();
 FILLER_ASAP7_75t_R FILLER_0_166_1315 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_1317 ();
 FILLER_ASAP7_75t_R FILLER_0_166_1321 ();
 FILLER_ASAP7_75t_R FILLER_0_166_1326 ();
 FILLER_ASAP7_75t_R FILLER_0_166_1333 ();
 FILLER_ASAP7_75t_R FILLER_0_166_1340 ();
 FILLER_ASAP7_75t_R FILLER_0_166_1347 ();
 FILLER_ASAP7_75t_R FILLER_0_166_1355 ();
 FILLER_ASAP7_75t_R FILLER_0_166_1362 ();
 FILLER_ASAP7_75t_R FILLER_0_166_1367 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166_1369 ();
 FILLER_ASAP7_75t_R FILLER_0_166_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_167_2 ();
 FILLER_ASAP7_75t_R FILLER_0_167_25 ();
 FILLER_ASAP7_75t_R FILLER_0_167_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_35 ();
 FILLER_ASAP7_75t_R FILLER_0_167_41 ();
 DECAPx2_ASAP7_75t_R FILLER_0_167_49 ();
 FILLER_ASAP7_75t_R FILLER_0_167_65 ();
 FILLER_ASAP7_75t_R FILLER_0_167_73 ();
 FILLER_ASAP7_75t_R FILLER_0_167_81 ();
 FILLER_ASAP7_75t_R FILLER_0_167_88 ();
 FILLER_ASAP7_75t_R FILLER_0_167_95 ();
 FILLER_ASAP7_75t_R FILLER_0_167_100 ();
 DECAPx6_ASAP7_75t_R FILLER_0_167_113 ();
 DECAPx1_ASAP7_75t_R FILLER_0_167_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_131 ();
 DECAPx2_ASAP7_75t_R FILLER_0_167_144 ();
 FILLER_ASAP7_75t_R FILLER_0_167_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_152 ();
 DECAPx1_ASAP7_75t_R FILLER_0_167_164 ();
 DECAPx1_ASAP7_75t_R FILLER_0_167_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_175 ();
 DECAPx2_ASAP7_75t_R FILLER_0_167_182 ();
 FILLER_ASAP7_75t_R FILLER_0_167_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_190 ();
 DECAPx2_ASAP7_75t_R FILLER_0_167_212 ();
 FILLER_ASAP7_75t_R FILLER_0_167_218 ();
 FILLER_ASAP7_75t_R FILLER_0_167_232 ();
 DECAPx10_ASAP7_75t_R FILLER_0_167_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_267 ();
 DECAPx4_ASAP7_75t_R FILLER_0_167_274 ();
 DECAPx1_ASAP7_75t_R FILLER_0_167_290 ();
 DECAPx1_ASAP7_75t_R FILLER_0_167_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_306 ();
 DECAPx6_ASAP7_75t_R FILLER_0_167_313 ();
 DECAPx2_ASAP7_75t_R FILLER_0_167_327 ();
 FILLER_ASAP7_75t_R FILLER_0_167_339 ();
 DECAPx2_ASAP7_75t_R FILLER_0_167_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_353 ();
 FILLER_ASAP7_75t_R FILLER_0_167_358 ();
 FILLER_ASAP7_75t_R FILLER_0_167_366 ();
 FILLER_ASAP7_75t_R FILLER_0_167_374 ();
 FILLER_ASAP7_75t_R FILLER_0_167_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_386 ();
 FILLER_ASAP7_75t_R FILLER_0_167_393 ();
 DECAPx1_ASAP7_75t_R FILLER_0_167_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_405 ();
 DECAPx6_ASAP7_75t_R FILLER_0_167_416 ();
 FILLER_ASAP7_75t_R FILLER_0_167_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_432 ();
 DECAPx1_ASAP7_75t_R FILLER_0_167_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_443 ();
 DECAPx4_ASAP7_75t_R FILLER_0_167_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_460 ();
 FILLER_ASAP7_75t_R FILLER_0_167_467 ();
 FILLER_ASAP7_75t_R FILLER_0_167_472 ();
 DECAPx1_ASAP7_75t_R FILLER_0_167_477 ();
 DECAPx6_ASAP7_75t_R FILLER_0_167_484 ();
 DECAPx2_ASAP7_75t_R FILLER_0_167_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_504 ();
 DECAPx4_ASAP7_75t_R FILLER_0_167_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_521 ();
 DECAPx10_ASAP7_75t_R FILLER_0_167_525 ();
 DECAPx10_ASAP7_75t_R FILLER_0_167_547 ();
 DECAPx10_ASAP7_75t_R FILLER_0_167_569 ();
 DECAPx6_ASAP7_75t_R FILLER_0_167_591 ();
 FILLER_ASAP7_75t_R FILLER_0_167_605 ();
 DECAPx4_ASAP7_75t_R FILLER_0_167_613 ();
 FILLER_ASAP7_75t_R FILLER_0_167_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_625 ();
 DECAPx4_ASAP7_75t_R FILLER_0_167_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_639 ();
 FILLER_ASAP7_75t_R FILLER_0_167_646 ();
 FILLER_ASAP7_75t_R FILLER_0_167_658 ();
 FILLER_ASAP7_75t_R FILLER_0_167_666 ();
 DECAPx2_ASAP7_75t_R FILLER_0_167_671 ();
 DECAPx10_ASAP7_75t_R FILLER_0_167_698 ();
 FILLER_ASAP7_75t_R FILLER_0_167_720 ();
 DECAPx4_ASAP7_75t_R FILLER_0_167_728 ();
 FILLER_ASAP7_75t_R FILLER_0_167_738 ();
 DECAPx4_ASAP7_75t_R FILLER_0_167_746 ();
 FILLER_ASAP7_75t_R FILLER_0_167_762 ();
 FILLER_ASAP7_75t_R FILLER_0_167_770 ();
 DECAPx2_ASAP7_75t_R FILLER_0_167_775 ();
 FILLER_ASAP7_75t_R FILLER_0_167_781 ();
 FILLER_ASAP7_75t_R FILLER_0_167_789 ();
 DECAPx6_ASAP7_75t_R FILLER_0_167_797 ();
 FILLER_ASAP7_75t_R FILLER_0_167_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_813 ();
 DECAPx2_ASAP7_75t_R FILLER_0_167_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_830 ();
 FILLER_ASAP7_75t_R FILLER_0_167_837 ();
 DECAPx4_ASAP7_75t_R FILLER_0_167_845 ();
 FILLER_ASAP7_75t_R FILLER_0_167_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_857 ();
 FILLER_ASAP7_75t_R FILLER_0_167_864 ();
 FILLER_ASAP7_75t_R FILLER_0_167_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_871 ();
 FILLER_ASAP7_75t_R FILLER_0_167_878 ();
 DECAPx2_ASAP7_75t_R FILLER_0_167_886 ();
 FILLER_ASAP7_75t_R FILLER_0_167_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_894 ();
 FILLER_ASAP7_75t_R FILLER_0_167_901 ();
 DECAPx2_ASAP7_75t_R FILLER_0_167_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_915 ();
 DECAPx2_ASAP7_75t_R FILLER_0_167_919 ();
 DECAPx2_ASAP7_75t_R FILLER_0_167_927 ();
 FILLER_ASAP7_75t_R FILLER_0_167_933 ();
 DECAPx2_ASAP7_75t_R FILLER_0_167_947 ();
 FILLER_ASAP7_75t_R FILLER_0_167_953 ();
 FILLER_ASAP7_75t_R FILLER_0_167_967 ();
 FILLER_ASAP7_75t_R FILLER_0_167_980 ();
 DECAPx1_ASAP7_75t_R FILLER_0_167_992 ();
 FILLER_ASAP7_75t_R FILLER_0_167_1002 ();
 DECAPx2_ASAP7_75t_R FILLER_0_167_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_1016 ();
 DECAPx2_ASAP7_75t_R FILLER_0_167_1023 ();
 FILLER_ASAP7_75t_R FILLER_0_167_1037 ();
 DECAPx1_ASAP7_75t_R FILLER_0_167_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_1055 ();
 FILLER_ASAP7_75t_R FILLER_0_167_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_1064 ();
 DECAPx2_ASAP7_75t_R FILLER_0_167_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_1079 ();
 FILLER_ASAP7_75t_R FILLER_0_167_1088 ();
 FILLER_ASAP7_75t_R FILLER_0_167_1098 ();
 DECAPx2_ASAP7_75t_R FILLER_0_167_1106 ();
 FILLER_ASAP7_75t_R FILLER_0_167_1112 ();
 DECAPx6_ASAP7_75t_R FILLER_0_167_1120 ();
 DECAPx2_ASAP7_75t_R FILLER_0_167_1134 ();
 FILLER_ASAP7_75t_R FILLER_0_167_1146 ();
 FILLER_ASAP7_75t_R FILLER_0_167_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_1154 ();
 FILLER_ASAP7_75t_R FILLER_0_167_1161 ();
 FILLER_ASAP7_75t_R FILLER_0_167_1169 ();
 DECAPx2_ASAP7_75t_R FILLER_0_167_1174 ();
 DECAPx1_ASAP7_75t_R FILLER_0_167_1201 ();
 DECAPx10_ASAP7_75t_R FILLER_0_167_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_0_167_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_0_167_1261 ();
 DECAPx6_ASAP7_75t_R FILLER_0_167_1283 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_1297 ();
 FILLER_ASAP7_75t_R FILLER_0_167_1319 ();
 DECAPx1_ASAP7_75t_R FILLER_0_167_1343 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167_1347 ();
 DECAPx2_ASAP7_75t_R FILLER_0_167_1353 ();
 FILLER_ASAP7_75t_R FILLER_0_167_1380 ();
 DECAPx1_ASAP7_75t_R FILLER_0_168_2 ();
 FILLER_ASAP7_75t_R FILLER_0_168_11 ();
 FILLER_ASAP7_75t_R FILLER_0_168_16 ();
 FILLER_ASAP7_75t_R FILLER_0_168_24 ();
 FILLER_ASAP7_75t_R FILLER_0_168_31 ();
 FILLER_ASAP7_75t_R FILLER_0_168_55 ();
 FILLER_ASAP7_75t_R FILLER_0_168_60 ();
 DECAPx1_ASAP7_75t_R FILLER_0_168_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_87 ();
 FILLER_ASAP7_75t_R FILLER_0_168_94 ();
 DECAPx1_ASAP7_75t_R FILLER_0_168_101 ();
 FILLER_ASAP7_75t_R FILLER_0_168_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_110 ();
 DECAPx6_ASAP7_75t_R FILLER_0_168_119 ();
 FILLER_ASAP7_75t_R FILLER_0_168_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_135 ();
 DECAPx6_ASAP7_75t_R FILLER_0_168_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_156 ();
 DECAPx2_ASAP7_75t_R FILLER_0_168_168 ();
 FILLER_ASAP7_75t_R FILLER_0_168_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_176 ();
 DECAPx1_ASAP7_75t_R FILLER_0_168_185 ();
 FILLER_ASAP7_75t_R FILLER_0_168_192 ();
 DECAPx2_ASAP7_75t_R FILLER_0_168_200 ();
 FILLER_ASAP7_75t_R FILLER_0_168_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_220 ();
 DECAPx10_ASAP7_75t_R FILLER_0_168_233 ();
 DECAPx4_ASAP7_75t_R FILLER_0_168_255 ();
 FILLER_ASAP7_75t_R FILLER_0_168_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_267 ();
 DECAPx2_ASAP7_75t_R FILLER_0_168_274 ();
 FILLER_ASAP7_75t_R FILLER_0_168_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_282 ();
 FILLER_ASAP7_75t_R FILLER_0_168_289 ();
 FILLER_ASAP7_75t_R FILLER_0_168_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_299 ();
 FILLER_ASAP7_75t_R FILLER_0_168_306 ();
 DECAPx1_ASAP7_75t_R FILLER_0_168_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_319 ();
 DECAPx1_ASAP7_75t_R FILLER_0_168_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_330 ();
 DECAPx1_ASAP7_75t_R FILLER_0_168_334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_168_344 ();
 DECAPx1_ASAP7_75t_R FILLER_0_168_372 ();
 FILLER_ASAP7_75t_R FILLER_0_168_382 ();
 FILLER_ASAP7_75t_R FILLER_0_168_390 ();
 FILLER_ASAP7_75t_R FILLER_0_168_400 ();
 DECAPx2_ASAP7_75t_R FILLER_0_168_408 ();
 FILLER_ASAP7_75t_R FILLER_0_168_414 ();
 DECAPx1_ASAP7_75t_R FILLER_0_168_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_426 ();
 FILLER_ASAP7_75t_R FILLER_0_168_433 ();
 FILLER_ASAP7_75t_R FILLER_0_168_442 ();
 FILLER_ASAP7_75t_R FILLER_0_168_447 ();
 FILLER_ASAP7_75t_R FILLER_0_168_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_461 ();
 FILLER_ASAP7_75t_R FILLER_0_168_464 ();
 DECAPx6_ASAP7_75t_R FILLER_0_168_474 ();
 FILLER_ASAP7_75t_R FILLER_0_168_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_490 ();
 FILLER_ASAP7_75t_R FILLER_0_168_497 ();
 DECAPx1_ASAP7_75t_R FILLER_0_168_502 ();
 FILLER_ASAP7_75t_R FILLER_0_168_509 ();
 FILLER_ASAP7_75t_R FILLER_0_168_518 ();
 FILLER_ASAP7_75t_R FILLER_0_168_526 ();
 DECAPx10_ASAP7_75t_R FILLER_0_168_534 ();
 FILLER_ASAP7_75t_R FILLER_0_168_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_558 ();
 DECAPx1_ASAP7_75t_R FILLER_0_168_567 ();
 DECAPx6_ASAP7_75t_R FILLER_0_168_581 ();
 FILLER_ASAP7_75t_R FILLER_0_168_595 ();
 FILLER_ASAP7_75t_R FILLER_0_168_603 ();
 DECAPx4_ASAP7_75t_R FILLER_0_168_612 ();
 FILLER_ASAP7_75t_R FILLER_0_168_630 ();
 DECAPx1_ASAP7_75t_R FILLER_0_168_638 ();
 FILLER_ASAP7_75t_R FILLER_0_168_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_650 ();
 DECAPx2_ASAP7_75t_R FILLER_0_168_654 ();
 DECAPx2_ASAP7_75t_R FILLER_0_168_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_673 ();
 FILLER_ASAP7_75t_R FILLER_0_168_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_168_689 ();
 FILLER_ASAP7_75t_R FILLER_0_168_727 ();
 FILLER_ASAP7_75t_R FILLER_0_168_735 ();
 FILLER_ASAP7_75t_R FILLER_0_168_743 ();
 DECAPx2_ASAP7_75t_R FILLER_0_168_755 ();
 FILLER_ASAP7_75t_R FILLER_0_168_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_783 ();
 FILLER_ASAP7_75t_R FILLER_0_168_789 ();
 FILLER_ASAP7_75t_R FILLER_0_168_797 ();
 DECAPx2_ASAP7_75t_R FILLER_0_168_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_811 ();
 FILLER_ASAP7_75t_R FILLER_0_168_818 ();
 DECAPx1_ASAP7_75t_R FILLER_0_168_826 ();
 FILLER_ASAP7_75t_R FILLER_0_168_838 ();
 DECAPx4_ASAP7_75t_R FILLER_0_168_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_856 ();
 FILLER_ASAP7_75t_R FILLER_0_168_863 ();
 DECAPx10_ASAP7_75t_R FILLER_0_168_871 ();
 DECAPx2_ASAP7_75t_R FILLER_0_168_904 ();
 DECAPx4_ASAP7_75t_R FILLER_0_168_921 ();
 FILLER_ASAP7_75t_R FILLER_0_168_931 ();
 DECAPx10_ASAP7_75t_R FILLER_0_168_954 ();
 DECAPx10_ASAP7_75t_R FILLER_0_168_976 ();
 FILLER_ASAP7_75t_R FILLER_0_168_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_1000 ();
 FILLER_ASAP7_75t_R FILLER_0_168_1023 ();
 DECAPx1_ASAP7_75t_R FILLER_0_168_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_1034 ();
 DECAPx4_ASAP7_75t_R FILLER_0_168_1046 ();
 FILLER_ASAP7_75t_R FILLER_0_168_1064 ();
 DECAPx2_ASAP7_75t_R FILLER_0_168_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_1078 ();
 DECAPx2_ASAP7_75t_R FILLER_0_168_1087 ();
 FILLER_ASAP7_75t_R FILLER_0_168_1093 ();
 DECAPx4_ASAP7_75t_R FILLER_0_168_1101 ();
 FILLER_ASAP7_75t_R FILLER_0_168_1122 ();
 DECAPx1_ASAP7_75t_R FILLER_0_168_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_1131 ();
 DECAPx4_ASAP7_75t_R FILLER_0_168_1138 ();
 DECAPx1_ASAP7_75t_R FILLER_0_168_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_1158 ();
 FILLER_ASAP7_75t_R FILLER_0_168_1170 ();
 DECAPx1_ASAP7_75t_R FILLER_0_168_1175 ();
 FILLER_ASAP7_75t_R FILLER_0_168_1182 ();
 FILLER_ASAP7_75t_R FILLER_0_168_1205 ();
 DECAPx10_ASAP7_75t_R FILLER_0_168_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_0_168_1239 ();
 FILLER_ASAP7_75t_R FILLER_0_168_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_0_168_1269 ();
 DECAPx6_ASAP7_75t_R FILLER_0_168_1291 ();
 FILLER_ASAP7_75t_R FILLER_0_168_1305 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_1307 ();
 FILLER_ASAP7_75t_R FILLER_0_168_1314 ();
 FILLER_ASAP7_75t_R FILLER_0_168_1321 ();
 DECAPx1_ASAP7_75t_R FILLER_0_168_1326 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_1330 ();
 FILLER_ASAP7_75t_R FILLER_0_168_1336 ();
 FILLER_ASAP7_75t_R FILLER_0_168_1343 ();
 FILLER_ASAP7_75t_R FILLER_0_168_1350 ();
 FILLER_ASAP7_75t_R FILLER_0_168_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_168_1364 ();
 FILLER_ASAP7_75t_R FILLER_0_168_1372 ();
 FILLER_ASAP7_75t_R FILLER_0_168_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_169_2 ();
 FILLER_ASAP7_75t_R FILLER_0_169_9 ();
 FILLER_ASAP7_75t_R FILLER_0_169_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_18 ();
 FILLER_ASAP7_75t_R FILLER_0_169_40 ();
 FILLER_ASAP7_75t_R FILLER_0_169_63 ();
 FILLER_ASAP7_75t_R FILLER_0_169_71 ();
 FILLER_ASAP7_75t_R FILLER_0_169_78 ();
 DECAPx1_ASAP7_75t_R FILLER_0_169_85 ();
 FILLER_ASAP7_75t_R FILLER_0_169_95 ();
 FILLER_ASAP7_75t_R FILLER_0_169_102 ();
 FILLER_ASAP7_75t_R FILLER_0_169_107 ();
 FILLER_ASAP7_75t_R FILLER_0_169_112 ();
 FILLER_ASAP7_75t_R FILLER_0_169_117 ();
 DECAPx4_ASAP7_75t_R FILLER_0_169_122 ();
 FILLER_ASAP7_75t_R FILLER_0_169_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_134 ();
 FILLER_ASAP7_75t_R FILLER_0_169_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_145 ();
 FILLER_ASAP7_75t_R FILLER_0_169_158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_169_170 ();
 FILLER_ASAP7_75t_R FILLER_0_169_192 ();
 FILLER_ASAP7_75t_R FILLER_0_169_199 ();
 DECAPx1_ASAP7_75t_R FILLER_0_169_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_215 ();
 FILLER_ASAP7_75t_R FILLER_0_169_222 ();
 DECAPx1_ASAP7_75t_R FILLER_0_169_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_240 ();
 DECAPx1_ASAP7_75t_R FILLER_0_169_244 ();
 DECAPx6_ASAP7_75t_R FILLER_0_169_258 ();
 DECAPx1_ASAP7_75t_R FILLER_0_169_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_279 ();
 FILLER_ASAP7_75t_R FILLER_0_169_286 ();
 DECAPx4_ASAP7_75t_R FILLER_0_169_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_169_308 ();
 DECAPx6_ASAP7_75t_R FILLER_0_169_330 ();
 DECAPx2_ASAP7_75t_R FILLER_0_169_344 ();
 DECAPx1_ASAP7_75t_R FILLER_0_169_356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_169_366 ();
 FILLER_ASAP7_75t_R FILLER_0_169_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_169_394 ();
 DECAPx2_ASAP7_75t_R FILLER_0_169_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_169_429 ();
 FILLER_ASAP7_75t_R FILLER_0_169_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_453 ();
 DECAPx2_ASAP7_75t_R FILLER_0_169_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_465 ();
 FILLER_ASAP7_75t_R FILLER_0_169_474 ();
 FILLER_ASAP7_75t_R FILLER_0_169_482 ();
 DECAPx2_ASAP7_75t_R FILLER_0_169_487 ();
 FILLER_ASAP7_75t_R FILLER_0_169_499 ();
 FILLER_ASAP7_75t_R FILLER_0_169_507 ();
 DECAPx4_ASAP7_75t_R FILLER_0_169_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_526 ();
 DECAPx2_ASAP7_75t_R FILLER_0_169_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_541 ();
 DECAPx1_ASAP7_75t_R FILLER_0_169_548 ();
 FILLER_ASAP7_75t_R FILLER_0_169_558 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_560 ();
 FILLER_ASAP7_75t_R FILLER_0_169_571 ();
 FILLER_ASAP7_75t_R FILLER_0_169_593 ();
 FILLER_ASAP7_75t_R FILLER_0_169_609 ();
 DECAPx2_ASAP7_75t_R FILLER_0_169_617 ();
 DECAPx1_ASAP7_75t_R FILLER_0_169_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_636 ();
 DECAPx10_ASAP7_75t_R FILLER_0_169_648 ();
 DECAPx6_ASAP7_75t_R FILLER_0_169_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_684 ();
 FILLER_ASAP7_75t_R FILLER_0_169_688 ();
 FILLER_ASAP7_75t_R FILLER_0_169_694 ();
 DECAPx10_ASAP7_75t_R FILLER_0_169_705 ();
 DECAPx2_ASAP7_75t_R FILLER_0_169_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_733 ();
 FILLER_ASAP7_75t_R FILLER_0_169_740 ();
 DECAPx2_ASAP7_75t_R FILLER_0_169_748 ();
 FILLER_ASAP7_75t_R FILLER_0_169_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_756 ();
 DECAPx2_ASAP7_75t_R FILLER_0_169_778 ();
 FILLER_ASAP7_75t_R FILLER_0_169_784 ();
 FILLER_ASAP7_75t_R FILLER_0_169_792 ();
 DECAPx1_ASAP7_75t_R FILLER_0_169_800 ();
 DECAPx2_ASAP7_75t_R FILLER_0_169_810 ();
 FILLER_ASAP7_75t_R FILLER_0_169_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_818 ();
 FILLER_ASAP7_75t_R FILLER_0_169_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_827 ();
 DECAPx2_ASAP7_75t_R FILLER_0_169_834 ();
 DECAPx10_ASAP7_75t_R FILLER_0_169_850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_169_872 ();
 DECAPx2_ASAP7_75t_R FILLER_0_169_894 ();
 FILLER_ASAP7_75t_R FILLER_0_169_900 ();
 FILLER_ASAP7_75t_R FILLER_0_169_923 ();
 FILLER_ASAP7_75t_R FILLER_0_169_927 ();
 DECAPx4_ASAP7_75t_R FILLER_0_169_935 ();
 FILLER_ASAP7_75t_R FILLER_0_169_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_947 ();
 FILLER_ASAP7_75t_R FILLER_0_169_951 ();
 DECAPx6_ASAP7_75t_R FILLER_0_169_965 ();
 DECAPx1_ASAP7_75t_R FILLER_0_169_979 ();
 DECAPx2_ASAP7_75t_R FILLER_0_169_995 ();
 DECAPx6_ASAP7_75t_R FILLER_0_169_1013 ();
 DECAPx1_ASAP7_75t_R FILLER_0_169_1027 ();
 FILLER_ASAP7_75t_R FILLER_0_169_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_1036 ();
 FILLER_ASAP7_75t_R FILLER_0_169_1047 ();
 DECAPx2_ASAP7_75t_R FILLER_0_169_1059 ();
 FILLER_ASAP7_75t_R FILLER_0_169_1065 ();
 DECAPx2_ASAP7_75t_R FILLER_0_169_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_1079 ();
 DECAPx10_ASAP7_75t_R FILLER_0_169_1086 ();
 DECAPx4_ASAP7_75t_R FILLER_0_169_1108 ();
 FILLER_ASAP7_75t_R FILLER_0_169_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_1120 ();
 DECAPx10_ASAP7_75t_R FILLER_0_169_1127 ();
 DECAPx4_ASAP7_75t_R FILLER_0_169_1149 ();
 FILLER_ASAP7_75t_R FILLER_0_169_1159 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_1161 ();
 FILLER_ASAP7_75t_R FILLER_0_169_1165 ();
 DECAPx4_ASAP7_75t_R FILLER_0_169_1175 ();
 FILLER_ASAP7_75t_R FILLER_0_169_1185 ();
 FILLER_ASAP7_75t_R FILLER_0_169_1192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_169_1197 ();
 FILLER_ASAP7_75t_R FILLER_0_169_1219 ();
 DECAPx6_ASAP7_75t_R FILLER_0_169_1233 ();
 DECAPx2_ASAP7_75t_R FILLER_0_169_1247 ();
 DECAPx6_ASAP7_75t_R FILLER_0_169_1274 ();
 DECAPx2_ASAP7_75t_R FILLER_0_169_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_1294 ();
 DECAPx2_ASAP7_75t_R FILLER_0_169_1317 ();
 DECAPx1_ASAP7_75t_R FILLER_0_169_1326 ();
 FILLER_ASAP7_75t_R FILLER_0_169_1333 ();
 FILLER_ASAP7_75t_R FILLER_0_169_1338 ();
 DECAPx1_ASAP7_75t_R FILLER_0_169_1345 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_1349 ();
 DECAPx1_ASAP7_75t_R FILLER_0_169_1355 ();
 FILLER_ASAP7_75t_R FILLER_0_169_1364 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169_1366 ();
 FILLER_ASAP7_75t_R FILLER_0_169_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_169_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_170_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_4 ();
 FILLER_ASAP7_75t_R FILLER_0_170_27 ();
 FILLER_ASAP7_75t_R FILLER_0_170_34 ();
 FILLER_ASAP7_75t_R FILLER_0_170_41 ();
 FILLER_ASAP7_75t_R FILLER_0_170_46 ();
 FILLER_ASAP7_75t_R FILLER_0_170_53 ();
 FILLER_ASAP7_75t_R FILLER_0_170_60 ();
 FILLER_ASAP7_75t_R FILLER_0_170_67 ();
 FILLER_ASAP7_75t_R FILLER_0_170_72 ();
 DECAPx1_ASAP7_75t_R FILLER_0_170_85 ();
 DECAPx2_ASAP7_75t_R FILLER_0_170_100 ();
 DECAPx10_ASAP7_75t_R FILLER_0_170_114 ();
 FILLER_ASAP7_75t_R FILLER_0_170_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_170_145 ();
 DECAPx4_ASAP7_75t_R FILLER_0_170_167 ();
 FILLER_ASAP7_75t_R FILLER_0_170_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_179 ();
 FILLER_ASAP7_75t_R FILLER_0_170_200 ();
 DECAPx1_ASAP7_75t_R FILLER_0_170_210 ();
 FILLER_ASAP7_75t_R FILLER_0_170_235 ();
 FILLER_ASAP7_75t_R FILLER_0_170_240 ();
 DECAPx1_ASAP7_75t_R FILLER_0_170_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_266 ();
 DECAPx4_ASAP7_75t_R FILLER_0_170_273 ();
 DECAPx6_ASAP7_75t_R FILLER_0_170_290 ();
 DECAPx6_ASAP7_75t_R FILLER_0_170_310 ();
 FILLER_ASAP7_75t_R FILLER_0_170_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_326 ();
 DECAPx4_ASAP7_75t_R FILLER_0_170_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_343 ();
 FILLER_ASAP7_75t_R FILLER_0_170_350 ();
 DECAPx6_ASAP7_75t_R FILLER_0_170_359 ();
 DECAPx2_ASAP7_75t_R FILLER_0_170_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_379 ();
 DECAPx1_ASAP7_75t_R FILLER_0_170_383 ();
 FILLER_ASAP7_75t_R FILLER_0_170_393 ();
 DECAPx2_ASAP7_75t_R FILLER_0_170_398 ();
 DECAPx1_ASAP7_75t_R FILLER_0_170_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_412 ();
 DECAPx2_ASAP7_75t_R FILLER_0_170_419 ();
 FILLER_ASAP7_75t_R FILLER_0_170_425 ();
 DECAPx10_ASAP7_75t_R FILLER_0_170_433 ();
 DECAPx2_ASAP7_75t_R FILLER_0_170_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_461 ();
 DECAPx1_ASAP7_75t_R FILLER_0_170_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_468 ();
 DECAPx1_ASAP7_75t_R FILLER_0_170_472 ();
 FILLER_ASAP7_75t_R FILLER_0_170_496 ();
 FILLER_ASAP7_75t_R FILLER_0_170_505 ();
 DECAPx6_ASAP7_75t_R FILLER_0_170_510 ();
 FILLER_ASAP7_75t_R FILLER_0_170_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_526 ();
 DECAPx2_ASAP7_75t_R FILLER_0_170_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_539 ();
 FILLER_ASAP7_75t_R FILLER_0_170_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_550 ();
 FILLER_ASAP7_75t_R FILLER_0_170_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_556 ();
 FILLER_ASAP7_75t_R FILLER_0_170_565 ();
 DECAPx6_ASAP7_75t_R FILLER_0_170_570 ();
 FILLER_ASAP7_75t_R FILLER_0_170_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_586 ();
 FILLER_ASAP7_75t_R FILLER_0_170_611 ();
 DECAPx1_ASAP7_75t_R FILLER_0_170_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_623 ();
 FILLER_ASAP7_75t_R FILLER_0_170_630 ();
 FILLER_ASAP7_75t_R FILLER_0_170_635 ();
 DECAPx2_ASAP7_75t_R FILLER_0_170_643 ();
 FILLER_ASAP7_75t_R FILLER_0_170_649 ();
 FILLER_ASAP7_75t_R FILLER_0_170_654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_170_662 ();
 FILLER_ASAP7_75t_R FILLER_0_170_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_678 ();
 FILLER_ASAP7_75t_R FILLER_0_170_688 ();
 FILLER_ASAP7_75t_R FILLER_0_170_699 ();
 DECAPx10_ASAP7_75t_R FILLER_0_170_722 ();
 DECAPx4_ASAP7_75t_R FILLER_0_170_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_754 ();
 FILLER_ASAP7_75t_R FILLER_0_170_760 ();
 DECAPx10_ASAP7_75t_R FILLER_0_170_765 ();
 DECAPx10_ASAP7_75t_R FILLER_0_170_787 ();
 DECAPx2_ASAP7_75t_R FILLER_0_170_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_815 ();
 DECAPx10_ASAP7_75t_R FILLER_0_170_822 ();
 DECAPx2_ASAP7_75t_R FILLER_0_170_844 ();
 FILLER_ASAP7_75t_R FILLER_0_170_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_852 ();
 DECAPx4_ASAP7_75t_R FILLER_0_170_865 ();
 FILLER_ASAP7_75t_R FILLER_0_170_881 ();
 FILLER_ASAP7_75t_R FILLER_0_170_895 ();
 DECAPx2_ASAP7_75t_R FILLER_0_170_903 ();
 DECAPx1_ASAP7_75t_R FILLER_0_170_917 ();
 DECAPx10_ASAP7_75t_R FILLER_0_170_924 ();
 DECAPx10_ASAP7_75t_R FILLER_0_170_946 ();
 DECAPx4_ASAP7_75t_R FILLER_0_170_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_978 ();
 FILLER_ASAP7_75t_R FILLER_0_170_991 ();
 FILLER_ASAP7_75t_R FILLER_0_170_1005 ();
 DECAPx6_ASAP7_75t_R FILLER_0_170_1013 ();
 FILLER_ASAP7_75t_R FILLER_0_170_1027 ();
 DECAPx1_ASAP7_75t_R FILLER_0_170_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_1041 ();
 DECAPx2_ASAP7_75t_R FILLER_0_170_1052 ();
 FILLER_ASAP7_75t_R FILLER_0_170_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_1060 ();
 DECAPx4_ASAP7_75t_R FILLER_0_170_1065 ();
 FILLER_ASAP7_75t_R FILLER_0_170_1075 ();
 DECAPx10_ASAP7_75t_R FILLER_0_170_1087 ();
 DECAPx10_ASAP7_75t_R FILLER_0_170_1109 ();
 FILLER_ASAP7_75t_R FILLER_0_170_1131 ();
 DECAPx2_ASAP7_75t_R FILLER_0_170_1145 ();
 DECAPx6_ASAP7_75t_R FILLER_0_170_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_1170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_170_1174 ();
 DECAPx6_ASAP7_75t_R FILLER_0_170_1196 ();
 DECAPx2_ASAP7_75t_R FILLER_0_170_1216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_170_1225 ();
 DECAPx6_ASAP7_75t_R FILLER_0_170_1247 ();
 FILLER_ASAP7_75t_R FILLER_0_170_1261 ();
 FILLER_ASAP7_75t_R FILLER_0_170_1269 ();
 FILLER_ASAP7_75t_R FILLER_0_170_1276 ();
 DECAPx6_ASAP7_75t_R FILLER_0_170_1281 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_1295 ();
 DECAPx6_ASAP7_75t_R FILLER_0_170_1316 ();
 FILLER_ASAP7_75t_R FILLER_0_170_1333 ();
 FILLER_ASAP7_75t_R FILLER_0_170_1338 ();
 DECAPx1_ASAP7_75t_R FILLER_0_170_1345 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170_1349 ();
 DECAPx1_ASAP7_75t_R FILLER_0_170_1355 ();
 DECAPx1_ASAP7_75t_R FILLER_0_170_1364 ();
 FILLER_ASAP7_75t_R FILLER_0_170_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_170_1380 ();
 DECAPx2_ASAP7_75t_R FILLER_0_171_2 ();
 FILLER_ASAP7_75t_R FILLER_0_171_29 ();
 FILLER_ASAP7_75t_R FILLER_0_171_37 ();
 FILLER_ASAP7_75t_R FILLER_0_171_45 ();
 FILLER_ASAP7_75t_R FILLER_0_171_52 ();
 FILLER_ASAP7_75t_R FILLER_0_171_60 ();
 FILLER_ASAP7_75t_R FILLER_0_171_68 ();
 FILLER_ASAP7_75t_R FILLER_0_171_75 ();
 FILLER_ASAP7_75t_R FILLER_0_171_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_82 ();
 DECAPx1_ASAP7_75t_R FILLER_0_171_89 ();
 FILLER_ASAP7_75t_R FILLER_0_171_101 ();
 FILLER_ASAP7_75t_R FILLER_0_171_111 ();
 DECAPx10_ASAP7_75t_R FILLER_0_171_116 ();
 FILLER_ASAP7_75t_R FILLER_0_171_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_140 ();
 FILLER_ASAP7_75t_R FILLER_0_171_153 ();
 FILLER_ASAP7_75t_R FILLER_0_171_166 ();
 DECAPx4_ASAP7_75t_R FILLER_0_171_171 ();
 DECAPx4_ASAP7_75t_R FILLER_0_171_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_202 ();
 FILLER_ASAP7_75t_R FILLER_0_171_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_215 ();
 DECAPx10_ASAP7_75t_R FILLER_0_171_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_241 ();
 FILLER_ASAP7_75t_R FILLER_0_171_250 ();
 DECAPx2_ASAP7_75t_R FILLER_0_171_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_268 ();
 DECAPx2_ASAP7_75t_R FILLER_0_171_276 ();
 DECAPx1_ASAP7_75t_R FILLER_0_171_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_292 ();
 DECAPx2_ASAP7_75t_R FILLER_0_171_299 ();
 DECAPx4_ASAP7_75t_R FILLER_0_171_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_321 ();
 FILLER_ASAP7_75t_R FILLER_0_171_328 ();
 FILLER_ASAP7_75t_R FILLER_0_171_338 ();
 DECAPx2_ASAP7_75t_R FILLER_0_171_346 ();
 FILLER_ASAP7_75t_R FILLER_0_171_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_362 ();
 FILLER_ASAP7_75t_R FILLER_0_171_369 ();
 DECAPx6_ASAP7_75t_R FILLER_0_171_377 ();
 FILLER_ASAP7_75t_R FILLER_0_171_391 ();
 FILLER_ASAP7_75t_R FILLER_0_171_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_403 ();
 FILLER_ASAP7_75t_R FILLER_0_171_409 ();
 DECAPx2_ASAP7_75t_R FILLER_0_171_417 ();
 FILLER_ASAP7_75t_R FILLER_0_171_423 ();
 FILLER_ASAP7_75t_R FILLER_0_171_433 ();
 DECAPx10_ASAP7_75t_R FILLER_0_171_441 ();
 DECAPx6_ASAP7_75t_R FILLER_0_171_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_477 ();
 DECAPx4_ASAP7_75t_R FILLER_0_171_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_494 ();
 DECAPx2_ASAP7_75t_R FILLER_0_171_501 ();
 FILLER_ASAP7_75t_R FILLER_0_171_515 ();
 FILLER_ASAP7_75t_R FILLER_0_171_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_525 ();
 FILLER_ASAP7_75t_R FILLER_0_171_532 ();
 DECAPx1_ASAP7_75t_R FILLER_0_171_541 ();
 FILLER_ASAP7_75t_R FILLER_0_171_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_553 ();
 DECAPx1_ASAP7_75t_R FILLER_0_171_560 ();
 DECAPx6_ASAP7_75t_R FILLER_0_171_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_584 ();
 DECAPx4_ASAP7_75t_R FILLER_0_171_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_601 ();
 FILLER_ASAP7_75t_R FILLER_0_171_624 ();
 DECAPx1_ASAP7_75t_R FILLER_0_171_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_636 ();
 DECAPx10_ASAP7_75t_R FILLER_0_171_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_679 ();
 DECAPx4_ASAP7_75t_R FILLER_0_171_689 ();
 FILLER_ASAP7_75t_R FILLER_0_171_702 ();
 DECAPx2_ASAP7_75t_R FILLER_0_171_710 ();
 FILLER_ASAP7_75t_R FILLER_0_171_719 ();
 DECAPx4_ASAP7_75t_R FILLER_0_171_742 ();
 FILLER_ASAP7_75t_R FILLER_0_171_752 ();
 DECAPx6_ASAP7_75t_R FILLER_0_171_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_780 ();
 DECAPx10_ASAP7_75t_R FILLER_0_171_803 ();
 DECAPx10_ASAP7_75t_R FILLER_0_171_825 ();
 DECAPx4_ASAP7_75t_R FILLER_0_171_847 ();
 DECAPx2_ASAP7_75t_R FILLER_0_171_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_875 ();
 FILLER_ASAP7_75t_R FILLER_0_171_888 ();
 FILLER_ASAP7_75t_R FILLER_0_171_893 ();
 FILLER_ASAP7_75t_R FILLER_0_171_906 ();
 DECAPx4_ASAP7_75t_R FILLER_0_171_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_924 ();
 DECAPx6_ASAP7_75t_R FILLER_0_171_927 ();
 FILLER_ASAP7_75t_R FILLER_0_171_953 ();
 DECAPx4_ASAP7_75t_R FILLER_0_171_967 ();
 FILLER_ASAP7_75t_R FILLER_0_171_977 ();
 DECAPx2_ASAP7_75t_R FILLER_0_171_984 ();
 DECAPx6_ASAP7_75t_R FILLER_0_171_996 ();
 FILLER_ASAP7_75t_R FILLER_0_171_1010 ();
 FILLER_ASAP7_75t_R FILLER_0_171_1022 ();
 DECAPx2_ASAP7_75t_R FILLER_0_171_1034 ();
 FILLER_ASAP7_75t_R FILLER_0_171_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_1042 ();
 FILLER_ASAP7_75t_R FILLER_0_171_1053 ();
 DECAPx6_ASAP7_75t_R FILLER_0_171_1063 ();
 DECAPx2_ASAP7_75t_R FILLER_0_171_1083 ();
 FILLER_ASAP7_75t_R FILLER_0_171_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_1091 ();
 FILLER_ASAP7_75t_R FILLER_0_171_1102 ();
 FILLER_ASAP7_75t_R FILLER_0_171_1110 ();
 FILLER_ASAP7_75t_R FILLER_0_171_1122 ();
 DECAPx1_ASAP7_75t_R FILLER_0_171_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_1134 ();
 FILLER_ASAP7_75t_R FILLER_0_171_1145 ();
 DECAPx1_ASAP7_75t_R FILLER_0_171_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_1157 ();
 DECAPx4_ASAP7_75t_R FILLER_0_171_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_1174 ();
 FILLER_ASAP7_75t_R FILLER_0_171_1181 ();
 DECAPx4_ASAP7_75t_R FILLER_0_171_1191 ();
 DECAPx1_ASAP7_75t_R FILLER_0_171_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_1215 ();
 FILLER_ASAP7_75t_R FILLER_0_171_1222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_171_1235 ();
 DECAPx10_ASAP7_75t_R FILLER_0_171_1257 ();
 DECAPx4_ASAP7_75t_R FILLER_0_171_1279 ();
 FILLER_ASAP7_75t_R FILLER_0_171_1289 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_1291 ();
 FILLER_ASAP7_75t_R FILLER_0_171_1295 ();
 DECAPx1_ASAP7_75t_R FILLER_0_171_1300 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_171_1310 ();
 DECAPx2_ASAP7_75t_R FILLER_0_171_1332 ();
 FILLER_ASAP7_75t_R FILLER_0_171_1338 ();
 FILLER_ASAP7_75t_R FILLER_0_171_1345 ();
 FILLER_ASAP7_75t_R FILLER_0_171_1352 ();
 FILLER_ASAP7_75t_R FILLER_0_171_1359 ();
 FILLER_ASAP7_75t_R FILLER_0_171_1366 ();
 FILLER_ASAP7_75t_R FILLER_0_171_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_171_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_172_2 ();
 FILLER_ASAP7_75t_R FILLER_0_172_9 ();
 FILLER_ASAP7_75t_R FILLER_0_172_16 ();
 DECAPx1_ASAP7_75t_R FILLER_0_172_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172_27 ();
 FILLER_ASAP7_75t_R FILLER_0_172_49 ();
 DECAPx2_ASAP7_75t_R FILLER_0_172_58 ();
 FILLER_ASAP7_75t_R FILLER_0_172_70 ();
 FILLER_ASAP7_75t_R FILLER_0_172_77 ();
 FILLER_ASAP7_75t_R FILLER_0_172_91 ();
 DECAPx1_ASAP7_75t_R FILLER_0_172_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172_102 ();
 FILLER_ASAP7_75t_R FILLER_0_172_109 ();
 DECAPx6_ASAP7_75t_R FILLER_0_172_114 ();
 FILLER_ASAP7_75t_R FILLER_0_172_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172_136 ();
 DECAPx2_ASAP7_75t_R FILLER_0_172_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172_151 ();
 FILLER_ASAP7_75t_R FILLER_0_172_155 ();
 FILLER_ASAP7_75t_R FILLER_0_172_165 ();
 DECAPx2_ASAP7_75t_R FILLER_0_172_170 ();
 FILLER_ASAP7_75t_R FILLER_0_172_176 ();
 DECAPx4_ASAP7_75t_R FILLER_0_172_183 ();
 FILLER_ASAP7_75t_R FILLER_0_172_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172_195 ();
 DECAPx6_ASAP7_75t_R FILLER_0_172_204 ();
 DECAPx6_ASAP7_75t_R FILLER_0_172_230 ();
 DECAPx1_ASAP7_75t_R FILLER_0_172_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172_248 ();
 DECAPx4_ASAP7_75t_R FILLER_0_172_254 ();
 FILLER_ASAP7_75t_R FILLER_0_172_269 ();
 DECAPx2_ASAP7_75t_R FILLER_0_172_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172_281 ();
 FILLER_ASAP7_75t_R FILLER_0_172_288 ();
 DECAPx1_ASAP7_75t_R FILLER_0_172_296 ();
 FILLER_ASAP7_75t_R FILLER_0_172_306 ();
 DECAPx2_ASAP7_75t_R FILLER_0_172_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172_321 ();
 FILLER_ASAP7_75t_R FILLER_0_172_329 ();
 DECAPx4_ASAP7_75t_R FILLER_0_172_337 ();
 FILLER_ASAP7_75t_R FILLER_0_172_347 ();
 DECAPx4_ASAP7_75t_R FILLER_0_172_355 ();
 FILLER_ASAP7_75t_R FILLER_0_172_365 ();
 FILLER_ASAP7_75t_R FILLER_0_172_373 ();
 FILLER_ASAP7_75t_R FILLER_0_172_382 ();
 FILLER_ASAP7_75t_R FILLER_0_172_390 ();
 DECAPx2_ASAP7_75t_R FILLER_0_172_399 ();
 FILLER_ASAP7_75t_R FILLER_0_172_405 ();
 FILLER_ASAP7_75t_R FILLER_0_172_412 ();
 DECAPx2_ASAP7_75t_R FILLER_0_172_420 ();
 FILLER_ASAP7_75t_R FILLER_0_172_426 ();
 FILLER_ASAP7_75t_R FILLER_0_172_434 ();
 DECAPx6_ASAP7_75t_R FILLER_0_172_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_172_456 ();
 DECAPx4_ASAP7_75t_R FILLER_0_172_464 ();
 FILLER_ASAP7_75t_R FILLER_0_172_480 ();
 DECAPx2_ASAP7_75t_R FILLER_0_172_487 ();
 FILLER_ASAP7_75t_R FILLER_0_172_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172_495 ();
 DECAPx2_ASAP7_75t_R FILLER_0_172_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172_508 ();
 DECAPx2_ASAP7_75t_R FILLER_0_172_512 ();
 FILLER_ASAP7_75t_R FILLER_0_172_518 ();
 FILLER_ASAP7_75t_R FILLER_0_172_527 ();
 DECAPx6_ASAP7_75t_R FILLER_0_172_537 ();
 FILLER_ASAP7_75t_R FILLER_0_172_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172_559 ();
 DECAPx6_ASAP7_75t_R FILLER_0_172_563 ();
 FILLER_ASAP7_75t_R FILLER_0_172_583 ();
 DECAPx2_ASAP7_75t_R FILLER_0_172_593 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172_599 ();
 FILLER_ASAP7_75t_R FILLER_0_172_610 ();
 FILLER_ASAP7_75t_R FILLER_0_172_618 ();
 FILLER_ASAP7_75t_R FILLER_0_172_627 ();
 DECAPx6_ASAP7_75t_R FILLER_0_172_635 ();
 DECAPx1_ASAP7_75t_R FILLER_0_172_649 ();
 DECAPx10_ASAP7_75t_R FILLER_0_172_659 ();
 FILLER_ASAP7_75t_R FILLER_0_172_681 ();
 DECAPx2_ASAP7_75t_R FILLER_0_172_686 ();
 FILLER_ASAP7_75t_R FILLER_0_172_692 ();
 DECAPx4_ASAP7_75t_R FILLER_0_172_697 ();
 FILLER_ASAP7_75t_R FILLER_0_172_707 ();
 DECAPx1_ASAP7_75t_R FILLER_0_172_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172_719 ();
 FILLER_ASAP7_75t_R FILLER_0_172_726 ();
 FILLER_ASAP7_75t_R FILLER_0_172_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172_733 ();
 DECAPx10_ASAP7_75t_R FILLER_0_172_756 ();
 FILLER_ASAP7_75t_R FILLER_0_172_784 ();
 DECAPx1_ASAP7_75t_R FILLER_0_172_789 ();
 DECAPx10_ASAP7_75t_R FILLER_0_172_814 ();
 DECAPx1_ASAP7_75t_R FILLER_0_172_836 ();
 FILLER_ASAP7_75t_R FILLER_0_172_852 ();
 FILLER_ASAP7_75t_R FILLER_0_172_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172_862 ();
 FILLER_ASAP7_75t_R FILLER_0_172_874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_172_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172_910 ();
 DECAPx4_ASAP7_75t_R FILLER_0_172_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172_942 ();
 DECAPx1_ASAP7_75t_R FILLER_0_172_954 ();
 FILLER_ASAP7_75t_R FILLER_0_172_979 ();
 FILLER_ASAP7_75t_R FILLER_0_172_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172_986 ();
 FILLER_ASAP7_75t_R FILLER_0_172_993 ();
 DECAPx2_ASAP7_75t_R FILLER_0_172_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172_1009 ();
 DECAPx2_ASAP7_75t_R FILLER_0_172_1021 ();
 DECAPx10_ASAP7_75t_R FILLER_0_172_1047 ();
 DECAPx4_ASAP7_75t_R FILLER_0_172_1069 ();
 FILLER_ASAP7_75t_R FILLER_0_172_1079 ();
 FILLER_ASAP7_75t_R FILLER_0_172_1091 ();
 FILLER_ASAP7_75t_R FILLER_0_172_1103 ();
 DECAPx4_ASAP7_75t_R FILLER_0_172_1111 ();
 FILLER_ASAP7_75t_R FILLER_0_172_1124 ();
 FILLER_ASAP7_75t_R FILLER_0_172_1132 ();
 DECAPx4_ASAP7_75t_R FILLER_0_172_1140 ();
 FILLER_ASAP7_75t_R FILLER_0_172_1150 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172_1152 ();
 FILLER_ASAP7_75t_R FILLER_0_172_1164 ();
 DECAPx1_ASAP7_75t_R FILLER_0_172_1172 ();
 DECAPx1_ASAP7_75t_R FILLER_0_172_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172_1185 ();
 DECAPx6_ASAP7_75t_R FILLER_0_172_1192 ();
 DECAPx1_ASAP7_75t_R FILLER_0_172_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172_1210 ();
 DECAPx2_ASAP7_75t_R FILLER_0_172_1222 ();
 DECAPx6_ASAP7_75t_R FILLER_0_172_1234 ();
 DECAPx2_ASAP7_75t_R FILLER_0_172_1248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_172_1274 ();
 DECAPx2_ASAP7_75t_R FILLER_0_172_1296 ();
 FILLER_ASAP7_75t_R FILLER_0_172_1302 ();
 FILLER_ASAP7_75t_R FILLER_0_172_1314 ();
 DECAPx1_ASAP7_75t_R FILLER_0_172_1338 ();
 FILLER_ASAP7_75t_R FILLER_0_172_1345 ();
 FILLER_ASAP7_75t_R FILLER_0_172_1350 ();
 FILLER_ASAP7_75t_R FILLER_0_172_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_172_1364 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172_1366 ();
 FILLER_ASAP7_75t_R FILLER_0_172_1372 ();
 FILLER_ASAP7_75t_R FILLER_0_172_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_173_2 ();
 FILLER_ASAP7_75t_R FILLER_0_173_9 ();
 DECAPx2_ASAP7_75t_R FILLER_0_173_16 ();
 FILLER_ASAP7_75t_R FILLER_0_173_27 ();
 DECAPx1_ASAP7_75t_R FILLER_0_173_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173_38 ();
 FILLER_ASAP7_75t_R FILLER_0_173_45 ();
 FILLER_ASAP7_75t_R FILLER_0_173_52 ();
 FILLER_ASAP7_75t_R FILLER_0_173_75 ();
 FILLER_ASAP7_75t_R FILLER_0_173_82 ();
 FILLER_ASAP7_75t_R FILLER_0_173_87 ();
 FILLER_ASAP7_75t_R FILLER_0_173_99 ();
 FILLER_ASAP7_75t_R FILLER_0_173_105 ();
 DECAPx2_ASAP7_75t_R FILLER_0_173_110 ();
 DECAPx2_ASAP7_75t_R FILLER_0_173_120 ();
 FILLER_ASAP7_75t_R FILLER_0_173_132 ();
 DECAPx6_ASAP7_75t_R FILLER_0_173_142 ();
 FILLER_ASAP7_75t_R FILLER_0_173_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173_158 ();
 DECAPx4_ASAP7_75t_R FILLER_0_173_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173_180 ();
 DECAPx2_ASAP7_75t_R FILLER_0_173_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173_192 ();
 FILLER_ASAP7_75t_R FILLER_0_173_201 ();
 FILLER_ASAP7_75t_R FILLER_0_173_213 ();
 DECAPx6_ASAP7_75t_R FILLER_0_173_220 ();
 FILLER_ASAP7_75t_R FILLER_0_173_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173_236 ();
 DECAPx2_ASAP7_75t_R FILLER_0_173_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173_281 ();
 FILLER_ASAP7_75t_R FILLER_0_173_289 ();
 DECAPx1_ASAP7_75t_R FILLER_0_173_301 ();
 DECAPx2_ASAP7_75t_R FILLER_0_173_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173_317 ();
 DECAPx1_ASAP7_75t_R FILLER_0_173_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173_328 ();
 DECAPx6_ASAP7_75t_R FILLER_0_173_335 ();
 DECAPx1_ASAP7_75t_R FILLER_0_173_349 ();
 DECAPx2_ASAP7_75t_R FILLER_0_173_359 ();
 FILLER_ASAP7_75t_R FILLER_0_173_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173_367 ();
 DECAPx4_ASAP7_75t_R FILLER_0_173_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173_381 ();
 FILLER_ASAP7_75t_R FILLER_0_173_387 ();
 FILLER_ASAP7_75t_R FILLER_0_173_409 ();
 FILLER_ASAP7_75t_R FILLER_0_173_437 ();
 DECAPx2_ASAP7_75t_R FILLER_0_173_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173_451 ();
 DECAPx2_ASAP7_75t_R FILLER_0_173_462 ();
 FILLER_ASAP7_75t_R FILLER_0_173_468 ();
 DECAPx1_ASAP7_75t_R FILLER_0_173_480 ();
 FILLER_ASAP7_75t_R FILLER_0_173_490 ();
 DECAPx1_ASAP7_75t_R FILLER_0_173_499 ();
 FILLER_ASAP7_75t_R FILLER_0_173_511 ();
 DECAPx2_ASAP7_75t_R FILLER_0_173_519 ();
 FILLER_ASAP7_75t_R FILLER_0_173_525 ();
 FILLER_ASAP7_75t_R FILLER_0_173_533 ();
 DECAPx6_ASAP7_75t_R FILLER_0_173_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173_552 ();
 DECAPx4_ASAP7_75t_R FILLER_0_173_567 ();
 FILLER_ASAP7_75t_R FILLER_0_173_583 ();
 FILLER_ASAP7_75t_R FILLER_0_173_591 ();
 DECAPx6_ASAP7_75t_R FILLER_0_173_599 ();
 FILLER_ASAP7_75t_R FILLER_0_173_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173_615 ();
 DECAPx1_ASAP7_75t_R FILLER_0_173_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173_628 ();
 DECAPx2_ASAP7_75t_R FILLER_0_173_632 ();
 FILLER_ASAP7_75t_R FILLER_0_173_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_173_647 ();
 DECAPx6_ASAP7_75t_R FILLER_0_173_669 ();
 FILLER_ASAP7_75t_R FILLER_0_173_683 ();
 FILLER_ASAP7_75t_R FILLER_0_173_691 ();
 FILLER_ASAP7_75t_R FILLER_0_173_699 ();
 DECAPx10_ASAP7_75t_R FILLER_0_173_707 ();
 DECAPx6_ASAP7_75t_R FILLER_0_173_729 ();
 DECAPx2_ASAP7_75t_R FILLER_0_173_743 ();
 FILLER_ASAP7_75t_R FILLER_0_173_752 ();
 FILLER_ASAP7_75t_R FILLER_0_173_766 ();
 FILLER_ASAP7_75t_R FILLER_0_173_780 ();
 FILLER_ASAP7_75t_R FILLER_0_173_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173_790 ();
 DECAPx2_ASAP7_75t_R FILLER_0_173_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173_804 ();
 FILLER_ASAP7_75t_R FILLER_0_173_811 ();
 DECAPx6_ASAP7_75t_R FILLER_0_173_816 ();
 FILLER_ASAP7_75t_R FILLER_0_173_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173_832 ();
 FILLER_ASAP7_75t_R FILLER_0_173_855 ();
 DECAPx2_ASAP7_75t_R FILLER_0_173_863 ();
 FILLER_ASAP7_75t_R FILLER_0_173_877 ();
 FILLER_ASAP7_75t_R FILLER_0_173_891 ();
 DECAPx2_ASAP7_75t_R FILLER_0_173_904 ();
 FILLER_ASAP7_75t_R FILLER_0_173_918 ();
 FILLER_ASAP7_75t_R FILLER_0_173_923 ();
 DECAPx2_ASAP7_75t_R FILLER_0_173_927 ();
 FILLER_ASAP7_75t_R FILLER_0_173_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173_935 ();
 FILLER_ASAP7_75t_R FILLER_0_173_942 ();
 DECAPx2_ASAP7_75t_R FILLER_0_173_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173_962 ();
 DECAPx1_ASAP7_75t_R FILLER_0_173_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173_975 ();
 DECAPx10_ASAP7_75t_R FILLER_0_173_997 ();
 DECAPx4_ASAP7_75t_R FILLER_0_173_1019 ();
 DECAPx10_ASAP7_75t_R FILLER_0_173_1039 ();
 FILLER_ASAP7_75t_R FILLER_0_173_1069 ();
 DECAPx2_ASAP7_75t_R FILLER_0_173_1077 ();
 FILLER_ASAP7_75t_R FILLER_0_173_1083 ();
 DECAPx4_ASAP7_75t_R FILLER_0_173_1091 ();
 FILLER_ASAP7_75t_R FILLER_0_173_1101 ();
 DECAPx10_ASAP7_75t_R FILLER_0_173_1109 ();
 DECAPx4_ASAP7_75t_R FILLER_0_173_1131 ();
 FILLER_ASAP7_75t_R FILLER_0_173_1141 ();
 FILLER_ASAP7_75t_R FILLER_0_173_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173_1151 ();
 DECAPx1_ASAP7_75t_R FILLER_0_173_1157 ();
 FILLER_ASAP7_75t_R FILLER_0_173_1167 ();
 DECAPx2_ASAP7_75t_R FILLER_0_173_1175 ();
 FILLER_ASAP7_75t_R FILLER_0_173_1181 ();
 DECAPx2_ASAP7_75t_R FILLER_0_173_1188 ();
 FILLER_ASAP7_75t_R FILLER_0_173_1194 ();
 FILLER_ASAP7_75t_R FILLER_0_173_1202 ();
 FILLER_ASAP7_75t_R FILLER_0_173_1210 ();
 DECAPx2_ASAP7_75t_R FILLER_0_173_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173_1225 ();
 FILLER_ASAP7_75t_R FILLER_0_173_1242 ();
 DECAPx10_ASAP7_75t_R FILLER_0_173_1264 ();
 DECAPx4_ASAP7_75t_R FILLER_0_173_1286 ();
 DECAPx6_ASAP7_75t_R FILLER_0_173_1302 ();
 FILLER_ASAP7_75t_R FILLER_0_173_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_173_1321 ();
 DECAPx4_ASAP7_75t_R FILLER_0_173_1343 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173_1353 ();
 FILLER_ASAP7_75t_R FILLER_0_173_1359 ();
 FILLER_ASAP7_75t_R FILLER_0_173_1366 ();
 FILLER_ASAP7_75t_R FILLER_0_173_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_173_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_174_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_174_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_29 ();
 FILLER_ASAP7_75t_R FILLER_0_174_36 ();
 FILLER_ASAP7_75t_R FILLER_0_174_59 ();
 FILLER_ASAP7_75t_R FILLER_0_174_66 ();
 FILLER_ASAP7_75t_R FILLER_0_174_73 ();
 FILLER_ASAP7_75t_R FILLER_0_174_80 ();
 FILLER_ASAP7_75t_R FILLER_0_174_87 ();
 FILLER_ASAP7_75t_R FILLER_0_174_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_96 ();
 DECAPx2_ASAP7_75t_R FILLER_0_174_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_115 ();
 DECAPx2_ASAP7_75t_R FILLER_0_174_122 ();
 FILLER_ASAP7_75t_R FILLER_0_174_128 ();
 DECAPx1_ASAP7_75t_R FILLER_0_174_135 ();
 DECAPx6_ASAP7_75t_R FILLER_0_174_145 ();
 DECAPx2_ASAP7_75t_R FILLER_0_174_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_165 ();
 FILLER_ASAP7_75t_R FILLER_0_174_169 ();
 DECAPx1_ASAP7_75t_R FILLER_0_174_179 ();
 FILLER_ASAP7_75t_R FILLER_0_174_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_195 ();
 DECAPx10_ASAP7_75t_R FILLER_0_174_204 ();
 DECAPx1_ASAP7_75t_R FILLER_0_174_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_230 ();
 FILLER_ASAP7_75t_R FILLER_0_174_252 ();
 DECAPx2_ASAP7_75t_R FILLER_0_174_265 ();
 FILLER_ASAP7_75t_R FILLER_0_174_271 ();
 FILLER_ASAP7_75t_R FILLER_0_174_279 ();
 DECAPx2_ASAP7_75t_R FILLER_0_174_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_293 ();
 FILLER_ASAP7_75t_R FILLER_0_174_300 ();
 FILLER_ASAP7_75t_R FILLER_0_174_307 ();
 DECAPx2_ASAP7_75t_R FILLER_0_174_313 ();
 FILLER_ASAP7_75t_R FILLER_0_174_319 ();
 FILLER_ASAP7_75t_R FILLER_0_174_328 ();
 FILLER_ASAP7_75t_R FILLER_0_174_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_339 ();
 DECAPx1_ASAP7_75t_R FILLER_0_174_346 ();
 DECAPx6_ASAP7_75t_R FILLER_0_174_370 ();
 FILLER_ASAP7_75t_R FILLER_0_174_390 ();
 DECAPx1_ASAP7_75t_R FILLER_0_174_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_399 ();
 FILLER_ASAP7_75t_R FILLER_0_174_406 ();
 FILLER_ASAP7_75t_R FILLER_0_174_414 ();
 FILLER_ASAP7_75t_R FILLER_0_174_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_424 ();
 FILLER_ASAP7_75t_R FILLER_0_174_431 ();
 FILLER_ASAP7_75t_R FILLER_0_174_439 ();
 DECAPx4_ASAP7_75t_R FILLER_0_174_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_454 ();
 FILLER_ASAP7_75t_R FILLER_0_174_460 ();
 FILLER_ASAP7_75t_R FILLER_0_174_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_466 ();
 FILLER_ASAP7_75t_R FILLER_0_174_477 ();
 FILLER_ASAP7_75t_R FILLER_0_174_484 ();
 DECAPx2_ASAP7_75t_R FILLER_0_174_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_502 ();
 FILLER_ASAP7_75t_R FILLER_0_174_509 ();
 FILLER_ASAP7_75t_R FILLER_0_174_517 ();
 DECAPx2_ASAP7_75t_R FILLER_0_174_525 ();
 FILLER_ASAP7_75t_R FILLER_0_174_538 ();
 DECAPx1_ASAP7_75t_R FILLER_0_174_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_550 ();
 DECAPx2_ASAP7_75t_R FILLER_0_174_561 ();
 FILLER_ASAP7_75t_R FILLER_0_174_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_569 ();
 DECAPx6_ASAP7_75t_R FILLER_0_174_580 ();
 DECAPx1_ASAP7_75t_R FILLER_0_174_594 ();
 FILLER_ASAP7_75t_R FILLER_0_174_606 ();
 DECAPx4_ASAP7_75t_R FILLER_0_174_614 ();
 FILLER_ASAP7_75t_R FILLER_0_174_628 ();
 FILLER_ASAP7_75t_R FILLER_0_174_636 ();
 FILLER_ASAP7_75t_R FILLER_0_174_646 ();
 FILLER_ASAP7_75t_R FILLER_0_174_654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_174_662 ();
 DECAPx4_ASAP7_75t_R FILLER_0_174_687 ();
 FILLER_ASAP7_75t_R FILLER_0_174_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_699 ();
 DECAPx2_ASAP7_75t_R FILLER_0_174_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_174_733 ();
 DECAPx2_ASAP7_75t_R FILLER_0_174_755 ();
 FILLER_ASAP7_75t_R FILLER_0_174_773 ();
 FILLER_ASAP7_75t_R FILLER_0_174_787 ();
 DECAPx2_ASAP7_75t_R FILLER_0_174_795 ();
 FILLER_ASAP7_75t_R FILLER_0_174_801 ();
 DECAPx4_ASAP7_75t_R FILLER_0_174_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_834 ();
 FILLER_ASAP7_75t_R FILLER_0_174_857 ();
 FILLER_ASAP7_75t_R FILLER_0_174_875 ();
 DECAPx6_ASAP7_75t_R FILLER_0_174_880 ();
 FILLER_ASAP7_75t_R FILLER_0_174_894 ();
 DECAPx1_ASAP7_75t_R FILLER_0_174_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_906 ();
 DECAPx2_ASAP7_75t_R FILLER_0_174_928 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_934 ();
 DECAPx1_ASAP7_75t_R FILLER_0_174_957 ();
 DECAPx2_ASAP7_75t_R FILLER_0_174_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_989 ();
 DECAPx2_ASAP7_75t_R FILLER_0_174_998 ();
 DECAPx2_ASAP7_75t_R FILLER_0_174_1025 ();
 DECAPx6_ASAP7_75t_R FILLER_0_174_1041 ();
 DECAPx4_ASAP7_75t_R FILLER_0_174_1067 ();
 FILLER_ASAP7_75t_R FILLER_0_174_1077 ();
 FILLER_ASAP7_75t_R FILLER_0_174_1085 ();
 FILLER_ASAP7_75t_R FILLER_0_174_1093 ();
 FILLER_ASAP7_75t_R FILLER_0_174_1101 ();
 DECAPx2_ASAP7_75t_R FILLER_0_174_1109 ();
 FILLER_ASAP7_75t_R FILLER_0_174_1115 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_1117 ();
 FILLER_ASAP7_75t_R FILLER_0_174_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_1126 ();
 FILLER_ASAP7_75t_R FILLER_0_174_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_1135 ();
 FILLER_ASAP7_75t_R FILLER_0_174_1142 ();
 DECAPx4_ASAP7_75t_R FILLER_0_174_1150 ();
 FILLER_ASAP7_75t_R FILLER_0_174_1160 ();
 DECAPx4_ASAP7_75t_R FILLER_0_174_1173 ();
 FILLER_ASAP7_75t_R FILLER_0_174_1189 ();
 FILLER_ASAP7_75t_R FILLER_0_174_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_1198 ();
 FILLER_ASAP7_75t_R FILLER_0_174_1205 ();
 DECAPx2_ASAP7_75t_R FILLER_0_174_1212 ();
 FILLER_ASAP7_75t_R FILLER_0_174_1218 ();
 DECAPx6_ASAP7_75t_R FILLER_0_174_1226 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_1240 ();
 FILLER_ASAP7_75t_R FILLER_0_174_1257 ();
 DECAPx10_ASAP7_75t_R FILLER_0_174_1269 ();
 DECAPx10_ASAP7_75t_R FILLER_0_174_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_0_174_1313 ();
 DECAPx6_ASAP7_75t_R FILLER_0_174_1335 ();
 FILLER_ASAP7_75t_R FILLER_0_174_1349 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_1351 ();
 FILLER_ASAP7_75t_R FILLER_0_174_1356 ();
 DECAPx1_ASAP7_75t_R FILLER_0_174_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174_1367 ();
 FILLER_ASAP7_75t_R FILLER_0_174_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_174_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_175_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_175_4 ();
 FILLER_ASAP7_75t_R FILLER_0_175_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_175_28 ();
 FILLER_ASAP7_75t_R FILLER_0_175_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_175_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_175_44 ();
 FILLER_ASAP7_75t_R FILLER_0_175_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_175_58 ();
 FILLER_ASAP7_75t_R FILLER_0_175_65 ();
 FILLER_ASAP7_75t_R FILLER_0_175_72 ();
 FILLER_ASAP7_75t_R FILLER_0_175_79 ();
 FILLER_ASAP7_75t_R FILLER_0_175_86 ();
 DECAPx1_ASAP7_75t_R FILLER_0_175_93 ();
 DECAPx1_ASAP7_75t_R FILLER_0_175_109 ();
 FILLER_ASAP7_75t_R FILLER_0_175_119 ();
 DECAPx10_ASAP7_75t_R FILLER_0_175_127 ();
 DECAPx4_ASAP7_75t_R FILLER_0_175_149 ();
 FILLER_ASAP7_75t_R FILLER_0_175_159 ();
 DECAPx4_ASAP7_75t_R FILLER_0_175_169 ();
 FILLER_ASAP7_75t_R FILLER_0_175_191 ();
 FILLER_ASAP7_75t_R FILLER_0_175_196 ();
 DECAPx10_ASAP7_75t_R FILLER_0_175_204 ();
 FILLER_ASAP7_75t_R FILLER_0_175_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_175_228 ();
 FILLER_ASAP7_75t_R FILLER_0_175_237 ();
 DECAPx2_ASAP7_75t_R FILLER_0_175_242 ();
 DECAPx6_ASAP7_75t_R FILLER_0_175_260 ();
 FILLER_ASAP7_75t_R FILLER_0_175_280 ();
 DECAPx2_ASAP7_75t_R FILLER_0_175_288 ();
 FILLER_ASAP7_75t_R FILLER_0_175_294 ();
 DECAPx6_ASAP7_75t_R FILLER_0_175_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_175_316 ();
 DECAPx2_ASAP7_75t_R FILLER_0_175_323 ();
 FILLER_ASAP7_75t_R FILLER_0_175_335 ();
 DECAPx2_ASAP7_75t_R FILLER_0_175_340 ();
 FILLER_ASAP7_75t_R FILLER_0_175_346 ();
 FILLER_ASAP7_75t_R FILLER_0_175_354 ();
 DECAPx1_ASAP7_75t_R FILLER_0_175_359 ();
 FILLER_ASAP7_75t_R FILLER_0_175_369 ();
 DECAPx6_ASAP7_75t_R FILLER_0_175_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_175_391 ();
 DECAPx1_ASAP7_75t_R FILLER_0_175_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_175_402 ();
 DECAPx2_ASAP7_75t_R FILLER_0_175_410 ();
 FILLER_ASAP7_75t_R FILLER_0_175_416 ();
 FILLER_ASAP7_75t_R FILLER_0_175_424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_175_433 ();
 DECAPx6_ASAP7_75t_R FILLER_0_175_467 ();
 DECAPx1_ASAP7_75t_R FILLER_0_175_481 ();
 FILLER_ASAP7_75t_R FILLER_0_175_490 ();
 FILLER_ASAP7_75t_R FILLER_0_175_499 ();
 FILLER_ASAP7_75t_R FILLER_0_175_509 ();
 FILLER_ASAP7_75t_R FILLER_0_175_521 ();
 FILLER_ASAP7_75t_R FILLER_0_175_529 ();
 DECAPx1_ASAP7_75t_R FILLER_0_175_536 ();
 FILLER_ASAP7_75t_R FILLER_0_175_548 ();
 DECAPx1_ASAP7_75t_R FILLER_0_175_553 ();
 FILLER_ASAP7_75t_R FILLER_0_175_567 ();
 DECAPx10_ASAP7_75t_R FILLER_0_175_579 ();
 DECAPx6_ASAP7_75t_R FILLER_0_175_607 ();
 FILLER_ASAP7_75t_R FILLER_0_175_621 ();
 FILLER_ASAP7_75t_R FILLER_0_175_629 ();
 DECAPx2_ASAP7_75t_R FILLER_0_175_638 ();
 DECAPx1_ASAP7_75t_R FILLER_0_175_650 ();
 FILLER_ASAP7_75t_R FILLER_0_175_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_175_664 ();
 DECAPx2_ASAP7_75t_R FILLER_0_175_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_175_677 ();
 DECAPx2_ASAP7_75t_R FILLER_0_175_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_175_690 ();
 FILLER_ASAP7_75t_R FILLER_0_175_713 ();
 DECAPx6_ASAP7_75t_R FILLER_0_175_718 ();
 FILLER_ASAP7_75t_R FILLER_0_175_732 ();
 FILLER_ASAP7_75t_R FILLER_0_175_738 ();
 DECAPx1_ASAP7_75t_R FILLER_0_175_748 ();
 DECAPx6_ASAP7_75t_R FILLER_0_175_764 ();
 DECAPx2_ASAP7_75t_R FILLER_0_175_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_175_784 ();
 FILLER_ASAP7_75t_R FILLER_0_175_795 ();
 FILLER_ASAP7_75t_R FILLER_0_175_807 ();
 FILLER_ASAP7_75t_R FILLER_0_175_815 ();
 FILLER_ASAP7_75t_R FILLER_0_175_823 ();
 DECAPx2_ASAP7_75t_R FILLER_0_175_828 ();
 FILLER_ASAP7_75t_R FILLER_0_175_834 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_175_836 ();
 DECAPx2_ASAP7_75t_R FILLER_0_175_840 ();
 FILLER_ASAP7_75t_R FILLER_0_175_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_175_848 ();
 FILLER_ASAP7_75t_R FILLER_0_175_854 ();
 FILLER_ASAP7_75t_R FILLER_0_175_866 ();
 FILLER_ASAP7_75t_R FILLER_0_175_871 ();
 FILLER_ASAP7_75t_R FILLER_0_175_876 ();
 DECAPx2_ASAP7_75t_R FILLER_0_175_908 ();
 FILLER_ASAP7_75t_R FILLER_0_175_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_175_924 ();
 DECAPx2_ASAP7_75t_R FILLER_0_175_927 ();
 DECAPx2_ASAP7_75t_R FILLER_0_175_955 ();
 FILLER_ASAP7_75t_R FILLER_0_175_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_175_963 ();
 DECAPx4_ASAP7_75t_R FILLER_0_175_972 ();
 FILLER_ASAP7_75t_R FILLER_0_175_994 ();
 FILLER_ASAP7_75t_R FILLER_0_175_999 ();
 FILLER_ASAP7_75t_R FILLER_0_175_1009 ();
 DECAPx2_ASAP7_75t_R FILLER_0_175_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_175_1023 ();
 DECAPx2_ASAP7_75t_R FILLER_0_175_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_175_1036 ();
 FILLER_ASAP7_75t_R FILLER_0_175_1040 ();
 DECAPx2_ASAP7_75t_R FILLER_0_175_1052 ();
 FILLER_ASAP7_75t_R FILLER_0_175_1058 ();
 DECAPx4_ASAP7_75t_R FILLER_0_175_1066 ();
 FILLER_ASAP7_75t_R FILLER_0_175_1076 ();
 FILLER_ASAP7_75t_R FILLER_0_175_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_175_1086 ();
 DECAPx2_ASAP7_75t_R FILLER_0_175_1093 ();
 FILLER_ASAP7_75t_R FILLER_0_175_1099 ();
 FILLER_ASAP7_75t_R FILLER_0_175_1112 ();
 FILLER_ASAP7_75t_R FILLER_0_175_1120 ();
 FILLER_ASAP7_75t_R FILLER_0_175_1128 ();
 FILLER_ASAP7_75t_R FILLER_0_175_1136 ();
 DECAPx1_ASAP7_75t_R FILLER_0_175_1144 ();
 FILLER_ASAP7_75t_R FILLER_0_175_1170 ();
 FILLER_ASAP7_75t_R FILLER_0_175_1177 ();
 FILLER_ASAP7_75t_R FILLER_0_175_1184 ();
 FILLER_ASAP7_75t_R FILLER_0_175_1192 ();
 FILLER_ASAP7_75t_R FILLER_0_175_1199 ();
 FILLER_ASAP7_75t_R FILLER_0_175_1207 ();
 FILLER_ASAP7_75t_R FILLER_0_175_1216 ();
 FILLER_ASAP7_75t_R FILLER_0_175_1224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_175_1232 ();
 DECAPx2_ASAP7_75t_R FILLER_0_175_1254 ();
 FILLER_ASAP7_75t_R FILLER_0_175_1260 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_175_1262 ();
 FILLER_ASAP7_75t_R FILLER_0_175_1269 ();
 FILLER_ASAP7_75t_R FILLER_0_175_1277 ();
 DECAPx10_ASAP7_75t_R FILLER_0_175_1285 ();
 DECAPx10_ASAP7_75t_R FILLER_0_175_1307 ();
 DECAPx10_ASAP7_75t_R FILLER_0_175_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_0_175_1351 ();
 FILLER_ASAP7_75t_R FILLER_0_175_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_175_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_176_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_4 ();
 FILLER_ASAP7_75t_R FILLER_0_176_8 ();
 DECAPx1_ASAP7_75t_R FILLER_0_176_15 ();
 FILLER_ASAP7_75t_R FILLER_0_176_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_27 ();
 FILLER_ASAP7_75t_R FILLER_0_176_49 ();
 FILLER_ASAP7_75t_R FILLER_0_176_56 ();
 FILLER_ASAP7_75t_R FILLER_0_176_63 ();
 DECAPx1_ASAP7_75t_R FILLER_0_176_70 ();
 DECAPx1_ASAP7_75t_R FILLER_0_176_79 ();
 FILLER_ASAP7_75t_R FILLER_0_176_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_93 ();
 FILLER_ASAP7_75t_R FILLER_0_176_105 ();
 DECAPx1_ASAP7_75t_R FILLER_0_176_117 ();
 DECAPx1_ASAP7_75t_R FILLER_0_176_129 ();
 DECAPx6_ASAP7_75t_R FILLER_0_176_137 ();
 FILLER_ASAP7_75t_R FILLER_0_176_151 ();
 DECAPx6_ASAP7_75t_R FILLER_0_176_174 ();
 FILLER_ASAP7_75t_R FILLER_0_176_188 ();
 FILLER_ASAP7_75t_R FILLER_0_176_211 ();
 DECAPx1_ASAP7_75t_R FILLER_0_176_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_229 ();
 DECAPx2_ASAP7_75t_R FILLER_0_176_238 ();
 FILLER_ASAP7_75t_R FILLER_0_176_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_246 ();
 DECAPx4_ASAP7_75t_R FILLER_0_176_259 ();
 FILLER_ASAP7_75t_R FILLER_0_176_269 ();
 DECAPx1_ASAP7_75t_R FILLER_0_176_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_281 ();
 DECAPx4_ASAP7_75t_R FILLER_0_176_304 ();
 FILLER_ASAP7_75t_R FILLER_0_176_320 ();
 FILLER_ASAP7_75t_R FILLER_0_176_328 ();
 FILLER_ASAP7_75t_R FILLER_0_176_336 ();
 FILLER_ASAP7_75t_R FILLER_0_176_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_348 ();
 DECAPx2_ASAP7_75t_R FILLER_0_176_355 ();
 FILLER_ASAP7_75t_R FILLER_0_176_361 ();
 FILLER_ASAP7_75t_R FILLER_0_176_369 ();
 DECAPx2_ASAP7_75t_R FILLER_0_176_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_385 ();
 DECAPx1_ASAP7_75t_R FILLER_0_176_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_396 ();
 FILLER_ASAP7_75t_R FILLER_0_176_403 ();
 FILLER_ASAP7_75t_R FILLER_0_176_411 ();
 DECAPx2_ASAP7_75t_R FILLER_0_176_421 ();
 DECAPx1_ASAP7_75t_R FILLER_0_176_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_437 ();
 FILLER_ASAP7_75t_R FILLER_0_176_441 ();
 DECAPx4_ASAP7_75t_R FILLER_0_176_449 ();
 FILLER_ASAP7_75t_R FILLER_0_176_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_461 ();
 DECAPx1_ASAP7_75t_R FILLER_0_176_464 ();
 FILLER_ASAP7_75t_R FILLER_0_176_478 ();
 FILLER_ASAP7_75t_R FILLER_0_176_490 ();
 FILLER_ASAP7_75t_R FILLER_0_176_496 ();
 DECAPx1_ASAP7_75t_R FILLER_0_176_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_512 ();
 FILLER_ASAP7_75t_R FILLER_0_176_523 ();
 DECAPx1_ASAP7_75t_R FILLER_0_176_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_534 ();
 DECAPx2_ASAP7_75t_R FILLER_0_176_541 ();
 DECAPx2_ASAP7_75t_R FILLER_0_176_553 ();
 FILLER_ASAP7_75t_R FILLER_0_176_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_561 ();
 DECAPx4_ASAP7_75t_R FILLER_0_176_572 ();
 FILLER_ASAP7_75t_R FILLER_0_176_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_584 ();
 DECAPx4_ASAP7_75t_R FILLER_0_176_588 ();
 FILLER_ASAP7_75t_R FILLER_0_176_604 ();
 FILLER_ASAP7_75t_R FILLER_0_176_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_614 ();
 FILLER_ASAP7_75t_R FILLER_0_176_622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_176_630 ();
 FILLER_ASAP7_75t_R FILLER_0_176_652 ();
 FILLER_ASAP7_75t_R FILLER_0_176_660 ();
 FILLER_ASAP7_75t_R FILLER_0_176_682 ();
 FILLER_ASAP7_75t_R FILLER_0_176_694 ();
 FILLER_ASAP7_75t_R FILLER_0_176_702 ();
 DECAPx10_ASAP7_75t_R FILLER_0_176_710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_176_743 ();
 DECAPx2_ASAP7_75t_R FILLER_0_176_765 ();
 FILLER_ASAP7_75t_R FILLER_0_176_771 ();
 DECAPx1_ASAP7_75t_R FILLER_0_176_777 ();
 FILLER_ASAP7_75t_R FILLER_0_176_791 ();
 FILLER_ASAP7_75t_R FILLER_0_176_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_799 ();
 FILLER_ASAP7_75t_R FILLER_0_176_818 ();
 FILLER_ASAP7_75t_R FILLER_0_176_826 ();
 FILLER_ASAP7_75t_R FILLER_0_176_834 ();
 DECAPx1_ASAP7_75t_R FILLER_0_176_842 ();
 DECAPx1_ASAP7_75t_R FILLER_0_176_851 ();
 DECAPx10_ASAP7_75t_R FILLER_0_176_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_889 ();
 FILLER_ASAP7_75t_R FILLER_0_176_928 ();
 DECAPx1_ASAP7_75t_R FILLER_0_176_936 ();
 FILLER_ASAP7_75t_R FILLER_0_176_952 ();
 FILLER_ASAP7_75t_R FILLER_0_176_968 ();
 FILLER_ASAP7_75t_R FILLER_0_176_978 ();
 DECAPx2_ASAP7_75t_R FILLER_0_176_987 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_993 ();
 DECAPx1_ASAP7_75t_R FILLER_0_176_1006 ();
 FILLER_ASAP7_75t_R FILLER_0_176_1015 ();
 DECAPx2_ASAP7_75t_R FILLER_0_176_1020 ();
 FILLER_ASAP7_75t_R FILLER_0_176_1029 ();
 FILLER_ASAP7_75t_R FILLER_0_176_1037 ();
 DECAPx1_ASAP7_75t_R FILLER_0_176_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_1049 ();
 FILLER_ASAP7_75t_R FILLER_0_176_1058 ();
 DECAPx4_ASAP7_75t_R FILLER_0_176_1066 ();
 FILLER_ASAP7_75t_R FILLER_0_176_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_0_176_1090 ();
 FILLER_ASAP7_75t_R FILLER_0_176_1096 ();
 DECAPx4_ASAP7_75t_R FILLER_0_176_1104 ();
 FILLER_ASAP7_75t_R FILLER_0_176_1114 ();
 FILLER_ASAP7_75t_R FILLER_0_176_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_1130 ();
 DECAPx4_ASAP7_75t_R FILLER_0_176_1137 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_1147 ();
 FILLER_ASAP7_75t_R FILLER_0_176_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_1156 ();
 FILLER_ASAP7_75t_R FILLER_0_176_1163 ();
 FILLER_ASAP7_75t_R FILLER_0_176_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_1173 ();
 FILLER_ASAP7_75t_R FILLER_0_176_1180 ();
 DECAPx1_ASAP7_75t_R FILLER_0_176_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_1194 ();
 DECAPx1_ASAP7_75t_R FILLER_0_176_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_1209 ();
 DECAPx1_ASAP7_75t_R FILLER_0_176_1216 ();
 DECAPx1_ASAP7_75t_R FILLER_0_176_1226 ();
 DECAPx1_ASAP7_75t_R FILLER_0_176_1236 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176_1240 ();
 FILLER_ASAP7_75t_R FILLER_0_176_1247 ();
 DECAPx2_ASAP7_75t_R FILLER_0_176_1255 ();
 FILLER_ASAP7_75t_R FILLER_0_176_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_0_176_1269 ();
 DECAPx10_ASAP7_75t_R FILLER_0_176_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_0_176_1313 ();
 DECAPx10_ASAP7_75t_R FILLER_0_176_1335 ();
 DECAPx6_ASAP7_75t_R FILLER_0_176_1357 ();
 DECAPx1_ASAP7_75t_R FILLER_0_176_1371 ();
 FILLER_ASAP7_75t_R FILLER_0_176_1380 ();
 DECAPx2_ASAP7_75t_R FILLER_0_177_2 ();
 FILLER_ASAP7_75t_R FILLER_0_177_14 ();
 FILLER_ASAP7_75t_R FILLER_0_177_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_24 ();
 FILLER_ASAP7_75t_R FILLER_0_177_28 ();
 FILLER_ASAP7_75t_R FILLER_0_177_51 ();
 FILLER_ASAP7_75t_R FILLER_0_177_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_58 ();
 FILLER_ASAP7_75t_R FILLER_0_177_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_71 ();
 FILLER_ASAP7_75t_R FILLER_0_177_75 ();
 FILLER_ASAP7_75t_R FILLER_0_177_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_90 ();
 FILLER_ASAP7_75t_R FILLER_0_177_97 ();
 DECAPx1_ASAP7_75t_R FILLER_0_177_105 ();
 FILLER_ASAP7_75t_R FILLER_0_177_115 ();
 DECAPx4_ASAP7_75t_R FILLER_0_177_125 ();
 FILLER_ASAP7_75t_R FILLER_0_177_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_137 ();
 DECAPx1_ASAP7_75t_R FILLER_0_177_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_154 ();
 FILLER_ASAP7_75t_R FILLER_0_177_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_160 ();
 FILLER_ASAP7_75t_R FILLER_0_177_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_166 ();
 DECAPx2_ASAP7_75t_R FILLER_0_177_175 ();
 FILLER_ASAP7_75t_R FILLER_0_177_187 ();
 DECAPx1_ASAP7_75t_R FILLER_0_177_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_199 ();
 FILLER_ASAP7_75t_R FILLER_0_177_212 ();
 FILLER_ASAP7_75t_R FILLER_0_177_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_228 ();
 DECAPx2_ASAP7_75t_R FILLER_0_177_235 ();
 FILLER_ASAP7_75t_R FILLER_0_177_241 ();
 FILLER_ASAP7_75t_R FILLER_0_177_248 ();
 FILLER_ASAP7_75t_R FILLER_0_177_253 ();
 DECAPx1_ASAP7_75t_R FILLER_0_177_276 ();
 DECAPx6_ASAP7_75t_R FILLER_0_177_290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_177_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_310 ();
 DECAPx1_ASAP7_75t_R FILLER_0_177_321 ();
 DECAPx10_ASAP7_75t_R FILLER_0_177_332 ();
 FILLER_ASAP7_75t_R FILLER_0_177_354 ();
 FILLER_ASAP7_75t_R FILLER_0_177_378 ();
 FILLER_ASAP7_75t_R FILLER_0_177_386 ();
 DECAPx2_ASAP7_75t_R FILLER_0_177_408 ();
 FILLER_ASAP7_75t_R FILLER_0_177_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_177_444 ();
 FILLER_ASAP7_75t_R FILLER_0_177_458 ();
 FILLER_ASAP7_75t_R FILLER_0_177_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_468 ();
 FILLER_ASAP7_75t_R FILLER_0_177_474 ();
 DECAPx1_ASAP7_75t_R FILLER_0_177_486 ();
 FILLER_ASAP7_75t_R FILLER_0_177_495 ();
 FILLER_ASAP7_75t_R FILLER_0_177_521 ();
 FILLER_ASAP7_75t_R FILLER_0_177_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_535 ();
 FILLER_ASAP7_75t_R FILLER_0_177_542 ();
 DECAPx4_ASAP7_75t_R FILLER_0_177_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_559 ();
 DECAPx2_ASAP7_75t_R FILLER_0_177_566 ();
 DECAPx1_ASAP7_75t_R FILLER_0_177_578 ();
 DECAPx2_ASAP7_75t_R FILLER_0_177_589 ();
 FILLER_ASAP7_75t_R FILLER_0_177_595 ();
 FILLER_ASAP7_75t_R FILLER_0_177_603 ();
 FILLER_ASAP7_75t_R FILLER_0_177_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_615 ();
 FILLER_ASAP7_75t_R FILLER_0_177_619 ();
 FILLER_ASAP7_75t_R FILLER_0_177_629 ();
 DECAPx4_ASAP7_75t_R FILLER_0_177_639 ();
 FILLER_ASAP7_75t_R FILLER_0_177_649 ();
 DECAPx10_ASAP7_75t_R FILLER_0_177_657 ();
 DECAPx2_ASAP7_75t_R FILLER_0_177_679 ();
 FILLER_ASAP7_75t_R FILLER_0_177_691 ();
 FILLER_ASAP7_75t_R FILLER_0_177_699 ();
 DECAPx4_ASAP7_75t_R FILLER_0_177_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_717 ();
 FILLER_ASAP7_75t_R FILLER_0_177_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_723 ();
 DECAPx2_ASAP7_75t_R FILLER_0_177_731 ();
 FILLER_ASAP7_75t_R FILLER_0_177_744 ();
 DECAPx2_ASAP7_75t_R FILLER_0_177_749 ();
 FILLER_ASAP7_75t_R FILLER_0_177_755 ();
 FILLER_ASAP7_75t_R FILLER_0_177_769 ();
 DECAPx2_ASAP7_75t_R FILLER_0_177_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_787 ();
 FILLER_ASAP7_75t_R FILLER_0_177_798 ();
 FILLER_ASAP7_75t_R FILLER_0_177_810 ();
 FILLER_ASAP7_75t_R FILLER_0_177_822 ();
 DECAPx2_ASAP7_75t_R FILLER_0_177_834 ();
 DECAPx2_ASAP7_75t_R FILLER_0_177_850 ();
 FILLER_ASAP7_75t_R FILLER_0_177_862 ();
 FILLER_ASAP7_75t_R FILLER_0_177_870 ();
 FILLER_ASAP7_75t_R FILLER_0_177_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_880 ();
 FILLER_ASAP7_75t_R FILLER_0_177_884 ();
 DECAPx1_ASAP7_75t_R FILLER_0_177_892 ();
 FILLER_ASAP7_75t_R FILLER_0_177_906 ();
 FILLER_ASAP7_75t_R FILLER_0_177_918 ();
 FILLER_ASAP7_75t_R FILLER_0_177_923 ();
 FILLER_ASAP7_75t_R FILLER_0_177_927 ();
 FILLER_ASAP7_75t_R FILLER_0_177_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_951 ();
 DECAPx2_ASAP7_75t_R FILLER_0_177_955 ();
 DECAPx1_ASAP7_75t_R FILLER_0_177_972 ();
 FILLER_ASAP7_75t_R FILLER_0_177_988 ();
 DECAPx2_ASAP7_75t_R FILLER_0_177_1002 ();
 FILLER_ASAP7_75t_R FILLER_0_177_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_1010 ();
 DECAPx4_ASAP7_75t_R FILLER_0_177_1017 ();
 FILLER_ASAP7_75t_R FILLER_0_177_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_1029 ();
 DECAPx6_ASAP7_75t_R FILLER_0_177_1050 ();
 DECAPx2_ASAP7_75t_R FILLER_0_177_1064 ();
 FILLER_ASAP7_75t_R FILLER_0_177_1077 ();
 DECAPx10_ASAP7_75t_R FILLER_0_177_1085 ();
 FILLER_ASAP7_75t_R FILLER_0_177_1107 ();
 DECAPx10_ASAP7_75t_R FILLER_0_177_1112 ();
 DECAPx4_ASAP7_75t_R FILLER_0_177_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_1144 ();
 FILLER_ASAP7_75t_R FILLER_0_177_1151 ();
 DECAPx2_ASAP7_75t_R FILLER_0_177_1159 ();
 FILLER_ASAP7_75t_R FILLER_0_177_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_1167 ();
 DECAPx2_ASAP7_75t_R FILLER_0_177_1174 ();
 FILLER_ASAP7_75t_R FILLER_0_177_1185 ();
 FILLER_ASAP7_75t_R FILLER_0_177_1207 ();
 DECAPx2_ASAP7_75t_R FILLER_0_177_1219 ();
 DECAPx2_ASAP7_75t_R FILLER_0_177_1231 ();
 FILLER_ASAP7_75t_R FILLER_0_177_1237 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_1239 ();
 DECAPx2_ASAP7_75t_R FILLER_0_177_1246 ();
 FILLER_ASAP7_75t_R FILLER_0_177_1252 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_1254 ();
 DECAPx2_ASAP7_75t_R FILLER_0_177_1261 ();
 FILLER_ASAP7_75t_R FILLER_0_177_1273 ();
 DECAPx10_ASAP7_75t_R FILLER_0_177_1281 ();
 DECAPx10_ASAP7_75t_R FILLER_0_177_1303 ();
 DECAPx10_ASAP7_75t_R FILLER_0_177_1325 ();
 DECAPx10_ASAP7_75t_R FILLER_0_177_1347 ();
 DECAPx4_ASAP7_75t_R FILLER_0_177_1369 ();
 FILLER_ASAP7_75t_R FILLER_0_177_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177_1381 ();
 DECAPx1_ASAP7_75t_R FILLER_0_178_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_6 ();
 FILLER_ASAP7_75t_R FILLER_0_178_28 ();
 FILLER_ASAP7_75t_R FILLER_0_178_36 ();
 FILLER_ASAP7_75t_R FILLER_0_178_43 ();
 DECAPx1_ASAP7_75t_R FILLER_0_178_50 ();
 FILLER_ASAP7_75t_R FILLER_0_178_76 ();
 DECAPx4_ASAP7_75t_R FILLER_0_178_81 ();
 FILLER_ASAP7_75t_R FILLER_0_178_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_93 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_103 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_125 ();
 DECAPx6_ASAP7_75t_R FILLER_0_178_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_161 ();
 FILLER_ASAP7_75t_R FILLER_0_178_173 ();
 DECAPx1_ASAP7_75t_R FILLER_0_178_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_185 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_213 ();
 DECAPx1_ASAP7_75t_R FILLER_0_178_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_230 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_237 ();
 FILLER_ASAP7_75t_R FILLER_0_178_243 ();
 FILLER_ASAP7_75t_R FILLER_0_178_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_251 ();
 FILLER_ASAP7_75t_R FILLER_0_178_278 ();
 DECAPx1_ASAP7_75t_R FILLER_0_178_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_294 ();
 FILLER_ASAP7_75t_R FILLER_0_178_300 ();
 FILLER_ASAP7_75t_R FILLER_0_178_312 ();
 DECAPx1_ASAP7_75t_R FILLER_0_178_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_340 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_351 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_373 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_395 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_417 ();
 FILLER_ASAP7_75t_R FILLER_0_178_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_425 ();
 DECAPx4_ASAP7_75t_R FILLER_0_178_436 ();
 FILLER_ASAP7_75t_R FILLER_0_178_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_448 ();
 FILLER_ASAP7_75t_R FILLER_0_178_452 ();
 FILLER_ASAP7_75t_R FILLER_0_178_460 ();
 FILLER_ASAP7_75t_R FILLER_0_178_464 ();
 FILLER_ASAP7_75t_R FILLER_0_178_472 ();
 FILLER_ASAP7_75t_R FILLER_0_178_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_486 ();
 FILLER_ASAP7_75t_R FILLER_0_178_497 ();
 FILLER_ASAP7_75t_R FILLER_0_178_521 ();
 FILLER_ASAP7_75t_R FILLER_0_178_533 ();
 FILLER_ASAP7_75t_R FILLER_0_178_540 ();
 FILLER_ASAP7_75t_R FILLER_0_178_550 ();
 FILLER_ASAP7_75t_R FILLER_0_178_559 ();
 FILLER_ASAP7_75t_R FILLER_0_178_566 ();
 FILLER_ASAP7_75t_R FILLER_0_178_574 ();
 FILLER_ASAP7_75t_R FILLER_0_178_582 ();
 DECAPx6_ASAP7_75t_R FILLER_0_178_590 ();
 FILLER_ASAP7_75t_R FILLER_0_178_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_606 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_610 ();
 FILLER_ASAP7_75t_R FILLER_0_178_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_618 ();
 DECAPx1_ASAP7_75t_R FILLER_0_178_622 ();
 DECAPx1_ASAP7_75t_R FILLER_0_178_632 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_642 ();
 FILLER_ASAP7_75t_R FILLER_0_178_648 ();
 DECAPx6_ASAP7_75t_R FILLER_0_178_656 ();
 DECAPx4_ASAP7_75t_R FILLER_0_178_673 ();
 FILLER_ASAP7_75t_R FILLER_0_178_683 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_692 ();
 FILLER_ASAP7_75t_R FILLER_0_178_701 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_709 ();
 FILLER_ASAP7_75t_R FILLER_0_178_725 ();
 FILLER_ASAP7_75t_R FILLER_0_178_733 ();
 DECAPx6_ASAP7_75t_R FILLER_0_178_741 ();
 FILLER_ASAP7_75t_R FILLER_0_178_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_769 ();
 FILLER_ASAP7_75t_R FILLER_0_178_780 ();
 FILLER_ASAP7_75t_R FILLER_0_178_787 ();
 FILLER_ASAP7_75t_R FILLER_0_178_801 ();
 FILLER_ASAP7_75t_R FILLER_0_178_821 ();
 FILLER_ASAP7_75t_R FILLER_0_178_833 ();
 FILLER_ASAP7_75t_R FILLER_0_178_845 ();
 DECAPx1_ASAP7_75t_R FILLER_0_178_857 ();
 FILLER_ASAP7_75t_R FILLER_0_178_869 ();
 FILLER_ASAP7_75t_R FILLER_0_178_877 ();
 DECAPx1_ASAP7_75t_R FILLER_0_178_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_895 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_902 ();
 FILLER_ASAP7_75t_R FILLER_0_178_914 ();
 FILLER_ASAP7_75t_R FILLER_0_178_936 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_948 ();
 FILLER_ASAP7_75t_R FILLER_0_178_970 ();
 FILLER_ASAP7_75t_R FILLER_0_178_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_998 ();
 DECAPx6_ASAP7_75t_R FILLER_0_178_1020 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_1034 ();
 FILLER_ASAP7_75t_R FILLER_0_178_1041 ();
 FILLER_ASAP7_75t_R FILLER_0_178_1049 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1057 ();
 FILLER_ASAP7_75t_R FILLER_0_178_1079 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_1081 ();
 DECAPx6_ASAP7_75t_R FILLER_0_178_1088 ();
 FILLER_ASAP7_75t_R FILLER_0_178_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_1104 ();
 FILLER_ASAP7_75t_R FILLER_0_178_1111 ();
 DECAPx1_ASAP7_75t_R FILLER_0_178_1119 ();
 DECAPx6_ASAP7_75t_R FILLER_0_178_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_1143 ();
 DECAPx4_ASAP7_75t_R FILLER_0_178_1150 ();
 FILLER_ASAP7_75t_R FILLER_0_178_1166 ();
 FILLER_ASAP7_75t_R FILLER_0_178_1175 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_1181 ();
 FILLER_ASAP7_75t_R FILLER_0_178_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_1189 ();
 DECAPx6_ASAP7_75t_R FILLER_0_178_1196 ();
 FILLER_ASAP7_75t_R FILLER_0_178_1210 ();
 FILLER_ASAP7_75t_R FILLER_0_178_1222 ();
 FILLER_ASAP7_75t_R FILLER_0_178_1227 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_1235 ();
 FILLER_ASAP7_75t_R FILLER_0_178_1241 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_1243 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_1250 ();
 FILLER_ASAP7_75t_R FILLER_0_178_1256 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_1258 ();
 DECAPx1_ASAP7_75t_R FILLER_0_178_1265 ();
 FILLER_ASAP7_75t_R FILLER_0_178_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1305 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1327 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1349 ();
 DECAPx4_ASAP7_75t_R FILLER_0_178_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178_1381 ();
 DECAPx1_ASAP7_75t_R FILLER_0_179_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_6 ();
 FILLER_ASAP7_75t_R FILLER_0_179_12 ();
 FILLER_ASAP7_75t_R FILLER_0_179_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_26 ();
 FILLER_ASAP7_75t_R FILLER_0_179_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_179_55 ();
 DECAPx2_ASAP7_75t_R FILLER_0_179_64 ();
 FILLER_ASAP7_75t_R FILLER_0_179_82 ();
 DECAPx1_ASAP7_75t_R FILLER_0_179_87 ();
 FILLER_ASAP7_75t_R FILLER_0_179_101 ();
 FILLER_ASAP7_75t_R FILLER_0_179_113 ();
 DECAPx1_ASAP7_75t_R FILLER_0_179_118 ();
 FILLER_ASAP7_75t_R FILLER_0_179_130 ();
 DECAPx1_ASAP7_75t_R FILLER_0_179_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_148 ();
 FILLER_ASAP7_75t_R FILLER_0_179_159 ();
 DECAPx6_ASAP7_75t_R FILLER_0_179_172 ();
 FILLER_ASAP7_75t_R FILLER_0_179_186 ();
 DECAPx1_ASAP7_75t_R FILLER_0_179_191 ();
 DECAPx1_ASAP7_75t_R FILLER_0_179_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_221 ();
 FILLER_ASAP7_75t_R FILLER_0_179_227 ();
 DECAPx1_ASAP7_75t_R FILLER_0_179_239 ();
 FILLER_ASAP7_75t_R FILLER_0_179_248 ();
 FILLER_ASAP7_75t_R FILLER_0_179_274 ();
 DECAPx2_ASAP7_75t_R FILLER_0_179_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_292 ();
 FILLER_ASAP7_75t_R FILLER_0_179_303 ();
 DECAPx1_ASAP7_75t_R FILLER_0_179_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_314 ();
 FILLER_ASAP7_75t_R FILLER_0_179_325 ();
 FILLER_ASAP7_75t_R FILLER_0_179_341 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_353 ();
 DECAPx6_ASAP7_75t_R FILLER_0_179_375 ();
 DECAPx2_ASAP7_75t_R FILLER_0_179_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_395 ();
 DECAPx6_ASAP7_75t_R FILLER_0_179_416 ();
 FILLER_ASAP7_75t_R FILLER_0_179_430 ();
 FILLER_ASAP7_75t_R FILLER_0_179_453 ();
 FILLER_ASAP7_75t_R FILLER_0_179_463 ();
 FILLER_ASAP7_75t_R FILLER_0_179_471 ();
 FILLER_ASAP7_75t_R FILLER_0_179_495 ();
 FILLER_ASAP7_75t_R FILLER_0_179_519 ();
 FILLER_ASAP7_75t_R FILLER_0_179_527 ();
 FILLER_ASAP7_75t_R FILLER_0_179_535 ();
 FILLER_ASAP7_75t_R FILLER_0_179_547 ();
 FILLER_ASAP7_75t_R FILLER_0_179_559 ();
 DECAPx1_ASAP7_75t_R FILLER_0_179_571 ();
 FILLER_ASAP7_75t_R FILLER_0_179_581 ();
 FILLER_ASAP7_75t_R FILLER_0_179_589 ();
 DECAPx2_ASAP7_75t_R FILLER_0_179_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_600 ();
 FILLER_ASAP7_75t_R FILLER_0_179_607 ();
 DECAPx2_ASAP7_75t_R FILLER_0_179_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_622 ();
 DECAPx4_ASAP7_75t_R FILLER_0_179_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_639 ();
 FILLER_ASAP7_75t_R FILLER_0_179_643 ();
 DECAPx1_ASAP7_75t_R FILLER_0_179_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_657 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_664 ();
 DECAPx1_ASAP7_75t_R FILLER_0_179_686 ();
 DECAPx6_ASAP7_75t_R FILLER_0_179_696 ();
 DECAPx2_ASAP7_75t_R FILLER_0_179_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_716 ();
 FILLER_ASAP7_75t_R FILLER_0_179_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_722 ();
 FILLER_ASAP7_75t_R FILLER_0_179_730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_739 ();
 DECAPx2_ASAP7_75t_R FILLER_0_179_761 ();
 FILLER_ASAP7_75t_R FILLER_0_179_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_769 ();
 DECAPx1_ASAP7_75t_R FILLER_0_179_775 ();
 FILLER_ASAP7_75t_R FILLER_0_179_789 ();
 FILLER_ASAP7_75t_R FILLER_0_179_801 ();
 FILLER_ASAP7_75t_R FILLER_0_179_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_815 ();
 FILLER_ASAP7_75t_R FILLER_0_179_826 ();
 FILLER_ASAP7_75t_R FILLER_0_179_838 ();
 FILLER_ASAP7_75t_R FILLER_0_179_850 ();
 FILLER_ASAP7_75t_R FILLER_0_179_862 ();
 FILLER_ASAP7_75t_R FILLER_0_179_870 ();
 FILLER_ASAP7_75t_R FILLER_0_179_878 ();
 FILLER_ASAP7_75t_R FILLER_0_179_886 ();
 FILLER_ASAP7_75t_R FILLER_0_179_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_893 ();
 DECAPx1_ASAP7_75t_R FILLER_0_179_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_908 ();
 DECAPx4_ASAP7_75t_R FILLER_0_179_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_924 ();
 DECAPx4_ASAP7_75t_R FILLER_0_179_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_937 ();
 DECAPx1_ASAP7_75t_R FILLER_0_179_944 ();
 FILLER_ASAP7_75t_R FILLER_0_179_954 ();
 FILLER_ASAP7_75t_R FILLER_0_179_962 ();
 DECAPx2_ASAP7_75t_R FILLER_0_179_970 ();
 FILLER_ASAP7_75t_R FILLER_0_179_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_978 ();
 FILLER_ASAP7_75t_R FILLER_0_179_991 ();
 DECAPx1_ASAP7_75t_R FILLER_0_179_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_1009 ();
 DECAPx4_ASAP7_75t_R FILLER_0_179_1015 ();
 FILLER_ASAP7_75t_R FILLER_0_179_1025 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_1027 ();
 DECAPx2_ASAP7_75t_R FILLER_0_179_1038 ();
 DECAPx2_ASAP7_75t_R FILLER_0_179_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_1057 ();
 DECAPx4_ASAP7_75t_R FILLER_0_179_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1081 ();
 FILLER_ASAP7_75t_R FILLER_0_179_1103 ();
 DECAPx2_ASAP7_75t_R FILLER_0_179_1111 ();
 FILLER_ASAP7_75t_R FILLER_0_179_1117 ();
 DECAPx2_ASAP7_75t_R FILLER_0_179_1125 ();
 FILLER_ASAP7_75t_R FILLER_0_179_1131 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1139 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1161 ();
 DECAPx1_ASAP7_75t_R FILLER_0_179_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_1187 ();
 FILLER_ASAP7_75t_R FILLER_0_179_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_1197 ();
 DECAPx4_ASAP7_75t_R FILLER_0_179_1204 ();
 FILLER_ASAP7_75t_R FILLER_0_179_1221 ();
 DECAPx6_ASAP7_75t_R FILLER_0_179_1229 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179_1243 ();
 FILLER_ASAP7_75t_R FILLER_0_179_1250 ();
 FILLER_ASAP7_75t_R FILLER_0_179_1258 ();
 DECAPx2_ASAP7_75t_R FILLER_0_179_1270 ();
 FILLER_ASAP7_75t_R FILLER_0_179_1276 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1284 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1306 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1328 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1350 ();
 DECAPx4_ASAP7_75t_R FILLER_0_179_1372 ();
 FILLER_ASAP7_75t_R FILLER_0_180_2 ();
 FILLER_ASAP7_75t_R FILLER_0_180_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_11 ();
 FILLER_ASAP7_75t_R FILLER_0_180_18 ();
 FILLER_ASAP7_75t_R FILLER_0_180_26 ();
 FILLER_ASAP7_75t_R FILLER_0_180_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_35 ();
 FILLER_ASAP7_75t_R FILLER_0_180_42 ();
 FILLER_ASAP7_75t_R FILLER_0_180_49 ();
 FILLER_ASAP7_75t_R FILLER_0_180_54 ();
 DECAPx6_ASAP7_75t_R FILLER_0_180_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_73 ();
 DECAPx2_ASAP7_75t_R FILLER_0_180_77 ();
 FILLER_ASAP7_75t_R FILLER_0_180_89 ();
 FILLER_ASAP7_75t_R FILLER_0_180_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_99 ();
 FILLER_ASAP7_75t_R FILLER_0_180_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_108 ();
 FILLER_ASAP7_75t_R FILLER_0_180_115 ();
 FILLER_ASAP7_75t_R FILLER_0_180_123 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_133 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_155 ();
 DECAPx4_ASAP7_75t_R FILLER_0_180_177 ();
 DECAPx2_ASAP7_75t_R FILLER_0_180_208 ();
 DECAPx1_ASAP7_75t_R FILLER_0_180_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_222 ();
 FILLER_ASAP7_75t_R FILLER_0_180_228 ();
 FILLER_ASAP7_75t_R FILLER_0_180_258 ();
 FILLER_ASAP7_75t_R FILLER_0_180_270 ();
 FILLER_ASAP7_75t_R FILLER_0_180_282 ();
 FILLER_ASAP7_75t_R FILLER_0_180_294 ();
 FILLER_ASAP7_75t_R FILLER_0_180_306 ();
 FILLER_ASAP7_75t_R FILLER_0_180_318 ();
 FILLER_ASAP7_75t_R FILLER_0_180_330 ();
 DECAPx4_ASAP7_75t_R FILLER_0_180_338 ();
 FILLER_ASAP7_75t_R FILLER_0_180_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_350 ();
 DECAPx2_ASAP7_75t_R FILLER_0_180_361 ();
 DECAPx2_ASAP7_75t_R FILLER_0_180_373 ();
 FILLER_ASAP7_75t_R FILLER_0_180_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_385 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_407 ();
 FILLER_ASAP7_75t_R FILLER_0_180_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_431 ();
 FILLER_ASAP7_75t_R FILLER_0_180_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_442 ();
 FILLER_ASAP7_75t_R FILLER_0_180_448 ();
 FILLER_ASAP7_75t_R FILLER_0_180_460 ();
 FILLER_ASAP7_75t_R FILLER_0_180_464 ();
 FILLER_ASAP7_75t_R FILLER_0_180_473 ();
 FILLER_ASAP7_75t_R FILLER_0_180_485 ();
 FILLER_ASAP7_75t_R FILLER_0_180_511 ();
 FILLER_ASAP7_75t_R FILLER_0_180_535 ();
 DECAPx1_ASAP7_75t_R FILLER_0_180_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_551 ();
 FILLER_ASAP7_75t_R FILLER_0_180_558 ();
 FILLER_ASAP7_75t_R FILLER_0_180_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_565 ();
 DECAPx2_ASAP7_75t_R FILLER_0_180_584 ();
 DECAPx1_ASAP7_75t_R FILLER_0_180_596 ();
 FILLER_ASAP7_75t_R FILLER_0_180_608 ();
 FILLER_ASAP7_75t_R FILLER_0_180_616 ();
 DECAPx6_ASAP7_75t_R FILLER_0_180_624 ();
 DECAPx1_ASAP7_75t_R FILLER_0_180_638 ();
 FILLER_ASAP7_75t_R FILLER_0_180_645 ();
 FILLER_ASAP7_75t_R FILLER_0_180_653 ();
 DECAPx4_ASAP7_75t_R FILLER_0_180_662 ();
 FILLER_ASAP7_75t_R FILLER_0_180_672 ();
 FILLER_ASAP7_75t_R FILLER_0_180_696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_707 ();
 FILLER_ASAP7_75t_R FILLER_0_180_740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_750 ();
 DECAPx4_ASAP7_75t_R FILLER_0_180_772 ();
 FILLER_ASAP7_75t_R FILLER_0_180_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_790 ();
 FILLER_ASAP7_75t_R FILLER_0_180_801 ();
 FILLER_ASAP7_75t_R FILLER_0_180_813 ();
 FILLER_ASAP7_75t_R FILLER_0_180_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_827 ();
 FILLER_ASAP7_75t_R FILLER_0_180_838 ();
 FILLER_ASAP7_75t_R FILLER_0_180_850 ();
 FILLER_ASAP7_75t_R FILLER_0_180_858 ();
 FILLER_ASAP7_75t_R FILLER_0_180_866 ();
 DECAPx6_ASAP7_75t_R FILLER_0_180_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_887 ();
 FILLER_ASAP7_75t_R FILLER_0_180_896 ();
 DECAPx2_ASAP7_75t_R FILLER_0_180_901 ();
 FILLER_ASAP7_75t_R FILLER_0_180_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_909 ();
 DECAPx1_ASAP7_75t_R FILLER_0_180_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_924 ();
 FILLER_ASAP7_75t_R FILLER_0_180_932 ();
 DECAPx1_ASAP7_75t_R FILLER_0_180_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_944 ();
 DECAPx1_ASAP7_75t_R FILLER_0_180_951 ();
 FILLER_ASAP7_75t_R FILLER_0_180_961 ();
 DECAPx1_ASAP7_75t_R FILLER_0_180_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_973 ();
 DECAPx2_ASAP7_75t_R FILLER_0_180_995 ();
 DECAPx6_ASAP7_75t_R FILLER_0_180_1009 ();
 DECAPx1_ASAP7_75t_R FILLER_0_180_1023 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_1027 ();
 FILLER_ASAP7_75t_R FILLER_0_180_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_1036 ();
 FILLER_ASAP7_75t_R FILLER_0_180_1043 ();
 DECAPx1_ASAP7_75t_R FILLER_0_180_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_1057 ();
 DECAPx2_ASAP7_75t_R FILLER_0_180_1068 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_0_180_1081 ();
 FILLER_ASAP7_75t_R FILLER_0_180_1087 ();
 DECAPx1_ASAP7_75t_R FILLER_0_180_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_1105 ();
 FILLER_ASAP7_75t_R FILLER_0_180_1113 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_1115 ();
 DECAPx4_ASAP7_75t_R FILLER_0_180_1127 ();
 FILLER_ASAP7_75t_R FILLER_0_180_1143 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_1145 ();
 FILLER_ASAP7_75t_R FILLER_0_180_1156 ();
 FILLER_ASAP7_75t_R FILLER_0_180_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_1166 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1173 ();
 DECAPx6_ASAP7_75t_R FILLER_0_180_1195 ();
 FILLER_ASAP7_75t_R FILLER_0_180_1209 ();
 DECAPx6_ASAP7_75t_R FILLER_0_180_1219 ();
 DECAPx2_ASAP7_75t_R FILLER_0_180_1233 ();
 DECAPx4_ASAP7_75t_R FILLER_0_180_1246 ();
 FILLER_ASAP7_75t_R FILLER_0_180_1256 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_1258 ();
 FILLER_ASAP7_75t_R FILLER_0_180_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_0_180_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1348 ();
 DECAPx4_ASAP7_75t_R FILLER_0_180_1370 ();
 FILLER_ASAP7_75t_R FILLER_0_180_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_181_2 ();
 FILLER_ASAP7_75t_R FILLER_0_181_9 ();
 FILLER_ASAP7_75t_R FILLER_0_181_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181_18 ();
 FILLER_ASAP7_75t_R FILLER_0_181_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181_43 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_47 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_69 ();
 FILLER_ASAP7_75t_R FILLER_0_181_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181_77 ();
 DECAPx4_ASAP7_75t_R FILLER_0_181_81 ();
 DECAPx4_ASAP7_75t_R FILLER_0_181_101 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181_123 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_134 ();
 DECAPx1_ASAP7_75t_R FILLER_0_181_156 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181_176 ();
 FILLER_ASAP7_75t_R FILLER_0_181_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181_185 ();
 FILLER_ASAP7_75t_R FILLER_0_181_196 ();
 FILLER_ASAP7_75t_R FILLER_0_181_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181_203 ();
 DECAPx6_ASAP7_75t_R FILLER_0_181_215 ();
 FILLER_ASAP7_75t_R FILLER_0_181_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181_231 ();
 FILLER_ASAP7_75t_R FILLER_0_181_250 ();
 FILLER_ASAP7_75t_R FILLER_0_181_262 ();
 FILLER_ASAP7_75t_R FILLER_0_181_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181_276 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_287 ();
 FILLER_ASAP7_75t_R FILLER_0_181_293 ();
 FILLER_ASAP7_75t_R FILLER_0_181_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181_307 ();
 FILLER_ASAP7_75t_R FILLER_0_181_318 ();
 FILLER_ASAP7_75t_R FILLER_0_181_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181_332 ();
 FILLER_ASAP7_75t_R FILLER_0_181_343 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_355 ();
 FILLER_ASAP7_75t_R FILLER_0_181_361 ();
 FILLER_ASAP7_75t_R FILLER_0_181_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181_387 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_394 ();
 FILLER_ASAP7_75t_R FILLER_0_181_406 ();
 FILLER_ASAP7_75t_R FILLER_0_181_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181_413 ();
 DECAPx6_ASAP7_75t_R FILLER_0_181_424 ();
 DECAPx1_ASAP7_75t_R FILLER_0_181_438 ();
 DECAPx1_ASAP7_75t_R FILLER_0_181_445 ();
 FILLER_ASAP7_75t_R FILLER_0_181_454 ();
 FILLER_ASAP7_75t_R FILLER_0_181_466 ();
 FILLER_ASAP7_75t_R FILLER_0_181_478 ();
 FILLER_ASAP7_75t_R FILLER_0_181_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181_495 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_520 ();
 FILLER_ASAP7_75t_R FILLER_0_181_536 ();
 FILLER_ASAP7_75t_R FILLER_0_181_548 ();
 FILLER_ASAP7_75t_R FILLER_0_181_560 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_576 ();
 FILLER_ASAP7_75t_R FILLER_0_181_582 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_592 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_604 ();
 FILLER_ASAP7_75t_R FILLER_0_181_610 ();
 FILLER_ASAP7_75t_R FILLER_0_181_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_626 ();
 FILLER_ASAP7_75t_R FILLER_0_181_648 ();
 FILLER_ASAP7_75t_R FILLER_0_181_656 ();
 DECAPx4_ASAP7_75t_R FILLER_0_181_664 ();
 FILLER_ASAP7_75t_R FILLER_0_181_674 ();
 DECAPx1_ASAP7_75t_R FILLER_0_181_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181_702 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_714 ();
 DECAPx6_ASAP7_75t_R FILLER_0_181_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181_750 ();
 FILLER_ASAP7_75t_R FILLER_0_181_758 ();
 FILLER_ASAP7_75t_R FILLER_0_181_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181_768 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_775 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_787 ();
 FILLER_ASAP7_75t_R FILLER_0_181_798 ();
 FILLER_ASAP7_75t_R FILLER_0_181_812 ();
 FILLER_ASAP7_75t_R FILLER_0_181_824 ();
 FILLER_ASAP7_75t_R FILLER_0_181_836 ();
 FILLER_ASAP7_75t_R FILLER_0_181_848 ();
 FILLER_ASAP7_75t_R FILLER_0_181_858 ();
 FILLER_ASAP7_75t_R FILLER_0_181_866 ();
 FILLER_ASAP7_75t_R FILLER_0_181_874 ();
 FILLER_ASAP7_75t_R FILLER_0_181_882 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_890 ();
 FILLER_ASAP7_75t_R FILLER_0_181_896 ();
 DECAPx4_ASAP7_75t_R FILLER_0_181_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181_916 ();
 FILLER_ASAP7_75t_R FILLER_0_181_923 ();
 DECAPx4_ASAP7_75t_R FILLER_0_181_927 ();
 DECAPx1_ASAP7_75t_R FILLER_0_181_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181_947 ();
 DECAPx1_ASAP7_75t_R FILLER_0_181_954 ();
 DECAPx6_ASAP7_75t_R FILLER_0_181_964 ();
 FILLER_ASAP7_75t_R FILLER_0_181_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181_980 ();
 FILLER_ASAP7_75t_R FILLER_0_181_991 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_996 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_1018 ();
 FILLER_ASAP7_75t_R FILLER_0_181_1024 ();
 DECAPx6_ASAP7_75t_R FILLER_0_181_1032 ();
 DECAPx1_ASAP7_75t_R FILLER_0_181_1046 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181_1059 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_1063 ();
 FILLER_ASAP7_75t_R FILLER_0_181_1069 ();
 FILLER_ASAP7_75t_R FILLER_0_181_1077 ();
 DECAPx4_ASAP7_75t_R FILLER_0_181_1085 ();
 FILLER_ASAP7_75t_R FILLER_0_181_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181_1097 ();
 FILLER_ASAP7_75t_R FILLER_0_181_1104 ();
 FILLER_ASAP7_75t_R FILLER_0_181_1113 ();
 FILLER_ASAP7_75t_R FILLER_0_181_1121 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_1128 ();
 DECAPx1_ASAP7_75t_R FILLER_0_181_1140 ();
 DECAPx4_ASAP7_75t_R FILLER_0_181_1150 ();
 DECAPx6_ASAP7_75t_R FILLER_0_181_1163 ();
 FILLER_ASAP7_75t_R FILLER_0_181_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181_1179 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_1192 ();
 FILLER_ASAP7_75t_R FILLER_0_181_1198 ();
 FILLER_ASAP7_75t_R FILLER_0_181_1206 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_1214 ();
 DECAPx6_ASAP7_75t_R FILLER_0_181_1227 ();
 DECAPx1_ASAP7_75t_R FILLER_0_181_1241 ();
 FILLER_ASAP7_75t_R FILLER_0_181_1251 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_1259 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181_1265 ();
 DECAPx1_ASAP7_75t_R FILLER_0_181_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1348 ();
 DECAPx4_ASAP7_75t_R FILLER_0_181_1370 ();
 FILLER_ASAP7_75t_R FILLER_0_181_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_182_2 ();
 FILLER_ASAP7_75t_R FILLER_0_182_25 ();
 DECAPx2_ASAP7_75t_R FILLER_0_182_32 ();
 FILLER_ASAP7_75t_R FILLER_0_182_41 ();
 FILLER_ASAP7_75t_R FILLER_0_182_46 ();
 DECAPx6_ASAP7_75t_R FILLER_0_182_51 ();
 DECAPx1_ASAP7_75t_R FILLER_0_182_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_69 ();
 DECAPx6_ASAP7_75t_R FILLER_0_182_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_94 ();
 FILLER_ASAP7_75t_R FILLER_0_182_98 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_120 ();
 DECAPx6_ASAP7_75t_R FILLER_0_182_142 ();
 DECAPx2_ASAP7_75t_R FILLER_0_182_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_162 ();
 DECAPx6_ASAP7_75t_R FILLER_0_182_166 ();
 FILLER_ASAP7_75t_R FILLER_0_182_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_182 ();
 FILLER_ASAP7_75t_R FILLER_0_182_193 ();
 DECAPx2_ASAP7_75t_R FILLER_0_182_198 ();
 FILLER_ASAP7_75t_R FILLER_0_182_204 ();
 DECAPx1_ASAP7_75t_R FILLER_0_182_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_218 ();
 FILLER_ASAP7_75t_R FILLER_0_182_225 ();
 DECAPx2_ASAP7_75t_R FILLER_0_182_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_243 ();
 DECAPx1_ASAP7_75t_R FILLER_0_182_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_258 ();
 FILLER_ASAP7_75t_R FILLER_0_182_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_271 ();
 FILLER_ASAP7_75t_R FILLER_0_182_282 ();
 DECAPx4_ASAP7_75t_R FILLER_0_182_291 ();
 FILLER_ASAP7_75t_R FILLER_0_182_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_303 ();
 DECAPx6_ASAP7_75t_R FILLER_0_182_311 ();
 DECAPx1_ASAP7_75t_R FILLER_0_182_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_329 ();
 FILLER_ASAP7_75t_R FILLER_0_182_342 ();
 DECAPx2_ASAP7_75t_R FILLER_0_182_358 ();
 FILLER_ASAP7_75t_R FILLER_0_182_364 ();
 DECAPx2_ASAP7_75t_R FILLER_0_182_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_378 ();
 FILLER_ASAP7_75t_R FILLER_0_182_385 ();
 FILLER_ASAP7_75t_R FILLER_0_182_394 ();
 FILLER_ASAP7_75t_R FILLER_0_182_403 ();
 FILLER_ASAP7_75t_R FILLER_0_182_413 ();
 DECAPx1_ASAP7_75t_R FILLER_0_182_421 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_428 ();
 FILLER_ASAP7_75t_R FILLER_0_182_460 ();
 DECAPx2_ASAP7_75t_R FILLER_0_182_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_470 ();
 FILLER_ASAP7_75t_R FILLER_0_182_481 ();
 FILLER_ASAP7_75t_R FILLER_0_182_511 ();
 FILLER_ASAP7_75t_R FILLER_0_182_523 ();
 DECAPx1_ASAP7_75t_R FILLER_0_182_533 ();
 DECAPx1_ASAP7_75t_R FILLER_0_182_547 ();
 FILLER_ASAP7_75t_R FILLER_0_182_556 ();
 FILLER_ASAP7_75t_R FILLER_0_182_563 ();
 FILLER_ASAP7_75t_R FILLER_0_182_575 ();
 DECAPx1_ASAP7_75t_R FILLER_0_182_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_586 ();
 DECAPx1_ASAP7_75t_R FILLER_0_182_593 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_597 ();
 FILLER_ASAP7_75t_R FILLER_0_182_608 ();
 DECAPx4_ASAP7_75t_R FILLER_0_182_613 ();
 FILLER_ASAP7_75t_R FILLER_0_182_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_631 ();
 DECAPx2_ASAP7_75t_R FILLER_0_182_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_648 ();
 DECAPx6_ASAP7_75t_R FILLER_0_182_659 ();
 FILLER_ASAP7_75t_R FILLER_0_182_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_675 ();
 FILLER_ASAP7_75t_R FILLER_0_182_682 ();
 FILLER_ASAP7_75t_R FILLER_0_182_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_689 ();
 DECAPx1_ASAP7_75t_R FILLER_0_182_710 ();
 DECAPx6_ASAP7_75t_R FILLER_0_182_726 ();
 DECAPx1_ASAP7_75t_R FILLER_0_182_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_744 ();
 DECAPx2_ASAP7_75t_R FILLER_0_182_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_757 ();
 FILLER_ASAP7_75t_R FILLER_0_182_765 ();
 DECAPx1_ASAP7_75t_R FILLER_0_182_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_777 ();
 DECAPx2_ASAP7_75t_R FILLER_0_182_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_794 ();
 FILLER_ASAP7_75t_R FILLER_0_182_800 ();
 FILLER_ASAP7_75t_R FILLER_0_182_812 ();
 DECAPx2_ASAP7_75t_R FILLER_0_182_824 ();
 FILLER_ASAP7_75t_R FILLER_0_182_830 ();
 FILLER_ASAP7_75t_R FILLER_0_182_842 ();
 FILLER_ASAP7_75t_R FILLER_0_182_854 ();
 FILLER_ASAP7_75t_R FILLER_0_182_862 ();
 FILLER_ASAP7_75t_R FILLER_0_182_870 ();
 FILLER_ASAP7_75t_R FILLER_0_182_882 ();
 DECAPx1_ASAP7_75t_R FILLER_0_182_890 ();
 FILLER_ASAP7_75t_R FILLER_0_182_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_916 ();
 FILLER_ASAP7_75t_R FILLER_0_182_938 ();
 DECAPx4_ASAP7_75t_R FILLER_0_182_951 ();
 FILLER_ASAP7_75t_R FILLER_0_182_961 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_963 ();
 FILLER_ASAP7_75t_R FILLER_0_182_969 ();
 DECAPx2_ASAP7_75t_R FILLER_0_182_978 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_995 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_1039 ();
 DECAPx4_ASAP7_75t_R FILLER_0_182_1046 ();
 FILLER_ASAP7_75t_R FILLER_0_182_1056 ();
 FILLER_ASAP7_75t_R FILLER_0_182_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_1066 ();
 DECAPx1_ASAP7_75t_R FILLER_0_182_1073 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1083 ();
 FILLER_ASAP7_75t_R FILLER_0_182_1105 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_1107 ();
 DECAPx2_ASAP7_75t_R FILLER_0_182_1115 ();
 FILLER_ASAP7_75t_R FILLER_0_182_1121 ();
 DECAPx4_ASAP7_75t_R FILLER_0_182_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_1140 ();
 FILLER_ASAP7_75t_R FILLER_0_182_1147 ();
 DECAPx1_ASAP7_75t_R FILLER_0_182_1155 ();
 DECAPx1_ASAP7_75t_R FILLER_0_182_1166 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_1170 ();
 DECAPx6_ASAP7_75t_R FILLER_0_182_1177 ();
 FILLER_ASAP7_75t_R FILLER_0_182_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_1193 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1205 ();
 FILLER_ASAP7_75t_R FILLER_0_182_1227 ();
 FILLER_ASAP7_75t_R FILLER_0_182_1235 ();
 FILLER_ASAP7_75t_R FILLER_0_182_1243 ();
 FILLER_ASAP7_75t_R FILLER_0_182_1253 ();
 FILLER_ASAP7_75t_R FILLER_0_182_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1269 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1313 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1335 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_182_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_183_2 ();
 FILLER_ASAP7_75t_R FILLER_0_183_7 ();
 FILLER_ASAP7_75t_R FILLER_0_183_14 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_21 ();
 FILLER_ASAP7_75t_R FILLER_0_183_33 ();
 FILLER_ASAP7_75t_R FILLER_0_183_38 ();
 FILLER_ASAP7_75t_R FILLER_0_183_46 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_51 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_183_69 ();
 DECAPx6_ASAP7_75t_R FILLER_0_183_80 ();
 DECAPx1_ASAP7_75t_R FILLER_0_183_94 ();
 FILLER_ASAP7_75t_R FILLER_0_183_102 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_110 ();
 FILLER_ASAP7_75t_R FILLER_0_183_116 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_128 ();
 FILLER_ASAP7_75t_R FILLER_0_183_137 ();
 DECAPx1_ASAP7_75t_R FILLER_0_183_145 ();
 FILLER_ASAP7_75t_R FILLER_0_183_155 ();
 DECAPx6_ASAP7_75t_R FILLER_0_183_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_183_181 ();
 DECAPx6_ASAP7_75t_R FILLER_0_183_192 ();
 DECAPx1_ASAP7_75t_R FILLER_0_183_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_183_216 ();
 FILLER_ASAP7_75t_R FILLER_0_183_223 ();
 FILLER_ASAP7_75t_R FILLER_0_183_235 ();
 FILLER_ASAP7_75t_R FILLER_0_183_259 ();
 DECAPx1_ASAP7_75t_R FILLER_0_183_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_183_273 ();
 FILLER_ASAP7_75t_R FILLER_0_183_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_183_282 ();
 FILLER_ASAP7_75t_R FILLER_0_183_289 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_297 ();
 DECAPx6_ASAP7_75t_R FILLER_0_183_319 ();
 FILLER_ASAP7_75t_R FILLER_0_183_333 ();
 FILLER_ASAP7_75t_R FILLER_0_183_363 ();
 FILLER_ASAP7_75t_R FILLER_0_183_371 ();
 DECAPx1_ASAP7_75t_R FILLER_0_183_376 ();
 DECAPx4_ASAP7_75t_R FILLER_0_183_386 ();
 FILLER_ASAP7_75t_R FILLER_0_183_396 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_183_410 ();
 FILLER_ASAP7_75t_R FILLER_0_183_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_183_419 ();
 DECAPx6_ASAP7_75t_R FILLER_0_183_428 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_183_448 ();
 FILLER_ASAP7_75t_R FILLER_0_183_454 ();
 DECAPx1_ASAP7_75t_R FILLER_0_183_466 ();
 FILLER_ASAP7_75t_R FILLER_0_183_480 ();
 FILLER_ASAP7_75t_R FILLER_0_183_485 ();
 FILLER_ASAP7_75t_R FILLER_0_183_513 ();
 FILLER_ASAP7_75t_R FILLER_0_183_521 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_183_539 ();
 FILLER_ASAP7_75t_R FILLER_0_183_545 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_553 ();
 FILLER_ASAP7_75t_R FILLER_0_183_564 ();
 DECAPx1_ASAP7_75t_R FILLER_0_183_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_183_576 ();
 DECAPx1_ASAP7_75t_R FILLER_0_183_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_183_586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_594 ();
 DECAPx6_ASAP7_75t_R FILLER_0_183_616 ();
 FILLER_ASAP7_75t_R FILLER_0_183_630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_638 ();
 DECAPx1_ASAP7_75t_R FILLER_0_183_660 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_183_691 ();
 FILLER_ASAP7_75t_R FILLER_0_183_695 ();
 DECAPx4_ASAP7_75t_R FILLER_0_183_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_183_710 ();
 DECAPx1_ASAP7_75t_R FILLER_0_183_721 ();
 FILLER_ASAP7_75t_R FILLER_0_183_735 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_745 ();
 FILLER_ASAP7_75t_R FILLER_0_183_751 ();
 DECAPx1_ASAP7_75t_R FILLER_0_183_763 ();
 FILLER_ASAP7_75t_R FILLER_0_183_773 ();
 FILLER_ASAP7_75t_R FILLER_0_183_781 ();
 DECAPx1_ASAP7_75t_R FILLER_0_183_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_183_793 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_806 ();
 FILLER_ASAP7_75t_R FILLER_0_183_812 ();
 DECAPx1_ASAP7_75t_R FILLER_0_183_824 ();
 FILLER_ASAP7_75t_R FILLER_0_183_838 ();
 FILLER_ASAP7_75t_R FILLER_0_183_850 ();
 FILLER_ASAP7_75t_R FILLER_0_183_860 ();
 FILLER_ASAP7_75t_R FILLER_0_183_868 ();
 FILLER_ASAP7_75t_R FILLER_0_183_876 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_884 ();
 DECAPx1_ASAP7_75t_R FILLER_0_183_902 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_916 ();
 FILLER_ASAP7_75t_R FILLER_0_183_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_183_924 ();
 FILLER_ASAP7_75t_R FILLER_0_183_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_183_929 ();
 FILLER_ASAP7_75t_R FILLER_0_183_937 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_183_948 ();
 DECAPx1_ASAP7_75t_R FILLER_0_183_965 ();
 DECAPx4_ASAP7_75t_R FILLER_0_183_972 ();
 FILLER_ASAP7_75t_R FILLER_0_183_982 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_991 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_183_997 ();
 FILLER_ASAP7_75t_R FILLER_0_183_1013 ();
 DECAPx6_ASAP7_75t_R FILLER_0_183_1025 ();
 FILLER_ASAP7_75t_R FILLER_0_183_1039 ();
 FILLER_ASAP7_75t_R FILLER_0_183_1044 ();
 FILLER_ASAP7_75t_R FILLER_0_183_1058 ();
 FILLER_ASAP7_75t_R FILLER_0_183_1066 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_1073 ();
 FILLER_ASAP7_75t_R FILLER_0_183_1087 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_183_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_0_183_1097 ();
 FILLER_ASAP7_75t_R FILLER_0_183_1113 ();
 FILLER_ASAP7_75t_R FILLER_0_183_1122 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_1130 ();
 FILLER_ASAP7_75t_R FILLER_0_183_1136 ();
 FILLER_ASAP7_75t_R FILLER_0_183_1144 ();
 FILLER_ASAP7_75t_R FILLER_0_183_1152 ();
 FILLER_ASAP7_75t_R FILLER_0_183_1160 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_1168 ();
 FILLER_ASAP7_75t_R FILLER_0_183_1180 ();
 FILLER_ASAP7_75t_R FILLER_0_183_1188 ();
 FILLER_ASAP7_75t_R FILLER_0_183_1196 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_1204 ();
 DECAPx4_ASAP7_75t_R FILLER_0_183_1216 ();
 FILLER_ASAP7_75t_R FILLER_0_183_1232 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1240 ();
 DECAPx6_ASAP7_75t_R FILLER_0_183_1262 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_1276 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_183_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1333 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1355 ();
 DECAPx1_ASAP7_75t_R FILLER_0_183_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_183_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_184_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_184_9 ();
 FILLER_ASAP7_75t_R FILLER_0_184_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_20 ();
 FILLER_ASAP7_75t_R FILLER_0_184_24 ();
 FILLER_ASAP7_75t_R FILLER_0_184_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_39 ();
 DECAPx4_ASAP7_75t_R FILLER_0_184_46 ();
 FILLER_ASAP7_75t_R FILLER_0_184_56 ();
 FILLER_ASAP7_75t_R FILLER_0_184_61 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_69 ();
 DECAPx1_ASAP7_75t_R FILLER_0_184_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_82 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_89 ();
 DECAPx6_ASAP7_75t_R FILLER_0_184_111 ();
 FILLER_ASAP7_75t_R FILLER_0_184_125 ();
 FILLER_ASAP7_75t_R FILLER_0_184_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_140 ();
 FILLER_ASAP7_75t_R FILLER_0_184_144 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_152 ();
 DECAPx6_ASAP7_75t_R FILLER_0_184_164 ();
 DECAPx1_ASAP7_75t_R FILLER_0_184_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_182 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_195 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_206 ();
 FILLER_ASAP7_75t_R FILLER_0_184_212 ();
 DECAPx1_ASAP7_75t_R FILLER_0_184_217 ();
 FILLER_ASAP7_75t_R FILLER_0_184_231 ();
 DECAPx1_ASAP7_75t_R FILLER_0_184_255 ();
 FILLER_ASAP7_75t_R FILLER_0_184_265 ();
 FILLER_ASAP7_75t_R FILLER_0_184_273 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_281 ();
 FILLER_ASAP7_75t_R FILLER_0_184_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_289 ();
 DECAPx1_ASAP7_75t_R FILLER_0_184_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_300 ();
 FILLER_ASAP7_75t_R FILLER_0_184_323 ();
 FILLER_ASAP7_75t_R FILLER_0_184_335 ();
 FILLER_ASAP7_75t_R FILLER_0_184_342 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_354 ();
 FILLER_ASAP7_75t_R FILLER_0_184_360 ();
 FILLER_ASAP7_75t_R FILLER_0_184_368 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_377 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_389 ();
 DECAPx1_ASAP7_75t_R FILLER_0_184_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_405 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_422 ();
 FILLER_ASAP7_75t_R FILLER_0_184_429 ();
 DECAPx6_ASAP7_75t_R FILLER_0_184_434 ();
 FILLER_ASAP7_75t_R FILLER_0_184_448 ();
 FILLER_ASAP7_75t_R FILLER_0_184_460 ();
 FILLER_ASAP7_75t_R FILLER_0_184_464 ();
 DECAPx1_ASAP7_75t_R FILLER_0_184_476 ();
 FILLER_ASAP7_75t_R FILLER_0_184_486 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_504 ();
 FILLER_ASAP7_75t_R FILLER_0_184_510 ();
 FILLER_ASAP7_75t_R FILLER_0_184_522 ();
 FILLER_ASAP7_75t_R FILLER_0_184_534 ();
 DECAPx1_ASAP7_75t_R FILLER_0_184_542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_184_552 ();
 DECAPx1_ASAP7_75t_R FILLER_0_184_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_565 ();
 FILLER_ASAP7_75t_R FILLER_0_184_576 ();
 FILLER_ASAP7_75t_R FILLER_0_184_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_586 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_594 ();
 FILLER_ASAP7_75t_R FILLER_0_184_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_602 ();
 DECAPx1_ASAP7_75t_R FILLER_0_184_609 ();
 FILLER_ASAP7_75t_R FILLER_0_184_619 ();
 FILLER_ASAP7_75t_R FILLER_0_184_627 ();
 FILLER_ASAP7_75t_R FILLER_0_184_635 ();
 DECAPx1_ASAP7_75t_R FILLER_0_184_643 ();
 DECAPx4_ASAP7_75t_R FILLER_0_184_653 ();
 FILLER_ASAP7_75t_R FILLER_0_184_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_665 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_669 ();
 DECAPx4_ASAP7_75t_R FILLER_0_184_691 ();
 FILLER_ASAP7_75t_R FILLER_0_184_711 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_723 ();
 FILLER_ASAP7_75t_R FILLER_0_184_739 ();
 FILLER_ASAP7_75t_R FILLER_0_184_747 ();
 DECAPx4_ASAP7_75t_R FILLER_0_184_755 ();
 FILLER_ASAP7_75t_R FILLER_0_184_765 ();
 FILLER_ASAP7_75t_R FILLER_0_184_774 ();
 DECAPx1_ASAP7_75t_R FILLER_0_184_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_786 ();
 FILLER_ASAP7_75t_R FILLER_0_184_799 ();
 FILLER_ASAP7_75t_R FILLER_0_184_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_809 ();
 FILLER_ASAP7_75t_R FILLER_0_184_820 ();
 FILLER_ASAP7_75t_R FILLER_0_184_832 ();
 FILLER_ASAP7_75t_R FILLER_0_184_844 ();
 FILLER_ASAP7_75t_R FILLER_0_184_856 ();
 FILLER_ASAP7_75t_R FILLER_0_184_864 ();
 FILLER_ASAP7_75t_R FILLER_0_184_879 ();
 DECAPx1_ASAP7_75t_R FILLER_0_184_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_895 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_901 ();
 FILLER_ASAP7_75t_R FILLER_0_184_907 ();
 FILLER_ASAP7_75t_R FILLER_0_184_915 ();
 FILLER_ASAP7_75t_R FILLER_0_184_922 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_935 ();
 FILLER_ASAP7_75t_R FILLER_0_184_942 ();
 FILLER_ASAP7_75t_R FILLER_0_184_950 ();
 FILLER_ASAP7_75t_R FILLER_0_184_962 ();
 FILLER_ASAP7_75t_R FILLER_0_184_970 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_978 ();
 FILLER_ASAP7_75t_R FILLER_0_184_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_995 ();
 FILLER_ASAP7_75t_R FILLER_0_184_1017 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_1019 ();
 FILLER_ASAP7_75t_R FILLER_0_184_1026 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_1038 ();
 FILLER_ASAP7_75t_R FILLER_0_184_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_1046 ();
 FILLER_ASAP7_75t_R FILLER_0_184_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_1060 ();
 DECAPx6_ASAP7_75t_R FILLER_0_184_1068 ();
 FILLER_ASAP7_75t_R FILLER_0_184_1082 ();
 DECAPx1_ASAP7_75t_R FILLER_0_184_1091 ();
 FILLER_ASAP7_75t_R FILLER_0_184_1101 ();
 DECAPx4_ASAP7_75t_R FILLER_0_184_1110 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_1131 ();
 FILLER_ASAP7_75t_R FILLER_0_184_1143 ();
 DECAPx4_ASAP7_75t_R FILLER_0_184_1156 ();
 DECAPx4_ASAP7_75t_R FILLER_0_184_1172 ();
 FILLER_ASAP7_75t_R FILLER_0_184_1182 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_1184 ();
 DECAPx1_ASAP7_75t_R FILLER_0_184_1191 ();
 FILLER_ASAP7_75t_R FILLER_0_184_1201 ();
 DECAPx4_ASAP7_75t_R FILLER_0_184_1214 ();
 FILLER_ASAP7_75t_R FILLER_0_184_1230 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_1232 ();
 DECAPx6_ASAP7_75t_R FILLER_0_184_1239 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_1253 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_1259 ();
 FILLER_ASAP7_75t_R FILLER_0_184_1266 ();
 DECAPx1_ASAP7_75t_R FILLER_0_184_1274 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1285 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1307 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1351 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_184_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184_1381 ();
 DECAPx1_ASAP7_75t_R FILLER_0_185_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_9 ();
 FILLER_ASAP7_75t_R FILLER_0_185_31 ();
 DECAPx4_ASAP7_75t_R FILLER_0_185_39 ();
 FILLER_ASAP7_75t_R FILLER_0_185_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_51 ();
 FILLER_ASAP7_75t_R FILLER_0_185_58 ();
 DECAPx6_ASAP7_75t_R FILLER_0_185_63 ();
 FILLER_ASAP7_75t_R FILLER_0_185_83 ();
 DECAPx4_ASAP7_75t_R FILLER_0_185_88 ();
 FILLER_ASAP7_75t_R FILLER_0_185_98 ();
 FILLER_ASAP7_75t_R FILLER_0_185_103 ();
 DECAPx4_ASAP7_75t_R FILLER_0_185_111 ();
 FILLER_ASAP7_75t_R FILLER_0_185_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_123 ();
 FILLER_ASAP7_75t_R FILLER_0_185_130 ();
 FILLER_ASAP7_75t_R FILLER_0_185_138 ();
 DECAPx1_ASAP7_75t_R FILLER_0_185_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_150 ();
 FILLER_ASAP7_75t_R FILLER_0_185_154 ();
 DECAPx6_ASAP7_75t_R FILLER_0_185_162 ();
 FILLER_ASAP7_75t_R FILLER_0_185_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_178 ();
 FILLER_ASAP7_75t_R FILLER_0_185_182 ();
 DECAPx4_ASAP7_75t_R FILLER_0_185_190 ();
 FILLER_ASAP7_75t_R FILLER_0_185_200 ();
 FILLER_ASAP7_75t_R FILLER_0_185_223 ();
 DECAPx4_ASAP7_75t_R FILLER_0_185_233 ();
 DECAPx1_ASAP7_75t_R FILLER_0_185_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_257 ();
 DECAPx1_ASAP7_75t_R FILLER_0_185_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_270 ();
 DECAPx2_ASAP7_75t_R FILLER_0_185_278 ();
 FILLER_ASAP7_75t_R FILLER_0_185_284 ();
 DECAPx1_ASAP7_75t_R FILLER_0_185_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_296 ();
 DECAPx4_ASAP7_75t_R FILLER_0_185_303 ();
 FILLER_ASAP7_75t_R FILLER_0_185_313 ();
 FILLER_ASAP7_75t_R FILLER_0_185_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_327 ();
 FILLER_ASAP7_75t_R FILLER_0_185_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_342 ();
 FILLER_ASAP7_75t_R FILLER_0_185_349 ();
 FILLER_ASAP7_75t_R FILLER_0_185_361 ();
 FILLER_ASAP7_75t_R FILLER_0_185_369 ();
 FILLER_ASAP7_75t_R FILLER_0_185_377 ();
 FILLER_ASAP7_75t_R FILLER_0_185_382 ();
 FILLER_ASAP7_75t_R FILLER_0_185_392 ();
 DECAPx4_ASAP7_75t_R FILLER_0_185_400 ();
 DECAPx1_ASAP7_75t_R FILLER_0_185_416 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_425 ();
 DECAPx2_ASAP7_75t_R FILLER_0_185_447 ();
 FILLER_ASAP7_75t_R FILLER_0_185_459 ();
 FILLER_ASAP7_75t_R FILLER_0_185_467 ();
 FILLER_ASAP7_75t_R FILLER_0_185_474 ();
 DECAPx1_ASAP7_75t_R FILLER_0_185_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_490 ();
 FILLER_ASAP7_75t_R FILLER_0_185_497 ();
 FILLER_ASAP7_75t_R FILLER_0_185_507 ();
 FILLER_ASAP7_75t_R FILLER_0_185_517 ();
 FILLER_ASAP7_75t_R FILLER_0_185_524 ();
 FILLER_ASAP7_75t_R FILLER_0_185_533 ();
 FILLER_ASAP7_75t_R FILLER_0_185_541 ();
 DECAPx6_ASAP7_75t_R FILLER_0_185_551 ();
 FILLER_ASAP7_75t_R FILLER_0_185_565 ();
 DECAPx4_ASAP7_75t_R FILLER_0_185_577 ();
 FILLER_ASAP7_75t_R FILLER_0_185_587 ();
 DECAPx4_ASAP7_75t_R FILLER_0_185_596 ();
 FILLER_ASAP7_75t_R FILLER_0_185_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_614 ();
 DECAPx2_ASAP7_75t_R FILLER_0_185_629 ();
 FILLER_ASAP7_75t_R FILLER_0_185_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_637 ();
 FILLER_ASAP7_75t_R FILLER_0_185_644 ();
 FILLER_ASAP7_75t_R FILLER_0_185_653 ();
 DECAPx4_ASAP7_75t_R FILLER_0_185_669 ();
 FILLER_ASAP7_75t_R FILLER_0_185_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_702 ();
 DECAPx2_ASAP7_75t_R FILLER_0_185_706 ();
 FILLER_ASAP7_75t_R FILLER_0_185_716 ();
 DECAPx1_ASAP7_75t_R FILLER_0_185_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_727 ();
 DECAPx2_ASAP7_75t_R FILLER_0_185_738 ();
 FILLER_ASAP7_75t_R FILLER_0_185_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_746 ();
 DECAPx2_ASAP7_75t_R FILLER_0_185_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_759 ();
 DECAPx6_ASAP7_75t_R FILLER_0_185_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_780 ();
 DECAPx2_ASAP7_75t_R FILLER_0_185_789 ();
 FILLER_ASAP7_75t_R FILLER_0_185_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_797 ();
 FILLER_ASAP7_75t_R FILLER_0_185_809 ();
 FILLER_ASAP7_75t_R FILLER_0_185_819 ();
 FILLER_ASAP7_75t_R FILLER_0_185_827 ();
 FILLER_ASAP7_75t_R FILLER_0_185_835 ();
 FILLER_ASAP7_75t_R FILLER_0_185_843 ();
 DECAPx2_ASAP7_75t_R FILLER_0_185_851 ();
 FILLER_ASAP7_75t_R FILLER_0_185_863 ();
 FILLER_ASAP7_75t_R FILLER_0_185_871 ();
 FILLER_ASAP7_75t_R FILLER_0_185_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_878 ();
 DECAPx2_ASAP7_75t_R FILLER_0_185_889 ();
 DECAPx2_ASAP7_75t_R FILLER_0_185_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_911 ();
 FILLER_ASAP7_75t_R FILLER_0_185_923 ();
 FILLER_ASAP7_75t_R FILLER_0_185_927 ();
 DECAPx2_ASAP7_75t_R FILLER_0_185_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_940 ();
 DECAPx2_ASAP7_75t_R FILLER_0_185_947 ();
 DECAPx4_ASAP7_75t_R FILLER_0_185_973 ();
 DECAPx4_ASAP7_75t_R FILLER_0_185_991 ();
 FILLER_ASAP7_75t_R FILLER_0_185_1006 ();
 DECAPx2_ASAP7_75t_R FILLER_0_185_1028 ();
 FILLER_ASAP7_75t_R FILLER_0_185_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_1036 ();
 FILLER_ASAP7_75t_R FILLER_0_185_1043 ();
 DECAPx6_ASAP7_75t_R FILLER_0_185_1051 ();
 FILLER_ASAP7_75t_R FILLER_0_185_1071 ();
 FILLER_ASAP7_75t_R FILLER_0_185_1083 ();
 DECAPx4_ASAP7_75t_R FILLER_0_185_1091 ();
 FILLER_ASAP7_75t_R FILLER_0_185_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_1103 ();
 FILLER_ASAP7_75t_R FILLER_0_185_1111 ();
 FILLER_ASAP7_75t_R FILLER_0_185_1120 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1130 ();
 FILLER_ASAP7_75t_R FILLER_0_185_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_1154 ();
 FILLER_ASAP7_75t_R FILLER_0_185_1161 ();
 DECAPx6_ASAP7_75t_R FILLER_0_185_1169 ();
 FILLER_ASAP7_75t_R FILLER_0_185_1183 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_1185 ();
 DECAPx4_ASAP7_75t_R FILLER_0_185_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_1203 ();
 DECAPx4_ASAP7_75t_R FILLER_0_185_1210 ();
 FILLER_ASAP7_75t_R FILLER_0_185_1220 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_1222 ();
 FILLER_ASAP7_75t_R FILLER_0_185_1229 ();
 DECAPx2_ASAP7_75t_R FILLER_0_185_1237 ();
 FILLER_ASAP7_75t_R FILLER_0_185_1249 ();
 FILLER_ASAP7_75t_R FILLER_0_185_1257 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_1259 ();
 FILLER_ASAP7_75t_R FILLER_0_185_1266 ();
 FILLER_ASAP7_75t_R FILLER_0_185_1274 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185_1276 ();
 FILLER_ASAP7_75t_R FILLER_0_185_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1354 ();
 DECAPx2_ASAP7_75t_R FILLER_0_185_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2 ();
 FILLER_ASAP7_75t_R FILLER_0_186_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_186_48 ();
 DECAPx4_ASAP7_75t_R FILLER_0_186_59 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_75 ();
 DECAPx1_ASAP7_75t_R FILLER_0_186_84 ();
 FILLER_ASAP7_75t_R FILLER_0_186_98 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_128 ();
 DECAPx1_ASAP7_75t_R FILLER_0_186_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_186_154 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_161 ();
 FILLER_ASAP7_75t_R FILLER_0_186_183 ();
 DECAPx6_ASAP7_75t_R FILLER_0_186_188 ();
 FILLER_ASAP7_75t_R FILLER_0_186_202 ();
 DECAPx4_ASAP7_75t_R FILLER_0_186_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_186_217 ();
 FILLER_ASAP7_75t_R FILLER_0_186_223 ();
 FILLER_ASAP7_75t_R FILLER_0_186_231 ();
 DECAPx1_ASAP7_75t_R FILLER_0_186_239 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_248 ();
 FILLER_ASAP7_75t_R FILLER_0_186_254 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_264 ();
 FILLER_ASAP7_75t_R FILLER_0_186_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_186_272 ();
 DECAPx1_ASAP7_75t_R FILLER_0_186_279 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_290 ();
 FILLER_ASAP7_75t_R FILLER_0_186_296 ();
 FILLER_ASAP7_75t_R FILLER_0_186_304 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_312 ();
 FILLER_ASAP7_75t_R FILLER_0_186_318 ();
 FILLER_ASAP7_75t_R FILLER_0_186_328 ();
 FILLER_ASAP7_75t_R FILLER_0_186_348 ();
 DECAPx1_ASAP7_75t_R FILLER_0_186_356 ();
 DECAPx1_ASAP7_75t_R FILLER_0_186_366 ();
 DECAPx4_ASAP7_75t_R FILLER_0_186_376 ();
 FILLER_ASAP7_75t_R FILLER_0_186_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_186_388 ();
 FILLER_ASAP7_75t_R FILLER_0_186_396 ();
 FILLER_ASAP7_75t_R FILLER_0_186_401 ();
 DECAPx1_ASAP7_75t_R FILLER_0_186_406 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_416 ();
 FILLER_ASAP7_75t_R FILLER_0_186_422 ();
 DECAPx6_ASAP7_75t_R FILLER_0_186_430 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_444 ();
 FILLER_ASAP7_75t_R FILLER_0_186_453 ();
 FILLER_ASAP7_75t_R FILLER_0_186_460 ();
 FILLER_ASAP7_75t_R FILLER_0_186_464 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_488 ();
 DECAPx1_ASAP7_75t_R FILLER_0_186_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_186_504 ();
 FILLER_ASAP7_75t_R FILLER_0_186_511 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_519 ();
 FILLER_ASAP7_75t_R FILLER_0_186_531 ();
 FILLER_ASAP7_75t_R FILLER_0_186_539 ();
 DECAPx6_ASAP7_75t_R FILLER_0_186_547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_186_561 ();
 FILLER_ASAP7_75t_R FILLER_0_186_575 ();
 FILLER_ASAP7_75t_R FILLER_0_186_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_186_582 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_186_595 ();
 FILLER_ASAP7_75t_R FILLER_0_186_602 ();
 DECAPx1_ASAP7_75t_R FILLER_0_186_610 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_186_623 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_630 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_657 ();
 DECAPx4_ASAP7_75t_R FILLER_0_186_679 ();
 FILLER_ASAP7_75t_R FILLER_0_186_689 ();
 FILLER_ASAP7_75t_R FILLER_0_186_697 ();
 FILLER_ASAP7_75t_R FILLER_0_186_711 ();
 FILLER_ASAP7_75t_R FILLER_0_186_716 ();
 FILLER_ASAP7_75t_R FILLER_0_186_728 ();
 DECAPx4_ASAP7_75t_R FILLER_0_186_742 ();
 FILLER_ASAP7_75t_R FILLER_0_186_752 ();
 FILLER_ASAP7_75t_R FILLER_0_186_762 ();
 FILLER_ASAP7_75t_R FILLER_0_186_774 ();
 FILLER_ASAP7_75t_R FILLER_0_186_782 ();
 DECAPx6_ASAP7_75t_R FILLER_0_186_790 ();
 FILLER_ASAP7_75t_R FILLER_0_186_811 ();
 FILLER_ASAP7_75t_R FILLER_0_186_819 ();
 FILLER_ASAP7_75t_R FILLER_0_186_827 ();
 DECAPx1_ASAP7_75t_R FILLER_0_186_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_186_841 ();
 FILLER_ASAP7_75t_R FILLER_0_186_852 ();
 FILLER_ASAP7_75t_R FILLER_0_186_860 ();
 FILLER_ASAP7_75t_R FILLER_0_186_868 ();
 FILLER_ASAP7_75t_R FILLER_0_186_876 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_186_890 ();
 FILLER_ASAP7_75t_R FILLER_0_186_901 ();
 FILLER_ASAP7_75t_R FILLER_0_186_913 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_186_926 ();
 FILLER_ASAP7_75t_R FILLER_0_186_933 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_941 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_963 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_186_969 ();
 DECAPx4_ASAP7_75t_R FILLER_0_186_992 ();
 DECAPx1_ASAP7_75t_R FILLER_0_186_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_186_1011 ();
 DECAPx6_ASAP7_75t_R FILLER_0_186_1018 ();
 DECAPx1_ASAP7_75t_R FILLER_0_186_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_186_1036 ();
 FILLER_ASAP7_75t_R FILLER_0_186_1042 ();
 DECAPx4_ASAP7_75t_R FILLER_0_186_1050 ();
 FILLER_ASAP7_75t_R FILLER_0_186_1060 ();
 FILLER_ASAP7_75t_R FILLER_0_186_1068 ();
 FILLER_ASAP7_75t_R FILLER_0_186_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1106 ();
 DECAPx6_ASAP7_75t_R FILLER_0_186_1128 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_1142 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_186_1148 ();
 FILLER_ASAP7_75t_R FILLER_0_186_1155 ();
 DECAPx4_ASAP7_75t_R FILLER_0_186_1167 ();
 FILLER_ASAP7_75t_R FILLER_0_186_1183 ();
 DECAPx4_ASAP7_75t_R FILLER_0_186_1191 ();
 FILLER_ASAP7_75t_R FILLER_0_186_1201 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_186_1203 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_1211 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_186_1217 ();
 FILLER_ASAP7_75t_R FILLER_0_186_1225 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_186_1227 ();
 DECAPx1_ASAP7_75t_R FILLER_0_186_1234 ();
 FILLER_ASAP7_75t_R FILLER_0_186_1249 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_186_1251 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_1263 ();
 FILLER_ASAP7_75t_R FILLER_0_186_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1305 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1327 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1349 ();
 DECAPx4_ASAP7_75t_R FILLER_0_186_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_186_1381 ();
 DECAPx6_ASAP7_75t_R FILLER_0_187_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_22 ();
 FILLER_ASAP7_75t_R FILLER_0_187_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_187_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_187_61 ();
 DECAPx2_ASAP7_75t_R FILLER_0_187_71 ();
 DECAPx6_ASAP7_75t_R FILLER_0_187_83 ();
 FILLER_ASAP7_75t_R FILLER_0_187_108 ();
 DECAPx4_ASAP7_75t_R FILLER_0_187_117 ();
 FILLER_ASAP7_75t_R FILLER_0_187_127 ();
 DECAPx6_ASAP7_75t_R FILLER_0_187_135 ();
 FILLER_ASAP7_75t_R FILLER_0_187_149 ();
 FILLER_ASAP7_75t_R FILLER_0_187_162 ();
 DECAPx4_ASAP7_75t_R FILLER_0_187_170 ();
 DECAPx2_ASAP7_75t_R FILLER_0_187_191 ();
 DECAPx2_ASAP7_75t_R FILLER_0_187_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_187_209 ();
 DECAPx1_ASAP7_75t_R FILLER_0_187_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_187_226 ();
 DECAPx6_ASAP7_75t_R FILLER_0_187_233 ();
 FILLER_ASAP7_75t_R FILLER_0_187_253 ();
 FILLER_ASAP7_75t_R FILLER_0_187_261 ();
 DECAPx2_ASAP7_75t_R FILLER_0_187_269 ();
 FILLER_ASAP7_75t_R FILLER_0_187_275 ();
 FILLER_ASAP7_75t_R FILLER_0_187_283 ();
 FILLER_ASAP7_75t_R FILLER_0_187_291 ();
 FILLER_ASAP7_75t_R FILLER_0_187_299 ();
 DECAPx4_ASAP7_75t_R FILLER_0_187_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_187_319 ();
 FILLER_ASAP7_75t_R FILLER_0_187_325 ();
 FILLER_ASAP7_75t_R FILLER_0_187_337 ();
 FILLER_ASAP7_75t_R FILLER_0_187_349 ();
 FILLER_ASAP7_75t_R FILLER_0_187_361 ();
 FILLER_ASAP7_75t_R FILLER_0_187_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_187_370 ();
 DECAPx6_ASAP7_75t_R FILLER_0_187_374 ();
 DECAPx2_ASAP7_75t_R FILLER_0_187_388 ();
 DECAPx1_ASAP7_75t_R FILLER_0_187_400 ();
 DECAPx1_ASAP7_75t_R FILLER_0_187_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_187_414 ();
 DECAPx1_ASAP7_75t_R FILLER_0_187_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_187_427 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_434 ();
 DECAPx1_ASAP7_75t_R FILLER_0_187_456 ();
 FILLER_ASAP7_75t_R FILLER_0_187_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_187_468 ();
 FILLER_ASAP7_75t_R FILLER_0_187_477 ();
 FILLER_ASAP7_75t_R FILLER_0_187_482 ();
 FILLER_ASAP7_75t_R FILLER_0_187_490 ();
 FILLER_ASAP7_75t_R FILLER_0_187_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_187_500 ();
 DECAPx2_ASAP7_75t_R FILLER_0_187_509 ();
 FILLER_ASAP7_75t_R FILLER_0_187_515 ();
 DECAPx2_ASAP7_75t_R FILLER_0_187_523 ();
 DECAPx6_ASAP7_75t_R FILLER_0_187_535 ();
 FILLER_ASAP7_75t_R FILLER_0_187_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_187_558 ();
 FILLER_ASAP7_75t_R FILLER_0_187_564 ();
 FILLER_ASAP7_75t_R FILLER_0_187_584 ();
 DECAPx2_ASAP7_75t_R FILLER_0_187_600 ();
 FILLER_ASAP7_75t_R FILLER_0_187_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_187_608 ();
 FILLER_ASAP7_75t_R FILLER_0_187_612 ();
 FILLER_ASAP7_75t_R FILLER_0_187_622 ();
 DECAPx1_ASAP7_75t_R FILLER_0_187_630 ();
 DECAPx2_ASAP7_75t_R FILLER_0_187_640 ();
 FILLER_ASAP7_75t_R FILLER_0_187_646 ();
 FILLER_ASAP7_75t_R FILLER_0_187_656 ();
 DECAPx2_ASAP7_75t_R FILLER_0_187_668 ();
 FILLER_ASAP7_75t_R FILLER_0_187_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_187_676 ();
 DECAPx4_ASAP7_75t_R FILLER_0_187_680 ();
 FILLER_ASAP7_75t_R FILLER_0_187_690 ();
 DECAPx1_ASAP7_75t_R FILLER_0_187_697 ();
 FILLER_ASAP7_75t_R FILLER_0_187_711 ();
 FILLER_ASAP7_75t_R FILLER_0_187_723 ();
 FILLER_ASAP7_75t_R FILLER_0_187_737 ();
 FILLER_ASAP7_75t_R FILLER_0_187_759 ();
 DECAPx1_ASAP7_75t_R FILLER_0_187_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_187_771 ();
 DECAPx6_ASAP7_75t_R FILLER_0_187_778 ();
 FILLER_ASAP7_75t_R FILLER_0_187_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_187_794 ();
 FILLER_ASAP7_75t_R FILLER_0_187_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_187_807 ();
 FILLER_ASAP7_75t_R FILLER_0_187_813 ();
 DECAPx2_ASAP7_75t_R FILLER_0_187_820 ();
 FILLER_ASAP7_75t_R FILLER_0_187_836 ();
 FILLER_ASAP7_75t_R FILLER_0_187_843 ();
 FILLER_ASAP7_75t_R FILLER_0_187_849 ();
 FILLER_ASAP7_75t_R FILLER_0_187_859 ();
 FILLER_ASAP7_75t_R FILLER_0_187_871 ();
 FILLER_ASAP7_75t_R FILLER_0_187_879 ();
 DECAPx1_ASAP7_75t_R FILLER_0_187_891 ();
 DECAPx2_ASAP7_75t_R FILLER_0_187_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_187_907 ();
 FILLER_ASAP7_75t_R FILLER_0_187_916 ();
 FILLER_ASAP7_75t_R FILLER_0_187_923 ();
 FILLER_ASAP7_75t_R FILLER_0_187_927 ();
 FILLER_ASAP7_75t_R FILLER_0_187_949 ();
 FILLER_ASAP7_75t_R FILLER_0_187_957 ();
 FILLER_ASAP7_75t_R FILLER_0_187_965 ();
 FILLER_ASAP7_75t_R FILLER_0_187_977 ();
 DECAPx1_ASAP7_75t_R FILLER_0_187_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_187_988 ();
 DECAPx6_ASAP7_75t_R FILLER_0_187_992 ();
 FILLER_ASAP7_75t_R FILLER_0_187_1016 ();
 FILLER_ASAP7_75t_R FILLER_0_187_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_187_1040 ();
 FILLER_ASAP7_75t_R FILLER_0_187_1046 ();
 FILLER_ASAP7_75t_R FILLER_0_187_1054 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_187_1084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1096 ();
 FILLER_ASAP7_75t_R FILLER_0_187_1118 ();
 FILLER_ASAP7_75t_R FILLER_0_187_1125 ();
 DECAPx2_ASAP7_75t_R FILLER_0_187_1133 ();
 FILLER_ASAP7_75t_R FILLER_0_187_1139 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1147 ();
 DECAPx1_ASAP7_75t_R FILLER_0_187_1169 ();
 FILLER_ASAP7_75t_R FILLER_0_187_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_187_1182 ();
 FILLER_ASAP7_75t_R FILLER_0_187_1189 ();
 DECAPx2_ASAP7_75t_R FILLER_0_187_1199 ();
 FILLER_ASAP7_75t_R FILLER_0_187_1208 ();
 DECAPx6_ASAP7_75t_R FILLER_0_187_1222 ();
 DECAPx2_ASAP7_75t_R FILLER_0_187_1236 ();
 FILLER_ASAP7_75t_R FILLER_0_187_1248 ();
 DECAPx1_ASAP7_75t_R FILLER_0_187_1257 ();
 FILLER_ASAP7_75t_R FILLER_0_187_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1281 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1303 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1325 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1347 ();
 DECAPx4_ASAP7_75t_R FILLER_0_187_1369 ();
 FILLER_ASAP7_75t_R FILLER_0_187_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_187_1381 ();
 DECAPx4_ASAP7_75t_R FILLER_0_188_2 ();
 FILLER_ASAP7_75t_R FILLER_0_188_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_14 ();
 DECAPx1_ASAP7_75t_R FILLER_0_188_31 ();
 FILLER_ASAP7_75t_R FILLER_0_188_41 ();
 FILLER_ASAP7_75t_R FILLER_0_188_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_51 ();
 DECAPx4_ASAP7_75t_R FILLER_0_188_58 ();
 DECAPx4_ASAP7_75t_R FILLER_0_188_79 ();
 DECAPx6_ASAP7_75t_R FILLER_0_188_95 ();
 FILLER_ASAP7_75t_R FILLER_0_188_109 ();
 DECAPx4_ASAP7_75t_R FILLER_0_188_118 ();
 FILLER_ASAP7_75t_R FILLER_0_188_128 ();
 DECAPx2_ASAP7_75t_R FILLER_0_188_136 ();
 FILLER_ASAP7_75t_R FILLER_0_188_142 ();
 FILLER_ASAP7_75t_R FILLER_0_188_150 ();
 DECAPx2_ASAP7_75t_R FILLER_0_188_158 ();
 DECAPx1_ASAP7_75t_R FILLER_0_188_170 ();
 FILLER_ASAP7_75t_R FILLER_0_188_180 ();
 DECAPx2_ASAP7_75t_R FILLER_0_188_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_201 ();
 FILLER_ASAP7_75t_R FILLER_0_188_229 ();
 DECAPx4_ASAP7_75t_R FILLER_0_188_238 ();
 FILLER_ASAP7_75t_R FILLER_0_188_248 ();
 DECAPx2_ASAP7_75t_R FILLER_0_188_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_264 ();
 DECAPx4_ASAP7_75t_R FILLER_0_188_273 ();
 FILLER_ASAP7_75t_R FILLER_0_188_289 ();
 FILLER_ASAP7_75t_R FILLER_0_188_297 ();
 FILLER_ASAP7_75t_R FILLER_0_188_305 ();
 DECAPx6_ASAP7_75t_R FILLER_0_188_313 ();
 FILLER_ASAP7_75t_R FILLER_0_188_337 ();
 FILLER_ASAP7_75t_R FILLER_0_188_345 ();
 FILLER_ASAP7_75t_R FILLER_0_188_357 ();
 FILLER_ASAP7_75t_R FILLER_0_188_365 ();
 FILLER_ASAP7_75t_R FILLER_0_188_373 ();
 FILLER_ASAP7_75t_R FILLER_0_188_381 ();
 FILLER_ASAP7_75t_R FILLER_0_188_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_391 ();
 DECAPx2_ASAP7_75t_R FILLER_0_188_395 ();
 FILLER_ASAP7_75t_R FILLER_0_188_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_403 ();
 FILLER_ASAP7_75t_R FILLER_0_188_411 ();
 FILLER_ASAP7_75t_R FILLER_0_188_420 ();
 FILLER_ASAP7_75t_R FILLER_0_188_430 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_438 ();
 FILLER_ASAP7_75t_R FILLER_0_188_460 ();
 DECAPx2_ASAP7_75t_R FILLER_0_188_464 ();
 FILLER_ASAP7_75t_R FILLER_0_188_470 ();
 FILLER_ASAP7_75t_R FILLER_0_188_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_480 ();
 DECAPx1_ASAP7_75t_R FILLER_0_188_487 ();
 DECAPx1_ASAP7_75t_R FILLER_0_188_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_502 ();
 FILLER_ASAP7_75t_R FILLER_0_188_509 ();
 DECAPx1_ASAP7_75t_R FILLER_0_188_517 ();
 DECAPx4_ASAP7_75t_R FILLER_0_188_524 ();
 FILLER_ASAP7_75t_R FILLER_0_188_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_542 ();
 FILLER_ASAP7_75t_R FILLER_0_188_549 ();
 DECAPx2_ASAP7_75t_R FILLER_0_188_559 ();
 FILLER_ASAP7_75t_R FILLER_0_188_565 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_577 ();
 DECAPx1_ASAP7_75t_R FILLER_0_188_599 ();
 FILLER_ASAP7_75t_R FILLER_0_188_611 ();
 DECAPx2_ASAP7_75t_R FILLER_0_188_621 ();
 FILLER_ASAP7_75t_R FILLER_0_188_633 ();
 DECAPx2_ASAP7_75t_R FILLER_0_188_641 ();
 FILLER_ASAP7_75t_R FILLER_0_188_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_649 ();
 DECAPx4_ASAP7_75t_R FILLER_0_188_656 ();
 FILLER_ASAP7_75t_R FILLER_0_188_672 ();
 DECAPx4_ASAP7_75t_R FILLER_0_188_680 ();
 FILLER_ASAP7_75t_R FILLER_0_188_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_692 ();
 FILLER_ASAP7_75t_R FILLER_0_188_700 ();
 FILLER_ASAP7_75t_R FILLER_0_188_708 ();
 DECAPx2_ASAP7_75t_R FILLER_0_188_715 ();
 FILLER_ASAP7_75t_R FILLER_0_188_721 ();
 FILLER_ASAP7_75t_R FILLER_0_188_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_735 ();
 FILLER_ASAP7_75t_R FILLER_0_188_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_748 ();
 FILLER_ASAP7_75t_R FILLER_0_188_756 ();
 FILLER_ASAP7_75t_R FILLER_0_188_764 ();
 DECAPx1_ASAP7_75t_R FILLER_0_188_772 ();
 FILLER_ASAP7_75t_R FILLER_0_188_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_785 ();
 FILLER_ASAP7_75t_R FILLER_0_188_791 ();
 DECAPx4_ASAP7_75t_R FILLER_0_188_803 ();
 FILLER_ASAP7_75t_R FILLER_0_188_819 ();
 DECAPx6_ASAP7_75t_R FILLER_0_188_841 ();
 DECAPx1_ASAP7_75t_R FILLER_0_188_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_859 ();
 FILLER_ASAP7_75t_R FILLER_0_188_865 ();
 FILLER_ASAP7_75t_R FILLER_0_188_872 ();
 FILLER_ASAP7_75t_R FILLER_0_188_881 ();
 FILLER_ASAP7_75t_R FILLER_0_188_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_891 ();
 DECAPx2_ASAP7_75t_R FILLER_0_188_902 ();
 FILLER_ASAP7_75t_R FILLER_0_188_908 ();
 DECAPx6_ASAP7_75t_R FILLER_0_188_916 ();
 DECAPx2_ASAP7_75t_R FILLER_0_188_930 ();
 FILLER_ASAP7_75t_R FILLER_0_188_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_945 ();
 FILLER_ASAP7_75t_R FILLER_0_188_958 ();
 DECAPx2_ASAP7_75t_R FILLER_0_188_966 ();
 DECAPx6_ASAP7_75t_R FILLER_0_188_978 ();
 DECAPx1_ASAP7_75t_R FILLER_0_188_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_996 ();
 DECAPx2_ASAP7_75t_R FILLER_0_188_1007 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_1013 ();
 DECAPx6_ASAP7_75t_R FILLER_0_188_1021 ();
 DECAPx1_ASAP7_75t_R FILLER_0_188_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_1039 ();
 FILLER_ASAP7_75t_R FILLER_0_188_1050 ();
 FILLER_ASAP7_75t_R FILLER_0_188_1062 ();
 FILLER_ASAP7_75t_R FILLER_0_188_1070 ();
 DECAPx2_ASAP7_75t_R FILLER_0_188_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_0_188_1095 ();
 FILLER_ASAP7_75t_R FILLER_0_188_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_1103 ();
 FILLER_ASAP7_75t_R FILLER_0_188_1110 ();
 DECAPx1_ASAP7_75t_R FILLER_0_188_1118 ();
 FILLER_ASAP7_75t_R FILLER_0_188_1128 ();
 DECAPx4_ASAP7_75t_R FILLER_0_188_1136 ();
 FILLER_ASAP7_75t_R FILLER_0_188_1146 ();
 FILLER_ASAP7_75t_R FILLER_0_188_1155 ();
 DECAPx4_ASAP7_75t_R FILLER_0_188_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_1173 ();
 DECAPx6_ASAP7_75t_R FILLER_0_188_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_188_1200 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_1202 ();
 FILLER_ASAP7_75t_R FILLER_0_188_1209 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_1211 ();
 DECAPx1_ASAP7_75t_R FILLER_0_188_1220 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_1224 ();
 DECAPx1_ASAP7_75t_R FILLER_0_188_1231 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_1235 ();
 DECAPx4_ASAP7_75t_R FILLER_0_188_1242 ();
 FILLER_ASAP7_75t_R FILLER_0_188_1252 ();
 DECAPx2_ASAP7_75t_R FILLER_0_188_1257 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188_1263 ();
 FILLER_ASAP7_75t_R FILLER_0_188_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1346 ();
 DECAPx6_ASAP7_75t_R FILLER_0_188_1368 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_8 ();
 FILLER_ASAP7_75t_R FILLER_0_189_15 ();
 FILLER_ASAP7_75t_R FILLER_0_189_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_25 ();
 FILLER_ASAP7_75t_R FILLER_0_189_32 ();
 FILLER_ASAP7_75t_R FILLER_0_189_40 ();
 DECAPx1_ASAP7_75t_R FILLER_0_189_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_51 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_58 ();
 FILLER_ASAP7_75t_R FILLER_0_189_64 ();
 FILLER_ASAP7_75t_R FILLER_0_189_69 ();
 DECAPx4_ASAP7_75t_R FILLER_0_189_77 ();
 FILLER_ASAP7_75t_R FILLER_0_189_87 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_101 ();
 DECAPx1_ASAP7_75t_R FILLER_0_189_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_112 ();
 FILLER_ASAP7_75t_R FILLER_0_189_119 ();
 FILLER_ASAP7_75t_R FILLER_0_189_127 ();
 DECAPx4_ASAP7_75t_R FILLER_0_189_135 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_156 ();
 FILLER_ASAP7_75t_R FILLER_0_189_178 ();
 FILLER_ASAP7_75t_R FILLER_0_189_186 ();
 DECAPx1_ASAP7_75t_R FILLER_0_189_193 ();
 DECAPx6_ASAP7_75t_R FILLER_0_189_208 ();
 FILLER_ASAP7_75t_R FILLER_0_189_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_224 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_233 ();
 FILLER_ASAP7_75t_R FILLER_0_189_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_241 ();
 FILLER_ASAP7_75t_R FILLER_0_189_248 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_256 ();
 FILLER_ASAP7_75t_R FILLER_0_189_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_264 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_271 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_283 ();
 DECAPx4_ASAP7_75t_R FILLER_0_189_305 ();
 DECAPx1_ASAP7_75t_R FILLER_0_189_321 ();
 DECAPx1_ASAP7_75t_R FILLER_0_189_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_335 ();
 FILLER_ASAP7_75t_R FILLER_0_189_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_348 ();
 DECAPx6_ASAP7_75t_R FILLER_0_189_356 ();
 DECAPx1_ASAP7_75t_R FILLER_0_189_378 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_388 ();
 FILLER_ASAP7_75t_R FILLER_0_189_400 ();
 DECAPx1_ASAP7_75t_R FILLER_0_189_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_412 ();
 FILLER_ASAP7_75t_R FILLER_0_189_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_421 ();
 FILLER_ASAP7_75t_R FILLER_0_189_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_430 ();
 DECAPx6_ASAP7_75t_R FILLER_0_189_437 ();
 FILLER_ASAP7_75t_R FILLER_0_189_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_453 ();
 FILLER_ASAP7_75t_R FILLER_0_189_464 ();
 DECAPx1_ASAP7_75t_R FILLER_0_189_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_476 ();
 FILLER_ASAP7_75t_R FILLER_0_189_483 ();
 DECAPx1_ASAP7_75t_R FILLER_0_189_491 ();
 DECAPx1_ASAP7_75t_R FILLER_0_189_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_505 ();
 FILLER_ASAP7_75t_R FILLER_0_189_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_515 ();
 DECAPx1_ASAP7_75t_R FILLER_0_189_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_526 ();
 FILLER_ASAP7_75t_R FILLER_0_189_533 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_543 ();
 DECAPx4_ASAP7_75t_R FILLER_0_189_565 ();
 FILLER_ASAP7_75t_R FILLER_0_189_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_577 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_584 ();
 FILLER_ASAP7_75t_R FILLER_0_189_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_592 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_599 ();
 FILLER_ASAP7_75t_R FILLER_0_189_611 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_619 ();
 FILLER_ASAP7_75t_R FILLER_0_189_625 ();
 DECAPx6_ASAP7_75t_R FILLER_0_189_633 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_653 ();
 DECAPx6_ASAP7_75t_R FILLER_0_189_675 ();
 FILLER_ASAP7_75t_R FILLER_0_189_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_691 ();
 FILLER_ASAP7_75t_R FILLER_0_189_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_699 ();
 FILLER_ASAP7_75t_R FILLER_0_189_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_722 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_733 ();
 FILLER_ASAP7_75t_R FILLER_0_189_739 ();
 FILLER_ASAP7_75t_R FILLER_0_189_751 ();
 DECAPx4_ASAP7_75t_R FILLER_0_189_758 ();
 FILLER_ASAP7_75t_R FILLER_0_189_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_770 ();
 DECAPx6_ASAP7_75t_R FILLER_0_189_781 ();
 DECAPx1_ASAP7_75t_R FILLER_0_189_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_799 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_811 ();
 DECAPx1_ASAP7_75t_R FILLER_0_189_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_826 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_833 ();
 FILLER_ASAP7_75t_R FILLER_0_189_844 ();
 DECAPx4_ASAP7_75t_R FILLER_0_189_849 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_865 ();
 FILLER_ASAP7_75t_R FILLER_0_189_871 ();
 FILLER_ASAP7_75t_R FILLER_0_189_879 ();
 DECAPx1_ASAP7_75t_R FILLER_0_189_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_891 ();
 FILLER_ASAP7_75t_R FILLER_0_189_900 ();
 DECAPx1_ASAP7_75t_R FILLER_0_189_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_911 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_924 ();
 DECAPx6_ASAP7_75t_R FILLER_0_189_927 ();
 DECAPx1_ASAP7_75t_R FILLER_0_189_941 ();
 FILLER_ASAP7_75t_R FILLER_0_189_951 ();
 FILLER_ASAP7_75t_R FILLER_0_189_959 ();
 FILLER_ASAP7_75t_R FILLER_0_189_971 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_976 ();
 DECAPx1_ASAP7_75t_R FILLER_0_189_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_1002 ();
 FILLER_ASAP7_75t_R FILLER_0_189_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_1011 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_1022 ();
 FILLER_ASAP7_75t_R FILLER_0_189_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_1030 ();
 DECAPx1_ASAP7_75t_R FILLER_0_189_1037 ();
 FILLER_ASAP7_75t_R FILLER_0_189_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_1053 ();
 FILLER_ASAP7_75t_R FILLER_0_189_1064 ();
 FILLER_ASAP7_75t_R FILLER_0_189_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_1076 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_1083 ();
 FILLER_ASAP7_75t_R FILLER_0_189_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_1091 ();
 FILLER_ASAP7_75t_R FILLER_0_189_1098 ();
 DECAPx1_ASAP7_75t_R FILLER_0_189_1105 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_1117 ();
 FILLER_ASAP7_75t_R FILLER_0_189_1123 ();
 FILLER_ASAP7_75t_R FILLER_0_189_1131 ();
 FILLER_ASAP7_75t_R FILLER_0_189_1139 ();
 FILLER_ASAP7_75t_R FILLER_0_189_1148 ();
 FILLER_ASAP7_75t_R FILLER_0_189_1156 ();
 DECAPx6_ASAP7_75t_R FILLER_0_189_1161 ();
 FILLER_ASAP7_75t_R FILLER_0_189_1175 ();
 DECAPx6_ASAP7_75t_R FILLER_0_189_1185 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_1199 ();
 DECAPx1_ASAP7_75t_R FILLER_0_189_1210 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189_1225 ();
 FILLER_ASAP7_75t_R FILLER_0_189_1232 ();
 DECAPx1_ASAP7_75t_R FILLER_0_189_1246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_189_1366 ();
 FILLER_ASAP7_75t_R FILLER_0_189_1380 ();
 DECAPx1_ASAP7_75t_R FILLER_0_190_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_6 ();
 DECAPx2_ASAP7_75t_R FILLER_0_190_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_19 ();
 DECAPx2_ASAP7_75t_R FILLER_0_190_27 ();
 FILLER_ASAP7_75t_R FILLER_0_190_33 ();
 FILLER_ASAP7_75t_R FILLER_0_190_40 ();
 FILLER_ASAP7_75t_R FILLER_0_190_48 ();
 DECAPx4_ASAP7_75t_R FILLER_0_190_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_66 ();
 FILLER_ASAP7_75t_R FILLER_0_190_73 ();
 DECAPx2_ASAP7_75t_R FILLER_0_190_81 ();
 DECAPx4_ASAP7_75t_R FILLER_0_190_93 ();
 FILLER_ASAP7_75t_R FILLER_0_190_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_105 ();
 DECAPx10_ASAP7_75t_R FILLER_0_190_112 ();
 DECAPx2_ASAP7_75t_R FILLER_0_190_134 ();
 FILLER_ASAP7_75t_R FILLER_0_190_146 ();
 FILLER_ASAP7_75t_R FILLER_0_190_154 ();
 FILLER_ASAP7_75t_R FILLER_0_190_162 ();
 FILLER_ASAP7_75t_R FILLER_0_190_170 ();
 DECAPx2_ASAP7_75t_R FILLER_0_190_180 ();
 FILLER_ASAP7_75t_R FILLER_0_190_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_188 ();
 FILLER_ASAP7_75t_R FILLER_0_190_197 ();
 DECAPx6_ASAP7_75t_R FILLER_0_190_205 ();
 DECAPx1_ASAP7_75t_R FILLER_0_190_219 ();
 DECAPx4_ASAP7_75t_R FILLER_0_190_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_239 ();
 FILLER_ASAP7_75t_R FILLER_0_190_246 ();
 FILLER_ASAP7_75t_R FILLER_0_190_254 ();
 DECAPx1_ASAP7_75t_R FILLER_0_190_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_266 ();
 DECAPx1_ASAP7_75t_R FILLER_0_190_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_279 ();
 FILLER_ASAP7_75t_R FILLER_0_190_287 ();
 DECAPx2_ASAP7_75t_R FILLER_0_190_296 ();
 FILLER_ASAP7_75t_R FILLER_0_190_305 ();
 DECAPx4_ASAP7_75t_R FILLER_0_190_314 ();
 FILLER_ASAP7_75t_R FILLER_0_190_324 ();
 FILLER_ASAP7_75t_R FILLER_0_190_329 ();
 FILLER_ASAP7_75t_R FILLER_0_190_337 ();
 FILLER_ASAP7_75t_R FILLER_0_190_349 ();
 DECAPx2_ASAP7_75t_R FILLER_0_190_356 ();
 FILLER_ASAP7_75t_R FILLER_0_190_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_364 ();
 FILLER_ASAP7_75t_R FILLER_0_190_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_373 ();
 DECAPx1_ASAP7_75t_R FILLER_0_190_380 ();
 FILLER_ASAP7_75t_R FILLER_0_190_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_394 ();
 DECAPx1_ASAP7_75t_R FILLER_0_190_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_405 ();
 FILLER_ASAP7_75t_R FILLER_0_190_409 ();
 DECAPx2_ASAP7_75t_R FILLER_0_190_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_423 ();
 DECAPx10_ASAP7_75t_R FILLER_0_190_431 ();
 DECAPx2_ASAP7_75t_R FILLER_0_190_453 ();
 FILLER_ASAP7_75t_R FILLER_0_190_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_461 ();
 FILLER_ASAP7_75t_R FILLER_0_190_464 ();
 FILLER_ASAP7_75t_R FILLER_0_190_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_477 ();
 DECAPx1_ASAP7_75t_R FILLER_0_190_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_485 ();
 FILLER_ASAP7_75t_R FILLER_0_190_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_495 ();
 DECAPx4_ASAP7_75t_R FILLER_0_190_502 ();
 FILLER_ASAP7_75t_R FILLER_0_190_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_514 ();
 FILLER_ASAP7_75t_R FILLER_0_190_521 ();
 DECAPx2_ASAP7_75t_R FILLER_0_190_526 ();
 FILLER_ASAP7_75t_R FILLER_0_190_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_534 ();
 FILLER_ASAP7_75t_R FILLER_0_190_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_540 ();
 FILLER_ASAP7_75t_R FILLER_0_190_544 ();
 DECAPx6_ASAP7_75t_R FILLER_0_190_552 ();
 DECAPx2_ASAP7_75t_R FILLER_0_190_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_572 ();
 FILLER_ASAP7_75t_R FILLER_0_190_583 ();
 DECAPx6_ASAP7_75t_R FILLER_0_190_591 ();
 DECAPx1_ASAP7_75t_R FILLER_0_190_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_609 ();
 FILLER_ASAP7_75t_R FILLER_0_190_618 ();
 DECAPx4_ASAP7_75t_R FILLER_0_190_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_190_658 ();
 DECAPx2_ASAP7_75t_R FILLER_0_190_680 ();
 FILLER_ASAP7_75t_R FILLER_0_190_686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_190_708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_190_730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_190_752 ();
 FILLER_ASAP7_75t_R FILLER_0_190_766 ();
 FILLER_ASAP7_75t_R FILLER_0_190_775 ();
 FILLER_ASAP7_75t_R FILLER_0_190_783 ();
 FILLER_ASAP7_75t_R FILLER_0_190_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_794 ();
 FILLER_ASAP7_75t_R FILLER_0_190_805 ();
 FILLER_ASAP7_75t_R FILLER_0_190_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_815 ();
 FILLER_ASAP7_75t_R FILLER_0_190_819 ();
 FILLER_ASAP7_75t_R FILLER_0_190_841 ();
 DECAPx2_ASAP7_75t_R FILLER_0_190_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_855 ();
 FILLER_ASAP7_75t_R FILLER_0_190_864 ();
 DECAPx4_ASAP7_75t_R FILLER_0_190_872 ();
 FILLER_ASAP7_75t_R FILLER_0_190_888 ();
 FILLER_ASAP7_75t_R FILLER_0_190_901 ();
 FILLER_ASAP7_75t_R FILLER_0_190_913 ();
 FILLER_ASAP7_75t_R FILLER_0_190_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_190_938 ();
 FILLER_ASAP7_75t_R FILLER_0_190_960 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_962 ();
 DECAPx4_ASAP7_75t_R FILLER_0_190_969 ();
 FILLER_ASAP7_75t_R FILLER_0_190_1000 ();
 DECAPx4_ASAP7_75t_R FILLER_0_190_1012 ();
 FILLER_ASAP7_75t_R FILLER_0_190_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_1024 ();
 FILLER_ASAP7_75t_R FILLER_0_190_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_1032 ();
 FILLER_ASAP7_75t_R FILLER_0_190_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_1045 ();
 FILLER_ASAP7_75t_R FILLER_0_190_1056 ();
 DECAPx10_ASAP7_75t_R FILLER_0_190_1064 ();
 FILLER_ASAP7_75t_R FILLER_0_190_1086 ();
 FILLER_ASAP7_75t_R FILLER_0_190_1095 ();
 DECAPx2_ASAP7_75t_R FILLER_0_190_1103 ();
 DECAPx1_ASAP7_75t_R FILLER_0_190_1115 ();
 FILLER_ASAP7_75t_R FILLER_0_190_1125 ();
 DECAPx6_ASAP7_75t_R FILLER_0_190_1130 ();
 DECAPx6_ASAP7_75t_R FILLER_0_190_1154 ();
 DECAPx1_ASAP7_75t_R FILLER_0_190_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190_1172 ();
 FILLER_ASAP7_75t_R FILLER_0_190_1178 ();
 FILLER_ASAP7_75t_R FILLER_0_190_1188 ();
 DECAPx10_ASAP7_75t_R FILLER_0_190_1200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_190_1222 ();
 DECAPx6_ASAP7_75t_R FILLER_0_190_1250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_190_1280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_190_1302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_190_1324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_190_1346 ();
 DECAPx6_ASAP7_75t_R FILLER_0_190_1368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_191_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_191_24 ();
 DECAPx2_ASAP7_75t_R FILLER_0_191_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_40 ();
 DECAPx1_ASAP7_75t_R FILLER_0_191_47 ();
 DECAPx10_ASAP7_75t_R FILLER_0_191_57 ();
 DECAPx2_ASAP7_75t_R FILLER_0_191_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_85 ();
 DECAPx6_ASAP7_75t_R FILLER_0_191_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_106 ();
 FILLER_ASAP7_75t_R FILLER_0_191_113 ();
 DECAPx4_ASAP7_75t_R FILLER_0_191_121 ();
 DECAPx2_ASAP7_75t_R FILLER_0_191_137 ();
 DECAPx1_ASAP7_75t_R FILLER_0_191_146 ();
 DECAPx2_ASAP7_75t_R FILLER_0_191_156 ();
 FILLER_ASAP7_75t_R FILLER_0_191_168 ();
 DECAPx6_ASAP7_75t_R FILLER_0_191_176 ();
 DECAPx2_ASAP7_75t_R FILLER_0_191_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_196 ();
 FILLER_ASAP7_75t_R FILLER_0_191_203 ();
 DECAPx10_ASAP7_75t_R FILLER_0_191_208 ();
 DECAPx2_ASAP7_75t_R FILLER_0_191_230 ();
 FILLER_ASAP7_75t_R FILLER_0_191_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_238 ();
 DECAPx1_ASAP7_75t_R FILLER_0_191_249 ();
 DECAPx6_ASAP7_75t_R FILLER_0_191_273 ();
 DECAPx6_ASAP7_75t_R FILLER_0_191_307 ();
 FILLER_ASAP7_75t_R FILLER_0_191_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_323 ();
 DECAPx2_ASAP7_75t_R FILLER_0_191_330 ();
 FILLER_ASAP7_75t_R FILLER_0_191_346 ();
 DECAPx2_ASAP7_75t_R FILLER_0_191_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_359 ();
 DECAPx1_ASAP7_75t_R FILLER_0_191_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_370 ();
 DECAPx6_ASAP7_75t_R FILLER_0_191_379 ();
 DECAPx1_ASAP7_75t_R FILLER_0_191_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_397 ();
 DECAPx2_ASAP7_75t_R FILLER_0_191_404 ();
 FILLER_ASAP7_75t_R FILLER_0_191_416 ();
 FILLER_ASAP7_75t_R FILLER_0_191_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_191_433 ();
 DECAPx2_ASAP7_75t_R FILLER_0_191_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_461 ();
 DECAPx2_ASAP7_75t_R FILLER_0_191_468 ();
 DECAPx2_ASAP7_75t_R FILLER_0_191_480 ();
 FILLER_ASAP7_75t_R FILLER_0_191_492 ();
 FILLER_ASAP7_75t_R FILLER_0_191_500 ();
 DECAPx2_ASAP7_75t_R FILLER_0_191_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_511 ();
 FILLER_ASAP7_75t_R FILLER_0_191_515 ();
 DECAPx1_ASAP7_75t_R FILLER_0_191_525 ();
 DECAPx2_ASAP7_75t_R FILLER_0_191_537 ();
 FILLER_ASAP7_75t_R FILLER_0_191_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_545 ();
 DECAPx1_ASAP7_75t_R FILLER_0_191_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_558 ();
 FILLER_ASAP7_75t_R FILLER_0_191_562 ();
 FILLER_ASAP7_75t_R FILLER_0_191_570 ();
 DECAPx2_ASAP7_75t_R FILLER_0_191_575 ();
 FILLER_ASAP7_75t_R FILLER_0_191_589 ();
 FILLER_ASAP7_75t_R FILLER_0_191_598 ();
 FILLER_ASAP7_75t_R FILLER_0_191_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_608 ();
 DECAPx6_ASAP7_75t_R FILLER_0_191_615 ();
 FILLER_ASAP7_75t_R FILLER_0_191_629 ();
 FILLER_ASAP7_75t_R FILLER_0_191_634 ();
 FILLER_ASAP7_75t_R FILLER_0_191_642 ();
 FILLER_ASAP7_75t_R FILLER_0_191_650 ();
 FILLER_ASAP7_75t_R FILLER_0_191_658 ();
 DECAPx10_ASAP7_75t_R FILLER_0_191_666 ();
 FILLER_ASAP7_75t_R FILLER_0_191_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_700 ();
 FILLER_ASAP7_75t_R FILLER_0_191_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_713 ();
 FILLER_ASAP7_75t_R FILLER_0_191_724 ();
 FILLER_ASAP7_75t_R FILLER_0_191_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_738 ();
 FILLER_ASAP7_75t_R FILLER_0_191_759 ();
 FILLER_ASAP7_75t_R FILLER_0_191_768 ();
 FILLER_ASAP7_75t_R FILLER_0_191_775 ();
 DECAPx2_ASAP7_75t_R FILLER_0_191_787 ();
 FILLER_ASAP7_75t_R FILLER_0_191_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_795 ();
 DECAPx6_ASAP7_75t_R FILLER_0_191_806 ();
 FILLER_ASAP7_75t_R FILLER_0_191_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_822 ();
 DECAPx4_ASAP7_75t_R FILLER_0_191_833 ();
 DECAPx2_ASAP7_75t_R FILLER_0_191_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_856 ();
 FILLER_ASAP7_75t_R FILLER_0_191_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_865 ();
 FILLER_ASAP7_75t_R FILLER_0_191_874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_191_882 ();
 DECAPx2_ASAP7_75t_R FILLER_0_191_904 ();
 FILLER_ASAP7_75t_R FILLER_0_191_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_912 ();
 DECAPx2_ASAP7_75t_R FILLER_0_191_919 ();
 FILLER_ASAP7_75t_R FILLER_0_191_927 ();
 FILLER_ASAP7_75t_R FILLER_0_191_935 ();
 FILLER_ASAP7_75t_R FILLER_0_191_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_944 ();
 FILLER_ASAP7_75t_R FILLER_0_191_951 ();
 DECAPx2_ASAP7_75t_R FILLER_0_191_959 ();
 FILLER_ASAP7_75t_R FILLER_0_191_965 ();
 FILLER_ASAP7_75t_R FILLER_0_191_973 ();
 FILLER_ASAP7_75t_R FILLER_0_191_981 ();
 DECAPx10_ASAP7_75t_R FILLER_0_191_986 ();
 FILLER_ASAP7_75t_R FILLER_0_191_1008 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_1010 ();
 FILLER_ASAP7_75t_R FILLER_0_191_1021 ();
 FILLER_ASAP7_75t_R FILLER_0_191_1033 ();
 FILLER_ASAP7_75t_R FILLER_0_191_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_1047 ();
 DECAPx2_ASAP7_75t_R FILLER_0_191_1058 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_1064 ();
 DECAPx10_ASAP7_75t_R FILLER_0_191_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_1093 ();
 DECAPx1_ASAP7_75t_R FILLER_0_191_1104 ();
 FILLER_ASAP7_75t_R FILLER_0_191_1114 ();
 FILLER_ASAP7_75t_R FILLER_0_191_1127 ();
 DECAPx4_ASAP7_75t_R FILLER_0_191_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_1145 ();
 DECAPx1_ASAP7_75t_R FILLER_0_191_1152 ();
 FILLER_ASAP7_75t_R FILLER_0_191_1162 ();
 FILLER_ASAP7_75t_R FILLER_0_191_1174 ();
 DECAPx2_ASAP7_75t_R FILLER_0_191_1181 ();
 FILLER_ASAP7_75t_R FILLER_0_191_1193 ();
 FILLER_ASAP7_75t_R FILLER_0_191_1198 ();
 DECAPx2_ASAP7_75t_R FILLER_0_191_1203 ();
 FILLER_ASAP7_75t_R FILLER_0_191_1209 ();
 FILLER_ASAP7_75t_R FILLER_0_191_1221 ();
 DECAPx6_ASAP7_75t_R FILLER_0_191_1229 ();
 DECAPx1_ASAP7_75t_R FILLER_0_191_1243 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191_1247 ();
 FILLER_ASAP7_75t_R FILLER_0_191_1260 ();
 FILLER_ASAP7_75t_R FILLER_0_191_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_0_191_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_191_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_191_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_191_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_191_1366 ();
 FILLER_ASAP7_75t_R FILLER_0_191_1380 ();
 DECAPx4_ASAP7_75t_R FILLER_0_192_2 ();
 FILLER_ASAP7_75t_R FILLER_0_192_12 ();
 DECAPx1_ASAP7_75t_R FILLER_0_192_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_24 ();
 DECAPx1_ASAP7_75t_R FILLER_0_192_31 ();
 FILLER_ASAP7_75t_R FILLER_0_192_41 ();
 DECAPx1_ASAP7_75t_R FILLER_0_192_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_53 ();
 FILLER_ASAP7_75t_R FILLER_0_192_60 ();
 DECAPx1_ASAP7_75t_R FILLER_0_192_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_72 ();
 DECAPx4_ASAP7_75t_R FILLER_0_192_83 ();
 DECAPx4_ASAP7_75t_R FILLER_0_192_99 ();
 FILLER_ASAP7_75t_R FILLER_0_192_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_111 ();
 FILLER_ASAP7_75t_R FILLER_0_192_118 ();
 DECAPx1_ASAP7_75t_R FILLER_0_192_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_130 ();
 DECAPx6_ASAP7_75t_R FILLER_0_192_137 ();
 FILLER_ASAP7_75t_R FILLER_0_192_151 ();
 DECAPx4_ASAP7_75t_R FILLER_0_192_159 ();
 FILLER_ASAP7_75t_R FILLER_0_192_169 ();
 DECAPx6_ASAP7_75t_R FILLER_0_192_177 ();
 DECAPx1_ASAP7_75t_R FILLER_0_192_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_195 ();
 FILLER_ASAP7_75t_R FILLER_0_192_202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_192_210 ();
 DECAPx4_ASAP7_75t_R FILLER_0_192_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_192_257 ();
 DECAPx2_ASAP7_75t_R FILLER_0_192_279 ();
 FILLER_ASAP7_75t_R FILLER_0_192_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_287 ();
 DECAPx1_ASAP7_75t_R FILLER_0_192_294 ();
 DECAPx4_ASAP7_75t_R FILLER_0_192_304 ();
 FILLER_ASAP7_75t_R FILLER_0_192_320 ();
 DECAPx4_ASAP7_75t_R FILLER_0_192_332 ();
 DECAPx2_ASAP7_75t_R FILLER_0_192_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_354 ();
 DECAPx4_ASAP7_75t_R FILLER_0_192_361 ();
 DECAPx1_ASAP7_75t_R FILLER_0_192_377 ();
 DECAPx2_ASAP7_75t_R FILLER_0_192_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_394 ();
 FILLER_ASAP7_75t_R FILLER_0_192_402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_192_412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_192_434 ();
 DECAPx2_ASAP7_75t_R FILLER_0_192_456 ();
 DECAPx6_ASAP7_75t_R FILLER_0_192_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_478 ();
 FILLER_ASAP7_75t_R FILLER_0_192_485 ();
 DECAPx10_ASAP7_75t_R FILLER_0_192_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_515 ();
 FILLER_ASAP7_75t_R FILLER_0_192_519 ();
 DECAPx4_ASAP7_75t_R FILLER_0_192_527 ();
 FILLER_ASAP7_75t_R FILLER_0_192_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_539 ();
 FILLER_ASAP7_75t_R FILLER_0_192_543 ();
 DECAPx2_ASAP7_75t_R FILLER_0_192_551 ();
 DECAPx2_ASAP7_75t_R FILLER_0_192_563 ();
 FILLER_ASAP7_75t_R FILLER_0_192_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_571 ();
 DECAPx1_ASAP7_75t_R FILLER_0_192_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_596 ();
 DECAPx2_ASAP7_75t_R FILLER_0_192_606 ();
 FILLER_ASAP7_75t_R FILLER_0_192_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_614 ();
 DECAPx1_ASAP7_75t_R FILLER_0_192_621 ();
 FILLER_ASAP7_75t_R FILLER_0_192_633 ();
 DECAPx1_ASAP7_75t_R FILLER_0_192_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_645 ();
 DECAPx1_ASAP7_75t_R FILLER_0_192_652 ();
 FILLER_ASAP7_75t_R FILLER_0_192_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_664 ();
 DECAPx6_ASAP7_75t_R FILLER_0_192_668 ();
 FILLER_ASAP7_75t_R FILLER_0_192_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_684 ();
 FILLER_ASAP7_75t_R FILLER_0_192_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_699 ();
 FILLER_ASAP7_75t_R FILLER_0_192_710 ();
 DECAPx1_ASAP7_75t_R FILLER_0_192_722 ();
 FILLER_ASAP7_75t_R FILLER_0_192_736 ();
 FILLER_ASAP7_75t_R FILLER_0_192_745 ();
 FILLER_ASAP7_75t_R FILLER_0_192_754 ();
 FILLER_ASAP7_75t_R FILLER_0_192_763 ();
 DECAPx1_ASAP7_75t_R FILLER_0_192_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_775 ();
 FILLER_ASAP7_75t_R FILLER_0_192_786 ();
 DECAPx4_ASAP7_75t_R FILLER_0_192_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_804 ();
 FILLER_ASAP7_75t_R FILLER_0_192_817 ();
 FILLER_ASAP7_75t_R FILLER_0_192_825 ();
 DECAPx10_ASAP7_75t_R FILLER_0_192_833 ();
 DECAPx2_ASAP7_75t_R FILLER_0_192_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_861 ();
 DECAPx4_ASAP7_75t_R FILLER_0_192_869 ();
 FILLER_ASAP7_75t_R FILLER_0_192_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_881 ();
 FILLER_ASAP7_75t_R FILLER_0_192_888 ();
 DECAPx4_ASAP7_75t_R FILLER_0_192_902 ();
 FILLER_ASAP7_75t_R FILLER_0_192_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_914 ();
 FILLER_ASAP7_75t_R FILLER_0_192_921 ();
 FILLER_ASAP7_75t_R FILLER_0_192_929 ();
 DECAPx2_ASAP7_75t_R FILLER_0_192_942 ();
 FILLER_ASAP7_75t_R FILLER_0_192_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_950 ();
 DECAPx2_ASAP7_75t_R FILLER_0_192_962 ();
 FILLER_ASAP7_75t_R FILLER_0_192_968 ();
 FILLER_ASAP7_75t_R FILLER_0_192_976 ();
 DECAPx4_ASAP7_75t_R FILLER_0_192_984 ();
 FILLER_ASAP7_75t_R FILLER_0_192_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_1006 ();
 DECAPx1_ASAP7_75t_R FILLER_0_192_1017 ();
 FILLER_ASAP7_75t_R FILLER_0_192_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_1033 ();
 DECAPx1_ASAP7_75t_R FILLER_0_192_1044 ();
 DECAPx10_ASAP7_75t_R FILLER_0_192_1058 ();
 FILLER_ASAP7_75t_R FILLER_0_192_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_1082 ();
 FILLER_ASAP7_75t_R FILLER_0_192_1093 ();
 DECAPx2_ASAP7_75t_R FILLER_0_192_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_1107 ();
 DECAPx1_ASAP7_75t_R FILLER_0_192_1118 ();
 FILLER_ASAP7_75t_R FILLER_0_192_1132 ();
 FILLER_ASAP7_75t_R FILLER_0_192_1141 ();
 FILLER_ASAP7_75t_R FILLER_0_192_1149 ();
 FILLER_ASAP7_75t_R FILLER_0_192_1163 ();
 FILLER_ASAP7_75t_R FILLER_0_192_1173 ();
 DECAPx1_ASAP7_75t_R FILLER_0_192_1181 ();
 FILLER_ASAP7_75t_R FILLER_0_192_1191 ();
 FILLER_ASAP7_75t_R FILLER_0_192_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192_1201 ();
 FILLER_ASAP7_75t_R FILLER_0_192_1208 ();
 DECAPx2_ASAP7_75t_R FILLER_0_192_1220 ();
 FILLER_ASAP7_75t_R FILLER_0_192_1232 ();
 FILLER_ASAP7_75t_R FILLER_0_192_1239 ();
 DECAPx4_ASAP7_75t_R FILLER_0_192_1246 ();
 FILLER_ASAP7_75t_R FILLER_0_192_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_192_1264 ();
 DECAPx10_ASAP7_75t_R FILLER_0_192_1286 ();
 DECAPx10_ASAP7_75t_R FILLER_0_192_1308 ();
 DECAPx10_ASAP7_75t_R FILLER_0_192_1330 ();
 DECAPx10_ASAP7_75t_R FILLER_0_192_1352 ();
 DECAPx2_ASAP7_75t_R FILLER_0_192_1374 ();
 FILLER_ASAP7_75t_R FILLER_0_192_1380 ();
 DECAPx4_ASAP7_75t_R FILLER_0_193_2 ();
 FILLER_ASAP7_75t_R FILLER_0_193_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_14 ();
 FILLER_ASAP7_75t_R FILLER_0_193_21 ();
 DECAPx2_ASAP7_75t_R FILLER_0_193_29 ();
 FILLER_ASAP7_75t_R FILLER_0_193_35 ();
 FILLER_ASAP7_75t_R FILLER_0_193_43 ();
 FILLER_ASAP7_75t_R FILLER_0_193_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_53 ();
 FILLER_ASAP7_75t_R FILLER_0_193_60 ();
 DECAPx2_ASAP7_75t_R FILLER_0_193_68 ();
 DECAPx2_ASAP7_75t_R FILLER_0_193_80 ();
 DECAPx6_ASAP7_75t_R FILLER_0_193_92 ();
 DECAPx1_ASAP7_75t_R FILLER_0_193_106 ();
 FILLER_ASAP7_75t_R FILLER_0_193_116 ();
 DECAPx2_ASAP7_75t_R FILLER_0_193_124 ();
 FILLER_ASAP7_75t_R FILLER_0_193_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_132 ();
 FILLER_ASAP7_75t_R FILLER_0_193_139 ();
 DECAPx2_ASAP7_75t_R FILLER_0_193_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_153 ();
 FILLER_ASAP7_75t_R FILLER_0_193_160 ();
 DECAPx4_ASAP7_75t_R FILLER_0_193_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_178 ();
 FILLER_ASAP7_75t_R FILLER_0_193_185 ();
 DECAPx10_ASAP7_75t_R FILLER_0_193_194 ();
 DECAPx4_ASAP7_75t_R FILLER_0_193_216 ();
 FILLER_ASAP7_75t_R FILLER_0_193_234 ();
 DECAPx2_ASAP7_75t_R FILLER_0_193_243 ();
 FILLER_ASAP7_75t_R FILLER_0_193_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_251 ();
 DECAPx4_ASAP7_75t_R FILLER_0_193_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_265 ();
 DECAPx1_ASAP7_75t_R FILLER_0_193_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_276 ();
 DECAPx2_ASAP7_75t_R FILLER_0_193_283 ();
 FILLER_ASAP7_75t_R FILLER_0_193_295 ();
 FILLER_ASAP7_75t_R FILLER_0_193_303 ();
 FILLER_ASAP7_75t_R FILLER_0_193_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_313 ();
 FILLER_ASAP7_75t_R FILLER_0_193_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_322 ();
 FILLER_ASAP7_75t_R FILLER_0_193_331 ();
 FILLER_ASAP7_75t_R FILLER_0_193_336 ();
 FILLER_ASAP7_75t_R FILLER_0_193_348 ();
 DECAPx4_ASAP7_75t_R FILLER_0_193_357 ();
 DECAPx10_ASAP7_75t_R FILLER_0_193_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_395 ();
 DECAPx1_ASAP7_75t_R FILLER_0_193_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_406 ();
 DECAPx10_ASAP7_75t_R FILLER_0_193_410 ();
 DECAPx4_ASAP7_75t_R FILLER_0_193_432 ();
 FILLER_ASAP7_75t_R FILLER_0_193_442 ();
 DECAPx6_ASAP7_75t_R FILLER_0_193_450 ();
 FILLER_ASAP7_75t_R FILLER_0_193_470 ();
 FILLER_ASAP7_75t_R FILLER_0_193_478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_193_490 ();
 DECAPx1_ASAP7_75t_R FILLER_0_193_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_516 ();
 DECAPx2_ASAP7_75t_R FILLER_0_193_523 ();
 FILLER_ASAP7_75t_R FILLER_0_193_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_531 ();
 DECAPx2_ASAP7_75t_R FILLER_0_193_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_546 ();
 DECAPx2_ASAP7_75t_R FILLER_0_193_553 ();
 FILLER_ASAP7_75t_R FILLER_0_193_567 ();
 DECAPx4_ASAP7_75t_R FILLER_0_193_579 ();
 FILLER_ASAP7_75t_R FILLER_0_193_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_597 ();
 DECAPx4_ASAP7_75t_R FILLER_0_193_604 ();
 FILLER_ASAP7_75t_R FILLER_0_193_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_616 ();
 FILLER_ASAP7_75t_R FILLER_0_193_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_627 ();
 DECAPx2_ASAP7_75t_R FILLER_0_193_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_640 ();
 FILLER_ASAP7_75t_R FILLER_0_193_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_649 ();
 FILLER_ASAP7_75t_R FILLER_0_193_656 ();
 FILLER_ASAP7_75t_R FILLER_0_193_661 ();
 DECAPx6_ASAP7_75t_R FILLER_0_193_669 ();
 DECAPx1_ASAP7_75t_R FILLER_0_193_683 ();
 FILLER_ASAP7_75t_R FILLER_0_193_708 ();
 FILLER_ASAP7_75t_R FILLER_0_193_715 ();
 FILLER_ASAP7_75t_R FILLER_0_193_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_729 ();
 FILLER_ASAP7_75t_R FILLER_0_193_740 ();
 FILLER_ASAP7_75t_R FILLER_0_193_747 ();
 DECAPx4_ASAP7_75t_R FILLER_0_193_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_765 ();
 FILLER_ASAP7_75t_R FILLER_0_193_772 ();
 DECAPx2_ASAP7_75t_R FILLER_0_193_780 ();
 DECAPx1_ASAP7_75t_R FILLER_0_193_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_804 ();
 FILLER_ASAP7_75t_R FILLER_0_193_811 ();
 DECAPx10_ASAP7_75t_R FILLER_0_193_820 ();
 DECAPx1_ASAP7_75t_R FILLER_0_193_842 ();
 DECAPx6_ASAP7_75t_R FILLER_0_193_852 ();
 DECAPx1_ASAP7_75t_R FILLER_0_193_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_870 ();
 DECAPx1_ASAP7_75t_R FILLER_0_193_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_885 ();
 FILLER_ASAP7_75t_R FILLER_0_193_893 ();
 FILLER_ASAP7_75t_R FILLER_0_193_901 ();
 DECAPx1_ASAP7_75t_R FILLER_0_193_909 ();
 DECAPx2_ASAP7_75t_R FILLER_0_193_919 ();
 DECAPx1_ASAP7_75t_R FILLER_0_193_927 ();
 DECAPx4_ASAP7_75t_R FILLER_0_193_937 ();
 FILLER_ASAP7_75t_R FILLER_0_193_947 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_949 ();
 DECAPx2_ASAP7_75t_R FILLER_0_193_956 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_962 ();
 FILLER_ASAP7_75t_R FILLER_0_193_969 ();
 DECAPx4_ASAP7_75t_R FILLER_0_193_982 ();
 FILLER_ASAP7_75t_R FILLER_0_193_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_994 ();
 DECAPx2_ASAP7_75t_R FILLER_0_193_1005 ();
 DECAPx2_ASAP7_75t_R FILLER_0_193_1021 ();
 FILLER_ASAP7_75t_R FILLER_0_193_1027 ();
 FILLER_ASAP7_75t_R FILLER_0_193_1034 ();
 DECAPx2_ASAP7_75t_R FILLER_0_193_1041 ();
 FILLER_ASAP7_75t_R FILLER_0_193_1047 ();
 FILLER_ASAP7_75t_R FILLER_0_193_1059 ();
 FILLER_ASAP7_75t_R FILLER_0_193_1069 ();
 DECAPx6_ASAP7_75t_R FILLER_0_193_1078 ();
 DECAPx1_ASAP7_75t_R FILLER_0_193_1092 ();
 DECAPx1_ASAP7_75t_R FILLER_0_193_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_1106 ();
 FILLER_ASAP7_75t_R FILLER_0_193_1117 ();
 FILLER_ASAP7_75t_R FILLER_0_193_1129 ();
 FILLER_ASAP7_75t_R FILLER_0_193_1137 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_1139 ();
 FILLER_ASAP7_75t_R FILLER_0_193_1146 ();
 DECAPx1_ASAP7_75t_R FILLER_0_193_1159 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_1163 ();
 DECAPx2_ASAP7_75t_R FILLER_0_193_1170 ();
 FILLER_ASAP7_75t_R FILLER_0_193_1176 ();
 DECAPx2_ASAP7_75t_R FILLER_0_193_1184 ();
 FILLER_ASAP7_75t_R FILLER_0_193_1190 ();
 DECAPx2_ASAP7_75t_R FILLER_0_193_1200 ();
 FILLER_ASAP7_75t_R FILLER_0_193_1212 ();
 DECAPx1_ASAP7_75t_R FILLER_0_193_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_1223 ();
 DECAPx1_ASAP7_75t_R FILLER_0_193_1231 ();
 FILLER_ASAP7_75t_R FILLER_0_193_1245 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193_1247 ();
 DECAPx1_ASAP7_75t_R FILLER_0_193_1258 ();
 FILLER_ASAP7_75t_R FILLER_0_193_1268 ();
 FILLER_ASAP7_75t_R FILLER_0_193_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_0_193_1280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_193_1302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_193_1324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_193_1346 ();
 DECAPx6_ASAP7_75t_R FILLER_0_193_1368 ();
 DECAPx2_ASAP7_75t_R FILLER_0_194_2 ();
 FILLER_ASAP7_75t_R FILLER_0_194_13 ();
 FILLER_ASAP7_75t_R FILLER_0_194_22 ();
 DECAPx2_ASAP7_75t_R FILLER_0_194_29 ();
 FILLER_ASAP7_75t_R FILLER_0_194_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_37 ();
 DECAPx1_ASAP7_75t_R FILLER_0_194_44 ();
 FILLER_ASAP7_75t_R FILLER_0_194_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_56 ();
 DECAPx1_ASAP7_75t_R FILLER_0_194_63 ();
 DECAPx2_ASAP7_75t_R FILLER_0_194_73 ();
 FILLER_ASAP7_75t_R FILLER_0_194_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_81 ();
 FILLER_ASAP7_75t_R FILLER_0_194_88 ();
 FILLER_ASAP7_75t_R FILLER_0_194_96 ();
 DECAPx4_ASAP7_75t_R FILLER_0_194_104 ();
 FILLER_ASAP7_75t_R FILLER_0_194_114 ();
 FILLER_ASAP7_75t_R FILLER_0_194_122 ();
 DECAPx2_ASAP7_75t_R FILLER_0_194_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_135 ();
 DECAPx2_ASAP7_75t_R FILLER_0_194_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_148 ();
 DECAPx6_ASAP7_75t_R FILLER_0_194_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_169 ();
 DECAPx2_ASAP7_75t_R FILLER_0_194_176 ();
 FILLER_ASAP7_75t_R FILLER_0_194_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_184 ();
 DECAPx1_ASAP7_75t_R FILLER_0_194_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_194_199 ();
 DECAPx4_ASAP7_75t_R FILLER_0_194_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_231 ();
 FILLER_ASAP7_75t_R FILLER_0_194_240 ();
 FILLER_ASAP7_75t_R FILLER_0_194_248 ();
 DECAPx1_ASAP7_75t_R FILLER_0_194_256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_194_266 ();
 DECAPx1_ASAP7_75t_R FILLER_0_194_288 ();
 FILLER_ASAP7_75t_R FILLER_0_194_299 ();
 DECAPx4_ASAP7_75t_R FILLER_0_194_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_317 ();
 DECAPx6_ASAP7_75t_R FILLER_0_194_321 ();
 FILLER_ASAP7_75t_R FILLER_0_194_345 ();
 FILLER_ASAP7_75t_R FILLER_0_194_354 ();
 FILLER_ASAP7_75t_R FILLER_0_194_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_363 ();
 FILLER_ASAP7_75t_R FILLER_0_194_370 ();
 DECAPx6_ASAP7_75t_R FILLER_0_194_375 ();
 FILLER_ASAP7_75t_R FILLER_0_194_395 ();
 FILLER_ASAP7_75t_R FILLER_0_194_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_406 ();
 FILLER_ASAP7_75t_R FILLER_0_194_413 ();
 FILLER_ASAP7_75t_R FILLER_0_194_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_425 ();
 DECAPx1_ASAP7_75t_R FILLER_0_194_432 ();
 DECAPx1_ASAP7_75t_R FILLER_0_194_443 ();
 DECAPx4_ASAP7_75t_R FILLER_0_194_450 ();
 FILLER_ASAP7_75t_R FILLER_0_194_460 ();
 FILLER_ASAP7_75t_R FILLER_0_194_464 ();
 DECAPx2_ASAP7_75t_R FILLER_0_194_472 ();
 FILLER_ASAP7_75t_R FILLER_0_194_486 ();
 DECAPx2_ASAP7_75t_R FILLER_0_194_494 ();
 DECAPx2_ASAP7_75t_R FILLER_0_194_506 ();
 FILLER_ASAP7_75t_R FILLER_0_194_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_194_535 ();
 FILLER_ASAP7_75t_R FILLER_0_194_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_543 ();
 DECAPx4_ASAP7_75t_R FILLER_0_194_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_560 ();
 FILLER_ASAP7_75t_R FILLER_0_194_571 ();
 DECAPx1_ASAP7_75t_R FILLER_0_194_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_589 ();
 FILLER_ASAP7_75t_R FILLER_0_194_597 ();
 FILLER_ASAP7_75t_R FILLER_0_194_605 ();
 FILLER_ASAP7_75t_R FILLER_0_194_610 ();
 FILLER_ASAP7_75t_R FILLER_0_194_620 ();
 DECAPx2_ASAP7_75t_R FILLER_0_194_629 ();
 FILLER_ASAP7_75t_R FILLER_0_194_641 ();
 DECAPx1_ASAP7_75t_R FILLER_0_194_649 ();
 FILLER_ASAP7_75t_R FILLER_0_194_656 ();
 FILLER_ASAP7_75t_R FILLER_0_194_664 ();
 DECAPx6_ASAP7_75t_R FILLER_0_194_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_688 ();
 DECAPx4_ASAP7_75t_R FILLER_0_194_692 ();
 FILLER_ASAP7_75t_R FILLER_0_194_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_704 ();
 FILLER_ASAP7_75t_R FILLER_0_194_715 ();
 FILLER_ASAP7_75t_R FILLER_0_194_727 ();
 DECAPx2_ASAP7_75t_R FILLER_0_194_739 ();
 DECAPx4_ASAP7_75t_R FILLER_0_194_765 ();
 FILLER_ASAP7_75t_R FILLER_0_194_781 ();
 FILLER_ASAP7_75t_R FILLER_0_194_788 ();
 FILLER_ASAP7_75t_R FILLER_0_194_802 ();
 DECAPx6_ASAP7_75t_R FILLER_0_194_809 ();
 FILLER_ASAP7_75t_R FILLER_0_194_823 ();
 DECAPx1_ASAP7_75t_R FILLER_0_194_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_835 ();
 FILLER_ASAP7_75t_R FILLER_0_194_842 ();
 DECAPx1_ASAP7_75t_R FILLER_0_194_850 ();
 FILLER_ASAP7_75t_R FILLER_0_194_860 ();
 DECAPx1_ASAP7_75t_R FILLER_0_194_868 ();
 DECAPx1_ASAP7_75t_R FILLER_0_194_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_884 ();
 DECAPx6_ASAP7_75t_R FILLER_0_194_888 ();
 DECAPx2_ASAP7_75t_R FILLER_0_194_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_908 ();
 FILLER_ASAP7_75t_R FILLER_0_194_915 ();
 DECAPx10_ASAP7_75t_R FILLER_0_194_923 ();
 DECAPx10_ASAP7_75t_R FILLER_0_194_945 ();
 FILLER_ASAP7_75t_R FILLER_0_194_973 ();
 DECAPx6_ASAP7_75t_R FILLER_0_194_981 ();
 FILLER_ASAP7_75t_R FILLER_0_194_995 ();
 DECAPx4_ASAP7_75t_R FILLER_0_194_1001 ();
 FILLER_ASAP7_75t_R FILLER_0_194_1021 ();
 DECAPx1_ASAP7_75t_R FILLER_0_194_1029 ();
 DECAPx1_ASAP7_75t_R FILLER_0_194_1043 ();
 DECAPx1_ASAP7_75t_R FILLER_0_194_1057 ();
 FILLER_ASAP7_75t_R FILLER_0_194_1069 ();
 FILLER_ASAP7_75t_R FILLER_0_194_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_1079 ();
 FILLER_ASAP7_75t_R FILLER_0_194_1090 ();
 FILLER_ASAP7_75t_R FILLER_0_194_1099 ();
 FILLER_ASAP7_75t_R FILLER_0_194_1104 ();
 DECAPx2_ASAP7_75t_R FILLER_0_194_1112 ();
 FILLER_ASAP7_75t_R FILLER_0_194_1118 ();
 FILLER_ASAP7_75t_R FILLER_0_194_1130 ();
 DECAPx1_ASAP7_75t_R FILLER_0_194_1138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_194_1149 ();
 DECAPx10_ASAP7_75t_R FILLER_0_194_1171 ();
 FILLER_ASAP7_75t_R FILLER_0_194_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_1195 ();
 FILLER_ASAP7_75t_R FILLER_0_194_1202 ();
 FILLER_ASAP7_75t_R FILLER_0_194_1210 ();
 FILLER_ASAP7_75t_R FILLER_0_194_1218 ();
 DECAPx6_ASAP7_75t_R FILLER_0_194_1223 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_1237 ();
 DECAPx2_ASAP7_75t_R FILLER_0_194_1244 ();
 FILLER_ASAP7_75t_R FILLER_0_194_1250 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_1252 ();
 DECAPx2_ASAP7_75t_R FILLER_0_194_1258 ();
 FILLER_ASAP7_75t_R FILLER_0_194_1264 ();
 FILLER_ASAP7_75t_R FILLER_0_194_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_194_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_0_194_1301 ();
 DECAPx10_ASAP7_75t_R FILLER_0_194_1323 ();
 DECAPx10_ASAP7_75t_R FILLER_0_194_1345 ();
 DECAPx6_ASAP7_75t_R FILLER_0_194_1367 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_194_1381 ();
 DECAPx6_ASAP7_75t_R FILLER_0_195_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_195_16 ();
 DECAPx2_ASAP7_75t_R FILLER_0_195_26 ();
 FILLER_ASAP7_75t_R FILLER_0_195_32 ();
 DECAPx2_ASAP7_75t_R FILLER_0_195_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_46 ();
 DECAPx6_ASAP7_75t_R FILLER_0_195_58 ();
 DECAPx2_ASAP7_75t_R FILLER_0_195_72 ();
 DECAPx2_ASAP7_75t_R FILLER_0_195_84 ();
 FILLER_ASAP7_75t_R FILLER_0_195_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_92 ();
 DECAPx2_ASAP7_75t_R FILLER_0_195_104 ();
 FILLER_ASAP7_75t_R FILLER_0_195_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_112 ();
 DECAPx6_ASAP7_75t_R FILLER_0_195_119 ();
 DECAPx1_ASAP7_75t_R FILLER_0_195_133 ();
 DECAPx2_ASAP7_75t_R FILLER_0_195_143 ();
 DECAPx2_ASAP7_75t_R FILLER_0_195_159 ();
 FILLER_ASAP7_75t_R FILLER_0_195_165 ();
 FILLER_ASAP7_75t_R FILLER_0_195_173 ();
 FILLER_ASAP7_75t_R FILLER_0_195_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_183 ();
 FILLER_ASAP7_75t_R FILLER_0_195_195 ();
 DECAPx6_ASAP7_75t_R FILLER_0_195_203 ();
 DECAPx1_ASAP7_75t_R FILLER_0_195_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_221 ();
 FILLER_ASAP7_75t_R FILLER_0_195_232 ();
 FILLER_ASAP7_75t_R FILLER_0_195_237 ();
 FILLER_ASAP7_75t_R FILLER_0_195_245 ();
 FILLER_ASAP7_75t_R FILLER_0_195_253 ();
 FILLER_ASAP7_75t_R FILLER_0_195_261 ();
 FILLER_ASAP7_75t_R FILLER_0_195_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_273 ();
 DECAPx6_ASAP7_75t_R FILLER_0_195_280 ();
 DECAPx2_ASAP7_75t_R FILLER_0_195_294 ();
 DECAPx6_ASAP7_75t_R FILLER_0_195_308 ();
 DECAPx2_ASAP7_75t_R FILLER_0_195_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_328 ();
 DECAPx1_ASAP7_75t_R FILLER_0_195_336 ();
 FILLER_ASAP7_75t_R FILLER_0_195_345 ();
 FILLER_ASAP7_75t_R FILLER_0_195_352 ();
 FILLER_ASAP7_75t_R FILLER_0_195_360 ();
 DECAPx6_ASAP7_75t_R FILLER_0_195_372 ();
 DECAPx1_ASAP7_75t_R FILLER_0_195_386 ();
 DECAPx10_ASAP7_75t_R FILLER_0_195_396 ();
 FILLER_ASAP7_75t_R FILLER_0_195_421 ();
 DECAPx2_ASAP7_75t_R FILLER_0_195_429 ();
 FILLER_ASAP7_75t_R FILLER_0_195_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_437 ();
 DECAPx6_ASAP7_75t_R FILLER_0_195_444 ();
 DECAPx1_ASAP7_75t_R FILLER_0_195_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_462 ();
 FILLER_ASAP7_75t_R FILLER_0_195_469 ();
 FILLER_ASAP7_75t_R FILLER_0_195_477 ();
 FILLER_ASAP7_75t_R FILLER_0_195_486 ();
 FILLER_ASAP7_75t_R FILLER_0_195_494 ();
 FILLER_ASAP7_75t_R FILLER_0_195_502 ();
 DECAPx4_ASAP7_75t_R FILLER_0_195_511 ();
 DECAPx6_ASAP7_75t_R FILLER_0_195_527 ();
 FILLER_ASAP7_75t_R FILLER_0_195_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_543 ();
 DECAPx2_ASAP7_75t_R FILLER_0_195_550 ();
 FILLER_ASAP7_75t_R FILLER_0_195_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_558 ();
 FILLER_ASAP7_75t_R FILLER_0_195_564 ();
 DECAPx2_ASAP7_75t_R FILLER_0_195_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_577 ();
 DECAPx1_ASAP7_75t_R FILLER_0_195_584 ();
 DECAPx4_ASAP7_75t_R FILLER_0_195_591 ();
 FILLER_ASAP7_75t_R FILLER_0_195_607 ();
 FILLER_ASAP7_75t_R FILLER_0_195_615 ();
 FILLER_ASAP7_75t_R FILLER_0_195_624 ();
 DECAPx6_ASAP7_75t_R FILLER_0_195_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_645 ();
 FILLER_ASAP7_75t_R FILLER_0_195_654 ();
 FILLER_ASAP7_75t_R FILLER_0_195_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_195_667 ();
 DECAPx1_ASAP7_75t_R FILLER_0_195_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_693 ();
 FILLER_ASAP7_75t_R FILLER_0_195_697 ();
 DECAPx6_ASAP7_75t_R FILLER_0_195_705 ();
 FILLER_ASAP7_75t_R FILLER_0_195_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_721 ();
 FILLER_ASAP7_75t_R FILLER_0_195_732 ();
 DECAPx2_ASAP7_75t_R FILLER_0_195_740 ();
 DECAPx1_ASAP7_75t_R FILLER_0_195_756 ();
 FILLER_ASAP7_75t_R FILLER_0_195_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_784 ();
 DECAPx1_ASAP7_75t_R FILLER_0_195_792 ();
 DECAPx1_ASAP7_75t_R FILLER_0_195_803 ();
 DECAPx1_ASAP7_75t_R FILLER_0_195_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_817 ();
 FILLER_ASAP7_75t_R FILLER_0_195_824 ();
 DECAPx4_ASAP7_75t_R FILLER_0_195_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_842 ();
 DECAPx2_ASAP7_75t_R FILLER_0_195_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_855 ();
 DECAPx2_ASAP7_75t_R FILLER_0_195_864 ();
 FILLER_ASAP7_75t_R FILLER_0_195_870 ();
 FILLER_ASAP7_75t_R FILLER_0_195_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_880 ();
 DECAPx1_ASAP7_75t_R FILLER_0_195_887 ();
 DECAPx6_ASAP7_75t_R FILLER_0_195_898 ();
 DECAPx1_ASAP7_75t_R FILLER_0_195_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_916 ();
 FILLER_ASAP7_75t_R FILLER_0_195_923 ();
 DECAPx4_ASAP7_75t_R FILLER_0_195_927 ();
 FILLER_ASAP7_75t_R FILLER_0_195_937 ();
 DECAPx2_ASAP7_75t_R FILLER_0_195_945 ();
 DECAPx6_ASAP7_75t_R FILLER_0_195_957 ();
 DECAPx1_ASAP7_75t_R FILLER_0_195_971 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_975 ();
 FILLER_ASAP7_75t_R FILLER_0_195_982 ();
 DECAPx6_ASAP7_75t_R FILLER_0_195_987 ();
 FILLER_ASAP7_75t_R FILLER_0_195_1011 ();
 FILLER_ASAP7_75t_R FILLER_0_195_1023 ();
 FILLER_ASAP7_75t_R FILLER_0_195_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_1037 ();
 DECAPx1_ASAP7_75t_R FILLER_0_195_1048 ();
 FILLER_ASAP7_75t_R FILLER_0_195_1062 ();
 FILLER_ASAP7_75t_R FILLER_0_195_1070 ();
 FILLER_ASAP7_75t_R FILLER_0_195_1078 ();
 FILLER_ASAP7_75t_R FILLER_0_195_1086 ();
 FILLER_ASAP7_75t_R FILLER_0_195_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_1096 ();
 DECAPx1_ASAP7_75t_R FILLER_0_195_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_1107 ();
 FILLER_ASAP7_75t_R FILLER_0_195_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_1118 ();
 FILLER_ASAP7_75t_R FILLER_0_195_1129 ();
 FILLER_ASAP7_75t_R FILLER_0_195_1141 ();
 FILLER_ASAP7_75t_R FILLER_0_195_1148 ();
 DECAPx4_ASAP7_75t_R FILLER_0_195_1153 ();
 FILLER_ASAP7_75t_R FILLER_0_195_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_1165 ();
 FILLER_ASAP7_75t_R FILLER_0_195_1176 ();
 DECAPx4_ASAP7_75t_R FILLER_0_195_1184 ();
 FILLER_ASAP7_75t_R FILLER_0_195_1194 ();
 FILLER_ASAP7_75t_R FILLER_0_195_1202 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_1204 ();
 DECAPx6_ASAP7_75t_R FILLER_0_195_1211 ();
 FILLER_ASAP7_75t_R FILLER_0_195_1225 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_1227 ();
 FILLER_ASAP7_75t_R FILLER_0_195_1238 ();
 DECAPx4_ASAP7_75t_R FILLER_0_195_1246 ();
 FILLER_ASAP7_75t_R FILLER_0_195_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_1263 ();
 FILLER_ASAP7_75t_R FILLER_0_195_1270 ();
 FILLER_ASAP7_75t_R FILLER_0_195_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_0_195_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_0_195_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_0_195_1333 ();
 DECAPx10_ASAP7_75t_R FILLER_0_195_1355 ();
 DECAPx1_ASAP7_75t_R FILLER_0_195_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_195_1381 ();
 DECAPx6_ASAP7_75t_R FILLER_0_196_2 ();
 FILLER_ASAP7_75t_R FILLER_0_196_22 ();
 DECAPx1_ASAP7_75t_R FILLER_0_196_30 ();
 DECAPx2_ASAP7_75t_R FILLER_0_196_40 ();
 DECAPx2_ASAP7_75t_R FILLER_0_196_49 ();
 DECAPx2_ASAP7_75t_R FILLER_0_196_61 ();
 DECAPx10_ASAP7_75t_R FILLER_0_196_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_109 ();
 FILLER_ASAP7_75t_R FILLER_0_196_116 ();
 DECAPx4_ASAP7_75t_R FILLER_0_196_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_134 ();
 DECAPx6_ASAP7_75t_R FILLER_0_196_141 ();
 FILLER_ASAP7_75t_R FILLER_0_196_155 ();
 DECAPx2_ASAP7_75t_R FILLER_0_196_163 ();
 FILLER_ASAP7_75t_R FILLER_0_196_169 ();
 DECAPx1_ASAP7_75t_R FILLER_0_196_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_181 ();
 FILLER_ASAP7_75t_R FILLER_0_196_188 ();
 FILLER_ASAP7_75t_R FILLER_0_196_196 ();
 DECAPx10_ASAP7_75t_R FILLER_0_196_209 ();
 DECAPx10_ASAP7_75t_R FILLER_0_196_238 ();
 FILLER_ASAP7_75t_R FILLER_0_196_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_262 ();
 FILLER_ASAP7_75t_R FILLER_0_196_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_271 ();
 FILLER_ASAP7_75t_R FILLER_0_196_278 ();
 FILLER_ASAP7_75t_R FILLER_0_196_287 ();
 FILLER_ASAP7_75t_R FILLER_0_196_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_297 ();
 DECAPx1_ASAP7_75t_R FILLER_0_196_306 ();
 DECAPx1_ASAP7_75t_R FILLER_0_196_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_317 ();
 DECAPx2_ASAP7_75t_R FILLER_0_196_325 ();
 DECAPx4_ASAP7_75t_R FILLER_0_196_337 ();
 DECAPx2_ASAP7_75t_R FILLER_0_196_350 ();
 FILLER_ASAP7_75t_R FILLER_0_196_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_358 ();
 DECAPx2_ASAP7_75t_R FILLER_0_196_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_373 ();
 FILLER_ASAP7_75t_R FILLER_0_196_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_382 ();
 FILLER_ASAP7_75t_R FILLER_0_196_386 ();
 FILLER_ASAP7_75t_R FILLER_0_196_395 ();
 DECAPx1_ASAP7_75t_R FILLER_0_196_403 ();
 DECAPx2_ASAP7_75t_R FILLER_0_196_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_416 ();
 DECAPx10_ASAP7_75t_R FILLER_0_196_423 ();
 DECAPx6_ASAP7_75t_R FILLER_0_196_445 ();
 FILLER_ASAP7_75t_R FILLER_0_196_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_461 ();
 DECAPx2_ASAP7_75t_R FILLER_0_196_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_470 ();
 DECAPx4_ASAP7_75t_R FILLER_0_196_477 ();
 DECAPx2_ASAP7_75t_R FILLER_0_196_493 ();
 FILLER_ASAP7_75t_R FILLER_0_196_499 ();
 DECAPx2_ASAP7_75t_R FILLER_0_196_507 ();
 FILLER_ASAP7_75t_R FILLER_0_196_518 ();
 FILLER_ASAP7_75t_R FILLER_0_196_540 ();
 DECAPx10_ASAP7_75t_R FILLER_0_196_548 ();
 DECAPx4_ASAP7_75t_R FILLER_0_196_576 ();
 FILLER_ASAP7_75t_R FILLER_0_196_586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_196_595 ();
 FILLER_ASAP7_75t_R FILLER_0_196_617 ();
 DECAPx2_ASAP7_75t_R FILLER_0_196_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_631 ();
 DECAPx2_ASAP7_75t_R FILLER_0_196_639 ();
 FILLER_ASAP7_75t_R FILLER_0_196_645 ();
 DECAPx2_ASAP7_75t_R FILLER_0_196_654 ();
 FILLER_ASAP7_75t_R FILLER_0_196_660 ();
 DECAPx6_ASAP7_75t_R FILLER_0_196_670 ();
 FILLER_ASAP7_75t_R FILLER_0_196_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_686 ();
 FILLER_ASAP7_75t_R FILLER_0_196_707 ();
 FILLER_ASAP7_75t_R FILLER_0_196_715 ();
 DECAPx2_ASAP7_75t_R FILLER_0_196_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_733 ();
 DECAPx1_ASAP7_75t_R FILLER_0_196_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_744 ();
 FILLER_ASAP7_75t_R FILLER_0_196_751 ();
 DECAPx2_ASAP7_75t_R FILLER_0_196_760 ();
 FILLER_ASAP7_75t_R FILLER_0_196_772 ();
 FILLER_ASAP7_75t_R FILLER_0_196_785 ();
 FILLER_ASAP7_75t_R FILLER_0_196_797 ();
 FILLER_ASAP7_75t_R FILLER_0_196_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_804 ();
 DECAPx2_ASAP7_75t_R FILLER_0_196_815 ();
 DECAPx4_ASAP7_75t_R FILLER_0_196_832 ();
 FILLER_ASAP7_75t_R FILLER_0_196_848 ();
 FILLER_ASAP7_75t_R FILLER_0_196_855 ();
 FILLER_ASAP7_75t_R FILLER_0_196_877 ();
 FILLER_ASAP7_75t_R FILLER_0_196_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_885 ();
 FILLER_ASAP7_75t_R FILLER_0_196_895 ();
 DECAPx4_ASAP7_75t_R FILLER_0_196_903 ();
 FILLER_ASAP7_75t_R FILLER_0_196_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_915 ();
 FILLER_ASAP7_75t_R FILLER_0_196_922 ();
 DECAPx2_ASAP7_75t_R FILLER_0_196_934 ();
 FILLER_ASAP7_75t_R FILLER_0_196_940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_196_953 ();
 FILLER_ASAP7_75t_R FILLER_0_196_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_977 ();
 DECAPx6_ASAP7_75t_R FILLER_0_196_984 ();
 DECAPx1_ASAP7_75t_R FILLER_0_196_998 ();
 FILLER_ASAP7_75t_R FILLER_0_196_1012 ();
 FILLER_ASAP7_75t_R FILLER_0_196_1024 ();
 FILLER_ASAP7_75t_R FILLER_0_196_1036 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_1038 ();
 DECAPx1_ASAP7_75t_R FILLER_0_196_1049 ();
 FILLER_ASAP7_75t_R FILLER_0_196_1063 ();
 DECAPx2_ASAP7_75t_R FILLER_0_196_1072 ();
 FILLER_ASAP7_75t_R FILLER_0_196_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_1080 ();
 DECAPx6_ASAP7_75t_R FILLER_0_196_1087 ();
 FILLER_ASAP7_75t_R FILLER_0_196_1109 ();
 FILLER_ASAP7_75t_R FILLER_0_196_1116 ();
 FILLER_ASAP7_75t_R FILLER_0_196_1128 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_1130 ();
 FILLER_ASAP7_75t_R FILLER_0_196_1137 ();
 FILLER_ASAP7_75t_R FILLER_0_196_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_1149 ();
 DECAPx4_ASAP7_75t_R FILLER_0_196_1161 ();
 FILLER_ASAP7_75t_R FILLER_0_196_1171 ();
 DECAPx2_ASAP7_75t_R FILLER_0_196_1180 ();
 FILLER_ASAP7_75t_R FILLER_0_196_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_196_1195 ();
 DECAPx2_ASAP7_75t_R FILLER_0_196_1203 ();
 FILLER_ASAP7_75t_R FILLER_0_196_1216 ();
 FILLER_ASAP7_75t_R FILLER_0_196_1224 ();
 DECAPx2_ASAP7_75t_R FILLER_0_196_1232 ();
 FILLER_ASAP7_75t_R FILLER_0_196_1238 ();
 FILLER_ASAP7_75t_R FILLER_0_196_1246 ();
 FILLER_ASAP7_75t_R FILLER_0_196_1254 ();
 DECAPx4_ASAP7_75t_R FILLER_0_196_1262 ();
 FILLER_ASAP7_75t_R FILLER_0_196_1272 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_1274 ();
 DECAPx10_ASAP7_75t_R FILLER_0_196_1281 ();
 DECAPx10_ASAP7_75t_R FILLER_0_196_1303 ();
 DECAPx10_ASAP7_75t_R FILLER_0_196_1325 ();
 DECAPx10_ASAP7_75t_R FILLER_0_196_1347 ();
 DECAPx4_ASAP7_75t_R FILLER_0_196_1369 ();
 FILLER_ASAP7_75t_R FILLER_0_196_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_196_1381 ();
 DECAPx2_ASAP7_75t_R FILLER_0_197_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_197_14 ();
 FILLER_ASAP7_75t_R FILLER_0_197_29 ();
 FILLER_ASAP7_75t_R FILLER_0_197_51 ();
 DECAPx4_ASAP7_75t_R FILLER_0_197_59 ();
 FILLER_ASAP7_75t_R FILLER_0_197_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_71 ();
 DECAPx2_ASAP7_75t_R FILLER_0_197_78 ();
 FILLER_ASAP7_75t_R FILLER_0_197_84 ();
 FILLER_ASAP7_75t_R FILLER_0_197_92 ();
 DECAPx4_ASAP7_75t_R FILLER_0_197_100 ();
 DECAPx6_ASAP7_75t_R FILLER_0_197_116 ();
 DECAPx1_ASAP7_75t_R FILLER_0_197_130 ();
 DECAPx2_ASAP7_75t_R FILLER_0_197_145 ();
 FILLER_ASAP7_75t_R FILLER_0_197_157 ();
 DECAPx2_ASAP7_75t_R FILLER_0_197_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_171 ();
 FILLER_ASAP7_75t_R FILLER_0_197_175 ();
 FILLER_ASAP7_75t_R FILLER_0_197_182 ();
 DECAPx4_ASAP7_75t_R FILLER_0_197_192 ();
 FILLER_ASAP7_75t_R FILLER_0_197_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_204 ();
 DECAPx6_ASAP7_75t_R FILLER_0_197_211 ();
 DECAPx2_ASAP7_75t_R FILLER_0_197_225 ();
 DECAPx1_ASAP7_75t_R FILLER_0_197_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_242 ();
 DECAPx2_ASAP7_75t_R FILLER_0_197_249 ();
 FILLER_ASAP7_75t_R FILLER_0_197_255 ();
 FILLER_ASAP7_75t_R FILLER_0_197_264 ();
 DECAPx6_ASAP7_75t_R FILLER_0_197_272 ();
 FILLER_ASAP7_75t_R FILLER_0_197_286 ();
 DECAPx4_ASAP7_75t_R FILLER_0_197_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_318 ();
 DECAPx2_ASAP7_75t_R FILLER_0_197_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_331 ();
 FILLER_ASAP7_75t_R FILLER_0_197_338 ();
 DECAPx1_ASAP7_75t_R FILLER_0_197_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_347 ();
 DECAPx4_ASAP7_75t_R FILLER_0_197_355 ();
 FILLER_ASAP7_75t_R FILLER_0_197_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_367 ();
 DECAPx2_ASAP7_75t_R FILLER_0_197_374 ();
 FILLER_ASAP7_75t_R FILLER_0_197_388 ();
 FILLER_ASAP7_75t_R FILLER_0_197_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_398 ();
 DECAPx1_ASAP7_75t_R FILLER_0_197_407 ();
 FILLER_ASAP7_75t_R FILLER_0_197_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_420 ();
 DECAPx1_ASAP7_75t_R FILLER_0_197_427 ();
 DECAPx2_ASAP7_75t_R FILLER_0_197_437 ();
 FILLER_ASAP7_75t_R FILLER_0_197_443 ();
 FILLER_ASAP7_75t_R FILLER_0_197_451 ();
 DECAPx4_ASAP7_75t_R FILLER_0_197_458 ();
 FILLER_ASAP7_75t_R FILLER_0_197_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_470 ();
 DECAPx6_ASAP7_75t_R FILLER_0_197_477 ();
 DECAPx1_ASAP7_75t_R FILLER_0_197_491 ();
 FILLER_ASAP7_75t_R FILLER_0_197_501 ();
 DECAPx2_ASAP7_75t_R FILLER_0_197_511 ();
 FILLER_ASAP7_75t_R FILLER_0_197_517 ();
 DECAPx2_ASAP7_75t_R FILLER_0_197_525 ();
 FILLER_ASAP7_75t_R FILLER_0_197_537 ();
 FILLER_ASAP7_75t_R FILLER_0_197_545 ();
 DECAPx1_ASAP7_75t_R FILLER_0_197_553 ();
 FILLER_ASAP7_75t_R FILLER_0_197_567 ();
 DECAPx4_ASAP7_75t_R FILLER_0_197_575 ();
 FILLER_ASAP7_75t_R FILLER_0_197_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_587 ();
 FILLER_ASAP7_75t_R FILLER_0_197_594 ();
 DECAPx4_ASAP7_75t_R FILLER_0_197_602 ();
 FILLER_ASAP7_75t_R FILLER_0_197_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_614 ();
 DECAPx2_ASAP7_75t_R FILLER_0_197_621 ();
 FILLER_ASAP7_75t_R FILLER_0_197_627 ();
 FILLER_ASAP7_75t_R FILLER_0_197_635 ();
 FILLER_ASAP7_75t_R FILLER_0_197_643 ();
 FILLER_ASAP7_75t_R FILLER_0_197_651 ();
 DECAPx10_ASAP7_75t_R FILLER_0_197_661 ();
 DECAPx2_ASAP7_75t_R FILLER_0_197_683 ();
 FILLER_ASAP7_75t_R FILLER_0_197_689 ();
 DECAPx2_ASAP7_75t_R FILLER_0_197_701 ();
 DECAPx4_ASAP7_75t_R FILLER_0_197_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_728 ();
 FILLER_ASAP7_75t_R FILLER_0_197_740 ();
 DECAPx2_ASAP7_75t_R FILLER_0_197_748 ();
 DECAPx2_ASAP7_75t_R FILLER_0_197_764 ();
 FILLER_ASAP7_75t_R FILLER_0_197_770 ();
 DECAPx4_ASAP7_75t_R FILLER_0_197_782 ();
 FILLER_ASAP7_75t_R FILLER_0_197_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_794 ();
 FILLER_ASAP7_75t_R FILLER_0_197_801 ();
 DECAPx2_ASAP7_75t_R FILLER_0_197_813 ();
 FILLER_ASAP7_75t_R FILLER_0_197_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_821 ();
 FILLER_ASAP7_75t_R FILLER_0_197_827 ();
 DECAPx4_ASAP7_75t_R FILLER_0_197_834 ();
 DECAPx1_ASAP7_75t_R FILLER_0_197_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_854 ();
 DECAPx2_ASAP7_75t_R FILLER_0_197_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_867 ();
 FILLER_ASAP7_75t_R FILLER_0_197_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_880 ();
 DECAPx1_ASAP7_75t_R FILLER_0_197_889 ();
 FILLER_ASAP7_75t_R FILLER_0_197_900 ();
 DECAPx4_ASAP7_75t_R FILLER_0_197_913 ();
 FILLER_ASAP7_75t_R FILLER_0_197_923 ();
 DECAPx6_ASAP7_75t_R FILLER_0_197_927 ();
 FILLER_ASAP7_75t_R FILLER_0_197_941 ();
 DECAPx4_ASAP7_75t_R FILLER_0_197_949 ();
 FILLER_ASAP7_75t_R FILLER_0_197_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_961 ();
 FILLER_ASAP7_75t_R FILLER_0_197_965 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_967 ();
 DECAPx2_ASAP7_75t_R FILLER_0_197_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_980 ();
 DECAPx2_ASAP7_75t_R FILLER_0_197_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_994 ();
 FILLER_ASAP7_75t_R FILLER_0_197_999 ();
 DECAPx1_ASAP7_75t_R FILLER_0_197_1011 ();
 FILLER_ASAP7_75t_R FILLER_0_197_1020 ();
 DECAPx1_ASAP7_75t_R FILLER_0_197_1032 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_1036 ();
 FILLER_ASAP7_75t_R FILLER_0_197_1042 ();
 FILLER_ASAP7_75t_R FILLER_0_197_1054 ();
 FILLER_ASAP7_75t_R FILLER_0_197_1062 ();
 DECAPx1_ASAP7_75t_R FILLER_0_197_1069 ();
 DECAPx2_ASAP7_75t_R FILLER_0_197_1085 ();
 FILLER_ASAP7_75t_R FILLER_0_197_1091 ();
 FILLER_ASAP7_75t_R FILLER_0_197_1098 ();
 FILLER_ASAP7_75t_R FILLER_0_197_1108 ();
 DECAPx2_ASAP7_75t_R FILLER_0_197_1115 ();
 FILLER_ASAP7_75t_R FILLER_0_197_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_1123 ();
 DECAPx6_ASAP7_75t_R FILLER_0_197_1129 ();
 DECAPx1_ASAP7_75t_R FILLER_0_197_1153 ();
 FILLER_ASAP7_75t_R FILLER_0_197_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_1165 ();
 DECAPx10_ASAP7_75t_R FILLER_0_197_1172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_197_1194 ();
 DECAPx2_ASAP7_75t_R FILLER_0_197_1216 ();
 FILLER_ASAP7_75t_R FILLER_0_197_1228 ();
 DECAPx6_ASAP7_75t_R FILLER_0_197_1235 ();
 DECAPx1_ASAP7_75t_R FILLER_0_197_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_0_197_1259 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_197_1281 ();
 DECAPx10_ASAP7_75t_R FILLER_0_197_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_197_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_197_1332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_197_1354 ();
 DECAPx2_ASAP7_75t_R FILLER_0_197_1376 ();
 DECAPx2_ASAP7_75t_R FILLER_0_198_2 ();
 FILLER_ASAP7_75t_R FILLER_0_198_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_10 ();
 DECAPx2_ASAP7_75t_R FILLER_0_198_17 ();
 DECAPx4_ASAP7_75t_R FILLER_0_198_34 ();
 FILLER_ASAP7_75t_R FILLER_0_198_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_46 ();
 DECAPx2_ASAP7_75t_R FILLER_0_198_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_73 ();
 DECAPx2_ASAP7_75t_R FILLER_0_198_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_86 ();
 FILLER_ASAP7_75t_R FILLER_0_198_93 ();
 DECAPx4_ASAP7_75t_R FILLER_0_198_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_111 ();
 DECAPx1_ASAP7_75t_R FILLER_0_198_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_122 ();
 FILLER_ASAP7_75t_R FILLER_0_198_130 ();
 DECAPx6_ASAP7_75t_R FILLER_0_198_138 ();
 DECAPx1_ASAP7_75t_R FILLER_0_198_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_156 ();
 FILLER_ASAP7_75t_R FILLER_0_198_163 ();
 FILLER_ASAP7_75t_R FILLER_0_198_171 ();
 DECAPx1_ASAP7_75t_R FILLER_0_198_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_183 ();
 FILLER_ASAP7_75t_R FILLER_0_198_200 ();
 DECAPx6_ASAP7_75t_R FILLER_0_198_213 ();
 DECAPx2_ASAP7_75t_R FILLER_0_198_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_233 ();
 DECAPx1_ASAP7_75t_R FILLER_0_198_240 ();
 DECAPx2_ASAP7_75t_R FILLER_0_198_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_257 ();
 FILLER_ASAP7_75t_R FILLER_0_198_264 ();
 DECAPx1_ASAP7_75t_R FILLER_0_198_272 ();
 FILLER_ASAP7_75t_R FILLER_0_198_282 ();
 DECAPx2_ASAP7_75t_R FILLER_0_198_290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_198_302 ();
 DECAPx2_ASAP7_75t_R FILLER_0_198_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_330 ();
 FILLER_ASAP7_75t_R FILLER_0_198_337 ();
 DECAPx1_ASAP7_75t_R FILLER_0_198_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_349 ();
 DECAPx6_ASAP7_75t_R FILLER_0_198_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_370 ();
 FILLER_ASAP7_75t_R FILLER_0_198_377 ();
 DECAPx1_ASAP7_75t_R FILLER_0_198_385 ();
 FILLER_ASAP7_75t_R FILLER_0_198_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_394 ();
 DECAPx1_ASAP7_75t_R FILLER_0_198_401 ();
 FILLER_ASAP7_75t_R FILLER_0_198_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_410 ();
 DECAPx1_ASAP7_75t_R FILLER_0_198_417 ();
 DECAPx1_ASAP7_75t_R FILLER_0_198_429 ();
 DECAPx1_ASAP7_75t_R FILLER_0_198_444 ();
 FILLER_ASAP7_75t_R FILLER_0_198_454 ();
 FILLER_ASAP7_75t_R FILLER_0_198_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_461 ();
 DECAPx1_ASAP7_75t_R FILLER_0_198_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_468 ();
 DECAPx2_ASAP7_75t_R FILLER_0_198_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_482 ();
 FILLER_ASAP7_75t_R FILLER_0_198_489 ();
 DECAPx1_ASAP7_75t_R FILLER_0_198_497 ();
 DECAPx2_ASAP7_75t_R FILLER_0_198_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_513 ();
 DECAPx2_ASAP7_75t_R FILLER_0_198_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_526 ();
 DECAPx4_ASAP7_75t_R FILLER_0_198_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_543 ();
 FILLER_ASAP7_75t_R FILLER_0_198_551 ();
 FILLER_ASAP7_75t_R FILLER_0_198_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_561 ();
 DECAPx4_ASAP7_75t_R FILLER_0_198_567 ();
 FILLER_ASAP7_75t_R FILLER_0_198_580 ();
 FILLER_ASAP7_75t_R FILLER_0_198_588 ();
 DECAPx6_ASAP7_75t_R FILLER_0_198_596 ();
 DECAPx2_ASAP7_75t_R FILLER_0_198_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_616 ();
 FILLER_ASAP7_75t_R FILLER_0_198_623 ();
 FILLER_ASAP7_75t_R FILLER_0_198_631 ();
 DECAPx4_ASAP7_75t_R FILLER_0_198_639 ();
 FILLER_ASAP7_75t_R FILLER_0_198_655 ();
 DECAPx10_ASAP7_75t_R FILLER_0_198_660 ();
 DECAPx10_ASAP7_75t_R FILLER_0_198_682 ();
 FILLER_ASAP7_75t_R FILLER_0_198_704 ();
 FILLER_ASAP7_75t_R FILLER_0_198_712 ();
 DECAPx10_ASAP7_75t_R FILLER_0_198_717 ();
 DECAPx4_ASAP7_75t_R FILLER_0_198_739 ();
 FILLER_ASAP7_75t_R FILLER_0_198_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_751 ();
 FILLER_ASAP7_75t_R FILLER_0_198_758 ();
 FILLER_ASAP7_75t_R FILLER_0_198_766 ();
 FILLER_ASAP7_75t_R FILLER_0_198_774 ();
 DECAPx4_ASAP7_75t_R FILLER_0_198_781 ();
 DECAPx2_ASAP7_75t_R FILLER_0_198_801 ();
 FILLER_ASAP7_75t_R FILLER_0_198_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_809 ();
 DECAPx2_ASAP7_75t_R FILLER_0_198_816 ();
 DECAPx2_ASAP7_75t_R FILLER_0_198_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_834 ();
 FILLER_ASAP7_75t_R FILLER_0_198_841 ();
 DECAPx6_ASAP7_75t_R FILLER_0_198_853 ();
 DECAPx1_ASAP7_75t_R FILLER_0_198_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_871 ();
 FILLER_ASAP7_75t_R FILLER_0_198_877 ();
 DECAPx4_ASAP7_75t_R FILLER_0_198_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_895 ();
 FILLER_ASAP7_75t_R FILLER_0_198_906 ();
 FILLER_ASAP7_75t_R FILLER_0_198_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_198_923 ();
 DECAPx2_ASAP7_75t_R FILLER_0_198_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_957 ();
 FILLER_ASAP7_75t_R FILLER_0_198_964 ();
 FILLER_ASAP7_75t_R FILLER_0_198_972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_198_977 ();
 DECAPx10_ASAP7_75t_R FILLER_0_198_999 ();
 DECAPx1_ASAP7_75t_R FILLER_0_198_1021 ();
 FILLER_ASAP7_75t_R FILLER_0_198_1031 ();
 FILLER_ASAP7_75t_R FILLER_0_198_1053 ();
 DECAPx2_ASAP7_75t_R FILLER_0_198_1065 ();
 FILLER_ASAP7_75t_R FILLER_0_198_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_1073 ();
 FILLER_ASAP7_75t_R FILLER_0_198_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_0_198_1091 ();
 FILLER_ASAP7_75t_R FILLER_0_198_1109 ();
 FILLER_ASAP7_75t_R FILLER_0_198_1116 ();
 DECAPx4_ASAP7_75t_R FILLER_0_198_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_1134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_198_1145 ();
 DECAPx4_ASAP7_75t_R FILLER_0_198_1167 ();
 DECAPx4_ASAP7_75t_R FILLER_0_198_1183 ();
 FILLER_ASAP7_75t_R FILLER_0_198_1193 ();
 DECAPx2_ASAP7_75t_R FILLER_0_198_1201 ();
 FILLER_ASAP7_75t_R FILLER_0_198_1207 ();
 FILLER_ASAP7_75t_R FILLER_0_198_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_1221 ();
 FILLER_ASAP7_75t_R FILLER_0_198_1228 ();
 FILLER_ASAP7_75t_R FILLER_0_198_1236 ();
 DECAPx6_ASAP7_75t_R FILLER_0_198_1244 ();
 DECAPx2_ASAP7_75t_R FILLER_0_198_1258 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_1264 ();
 DECAPx1_ASAP7_75t_R FILLER_0_198_1271 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_198_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_0_198_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_198_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_198_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_198_1348 ();
 DECAPx4_ASAP7_75t_R FILLER_0_198_1370 ();
 FILLER_ASAP7_75t_R FILLER_0_198_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_199_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_199_24 ();
 FILLER_ASAP7_75t_R FILLER_0_199_38 ();
 FILLER_ASAP7_75t_R FILLER_0_199_50 ();
 DECAPx10_ASAP7_75t_R FILLER_0_199_62 ();
 FILLER_ASAP7_75t_R FILLER_0_199_84 ();
 FILLER_ASAP7_75t_R FILLER_0_199_91 ();
 DECAPx4_ASAP7_75t_R FILLER_0_199_99 ();
 FILLER_ASAP7_75t_R FILLER_0_199_109 ();
 FILLER_ASAP7_75t_R FILLER_0_199_115 ();
 FILLER_ASAP7_75t_R FILLER_0_199_125 ();
 FILLER_ASAP7_75t_R FILLER_0_199_133 ();
 FILLER_ASAP7_75t_R FILLER_0_199_141 ();
 DECAPx2_ASAP7_75t_R FILLER_0_199_149 ();
 FILLER_ASAP7_75t_R FILLER_0_199_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_199_157 ();
 FILLER_ASAP7_75t_R FILLER_0_199_169 ();
 DECAPx10_ASAP7_75t_R FILLER_0_199_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_199_197 ();
 DECAPx10_ASAP7_75t_R FILLER_0_199_204 ();
 DECAPx1_ASAP7_75t_R FILLER_0_199_236 ();
 FILLER_ASAP7_75t_R FILLER_0_199_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_199_248 ();
 FILLER_ASAP7_75t_R FILLER_0_199_255 ();
 DECAPx2_ASAP7_75t_R FILLER_0_199_264 ();
 DECAPx2_ASAP7_75t_R FILLER_0_199_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_199_283 ();
 DECAPx1_ASAP7_75t_R FILLER_0_199_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_199_296 ();
 FILLER_ASAP7_75t_R FILLER_0_199_303 ();
 FILLER_ASAP7_75t_R FILLER_0_199_311 ();
 DECAPx6_ASAP7_75t_R FILLER_0_199_319 ();
 DECAPx2_ASAP7_75t_R FILLER_0_199_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_199_347 ();
 DECAPx1_ASAP7_75t_R FILLER_0_199_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_199_364 ();
 DECAPx6_ASAP7_75t_R FILLER_0_199_386 ();
 FILLER_ASAP7_75t_R FILLER_0_199_406 ();
 DECAPx10_ASAP7_75t_R FILLER_0_199_414 ();
 DECAPx4_ASAP7_75t_R FILLER_0_199_436 ();
 FILLER_ASAP7_75t_R FILLER_0_199_446 ();
 DECAPx2_ASAP7_75t_R FILLER_0_199_468 ();
 FILLER_ASAP7_75t_R FILLER_0_199_482 ();
 DECAPx1_ASAP7_75t_R FILLER_0_199_490 ();
 DECAPx6_ASAP7_75t_R FILLER_0_199_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_199_511 ();
 FILLER_ASAP7_75t_R FILLER_0_199_518 ();
 DECAPx4_ASAP7_75t_R FILLER_0_199_526 ();
 DECAPx6_ASAP7_75t_R FILLER_0_199_546 ();
 DECAPx2_ASAP7_75t_R FILLER_0_199_560 ();
 FILLER_ASAP7_75t_R FILLER_0_199_594 ();
 DECAPx6_ASAP7_75t_R FILLER_0_199_603 ();
 DECAPx1_ASAP7_75t_R FILLER_0_199_617 ();
 DECAPx2_ASAP7_75t_R FILLER_0_199_629 ();
 FILLER_ASAP7_75t_R FILLER_0_199_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_199_637 ();
 FILLER_ASAP7_75t_R FILLER_0_199_645 ();
 FILLER_ASAP7_75t_R FILLER_0_199_650 ();
 DECAPx10_ASAP7_75t_R FILLER_0_199_658 ();
 DECAPx6_ASAP7_75t_R FILLER_0_199_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_199_694 ();
 DECAPx4_ASAP7_75t_R FILLER_0_199_698 ();
 FILLER_ASAP7_75t_R FILLER_0_199_708 ();
 DECAPx6_ASAP7_75t_R FILLER_0_199_716 ();
 DECAPx2_ASAP7_75t_R FILLER_0_199_730 ();
 FILLER_ASAP7_75t_R FILLER_0_199_742 ();
 DECAPx6_ASAP7_75t_R FILLER_0_199_750 ();
 DECAPx2_ASAP7_75t_R FILLER_0_199_770 ();
 DECAPx2_ASAP7_75t_R FILLER_0_199_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_199_794 ();
 DECAPx6_ASAP7_75t_R FILLER_0_199_798 ();
 DECAPx2_ASAP7_75t_R FILLER_0_199_812 ();
 DECAPx4_ASAP7_75t_R FILLER_0_199_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_199_839 ();
 FILLER_ASAP7_75t_R FILLER_0_199_846 ();
 FILLER_ASAP7_75t_R FILLER_0_199_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_199_856 ();
 DECAPx10_ASAP7_75t_R FILLER_0_199_863 ();
 FILLER_ASAP7_75t_R FILLER_0_199_892 ();
 FILLER_ASAP7_75t_R FILLER_0_199_901 ();
 FILLER_ASAP7_75t_R FILLER_0_199_909 ();
 DECAPx2_ASAP7_75t_R FILLER_0_199_919 ();
 DECAPx6_ASAP7_75t_R FILLER_0_199_927 ();
 DECAPx2_ASAP7_75t_R FILLER_0_199_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_199_950 ();
 FILLER_ASAP7_75t_R FILLER_0_199_962 ();
 FILLER_ASAP7_75t_R FILLER_0_199_969 ();
 FILLER_ASAP7_75t_R FILLER_0_199_978 ();
 DECAPx6_ASAP7_75t_R FILLER_0_199_1000 ();
 DECAPx1_ASAP7_75t_R FILLER_0_199_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_199_1018 ();
 FILLER_ASAP7_75t_R FILLER_0_199_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_199_1029 ();
 DECAPx1_ASAP7_75t_R FILLER_0_199_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_199_1044 ();
 DECAPx1_ASAP7_75t_R FILLER_0_199_1048 ();
 DECAPx1_ASAP7_75t_R FILLER_0_199_1058 ();
 DECAPx4_ASAP7_75t_R FILLER_0_199_1068 ();
 FILLER_ASAP7_75t_R FILLER_0_199_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_0_199_1097 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_199_1119 ();
 FILLER_ASAP7_75t_R FILLER_0_199_1126 ();
 FILLER_ASAP7_75t_R FILLER_0_199_1134 ();
 DECAPx6_ASAP7_75t_R FILLER_0_199_1142 ();
 DECAPx2_ASAP7_75t_R FILLER_0_199_1156 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_199_1162 ();
 FILLER_ASAP7_75t_R FILLER_0_199_1169 ();
 DECAPx2_ASAP7_75t_R FILLER_0_199_1178 ();
 FILLER_ASAP7_75t_R FILLER_0_199_1184 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_199_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_199_1195 ();
 DECAPx1_ASAP7_75t_R FILLER_0_199_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_199_1207 ();
 FILLER_ASAP7_75t_R FILLER_0_199_1213 ();
 DECAPx1_ASAP7_75t_R FILLER_0_199_1221 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_199_1225 ();
 FILLER_ASAP7_75t_R FILLER_0_199_1232 ();
 FILLER_ASAP7_75t_R FILLER_0_199_1240 ();
 FILLER_ASAP7_75t_R FILLER_0_199_1248 ();
 DECAPx2_ASAP7_75t_R FILLER_0_199_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_199_1267 ();
 FILLER_ASAP7_75t_R FILLER_0_199_1274 ();
 DECAPx10_ASAP7_75t_R FILLER_0_199_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_0_199_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_0_199_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_0_199_1353 ();
 DECAPx2_ASAP7_75t_R FILLER_0_199_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_199_1381 ();
 DECAPx2_ASAP7_75t_R FILLER_0_200_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_200_18 ();
 FILLER_ASAP7_75t_R FILLER_0_200_38 ();
 FILLER_ASAP7_75t_R FILLER_0_200_50 ();
 FILLER_ASAP7_75t_R FILLER_0_200_62 ();
 FILLER_ASAP7_75t_R FILLER_0_200_71 ();
 FILLER_ASAP7_75t_R FILLER_0_200_79 ();
 FILLER_ASAP7_75t_R FILLER_0_200_87 ();
 DECAPx4_ASAP7_75t_R FILLER_0_200_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_107 ();
 FILLER_ASAP7_75t_R FILLER_0_200_124 ();
 DECAPx2_ASAP7_75t_R FILLER_0_200_132 ();
 FILLER_ASAP7_75t_R FILLER_0_200_138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_200_146 ();
 FILLER_ASAP7_75t_R FILLER_0_200_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_154 ();
 DECAPx6_ASAP7_75t_R FILLER_0_200_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_175 ();
 FILLER_ASAP7_75t_R FILLER_0_200_182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_200_190 ();
 DECAPx4_ASAP7_75t_R FILLER_0_200_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_222 ();
 FILLER_ASAP7_75t_R FILLER_0_200_233 ();
 FILLER_ASAP7_75t_R FILLER_0_200_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_242 ();
 DECAPx2_ASAP7_75t_R FILLER_0_200_253 ();
 FILLER_ASAP7_75t_R FILLER_0_200_265 ();
 DECAPx2_ASAP7_75t_R FILLER_0_200_273 ();
 DECAPx10_ASAP7_75t_R FILLER_0_200_285 ();
 DECAPx4_ASAP7_75t_R FILLER_0_200_307 ();
 FILLER_ASAP7_75t_R FILLER_0_200_324 ();
 DECAPx4_ASAP7_75t_R FILLER_0_200_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_346 ();
 FILLER_ASAP7_75t_R FILLER_0_200_355 ();
 FILLER_ASAP7_75t_R FILLER_0_200_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_362 ();
 DECAPx1_ASAP7_75t_R FILLER_0_200_369 ();
 DECAPx1_ASAP7_75t_R FILLER_0_200_376 ();
 DECAPx1_ASAP7_75t_R FILLER_0_200_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_391 ();
 DECAPx1_ASAP7_75t_R FILLER_0_200_395 ();
 DECAPx2_ASAP7_75t_R FILLER_0_200_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_411 ();
 DECAPx10_ASAP7_75t_R FILLER_0_200_418 ();
 DECAPx1_ASAP7_75t_R FILLER_0_200_440 ();
 DECAPx4_ASAP7_75t_R FILLER_0_200_450 ();
 FILLER_ASAP7_75t_R FILLER_0_200_460 ();
 DECAPx2_ASAP7_75t_R FILLER_0_200_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_470 ();
 DECAPx2_ASAP7_75t_R FILLER_0_200_477 ();
 DECAPx10_ASAP7_75t_R FILLER_0_200_489 ();
 DECAPx1_ASAP7_75t_R FILLER_0_200_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_515 ();
 DECAPx1_ASAP7_75t_R FILLER_0_200_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_527 ();
 DECAPx1_ASAP7_75t_R FILLER_0_200_534 ();
 FILLER_ASAP7_75t_R FILLER_0_200_544 ();
 FILLER_ASAP7_75t_R FILLER_0_200_552 ();
 DECAPx2_ASAP7_75t_R FILLER_0_200_560 ();
 FILLER_ASAP7_75t_R FILLER_0_200_571 ();
 FILLER_ASAP7_75t_R FILLER_0_200_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_581 ();
 FILLER_ASAP7_75t_R FILLER_0_200_585 ();
 FILLER_ASAP7_75t_R FILLER_0_200_593 ();
 FILLER_ASAP7_75t_R FILLER_0_200_602 ();
 DECAPx10_ASAP7_75t_R FILLER_0_200_610 ();
 DECAPx2_ASAP7_75t_R FILLER_0_200_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_638 ();
 FILLER_ASAP7_75t_R FILLER_0_200_645 ();
 DECAPx4_ASAP7_75t_R FILLER_0_200_653 ();
 FILLER_ASAP7_75t_R FILLER_0_200_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_665 ();
 FILLER_ASAP7_75t_R FILLER_0_200_687 ();
 FILLER_ASAP7_75t_R FILLER_0_200_692 ();
 FILLER_ASAP7_75t_R FILLER_0_200_700 ();
 FILLER_ASAP7_75t_R FILLER_0_200_708 ();
 FILLER_ASAP7_75t_R FILLER_0_200_716 ();
 DECAPx2_ASAP7_75t_R FILLER_0_200_724 ();
 FILLER_ASAP7_75t_R FILLER_0_200_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_732 ();
 FILLER_ASAP7_75t_R FILLER_0_200_745 ();
 DECAPx1_ASAP7_75t_R FILLER_0_200_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_757 ();
 FILLER_ASAP7_75t_R FILLER_0_200_764 ();
 DECAPx2_ASAP7_75t_R FILLER_0_200_772 ();
 FILLER_ASAP7_75t_R FILLER_0_200_785 ();
 DECAPx4_ASAP7_75t_R FILLER_0_200_790 ();
 FILLER_ASAP7_75t_R FILLER_0_200_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_802 ();
 FILLER_ASAP7_75t_R FILLER_0_200_809 ();
 FILLER_ASAP7_75t_R FILLER_0_200_817 ();
 DECAPx6_ASAP7_75t_R FILLER_0_200_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_839 ();
 DECAPx4_ASAP7_75t_R FILLER_0_200_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_857 ();
 DECAPx4_ASAP7_75t_R FILLER_0_200_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_874 ();
 DECAPx6_ASAP7_75t_R FILLER_0_200_878 ();
 DECAPx1_ASAP7_75t_R FILLER_0_200_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_896 ();
 DECAPx2_ASAP7_75t_R FILLER_0_200_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_200_919 ();
 FILLER_ASAP7_75t_R FILLER_0_200_925 ();
 DECAPx1_ASAP7_75t_R FILLER_0_200_933 ();
 DECAPx1_ASAP7_75t_R FILLER_0_200_943 ();
 DECAPx2_ASAP7_75t_R FILLER_0_200_953 ();
 FILLER_ASAP7_75t_R FILLER_0_200_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_961 ();
 FILLER_ASAP7_75t_R FILLER_0_200_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_970 ();
 FILLER_ASAP7_75t_R FILLER_0_200_977 ();
 DECAPx10_ASAP7_75t_R FILLER_0_200_984 ();
 DECAPx2_ASAP7_75t_R FILLER_0_200_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_1012 ();
 FILLER_ASAP7_75t_R FILLER_0_200_1019 ();
 DECAPx2_ASAP7_75t_R FILLER_0_200_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_1033 ();
 DECAPx6_ASAP7_75t_R FILLER_0_200_1039 ();
 DECAPx1_ASAP7_75t_R FILLER_0_200_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_1057 ();
 FILLER_ASAP7_75t_R FILLER_0_200_1064 ();
 DECAPx2_ASAP7_75t_R FILLER_0_200_1072 ();
 FILLER_ASAP7_75t_R FILLER_0_200_1078 ();
 FILLER_ASAP7_75t_R FILLER_0_200_1086 ();
 DECAPx2_ASAP7_75t_R FILLER_0_200_1096 ();
 FILLER_ASAP7_75t_R FILLER_0_200_1102 ();
 DECAPx4_ASAP7_75t_R FILLER_0_200_1111 ();
 FILLER_ASAP7_75t_R FILLER_0_200_1127 ();
 DECAPx2_ASAP7_75t_R FILLER_0_200_1135 ();
 FILLER_ASAP7_75t_R FILLER_0_200_1147 ();
 FILLER_ASAP7_75t_R FILLER_0_200_1156 ();
 DECAPx4_ASAP7_75t_R FILLER_0_200_1164 ();
 FILLER_ASAP7_75t_R FILLER_0_200_1174 ();
 DECAPx1_ASAP7_75t_R FILLER_0_200_1182 ();
 FILLER_ASAP7_75t_R FILLER_0_200_1192 ();
 FILLER_ASAP7_75t_R FILLER_0_200_1200 ();
 DECAPx1_ASAP7_75t_R FILLER_0_200_1208 ();
 DECAPx2_ASAP7_75t_R FILLER_0_200_1218 ();
 FILLER_ASAP7_75t_R FILLER_0_200_1224 ();
 DECAPx6_ASAP7_75t_R FILLER_0_200_1231 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200_1245 ();
 FILLER_ASAP7_75t_R FILLER_0_200_1252 ();
 DECAPx6_ASAP7_75t_R FILLER_0_200_1258 ();
 FILLER_ASAP7_75t_R FILLER_0_200_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_200_1286 ();
 DECAPx10_ASAP7_75t_R FILLER_0_200_1308 ();
 DECAPx10_ASAP7_75t_R FILLER_0_200_1330 ();
 DECAPx10_ASAP7_75t_R FILLER_0_200_1352 ();
 DECAPx2_ASAP7_75t_R FILLER_0_200_1374 ();
 FILLER_ASAP7_75t_R FILLER_0_200_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_201_2 ();
 FILLER_ASAP7_75t_R FILLER_0_201_10 ();
 DECAPx4_ASAP7_75t_R FILLER_0_201_23 ();
 FILLER_ASAP7_75t_R FILLER_0_201_38 ();
 FILLER_ASAP7_75t_R FILLER_0_201_45 ();
 DECAPx4_ASAP7_75t_R FILLER_0_201_55 ();
 DECAPx1_ASAP7_75t_R FILLER_0_201_76 ();
 FILLER_ASAP7_75t_R FILLER_0_201_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_88 ();
 FILLER_ASAP7_75t_R FILLER_0_201_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_97 ();
 DECAPx2_ASAP7_75t_R FILLER_0_201_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_109 ();
 FILLER_ASAP7_75t_R FILLER_0_201_115 ();
 FILLER_ASAP7_75t_R FILLER_0_201_125 ();
 DECAPx10_ASAP7_75t_R FILLER_0_201_135 ();
 DECAPx6_ASAP7_75t_R FILLER_0_201_157 ();
 DECAPx2_ASAP7_75t_R FILLER_0_201_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_177 ();
 FILLER_ASAP7_75t_R FILLER_0_201_184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_201_192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_201_214 ();
 FILLER_ASAP7_75t_R FILLER_0_201_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_230 ();
 FILLER_ASAP7_75t_R FILLER_0_201_237 ();
 DECAPx4_ASAP7_75t_R FILLER_0_201_249 ();
 DECAPx10_ASAP7_75t_R FILLER_0_201_269 ();
 DECAPx10_ASAP7_75t_R FILLER_0_201_291 ();
 DECAPx6_ASAP7_75t_R FILLER_0_201_313 ();
 DECAPx1_ASAP7_75t_R FILLER_0_201_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_331 ();
 FILLER_ASAP7_75t_R FILLER_0_201_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_340 ();
 FILLER_ASAP7_75t_R FILLER_0_201_349 ();
 FILLER_ASAP7_75t_R FILLER_0_201_358 ();
 DECAPx6_ASAP7_75t_R FILLER_0_201_367 ();
 FILLER_ASAP7_75t_R FILLER_0_201_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_383 ();
 FILLER_ASAP7_75t_R FILLER_0_201_390 ();
 DECAPx6_ASAP7_75t_R FILLER_0_201_398 ();
 DECAPx1_ASAP7_75t_R FILLER_0_201_412 ();
 FILLER_ASAP7_75t_R FILLER_0_201_424 ();
 FILLER_ASAP7_75t_R FILLER_0_201_429 ();
 FILLER_ASAP7_75t_R FILLER_0_201_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_440 ();
 FILLER_ASAP7_75t_R FILLER_0_201_444 ();
 DECAPx6_ASAP7_75t_R FILLER_0_201_454 ();
 FILLER_ASAP7_75t_R FILLER_0_201_474 ();
 DECAPx1_ASAP7_75t_R FILLER_0_201_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_486 ();
 DECAPx2_ASAP7_75t_R FILLER_0_201_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_499 ();
 DECAPx4_ASAP7_75t_R FILLER_0_201_506 ();
 FILLER_ASAP7_75t_R FILLER_0_201_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_518 ();
 FILLER_ASAP7_75t_R FILLER_0_201_528 ();
 DECAPx6_ASAP7_75t_R FILLER_0_201_536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_201_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_554 ();
 DECAPx6_ASAP7_75t_R FILLER_0_201_561 ();
 FILLER_ASAP7_75t_R FILLER_0_201_582 ();
 DECAPx1_ASAP7_75t_R FILLER_0_201_592 ();
 FILLER_ASAP7_75t_R FILLER_0_201_599 ();
 FILLER_ASAP7_75t_R FILLER_0_201_609 ();
 DECAPx2_ASAP7_75t_R FILLER_0_201_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_623 ();
 FILLER_ASAP7_75t_R FILLER_0_201_630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_201_635 ();
 DECAPx6_ASAP7_75t_R FILLER_0_201_657 ();
 DECAPx1_ASAP7_75t_R FILLER_0_201_671 ();
 FILLER_ASAP7_75t_R FILLER_0_201_687 ();
 FILLER_ASAP7_75t_R FILLER_0_201_692 ();
 DECAPx1_ASAP7_75t_R FILLER_0_201_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_704 ();
 DECAPx10_ASAP7_75t_R FILLER_0_201_708 ();
 DECAPx2_ASAP7_75t_R FILLER_0_201_730 ();
 FILLER_ASAP7_75t_R FILLER_0_201_736 ();
 FILLER_ASAP7_75t_R FILLER_0_201_748 ();
 FILLER_ASAP7_75t_R FILLER_0_201_768 ();
 FILLER_ASAP7_75t_R FILLER_0_201_781 ();
 DECAPx4_ASAP7_75t_R FILLER_0_201_791 ();
 FILLER_ASAP7_75t_R FILLER_0_201_807 ();
 FILLER_ASAP7_75t_R FILLER_0_201_815 ();
 FILLER_ASAP7_75t_R FILLER_0_201_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_829 ();
 FILLER_ASAP7_75t_R FILLER_0_201_838 ();
 FILLER_ASAP7_75t_R FILLER_0_201_850 ();
 DECAPx6_ASAP7_75t_R FILLER_0_201_856 ();
 FILLER_ASAP7_75t_R FILLER_0_201_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_201_883 ();
 DECAPx2_ASAP7_75t_R FILLER_0_201_905 ();
 FILLER_ASAP7_75t_R FILLER_0_201_916 ();
 FILLER_ASAP7_75t_R FILLER_0_201_923 ();
 DECAPx4_ASAP7_75t_R FILLER_0_201_927 ();
 FILLER_ASAP7_75t_R FILLER_0_201_943 ();
 DECAPx6_ASAP7_75t_R FILLER_0_201_951 ();
 FILLER_ASAP7_75t_R FILLER_0_201_965 ();
 FILLER_ASAP7_75t_R FILLER_0_201_973 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_975 ();
 DECAPx2_ASAP7_75t_R FILLER_0_201_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_988 ();
 FILLER_ASAP7_75t_R FILLER_0_201_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_201_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_1024 ();
 FILLER_ASAP7_75t_R FILLER_0_201_1031 ();
 FILLER_ASAP7_75t_R FILLER_0_201_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_1045 ();
 DECAPx1_ASAP7_75t_R FILLER_0_201_1053 ();
 DECAPx1_ASAP7_75t_R FILLER_0_201_1063 ();
 DECAPx1_ASAP7_75t_R FILLER_0_201_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_1082 ();
 DECAPx2_ASAP7_75t_R FILLER_0_201_1089 ();
 FILLER_ASAP7_75t_R FILLER_0_201_1095 ();
 FILLER_ASAP7_75t_R FILLER_0_201_1100 ();
 FILLER_ASAP7_75t_R FILLER_0_201_1109 ();
 DECAPx2_ASAP7_75t_R FILLER_0_201_1118 ();
 FILLER_ASAP7_75t_R FILLER_0_201_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_1126 ();
 DECAPx6_ASAP7_75t_R FILLER_0_201_1133 ();
 DECAPx2_ASAP7_75t_R FILLER_0_201_1157 ();
 FILLER_ASAP7_75t_R FILLER_0_201_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_1165 ();
 DECAPx6_ASAP7_75t_R FILLER_0_201_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_1191 ();
 FILLER_ASAP7_75t_R FILLER_0_201_1198 ();
 FILLER_ASAP7_75t_R FILLER_0_201_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_1209 ();
 DECAPx4_ASAP7_75t_R FILLER_0_201_1217 ();
 FILLER_ASAP7_75t_R FILLER_0_201_1227 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_1229 ();
 DECAPx1_ASAP7_75t_R FILLER_0_201_1236 ();
 FILLER_ASAP7_75t_R FILLER_0_201_1246 ();
 FILLER_ASAP7_75t_R FILLER_0_201_1253 ();
 FILLER_ASAP7_75t_R FILLER_0_201_1261 ();
 DECAPx2_ASAP7_75t_R FILLER_0_201_1269 ();
 FILLER_ASAP7_75t_R FILLER_0_201_1275 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201_1277 ();
 DECAPx10_ASAP7_75t_R FILLER_0_201_1284 ();
 DECAPx10_ASAP7_75t_R FILLER_0_201_1306 ();
 DECAPx10_ASAP7_75t_R FILLER_0_201_1328 ();
 DECAPx10_ASAP7_75t_R FILLER_0_201_1350 ();
 DECAPx4_ASAP7_75t_R FILLER_0_201_1372 ();
 DECAPx2_ASAP7_75t_R FILLER_0_202_2 ();
 FILLER_ASAP7_75t_R FILLER_0_202_13 ();
 FILLER_ASAP7_75t_R FILLER_0_202_21 ();
 FILLER_ASAP7_75t_R FILLER_0_202_27 ();
 DECAPx4_ASAP7_75t_R FILLER_0_202_32 ();
 FILLER_ASAP7_75t_R FILLER_0_202_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_44 ();
 DECAPx2_ASAP7_75t_R FILLER_0_202_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_57 ();
 FILLER_ASAP7_75t_R FILLER_0_202_65 ();
 FILLER_ASAP7_75t_R FILLER_0_202_77 ();
 DECAPx2_ASAP7_75t_R FILLER_0_202_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_91 ();
 DECAPx10_ASAP7_75t_R FILLER_0_202_98 ();
 DECAPx4_ASAP7_75t_R FILLER_0_202_120 ();
 FILLER_ASAP7_75t_R FILLER_0_202_135 ();
 FILLER_ASAP7_75t_R FILLER_0_202_143 ();
 DECAPx4_ASAP7_75t_R FILLER_0_202_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_161 ();
 FILLER_ASAP7_75t_R FILLER_0_202_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_170 ();
 FILLER_ASAP7_75t_R FILLER_0_202_177 ();
 FILLER_ASAP7_75t_R FILLER_0_202_190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_202_199 ();
 FILLER_ASAP7_75t_R FILLER_0_202_221 ();
 FILLER_ASAP7_75t_R FILLER_0_202_233 ();
 FILLER_ASAP7_75t_R FILLER_0_202_242 ();
 FILLER_ASAP7_75t_R FILLER_0_202_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_256 ();
 DECAPx1_ASAP7_75t_R FILLER_0_202_279 ();
 FILLER_ASAP7_75t_R FILLER_0_202_286 ();
 DECAPx4_ASAP7_75t_R FILLER_0_202_298 ();
 FILLER_ASAP7_75t_R FILLER_0_202_314 ();
 FILLER_ASAP7_75t_R FILLER_0_202_322 ();
 FILLER_ASAP7_75t_R FILLER_0_202_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_332 ();
 FILLER_ASAP7_75t_R FILLER_0_202_339 ();
 DECAPx4_ASAP7_75t_R FILLER_0_202_344 ();
 DECAPx4_ASAP7_75t_R FILLER_0_202_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_370 ();
 DECAPx1_ASAP7_75t_R FILLER_0_202_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_390 ();
 FILLER_ASAP7_75t_R FILLER_0_202_397 ();
 DECAPx2_ASAP7_75t_R FILLER_0_202_405 ();
 FILLER_ASAP7_75t_R FILLER_0_202_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_413 ();
 FILLER_ASAP7_75t_R FILLER_0_202_417 ();
 DECAPx2_ASAP7_75t_R FILLER_0_202_427 ();
 FILLER_ASAP7_75t_R FILLER_0_202_433 ();
 DECAPx2_ASAP7_75t_R FILLER_0_202_441 ();
 DECAPx2_ASAP7_75t_R FILLER_0_202_453 ();
 FILLER_ASAP7_75t_R FILLER_0_202_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_461 ();
 FILLER_ASAP7_75t_R FILLER_0_202_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_466 ();
 FILLER_ASAP7_75t_R FILLER_0_202_489 ();
 DECAPx1_ASAP7_75t_R FILLER_0_202_497 ();
 DECAPx2_ASAP7_75t_R FILLER_0_202_509 ();
 FILLER_ASAP7_75t_R FILLER_0_202_515 ();
 DECAPx2_ASAP7_75t_R FILLER_0_202_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_529 ();
 DECAPx6_ASAP7_75t_R FILLER_0_202_536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_202_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_554 ();
 DECAPx1_ASAP7_75t_R FILLER_0_202_565 ();
 DECAPx1_ASAP7_75t_R FILLER_0_202_591 ();
 DECAPx4_ASAP7_75t_R FILLER_0_202_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_612 ();
 DECAPx6_ASAP7_75t_R FILLER_0_202_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_634 ();
 FILLER_ASAP7_75t_R FILLER_0_202_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_644 ();
 FILLER_ASAP7_75t_R FILLER_0_202_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_653 ();
 DECAPx6_ASAP7_75t_R FILLER_0_202_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_674 ();
 DECAPx6_ASAP7_75t_R FILLER_0_202_687 ();
 DECAPx2_ASAP7_75t_R FILLER_0_202_701 ();
 FILLER_ASAP7_75t_R FILLER_0_202_713 ();
 DECAPx10_ASAP7_75t_R FILLER_0_202_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_743 ();
 FILLER_ASAP7_75t_R FILLER_0_202_750 ();
 FILLER_ASAP7_75t_R FILLER_0_202_758 ();
 FILLER_ASAP7_75t_R FILLER_0_202_766 ();
 FILLER_ASAP7_75t_R FILLER_0_202_774 ();
 FILLER_ASAP7_75t_R FILLER_0_202_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_781 ();
 DECAPx6_ASAP7_75t_R FILLER_0_202_788 ();
 DECAPx2_ASAP7_75t_R FILLER_0_202_805 ();
 FILLER_ASAP7_75t_R FILLER_0_202_811 ();
 DECAPx10_ASAP7_75t_R FILLER_0_202_819 ();
 FILLER_ASAP7_75t_R FILLER_0_202_841 ();
 DECAPx2_ASAP7_75t_R FILLER_0_202_851 ();
 DECAPx2_ASAP7_75t_R FILLER_0_202_863 ();
 FILLER_ASAP7_75t_R FILLER_0_202_875 ();
 DECAPx4_ASAP7_75t_R FILLER_0_202_886 ();
 FILLER_ASAP7_75t_R FILLER_0_202_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_898 ();
 DECAPx1_ASAP7_75t_R FILLER_0_202_909 ();
 FILLER_ASAP7_75t_R FILLER_0_202_922 ();
 FILLER_ASAP7_75t_R FILLER_0_202_930 ();
 DECAPx6_ASAP7_75t_R FILLER_0_202_938 ();
 DECAPx2_ASAP7_75t_R FILLER_0_202_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_974 ();
 DECAPx2_ASAP7_75t_R FILLER_0_202_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_992 ();
 FILLER_ASAP7_75t_R FILLER_0_202_999 ();
 DECAPx10_ASAP7_75t_R FILLER_0_202_1009 ();
 FILLER_ASAP7_75t_R FILLER_0_202_1031 ();
 FILLER_ASAP7_75t_R FILLER_0_202_1039 ();
 FILLER_ASAP7_75t_R FILLER_0_202_1047 ();
 DECAPx1_ASAP7_75t_R FILLER_0_202_1055 ();
 FILLER_ASAP7_75t_R FILLER_0_202_1065 ();
 FILLER_ASAP7_75t_R FILLER_0_202_1073 ();
 DECAPx1_ASAP7_75t_R FILLER_0_202_1081 ();
 FILLER_ASAP7_75t_R FILLER_0_202_1095 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_1097 ();
 FILLER_ASAP7_75t_R FILLER_0_202_1104 ();
 DECAPx6_ASAP7_75t_R FILLER_0_202_1112 ();
 DECAPx1_ASAP7_75t_R FILLER_0_202_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_1130 ();
 FILLER_ASAP7_75t_R FILLER_0_202_1137 ();
 DECAPx2_ASAP7_75t_R FILLER_0_202_1142 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_1148 ();
 FILLER_ASAP7_75t_R FILLER_0_202_1155 ();
 DECAPx1_ASAP7_75t_R FILLER_0_202_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_1167 ();
 FILLER_ASAP7_75t_R FILLER_0_202_1174 ();
 DECAPx6_ASAP7_75t_R FILLER_0_202_1182 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_1196 ();
 FILLER_ASAP7_75t_R FILLER_0_202_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_1206 ();
 DECAPx1_ASAP7_75t_R FILLER_0_202_1213 ();
 DECAPx1_ASAP7_75t_R FILLER_0_202_1233 ();
 DECAPx2_ASAP7_75t_R FILLER_0_202_1243 ();
 FILLER_ASAP7_75t_R FILLER_0_202_1249 ();
 DECAPx1_ASAP7_75t_R FILLER_0_202_1259 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202_1263 ();
 DECAPx10_ASAP7_75t_R FILLER_0_202_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_202_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_202_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_202_1338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_202_1360 ();
 FILLER_ASAP7_75t_R FILLER_0_203_2 ();
 FILLER_ASAP7_75t_R FILLER_0_203_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_11 ();
 FILLER_ASAP7_75t_R FILLER_0_203_20 ();
 FILLER_ASAP7_75t_R FILLER_0_203_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_29 ();
 DECAPx2_ASAP7_75t_R FILLER_0_203_36 ();
 FILLER_ASAP7_75t_R FILLER_0_203_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_44 ();
 DECAPx4_ASAP7_75t_R FILLER_0_203_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_61 ();
 DECAPx1_ASAP7_75t_R FILLER_0_203_68 ();
 FILLER_ASAP7_75t_R FILLER_0_203_78 ();
 FILLER_ASAP7_75t_R FILLER_0_203_91 ();
 DECAPx2_ASAP7_75t_R FILLER_0_203_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_105 ();
 FILLER_ASAP7_75t_R FILLER_0_203_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_114 ();
 DECAPx1_ASAP7_75t_R FILLER_0_203_123 ();
 FILLER_ASAP7_75t_R FILLER_0_203_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_137 ();
 FILLER_ASAP7_75t_R FILLER_0_203_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_146 ();
 FILLER_ASAP7_75t_R FILLER_0_203_153 ();
 FILLER_ASAP7_75t_R FILLER_0_203_161 ();
 DECAPx1_ASAP7_75t_R FILLER_0_203_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_178 ();
 FILLER_ASAP7_75t_R FILLER_0_203_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_188 ();
 DECAPx6_ASAP7_75t_R FILLER_0_203_195 ();
 DECAPx2_ASAP7_75t_R FILLER_0_203_209 ();
 DECAPx10_ASAP7_75t_R FILLER_0_203_221 ();
 DECAPx4_ASAP7_75t_R FILLER_0_203_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_253 ();
 DECAPx6_ASAP7_75t_R FILLER_0_203_261 ();
 FILLER_ASAP7_75t_R FILLER_0_203_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_277 ();
 DECAPx2_ASAP7_75t_R FILLER_0_203_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_289 ();
 FILLER_ASAP7_75t_R FILLER_0_203_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_298 ();
 DECAPx6_ASAP7_75t_R FILLER_0_203_305 ();
 FILLER_ASAP7_75t_R FILLER_0_203_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_321 ();
 DECAPx2_ASAP7_75t_R FILLER_0_203_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_203_341 ();
 DECAPx10_ASAP7_75t_R FILLER_0_203_366 ();
 DECAPx1_ASAP7_75t_R FILLER_0_203_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_392 ();
 FILLER_ASAP7_75t_R FILLER_0_203_399 ();
 DECAPx10_ASAP7_75t_R FILLER_0_203_408 ();
 DECAPx10_ASAP7_75t_R FILLER_0_203_430 ();
 DECAPx6_ASAP7_75t_R FILLER_0_203_452 ();
 FILLER_ASAP7_75t_R FILLER_0_203_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_474 ();
 FILLER_ASAP7_75t_R FILLER_0_203_478 ();
 FILLER_ASAP7_75t_R FILLER_0_203_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_488 ();
 DECAPx1_ASAP7_75t_R FILLER_0_203_495 ();
 DECAPx2_ASAP7_75t_R FILLER_0_203_505 ();
 FILLER_ASAP7_75t_R FILLER_0_203_511 ();
 DECAPx1_ASAP7_75t_R FILLER_0_203_519 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_523 ();
 FILLER_ASAP7_75t_R FILLER_0_203_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_531 ();
 DECAPx1_ASAP7_75t_R FILLER_0_203_538 ();
 FILLER_ASAP7_75t_R FILLER_0_203_554 ();
 DECAPx4_ASAP7_75t_R FILLER_0_203_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_572 ();
 DECAPx2_ASAP7_75t_R FILLER_0_203_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_592 ();
 DECAPx2_ASAP7_75t_R FILLER_0_203_599 ();
 FILLER_ASAP7_75t_R FILLER_0_203_605 ();
 FILLER_ASAP7_75t_R FILLER_0_203_613 ();
 FILLER_ASAP7_75t_R FILLER_0_203_621 ();
 FILLER_ASAP7_75t_R FILLER_0_203_645 ();
 FILLER_ASAP7_75t_R FILLER_0_203_653 ();
 DECAPx6_ASAP7_75t_R FILLER_0_203_658 ();
 DECAPx1_ASAP7_75t_R FILLER_0_203_672 ();
 DECAPx6_ASAP7_75t_R FILLER_0_203_688 ();
 FILLER_ASAP7_75t_R FILLER_0_203_702 ();
 FILLER_ASAP7_75t_R FILLER_0_203_710 ();
 DECAPx2_ASAP7_75t_R FILLER_0_203_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_724 ();
 DECAPx6_ASAP7_75t_R FILLER_0_203_731 ();
 FILLER_ASAP7_75t_R FILLER_0_203_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_747 ();
 FILLER_ASAP7_75t_R FILLER_0_203_753 ();
 FILLER_ASAP7_75t_R FILLER_0_203_760 ();
 DECAPx6_ASAP7_75t_R FILLER_0_203_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_782 ();
 DECAPx6_ASAP7_75t_R FILLER_0_203_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_805 ();
 FILLER_ASAP7_75t_R FILLER_0_203_812 ();
 FILLER_ASAP7_75t_R FILLER_0_203_820 ();
 DECAPx2_ASAP7_75t_R FILLER_0_203_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_833 ();
 DECAPx1_ASAP7_75t_R FILLER_0_203_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_848 ();
 FILLER_ASAP7_75t_R FILLER_0_203_864 ();
 DECAPx2_ASAP7_75t_R FILLER_0_203_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_875 ();
 DECAPx2_ASAP7_75t_R FILLER_0_203_882 ();
 FILLER_ASAP7_75t_R FILLER_0_203_888 ();
 FILLER_ASAP7_75t_R FILLER_0_203_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_899 ();
 FILLER_ASAP7_75t_R FILLER_0_203_908 ();
 DECAPx2_ASAP7_75t_R FILLER_0_203_916 ();
 FILLER_ASAP7_75t_R FILLER_0_203_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_924 ();
 FILLER_ASAP7_75t_R FILLER_0_203_927 ();
 FILLER_ASAP7_75t_R FILLER_0_203_937 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_939 ();
 FILLER_ASAP7_75t_R FILLER_0_203_946 ();
 FILLER_ASAP7_75t_R FILLER_0_203_954 ();
 DECAPx6_ASAP7_75t_R FILLER_0_203_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_976 ();
 DECAPx6_ASAP7_75t_R FILLER_0_203_983 ();
 FILLER_ASAP7_75t_R FILLER_0_203_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_999 ();
 DECAPx10_ASAP7_75t_R FILLER_0_203_1006 ();
 DECAPx2_ASAP7_75t_R FILLER_0_203_1028 ();
 FILLER_ASAP7_75t_R FILLER_0_203_1034 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_1036 ();
 DECAPx1_ASAP7_75t_R FILLER_0_203_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_1053 ();
 FILLER_ASAP7_75t_R FILLER_0_203_1057 ();
 DECAPx4_ASAP7_75t_R FILLER_0_203_1065 ();
 DECAPx4_ASAP7_75t_R FILLER_0_203_1082 ();
 FILLER_ASAP7_75t_R FILLER_0_203_1092 ();
 FILLER_ASAP7_75t_R FILLER_0_203_1102 ();
 FILLER_ASAP7_75t_R FILLER_0_203_1110 ();
 DECAPx1_ASAP7_75t_R FILLER_0_203_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_1121 ();
 FILLER_ASAP7_75t_R FILLER_0_203_1128 ();
 FILLER_ASAP7_75t_R FILLER_0_203_1136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_203_1145 ();
 DECAPx6_ASAP7_75t_R FILLER_0_203_1167 ();
 FILLER_ASAP7_75t_R FILLER_0_203_1181 ();
 FILLER_ASAP7_75t_R FILLER_0_203_1193 ();
 DECAPx1_ASAP7_75t_R FILLER_0_203_1201 ();
 DECAPx4_ASAP7_75t_R FILLER_0_203_1210 ();
 FILLER_ASAP7_75t_R FILLER_0_203_1220 ();
 FILLER_ASAP7_75t_R FILLER_0_203_1233 ();
 DECAPx2_ASAP7_75t_R FILLER_0_203_1241 ();
 DECAPx2_ASAP7_75t_R FILLER_0_203_1253 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_1259 ();
 FILLER_ASAP7_75t_R FILLER_0_203_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_203_1275 ();
 DECAPx10_ASAP7_75t_R FILLER_0_203_1297 ();
 DECAPx10_ASAP7_75t_R FILLER_0_203_1319 ();
 DECAPx10_ASAP7_75t_R FILLER_0_203_1341 ();
 DECAPx6_ASAP7_75t_R FILLER_0_203_1363 ();
 DECAPx1_ASAP7_75t_R FILLER_0_203_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_204_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_204_4 ();
 DECAPx1_ASAP7_75t_R FILLER_0_204_11 ();
 DECAPx2_ASAP7_75t_R FILLER_0_204_21 ();
 FILLER_ASAP7_75t_R FILLER_0_204_27 ();
 FILLER_ASAP7_75t_R FILLER_0_204_35 ();
 FILLER_ASAP7_75t_R FILLER_0_204_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_204_45 ();
 DECAPx10_ASAP7_75t_R FILLER_0_204_52 ();
 DECAPx4_ASAP7_75t_R FILLER_0_204_74 ();
 FILLER_ASAP7_75t_R FILLER_0_204_84 ();
 DECAPx4_ASAP7_75t_R FILLER_0_204_92 ();
 FILLER_ASAP7_75t_R FILLER_0_204_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_204_104 ();
 DECAPx4_ASAP7_75t_R FILLER_0_204_115 ();
 FILLER_ASAP7_75t_R FILLER_0_204_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_204_139 ();
 DECAPx6_ASAP7_75t_R FILLER_0_204_143 ();
 DECAPx2_ASAP7_75t_R FILLER_0_204_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_204_163 ();
 DECAPx6_ASAP7_75t_R FILLER_0_204_170 ();
 DECAPx1_ASAP7_75t_R FILLER_0_204_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_204_188 ();
 DECAPx2_ASAP7_75t_R FILLER_0_204_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_204_198 ();
 DECAPx2_ASAP7_75t_R FILLER_0_204_202 ();
 FILLER_ASAP7_75t_R FILLER_0_204_208 ();
 DECAPx4_ASAP7_75t_R FILLER_0_204_221 ();
 FILLER_ASAP7_75t_R FILLER_0_204_238 ();
 FILLER_ASAP7_75t_R FILLER_0_204_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_204_245 ();
 FILLER_ASAP7_75t_R FILLER_0_204_249 ();
 DECAPx1_ASAP7_75t_R FILLER_0_204_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_204_261 ();
 DECAPx2_ASAP7_75t_R FILLER_0_204_268 ();
 FILLER_ASAP7_75t_R FILLER_0_204_274 ();
 FILLER_ASAP7_75t_R FILLER_0_204_282 ();
 FILLER_ASAP7_75t_R FILLER_0_204_290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_204_298 ();
 FILLER_ASAP7_75t_R FILLER_0_204_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_204_306 ();
 FILLER_ASAP7_75t_R FILLER_0_204_314 ();
 FILLER_ASAP7_75t_R FILLER_0_204_324 ();
 DECAPx2_ASAP7_75t_R FILLER_0_204_332 ();
 DECAPx4_ASAP7_75t_R FILLER_0_204_344 ();
 FILLER_ASAP7_75t_R FILLER_0_204_354 ();
 FILLER_ASAP7_75t_R FILLER_0_204_359 ();
 DECAPx1_ASAP7_75t_R FILLER_0_204_364 ();
 DECAPx10_ASAP7_75t_R FILLER_0_204_375 ();
 DECAPx6_ASAP7_75t_R FILLER_0_204_397 ();
 DECAPx2_ASAP7_75t_R FILLER_0_204_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_204_417 ();
 DECAPx4_ASAP7_75t_R FILLER_0_204_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_204_435 ();
 FILLER_ASAP7_75t_R FILLER_0_204_442 ();
 DECAPx4_ASAP7_75t_R FILLER_0_204_450 ();
 FILLER_ASAP7_75t_R FILLER_0_204_460 ();
 DECAPx10_ASAP7_75t_R FILLER_0_204_464 ();
 DECAPx6_ASAP7_75t_R FILLER_0_204_486 ();
 DECAPx2_ASAP7_75t_R FILLER_0_204_500 ();
 DECAPx2_ASAP7_75t_R FILLER_0_204_512 ();
 FILLER_ASAP7_75t_R FILLER_0_204_518 ();
 FILLER_ASAP7_75t_R FILLER_0_204_523 ();
 DECAPx2_ASAP7_75t_R FILLER_0_204_530 ();
 FILLER_ASAP7_75t_R FILLER_0_204_542 ();
 FILLER_ASAP7_75t_R FILLER_0_204_550 ();
 DECAPx6_ASAP7_75t_R FILLER_0_204_558 ();
 FILLER_ASAP7_75t_R FILLER_0_204_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_204_574 ();
 FILLER_ASAP7_75t_R FILLER_0_204_581 ();
 FILLER_ASAP7_75t_R FILLER_0_204_589 ();
 FILLER_ASAP7_75t_R FILLER_0_204_597 ();
 DECAPx1_ASAP7_75t_R FILLER_0_204_602 ();
 FILLER_ASAP7_75t_R FILLER_0_204_612 ();
 DECAPx1_ASAP7_75t_R FILLER_0_204_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_204_624 ();
 FILLER_ASAP7_75t_R FILLER_0_204_631 ();
 FILLER_ASAP7_75t_R FILLER_0_204_636 ();
 FILLER_ASAP7_75t_R FILLER_0_204_646 ();
 DECAPx10_ASAP7_75t_R FILLER_0_204_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_204_676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_204_689 ();
 FILLER_ASAP7_75t_R FILLER_0_204_711 ();
 FILLER_ASAP7_75t_R FILLER_0_204_719 ();
 FILLER_ASAP7_75t_R FILLER_0_204_724 ();
 DECAPx1_ASAP7_75t_R FILLER_0_204_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_204_740 ();
 DECAPx4_ASAP7_75t_R FILLER_0_204_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_204_757 ();
 FILLER_ASAP7_75t_R FILLER_0_204_768 ();
 FILLER_ASAP7_75t_R FILLER_0_204_780 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_204_782 ();
 DECAPx2_ASAP7_75t_R FILLER_0_204_789 ();
 DECAPx4_ASAP7_75t_R FILLER_0_204_804 ();
 DECAPx2_ASAP7_75t_R FILLER_0_204_820 ();
 DECAPx4_ASAP7_75t_R FILLER_0_204_832 ();
 DECAPx2_ASAP7_75t_R FILLER_0_204_848 ();
 FILLER_ASAP7_75t_R FILLER_0_204_854 ();
 FILLER_ASAP7_75t_R FILLER_0_204_862 ();
 FILLER_ASAP7_75t_R FILLER_0_204_874 ();
 FILLER_ASAP7_75t_R FILLER_0_204_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_204_890 ();
 DECAPx2_ASAP7_75t_R FILLER_0_204_914 ();
 FILLER_ASAP7_75t_R FILLER_0_204_926 ();
 FILLER_ASAP7_75t_R FILLER_0_204_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_204_936 ();
 DECAPx1_ASAP7_75t_R FILLER_0_204_943 ();
 FILLER_ASAP7_75t_R FILLER_0_204_954 ();
 DECAPx6_ASAP7_75t_R FILLER_0_204_962 ();
 DECAPx1_ASAP7_75t_R FILLER_0_204_976 ();
 DECAPx6_ASAP7_75t_R FILLER_0_204_986 ();
 FILLER_ASAP7_75t_R FILLER_0_204_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_204_1002 ();
 DECAPx4_ASAP7_75t_R FILLER_0_204_1009 ();
 FILLER_ASAP7_75t_R FILLER_0_204_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_204_1021 ();
 FILLER_ASAP7_75t_R FILLER_0_204_1029 ();
 FILLER_ASAP7_75t_R FILLER_0_204_1042 ();
 DECAPx2_ASAP7_75t_R FILLER_0_204_1049 ();
 FILLER_ASAP7_75t_R FILLER_0_204_1055 ();
 DECAPx4_ASAP7_75t_R FILLER_0_204_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_204_1077 ();
 FILLER_ASAP7_75t_R FILLER_0_204_1084 ();
 FILLER_ASAP7_75t_R FILLER_0_204_1091 ();
 DECAPx1_ASAP7_75t_R FILLER_0_204_1103 ();
 FILLER_ASAP7_75t_R FILLER_0_204_1117 ();
 FILLER_ASAP7_75t_R FILLER_0_204_1125 ();
 DECAPx6_ASAP7_75t_R FILLER_0_204_1130 ();
 FILLER_ASAP7_75t_R FILLER_0_204_1154 ();
 DECAPx10_ASAP7_75t_R FILLER_0_204_1166 ();
 FILLER_ASAP7_75t_R FILLER_0_204_1194 ();
 FILLER_ASAP7_75t_R FILLER_0_204_1202 ();
 FILLER_ASAP7_75t_R FILLER_0_204_1210 ();
 FILLER_ASAP7_75t_R FILLER_0_204_1218 ();
 FILLER_ASAP7_75t_R FILLER_0_204_1226 ();
 DECAPx2_ASAP7_75t_R FILLER_0_204_1234 ();
 FILLER_ASAP7_75t_R FILLER_0_204_1240 ();
 FILLER_ASAP7_75t_R FILLER_0_204_1248 ();
 DECAPx1_ASAP7_75t_R FILLER_0_204_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_204_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_0_204_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_204_1294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_204_1316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_204_1338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_204_1360 ();
 DECAPx1_ASAP7_75t_R FILLER_0_205_2 ();
 FILLER_ASAP7_75t_R FILLER_0_205_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_14 ();
 DECAPx1_ASAP7_75t_R FILLER_0_205_23 ();
 DECAPx1_ASAP7_75t_R FILLER_0_205_35 ();
 DECAPx1_ASAP7_75t_R FILLER_0_205_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_51 ();
 DECAPx1_ASAP7_75t_R FILLER_0_205_58 ();
 DECAPx2_ASAP7_75t_R FILLER_0_205_69 ();
 FILLER_ASAP7_75t_R FILLER_0_205_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_77 ();
 FILLER_ASAP7_75t_R FILLER_0_205_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_88 ();
 DECAPx4_ASAP7_75t_R FILLER_0_205_97 ();
 FILLER_ASAP7_75t_R FILLER_0_205_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_109 ();
 DECAPx10_ASAP7_75t_R FILLER_0_205_116 ();
 FILLER_ASAP7_75t_R FILLER_0_205_138 ();
 DECAPx6_ASAP7_75t_R FILLER_0_205_146 ();
 FILLER_ASAP7_75t_R FILLER_0_205_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_162 ();
 DECAPx4_ASAP7_75t_R FILLER_0_205_166 ();
 FILLER_ASAP7_75t_R FILLER_0_205_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_178 ();
 FILLER_ASAP7_75t_R FILLER_0_205_185 ();
 DECAPx4_ASAP7_75t_R FILLER_0_205_203 ();
 FILLER_ASAP7_75t_R FILLER_0_205_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_215 ();
 DECAPx4_ASAP7_75t_R FILLER_0_205_222 ();
 FILLER_ASAP7_75t_R FILLER_0_205_242 ();
 DECAPx1_ASAP7_75t_R FILLER_0_205_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_254 ();
 FILLER_ASAP7_75t_R FILLER_0_205_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_265 ();
 DECAPx1_ASAP7_75t_R FILLER_0_205_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_273 ();
 FILLER_ASAP7_75t_R FILLER_0_205_280 ();
 FILLER_ASAP7_75t_R FILLER_0_205_290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_205_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_305 ();
 FILLER_ASAP7_75t_R FILLER_0_205_312 ();
 DECAPx1_ASAP7_75t_R FILLER_0_205_317 ();
 FILLER_ASAP7_75t_R FILLER_0_205_341 ();
 DECAPx2_ASAP7_75t_R FILLER_0_205_349 ();
 FILLER_ASAP7_75t_R FILLER_0_205_355 ();
 DECAPx6_ASAP7_75t_R FILLER_0_205_363 ();
 DECAPx2_ASAP7_75t_R FILLER_0_205_377 ();
 FILLER_ASAP7_75t_R FILLER_0_205_389 ();
 DECAPx4_ASAP7_75t_R FILLER_0_205_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_407 ();
 DECAPx4_ASAP7_75t_R FILLER_0_205_416 ();
 FILLER_ASAP7_75t_R FILLER_0_205_426 ();
 FILLER_ASAP7_75t_R FILLER_0_205_434 ();
 FILLER_ASAP7_75t_R FILLER_0_205_442 ();
 DECAPx4_ASAP7_75t_R FILLER_0_205_451 ();
 FILLER_ASAP7_75t_R FILLER_0_205_461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_205_471 ();
 DECAPx4_ASAP7_75t_R FILLER_0_205_493 ();
 FILLER_ASAP7_75t_R FILLER_0_205_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_505 ();
 FILLER_ASAP7_75t_R FILLER_0_205_512 ();
 FILLER_ASAP7_75t_R FILLER_0_205_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_523 ();
 FILLER_ASAP7_75t_R FILLER_0_205_530 ();
 DECAPx4_ASAP7_75t_R FILLER_0_205_535 ();
 DECAPx6_ASAP7_75t_R FILLER_0_205_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_565 ();
 FILLER_ASAP7_75t_R FILLER_0_205_576 ();
 DECAPx4_ASAP7_75t_R FILLER_0_205_581 ();
 FILLER_ASAP7_75t_R FILLER_0_205_591 ();
 DECAPx4_ASAP7_75t_R FILLER_0_205_599 ();
 DECAPx2_ASAP7_75t_R FILLER_0_205_616 ();
 FILLER_ASAP7_75t_R FILLER_0_205_625 ();
 FILLER_ASAP7_75t_R FILLER_0_205_630 ();
 DECAPx1_ASAP7_75t_R FILLER_0_205_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_643 ();
 DECAPx4_ASAP7_75t_R FILLER_0_205_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_657 ();
 FILLER_ASAP7_75t_R FILLER_0_205_661 ();
 FILLER_ASAP7_75t_R FILLER_0_205_666 ();
 DECAPx1_ASAP7_75t_R FILLER_0_205_678 ();
 DECAPx6_ASAP7_75t_R FILLER_0_205_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_702 ();
 DECAPx2_ASAP7_75t_R FILLER_0_205_706 ();
 FILLER_ASAP7_75t_R FILLER_0_205_712 ();
 FILLER_ASAP7_75t_R FILLER_0_205_725 ();
 FILLER_ASAP7_75t_R FILLER_0_205_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_735 ();
 DECAPx1_ASAP7_75t_R FILLER_0_205_746 ();
 FILLER_ASAP7_75t_R FILLER_0_205_760 ();
 DECAPx10_ASAP7_75t_R FILLER_0_205_768 ();
 DECAPx4_ASAP7_75t_R FILLER_0_205_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_800 ();
 FILLER_ASAP7_75t_R FILLER_0_205_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_809 ();
 DECAPx6_ASAP7_75t_R FILLER_0_205_816 ();
 FILLER_ASAP7_75t_R FILLER_0_205_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_832 ();
 DECAPx4_ASAP7_75t_R FILLER_0_205_839 ();
 DECAPx2_ASAP7_75t_R FILLER_0_205_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_861 ();
 DECAPx1_ASAP7_75t_R FILLER_0_205_872 ();
 DECAPx4_ASAP7_75t_R FILLER_0_205_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_891 ();
 FILLER_ASAP7_75t_R FILLER_0_205_902 ();
 DECAPx6_ASAP7_75t_R FILLER_0_205_909 ();
 FILLER_ASAP7_75t_R FILLER_0_205_923 ();
 DECAPx10_ASAP7_75t_R FILLER_0_205_927 ();
 DECAPx6_ASAP7_75t_R FILLER_0_205_949 ();
 DECAPx1_ASAP7_75t_R FILLER_0_205_963 ();
 DECAPx2_ASAP7_75t_R FILLER_0_205_973 ();
 DECAPx10_ASAP7_75t_R FILLER_0_205_990 ();
 DECAPx2_ASAP7_75t_R FILLER_0_205_1012 ();
 FILLER_ASAP7_75t_R FILLER_0_205_1023 ();
 FILLER_ASAP7_75t_R FILLER_0_205_1043 ();
 FILLER_ASAP7_75t_R FILLER_0_205_1063 ();
 DECAPx2_ASAP7_75t_R FILLER_0_205_1071 ();
 FILLER_ASAP7_75t_R FILLER_0_205_1077 ();
 FILLER_ASAP7_75t_R FILLER_0_205_1085 ();
 FILLER_ASAP7_75t_R FILLER_0_205_1092 ();
 FILLER_ASAP7_75t_R FILLER_0_205_1104 ();
 FILLER_ASAP7_75t_R FILLER_0_205_1116 ();
 FILLER_ASAP7_75t_R FILLER_0_205_1128 ();
 FILLER_ASAP7_75t_R FILLER_0_205_1136 ();
 DECAPx1_ASAP7_75t_R FILLER_0_205_1144 ();
 FILLER_ASAP7_75t_R FILLER_0_205_1153 ();
 DECAPx1_ASAP7_75t_R FILLER_0_205_1161 ();
 FILLER_ASAP7_75t_R FILLER_0_205_1169 ();
 DECAPx1_ASAP7_75t_R FILLER_0_205_1182 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_205_1192 ();
 FILLER_ASAP7_75t_R FILLER_0_205_1216 ();
 DECAPx6_ASAP7_75t_R FILLER_0_205_1226 ();
 DECAPx1_ASAP7_75t_R FILLER_0_205_1240 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_1244 ();
 FILLER_ASAP7_75t_R FILLER_0_205_1251 ();
 DECAPx1_ASAP7_75t_R FILLER_0_205_1259 ();
 FILLER_ASAP7_75t_R FILLER_0_205_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_0_205_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_0_205_1301 ();
 DECAPx10_ASAP7_75t_R FILLER_0_205_1323 ();
 DECAPx10_ASAP7_75t_R FILLER_0_205_1345 ();
 DECAPx6_ASAP7_75t_R FILLER_0_205_1367 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_206_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_206_25 ();
 DECAPx1_ASAP7_75t_R FILLER_0_206_47 ();
 FILLER_ASAP7_75t_R FILLER_0_206_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_59 ();
 FILLER_ASAP7_75t_R FILLER_0_206_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_68 ();
 FILLER_ASAP7_75t_R FILLER_0_206_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_77 ();
 DECAPx1_ASAP7_75t_R FILLER_0_206_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_88 ();
 DECAPx4_ASAP7_75t_R FILLER_0_206_100 ();
 FILLER_ASAP7_75t_R FILLER_0_206_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_112 ();
 FILLER_ASAP7_75t_R FILLER_0_206_117 ();
 FILLER_ASAP7_75t_R FILLER_0_206_125 ();
 DECAPx2_ASAP7_75t_R FILLER_0_206_137 ();
 DECAPx4_ASAP7_75t_R FILLER_0_206_149 ();
 FILLER_ASAP7_75t_R FILLER_0_206_165 ();
 DECAPx2_ASAP7_75t_R FILLER_0_206_177 ();
 FILLER_ASAP7_75t_R FILLER_0_206_183 ();
 DECAPx2_ASAP7_75t_R FILLER_0_206_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_197 ();
 DECAPx10_ASAP7_75t_R FILLER_0_206_204 ();
 DECAPx4_ASAP7_75t_R FILLER_0_206_226 ();
 DECAPx1_ASAP7_75t_R FILLER_0_206_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_248 ();
 DECAPx4_ASAP7_75t_R FILLER_0_206_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_269 ();
 DECAPx1_ASAP7_75t_R FILLER_0_206_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_280 ();
 DECAPx2_ASAP7_75t_R FILLER_0_206_287 ();
 FILLER_ASAP7_75t_R FILLER_0_206_293 ();
 DECAPx2_ASAP7_75t_R FILLER_0_206_301 ();
 FILLER_ASAP7_75t_R FILLER_0_206_307 ();
 FILLER_ASAP7_75t_R FILLER_0_206_317 ();
 DECAPx2_ASAP7_75t_R FILLER_0_206_322 ();
 FILLER_ASAP7_75t_R FILLER_0_206_328 ();
 FILLER_ASAP7_75t_R FILLER_0_206_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_342 ();
 FILLER_ASAP7_75t_R FILLER_0_206_351 ();
 FILLER_ASAP7_75t_R FILLER_0_206_359 ();
 DECAPx2_ASAP7_75t_R FILLER_0_206_368 ();
 FILLER_ASAP7_75t_R FILLER_0_206_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_376 ();
 DECAPx4_ASAP7_75t_R FILLER_0_206_383 ();
 FILLER_ASAP7_75t_R FILLER_0_206_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_395 ();
 DECAPx2_ASAP7_75t_R FILLER_0_206_404 ();
 FILLER_ASAP7_75t_R FILLER_0_206_410 ();
 FILLER_ASAP7_75t_R FILLER_0_206_420 ();
 DECAPx2_ASAP7_75t_R FILLER_0_206_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_438 ();
 FILLER_ASAP7_75t_R FILLER_0_206_445 ();
 DECAPx2_ASAP7_75t_R FILLER_0_206_453 ();
 FILLER_ASAP7_75t_R FILLER_0_206_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_461 ();
 FILLER_ASAP7_75t_R FILLER_0_206_464 ();
 FILLER_ASAP7_75t_R FILLER_0_206_476 ();
 DECAPx6_ASAP7_75t_R FILLER_0_206_488 ();
 FILLER_ASAP7_75t_R FILLER_0_206_508 ();
 FILLER_ASAP7_75t_R FILLER_0_206_516 ();
 FILLER_ASAP7_75t_R FILLER_0_206_523 ();
 DECAPx10_ASAP7_75t_R FILLER_0_206_528 ();
 DECAPx6_ASAP7_75t_R FILLER_0_206_550 ();
 DECAPx1_ASAP7_75t_R FILLER_0_206_564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_206_571 ();
 DECAPx6_ASAP7_75t_R FILLER_0_206_593 ();
 DECAPx2_ASAP7_75t_R FILLER_0_206_607 ();
 DECAPx10_ASAP7_75t_R FILLER_0_206_620 ();
 DECAPx6_ASAP7_75t_R FILLER_0_206_642 ();
 DECAPx1_ASAP7_75t_R FILLER_0_206_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_660 ();
 DECAPx10_ASAP7_75t_R FILLER_0_206_667 ();
 DECAPx4_ASAP7_75t_R FILLER_0_206_689 ();
 FILLER_ASAP7_75t_R FILLER_0_206_699 ();
 FILLER_ASAP7_75t_R FILLER_0_206_707 ();
 DECAPx10_ASAP7_75t_R FILLER_0_206_712 ();
 DECAPx10_ASAP7_75t_R FILLER_0_206_734 ();
 DECAPx1_ASAP7_75t_R FILLER_0_206_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_760 ();
 DECAPx6_ASAP7_75t_R FILLER_0_206_771 ();
 DECAPx2_ASAP7_75t_R FILLER_0_206_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_797 ();
 FILLER_ASAP7_75t_R FILLER_0_206_808 ();
 FILLER_ASAP7_75t_R FILLER_0_206_820 ();
 FILLER_ASAP7_75t_R FILLER_0_206_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_829 ();
 DECAPx2_ASAP7_75t_R FILLER_0_206_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_846 ();
 FILLER_ASAP7_75t_R FILLER_0_206_853 ();
 DECAPx4_ASAP7_75t_R FILLER_0_206_861 ();
 FILLER_ASAP7_75t_R FILLER_0_206_877 ();
 FILLER_ASAP7_75t_R FILLER_0_206_886 ();
 FILLER_ASAP7_75t_R FILLER_0_206_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_895 ();
 FILLER_ASAP7_75t_R FILLER_0_206_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_905 ();
 FILLER_ASAP7_75t_R FILLER_0_206_916 ();
 FILLER_ASAP7_75t_R FILLER_0_206_923 ();
 FILLER_ASAP7_75t_R FILLER_0_206_931 ();
 DECAPx1_ASAP7_75t_R FILLER_0_206_939 ();
 DECAPx6_ASAP7_75t_R FILLER_0_206_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_967 ();
 FILLER_ASAP7_75t_R FILLER_0_206_979 ();
 DECAPx6_ASAP7_75t_R FILLER_0_206_987 ();
 DECAPx1_ASAP7_75t_R FILLER_0_206_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_1005 ();
 FILLER_ASAP7_75t_R FILLER_0_206_1027 ();
 FILLER_ASAP7_75t_R FILLER_0_206_1035 ();
 DECAPx2_ASAP7_75t_R FILLER_0_206_1047 ();
 FILLER_ASAP7_75t_R FILLER_0_206_1061 ();
 DECAPx1_ASAP7_75t_R FILLER_0_206_1068 ();
 FILLER_ASAP7_75t_R FILLER_0_206_1078 ();
 DECAPx1_ASAP7_75t_R FILLER_0_206_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_1090 ();
 FILLER_ASAP7_75t_R FILLER_0_206_1097 ();
 DECAPx2_ASAP7_75t_R FILLER_0_206_1109 ();
 FILLER_ASAP7_75t_R FILLER_0_206_1115 ();
 FILLER_ASAP7_75t_R FILLER_0_206_1124 ();
 FILLER_ASAP7_75t_R FILLER_0_206_1131 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_1133 ();
 FILLER_ASAP7_75t_R FILLER_0_206_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206_1142 ();
 DECAPx1_ASAP7_75t_R FILLER_0_206_1149 ();
 FILLER_ASAP7_75t_R FILLER_0_206_1163 ();
 FILLER_ASAP7_75t_R FILLER_0_206_1171 ();
 FILLER_ASAP7_75t_R FILLER_0_206_1181 ();
 DECAPx6_ASAP7_75t_R FILLER_0_206_1188 ();
 FILLER_ASAP7_75t_R FILLER_0_206_1202 ();
 DECAPx1_ASAP7_75t_R FILLER_0_206_1214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_206_1224 ();
 FILLER_ASAP7_75t_R FILLER_0_206_1252 ();
 FILLER_ASAP7_75t_R FILLER_0_206_1260 ();
 FILLER_ASAP7_75t_R FILLER_0_206_1274 ();
 DECAPx10_ASAP7_75t_R FILLER_0_206_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_206_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_206_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_206_1348 ();
 DECAPx4_ASAP7_75t_R FILLER_0_206_1370 ();
 FILLER_ASAP7_75t_R FILLER_0_206_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_207_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_4 ();
 FILLER_ASAP7_75t_R FILLER_0_207_8 ();
 FILLER_ASAP7_75t_R FILLER_0_207_15 ();
 DECAPx6_ASAP7_75t_R FILLER_0_207_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_36 ();
 FILLER_ASAP7_75t_R FILLER_0_207_47 ();
 DECAPx2_ASAP7_75t_R FILLER_0_207_57 ();
 FILLER_ASAP7_75t_R FILLER_0_207_63 ();
 DECAPx4_ASAP7_75t_R FILLER_0_207_71 ();
 FILLER_ASAP7_75t_R FILLER_0_207_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_83 ();
 FILLER_ASAP7_75t_R FILLER_0_207_90 ();
 DECAPx2_ASAP7_75t_R FILLER_0_207_98 ();
 FILLER_ASAP7_75t_R FILLER_0_207_104 ();
 DECAPx2_ASAP7_75t_R FILLER_0_207_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_117 ();
 FILLER_ASAP7_75t_R FILLER_0_207_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_126 ();
 DECAPx4_ASAP7_75t_R FILLER_0_207_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_143 ();
 DECAPx2_ASAP7_75t_R FILLER_0_207_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_156 ();
 DECAPx4_ASAP7_75t_R FILLER_0_207_169 ();
 FILLER_ASAP7_75t_R FILLER_0_207_179 ();
 FILLER_ASAP7_75t_R FILLER_0_207_187 ();
 DECAPx2_ASAP7_75t_R FILLER_0_207_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_199 ();
 DECAPx10_ASAP7_75t_R FILLER_0_207_210 ();
 DECAPx2_ASAP7_75t_R FILLER_0_207_232 ();
 DECAPx2_ASAP7_75t_R FILLER_0_207_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_251 ();
 FILLER_ASAP7_75t_R FILLER_0_207_255 ();
 DECAPx2_ASAP7_75t_R FILLER_0_207_263 ();
 DECAPx2_ASAP7_75t_R FILLER_0_207_275 ();
 FILLER_ASAP7_75t_R FILLER_0_207_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_283 ();
 DECAPx4_ASAP7_75t_R FILLER_0_207_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_314 ();
 DECAPx6_ASAP7_75t_R FILLER_0_207_321 ();
 DECAPx2_ASAP7_75t_R FILLER_0_207_335 ();
 DECAPx4_ASAP7_75t_R FILLER_0_207_347 ();
 FILLER_ASAP7_75t_R FILLER_0_207_357 ();
 DECAPx4_ASAP7_75t_R FILLER_0_207_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_375 ();
 FILLER_ASAP7_75t_R FILLER_0_207_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_384 ();
 FILLER_ASAP7_75t_R FILLER_0_207_388 ();
 DECAPx4_ASAP7_75t_R FILLER_0_207_393 ();
 FILLER_ASAP7_75t_R FILLER_0_207_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_405 ();
 FILLER_ASAP7_75t_R FILLER_0_207_412 ();
 DECAPx1_ASAP7_75t_R FILLER_0_207_420 ();
 DECAPx1_ASAP7_75t_R FILLER_0_207_427 ();
 DECAPx10_ASAP7_75t_R FILLER_0_207_437 ();
 FILLER_ASAP7_75t_R FILLER_0_207_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_461 ();
 DECAPx1_ASAP7_75t_R FILLER_0_207_470 ();
 DECAPx6_ASAP7_75t_R FILLER_0_207_495 ();
 FILLER_ASAP7_75t_R FILLER_0_207_516 ();
 DECAPx6_ASAP7_75t_R FILLER_0_207_521 ();
 DECAPx10_ASAP7_75t_R FILLER_0_207_541 ();
 FILLER_ASAP7_75t_R FILLER_0_207_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_565 ();
 FILLER_ASAP7_75t_R FILLER_0_207_572 ();
 DECAPx4_ASAP7_75t_R FILLER_0_207_595 ();
 DECAPx6_ASAP7_75t_R FILLER_0_207_617 ();
 DECAPx2_ASAP7_75t_R FILLER_0_207_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_637 ();
 DECAPx2_ASAP7_75t_R FILLER_0_207_644 ();
 FILLER_ASAP7_75t_R FILLER_0_207_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_652 ();
 FILLER_ASAP7_75t_R FILLER_0_207_659 ();
 DECAPx1_ASAP7_75t_R FILLER_0_207_667 ();
 FILLER_ASAP7_75t_R FILLER_0_207_677 ();
 DECAPx6_ASAP7_75t_R FILLER_0_207_685 ();
 DECAPx2_ASAP7_75t_R FILLER_0_207_699 ();
 DECAPx4_ASAP7_75t_R FILLER_0_207_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_721 ();
 DECAPx6_ASAP7_75t_R FILLER_0_207_730 ();
 DECAPx2_ASAP7_75t_R FILLER_0_207_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_750 ();
 FILLER_ASAP7_75t_R FILLER_0_207_755 ();
 DECAPx1_ASAP7_75t_R FILLER_0_207_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_769 ();
 FILLER_ASAP7_75t_R FILLER_0_207_780 ();
 DECAPx1_ASAP7_75t_R FILLER_0_207_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_795 ();
 DECAPx1_ASAP7_75t_R FILLER_0_207_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_810 ();
 FILLER_ASAP7_75t_R FILLER_0_207_831 ();
 FILLER_ASAP7_75t_R FILLER_0_207_841 ();
 FILLER_ASAP7_75t_R FILLER_0_207_850 ();
 DECAPx6_ASAP7_75t_R FILLER_0_207_859 ();
 DECAPx2_ASAP7_75t_R FILLER_0_207_880 ();
 FILLER_ASAP7_75t_R FILLER_0_207_886 ();
 FILLER_ASAP7_75t_R FILLER_0_207_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_902 ();
 FILLER_ASAP7_75t_R FILLER_0_207_908 ();
 DECAPx1_ASAP7_75t_R FILLER_0_207_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_924 ();
 DECAPx2_ASAP7_75t_R FILLER_0_207_927 ();
 DECAPx2_ASAP7_75t_R FILLER_0_207_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_945 ();
 FILLER_ASAP7_75t_R FILLER_0_207_950 ();
 DECAPx1_ASAP7_75t_R FILLER_0_207_964 ();
 FILLER_ASAP7_75t_R FILLER_0_207_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_976 ();
 DECAPx1_ASAP7_75t_R FILLER_0_207_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_987 ();
 DECAPx6_ASAP7_75t_R FILLER_0_207_994 ();
 DECAPx2_ASAP7_75t_R FILLER_0_207_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_1017 ();
 FILLER_ASAP7_75t_R FILLER_0_207_1024 ();
 FILLER_ASAP7_75t_R FILLER_0_207_1036 ();
 FILLER_ASAP7_75t_R FILLER_0_207_1044 ();
 FILLER_ASAP7_75t_R FILLER_0_207_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_1053 ();
 FILLER_ASAP7_75t_R FILLER_0_207_1064 ();
 FILLER_ASAP7_75t_R FILLER_0_207_1069 ();
 FILLER_ASAP7_75t_R FILLER_0_207_1077 ();
 FILLER_ASAP7_75t_R FILLER_0_207_1084 ();
 FILLER_ASAP7_75t_R FILLER_0_207_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_1093 ();
 DECAPx1_ASAP7_75t_R FILLER_0_207_1104 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_1108 ();
 FILLER_ASAP7_75t_R FILLER_0_207_1115 ();
 DECAPx1_ASAP7_75t_R FILLER_0_207_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_1127 ();
 DECAPx1_ASAP7_75t_R FILLER_0_207_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_1137 ();
 DECAPx2_ASAP7_75t_R FILLER_0_207_1143 ();
 FILLER_ASAP7_75t_R FILLER_0_207_1149 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_1151 ();
 DECAPx4_ASAP7_75t_R FILLER_0_207_1158 ();
 FILLER_ASAP7_75t_R FILLER_0_207_1168 ();
 DECAPx1_ASAP7_75t_R FILLER_0_207_1176 ();
 FILLER_ASAP7_75t_R FILLER_0_207_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_207_1193 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_1195 ();
 FILLER_ASAP7_75t_R FILLER_0_207_1202 ();
 DECAPx2_ASAP7_75t_R FILLER_0_207_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_1216 ();
 FILLER_ASAP7_75t_R FILLER_0_207_1222 ();
 DECAPx4_ASAP7_75t_R FILLER_0_207_1234 ();
 FILLER_ASAP7_75t_R FILLER_0_207_1244 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207_1246 ();
 FILLER_ASAP7_75t_R FILLER_0_207_1253 ();
 FILLER_ASAP7_75t_R FILLER_0_207_1260 ();
 DECAPx2_ASAP7_75t_R FILLER_0_207_1268 ();
 FILLER_ASAP7_75t_R FILLER_0_207_1274 ();
 DECAPx10_ASAP7_75t_R FILLER_0_207_1282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_207_1304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_207_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_207_1348 ();
 DECAPx4_ASAP7_75t_R FILLER_0_207_1370 ();
 FILLER_ASAP7_75t_R FILLER_0_207_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_208_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_208_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_19 ();
 FILLER_ASAP7_75t_R FILLER_0_208_26 ();
 DECAPx1_ASAP7_75t_R FILLER_0_208_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_38 ();
 FILLER_ASAP7_75t_R FILLER_0_208_45 ();
 FILLER_ASAP7_75t_R FILLER_0_208_50 ();
 DECAPx4_ASAP7_75t_R FILLER_0_208_60 ();
 FILLER_ASAP7_75t_R FILLER_0_208_70 ();
 FILLER_ASAP7_75t_R FILLER_0_208_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_80 ();
 DECAPx1_ASAP7_75t_R FILLER_0_208_84 ();
 DECAPx4_ASAP7_75t_R FILLER_0_208_91 ();
 FILLER_ASAP7_75t_R FILLER_0_208_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_103 ();
 FILLER_ASAP7_75t_R FILLER_0_208_109 ();
 FILLER_ASAP7_75t_R FILLER_0_208_123 ();
 DECAPx4_ASAP7_75t_R FILLER_0_208_130 ();
 FILLER_ASAP7_75t_R FILLER_0_208_148 ();
 DECAPx1_ASAP7_75t_R FILLER_0_208_156 ();
 FILLER_ASAP7_75t_R FILLER_0_208_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_168 ();
 FILLER_ASAP7_75t_R FILLER_0_208_177 ();
 DECAPx1_ASAP7_75t_R FILLER_0_208_186 ();
 FILLER_ASAP7_75t_R FILLER_0_208_195 ();
 FILLER_ASAP7_75t_R FILLER_0_208_203 ();
 DECAPx6_ASAP7_75t_R FILLER_0_208_211 ();
 FILLER_ASAP7_75t_R FILLER_0_208_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_227 ();
 FILLER_ASAP7_75t_R FILLER_0_208_238 ();
 FILLER_ASAP7_75t_R FILLER_0_208_248 ();
 DECAPx1_ASAP7_75t_R FILLER_0_208_253 ();
 DECAPx2_ASAP7_75t_R FILLER_0_208_263 ();
 FILLER_ASAP7_75t_R FILLER_0_208_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_277 ();
 FILLER_ASAP7_75t_R FILLER_0_208_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_286 ();
 DECAPx10_ASAP7_75t_R FILLER_0_208_295 ();
 DECAPx2_ASAP7_75t_R FILLER_0_208_317 ();
 FILLER_ASAP7_75t_R FILLER_0_208_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_325 ();
 DECAPx6_ASAP7_75t_R FILLER_0_208_336 ();
 DECAPx4_ASAP7_75t_R FILLER_0_208_356 ();
 DECAPx2_ASAP7_75t_R FILLER_0_208_372 ();
 FILLER_ASAP7_75t_R FILLER_0_208_378 ();
 FILLER_ASAP7_75t_R FILLER_0_208_386 ();
 DECAPx4_ASAP7_75t_R FILLER_0_208_396 ();
 FILLER_ASAP7_75t_R FILLER_0_208_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_408 ();
 DECAPx10_ASAP7_75t_R FILLER_0_208_415 ();
 DECAPx10_ASAP7_75t_R FILLER_0_208_437 ();
 FILLER_ASAP7_75t_R FILLER_0_208_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_461 ();
 DECAPx1_ASAP7_75t_R FILLER_0_208_464 ();
 FILLER_ASAP7_75t_R FILLER_0_208_476 ();
 DECAPx2_ASAP7_75t_R FILLER_0_208_481 ();
 FILLER_ASAP7_75t_R FILLER_0_208_498 ();
 FILLER_ASAP7_75t_R FILLER_0_208_522 ();
 FILLER_ASAP7_75t_R FILLER_0_208_536 ();
 FILLER_ASAP7_75t_R FILLER_0_208_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_550 ();
 DECAPx2_ASAP7_75t_R FILLER_0_208_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_567 ();
 FILLER_ASAP7_75t_R FILLER_0_208_574 ();
 DECAPx1_ASAP7_75t_R FILLER_0_208_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_592 ();
 DECAPx6_ASAP7_75t_R FILLER_0_208_596 ();
 DECAPx1_ASAP7_75t_R FILLER_0_208_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_614 ();
 FILLER_ASAP7_75t_R FILLER_0_208_637 ();
 DECAPx1_ASAP7_75t_R FILLER_0_208_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_664 ();
 DECAPx1_ASAP7_75t_R FILLER_0_208_668 ();
 FILLER_ASAP7_75t_R FILLER_0_208_678 ();
 DECAPx4_ASAP7_75t_R FILLER_0_208_688 ();
 FILLER_ASAP7_75t_R FILLER_0_208_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_700 ();
 FILLER_ASAP7_75t_R FILLER_0_208_707 ();
 FILLER_ASAP7_75t_R FILLER_0_208_719 ();
 FILLER_ASAP7_75t_R FILLER_0_208_733 ();
 DECAPx2_ASAP7_75t_R FILLER_0_208_741 ();
 FILLER_ASAP7_75t_R FILLER_0_208_747 ();
 DECAPx2_ASAP7_75t_R FILLER_0_208_757 ();
 FILLER_ASAP7_75t_R FILLER_0_208_763 ();
 DECAPx2_ASAP7_75t_R FILLER_0_208_771 ();
 FILLER_ASAP7_75t_R FILLER_0_208_777 ();
 FILLER_ASAP7_75t_R FILLER_0_208_785 ();
 DECAPx2_ASAP7_75t_R FILLER_0_208_793 ();
 FILLER_ASAP7_75t_R FILLER_0_208_809 ();
 DECAPx2_ASAP7_75t_R FILLER_0_208_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_827 ();
 FILLER_ASAP7_75t_R FILLER_0_208_838 ();
 FILLER_ASAP7_75t_R FILLER_0_208_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_847 ();
 FILLER_ASAP7_75t_R FILLER_0_208_856 ();
 DECAPx2_ASAP7_75t_R FILLER_0_208_865 ();
 FILLER_ASAP7_75t_R FILLER_0_208_871 ();
 DECAPx2_ASAP7_75t_R FILLER_0_208_880 ();
 DECAPx4_ASAP7_75t_R FILLER_0_208_898 ();
 FILLER_ASAP7_75t_R FILLER_0_208_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_910 ();
 DECAPx4_ASAP7_75t_R FILLER_0_208_915 ();
 FILLER_ASAP7_75t_R FILLER_0_208_925 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_927 ();
 FILLER_ASAP7_75t_R FILLER_0_208_934 ();
 FILLER_ASAP7_75t_R FILLER_0_208_942 ();
 DECAPx4_ASAP7_75t_R FILLER_0_208_954 ();
 DECAPx2_ASAP7_75t_R FILLER_0_208_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_976 ();
 FILLER_ASAP7_75t_R FILLER_0_208_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_985 ();
 DECAPx10_ASAP7_75t_R FILLER_0_208_992 ();
 FILLER_ASAP7_75t_R FILLER_0_208_1014 ();
 DECAPx2_ASAP7_75t_R FILLER_0_208_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_1032 ();
 FILLER_ASAP7_75t_R FILLER_0_208_1043 ();
 DECAPx2_ASAP7_75t_R FILLER_0_208_1056 ();
 FILLER_ASAP7_75t_R FILLER_0_208_1062 ();
 FILLER_ASAP7_75t_R FILLER_0_208_1070 ();
 DECAPx1_ASAP7_75t_R FILLER_0_208_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_1081 ();
 FILLER_ASAP7_75t_R FILLER_0_208_1110 ();
 DECAPx2_ASAP7_75t_R FILLER_0_208_1117 ();
 FILLER_ASAP7_75t_R FILLER_0_208_1133 ();
 FILLER_ASAP7_75t_R FILLER_0_208_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_1140 ();
 FILLER_ASAP7_75t_R FILLER_0_208_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_1149 ();
 FILLER_ASAP7_75t_R FILLER_0_208_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_1162 ();
 FILLER_ASAP7_75t_R FILLER_0_208_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_1171 ();
 FILLER_ASAP7_75t_R FILLER_0_208_1178 ();
 DECAPx2_ASAP7_75t_R FILLER_0_208_1191 ();
 DECAPx4_ASAP7_75t_R FILLER_0_208_1205 ();
 FILLER_ASAP7_75t_R FILLER_0_208_1221 ();
 DECAPx6_ASAP7_75t_R FILLER_0_208_1228 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_1242 ();
 FILLER_ASAP7_75t_R FILLER_0_208_1248 ();
 FILLER_ASAP7_75t_R FILLER_0_208_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_0_208_1269 ();
 DECAPx10_ASAP7_75t_R FILLER_0_208_1291 ();
 DECAPx10_ASAP7_75t_R FILLER_0_208_1313 ();
 DECAPx10_ASAP7_75t_R FILLER_0_208_1335 ();
 DECAPx10_ASAP7_75t_R FILLER_0_208_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_208_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_209_2 ();
 FILLER_ASAP7_75t_R FILLER_0_209_22 ();
 FILLER_ASAP7_75t_R FILLER_0_209_35 ();
 DECAPx1_ASAP7_75t_R FILLER_0_209_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_44 ();
 DECAPx10_ASAP7_75t_R FILLER_0_209_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_73 ();
 FILLER_ASAP7_75t_R FILLER_0_209_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_82 ();
 DECAPx2_ASAP7_75t_R FILLER_0_209_88 ();
 FILLER_ASAP7_75t_R FILLER_0_209_99 ();
 FILLER_ASAP7_75t_R FILLER_0_209_111 ();
 FILLER_ASAP7_75t_R FILLER_0_209_123 ();
 FILLER_ASAP7_75t_R FILLER_0_209_131 ();
 FILLER_ASAP7_75t_R FILLER_0_209_138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_209_147 ();
 DECAPx4_ASAP7_75t_R FILLER_0_209_169 ();
 FILLER_ASAP7_75t_R FILLER_0_209_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_181 ();
 FILLER_ASAP7_75t_R FILLER_0_209_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_189 ();
 DECAPx2_ASAP7_75t_R FILLER_0_209_196 ();
 FILLER_ASAP7_75t_R FILLER_0_209_202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_209_210 ();
 DECAPx2_ASAP7_75t_R FILLER_0_209_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_238 ();
 FILLER_ASAP7_75t_R FILLER_0_209_245 ();
 FILLER_ASAP7_75t_R FILLER_0_209_255 ();
 DECAPx2_ASAP7_75t_R FILLER_0_209_263 ();
 DECAPx1_ASAP7_75t_R FILLER_0_209_275 ();
 FILLER_ASAP7_75t_R FILLER_0_209_286 ();
 DECAPx1_ASAP7_75t_R FILLER_0_209_294 ();
 DECAPx1_ASAP7_75t_R FILLER_0_209_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_310 ();
 DECAPx2_ASAP7_75t_R FILLER_0_209_319 ();
 FILLER_ASAP7_75t_R FILLER_0_209_325 ();
 FILLER_ASAP7_75t_R FILLER_0_209_339 ();
 DECAPx6_ASAP7_75t_R FILLER_0_209_348 ();
 FILLER_ASAP7_75t_R FILLER_0_209_368 ();
 FILLER_ASAP7_75t_R FILLER_0_209_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_383 ();
 FILLER_ASAP7_75t_R FILLER_0_209_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_392 ();
 DECAPx2_ASAP7_75t_R FILLER_0_209_399 ();
 FILLER_ASAP7_75t_R FILLER_0_209_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_407 ();
 FILLER_ASAP7_75t_R FILLER_0_209_414 ();
 FILLER_ASAP7_75t_R FILLER_0_209_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_209_431 ();
 DECAPx6_ASAP7_75t_R FILLER_0_209_453 ();
 FILLER_ASAP7_75t_R FILLER_0_209_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_469 ();
 FILLER_ASAP7_75t_R FILLER_0_209_476 ();
 DECAPx4_ASAP7_75t_R FILLER_0_209_481 ();
 DECAPx2_ASAP7_75t_R FILLER_0_209_503 ();
 FILLER_ASAP7_75t_R FILLER_0_209_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_511 ();
 FILLER_ASAP7_75t_R FILLER_0_209_533 ();
 DECAPx1_ASAP7_75t_R FILLER_0_209_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_551 ();
 FILLER_ASAP7_75t_R FILLER_0_209_558 ();
 DECAPx1_ASAP7_75t_R FILLER_0_209_563 ();
 DECAPx2_ASAP7_75t_R FILLER_0_209_575 ();
 DECAPx10_ASAP7_75t_R FILLER_0_209_586 ();
 DECAPx2_ASAP7_75t_R FILLER_0_209_608 ();
 DECAPx1_ASAP7_75t_R FILLER_0_209_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_640 ();
 DECAPx6_ASAP7_75t_R FILLER_0_209_644 ();
 DECAPx1_ASAP7_75t_R FILLER_0_209_658 ();
 DECAPx2_ASAP7_75t_R FILLER_0_209_668 ();
 FILLER_ASAP7_75t_R FILLER_0_209_680 ();
 DECAPx10_ASAP7_75t_R FILLER_0_209_690 ();
 DECAPx4_ASAP7_75t_R FILLER_0_209_712 ();
 FILLER_ASAP7_75t_R FILLER_0_209_722 ();
 DECAPx6_ASAP7_75t_R FILLER_0_209_730 ();
 DECAPx1_ASAP7_75t_R FILLER_0_209_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_748 ();
 DECAPx2_ASAP7_75t_R FILLER_0_209_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_763 ();
 DECAPx1_ASAP7_75t_R FILLER_0_209_772 ();
 DECAPx1_ASAP7_75t_R FILLER_0_209_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_786 ();
 FILLER_ASAP7_75t_R FILLER_0_209_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_797 ();
 FILLER_ASAP7_75t_R FILLER_0_209_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_810 ();
 FILLER_ASAP7_75t_R FILLER_0_209_821 ();
 FILLER_ASAP7_75t_R FILLER_0_209_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_828 ();
 DECAPx1_ASAP7_75t_R FILLER_0_209_839 ();
 FILLER_ASAP7_75t_R FILLER_0_209_849 ();
 DECAPx4_ASAP7_75t_R FILLER_0_209_857 ();
 FILLER_ASAP7_75t_R FILLER_0_209_867 ();
 FILLER_ASAP7_75t_R FILLER_0_209_875 ();
 FILLER_ASAP7_75t_R FILLER_0_209_883 ();
 DECAPx6_ASAP7_75t_R FILLER_0_209_891 ();
 DECAPx1_ASAP7_75t_R FILLER_0_209_905 ();
 DECAPx2_ASAP7_75t_R FILLER_0_209_916 ();
 FILLER_ASAP7_75t_R FILLER_0_209_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_924 ();
 FILLER_ASAP7_75t_R FILLER_0_209_927 ();
 DECAPx1_ASAP7_75t_R FILLER_0_209_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_940 ();
 FILLER_ASAP7_75t_R FILLER_0_209_951 ();
 FILLER_ASAP7_75t_R FILLER_0_209_959 ();
 FILLER_ASAP7_75t_R FILLER_0_209_964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_209_972 ();
 FILLER_ASAP7_75t_R FILLER_0_209_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_988 ();
 FILLER_ASAP7_75t_R FILLER_0_209_1010 ();
 FILLER_ASAP7_75t_R FILLER_0_209_1016 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_1018 ();
 FILLER_ASAP7_75t_R FILLER_0_209_1029 ();
 FILLER_ASAP7_75t_R FILLER_0_209_1041 ();
 FILLER_ASAP7_75t_R FILLER_0_209_1049 ();
 DECAPx1_ASAP7_75t_R FILLER_0_209_1057 ();
 FILLER_ASAP7_75t_R FILLER_0_209_1067 ();
 DECAPx1_ASAP7_75t_R FILLER_0_209_1077 ();
 DECAPx2_ASAP7_75t_R FILLER_0_209_1091 ();
 FILLER_ASAP7_75t_R FILLER_0_209_1097 ();
 DECAPx1_ASAP7_75t_R FILLER_0_209_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_1113 ();
 DECAPx2_ASAP7_75t_R FILLER_0_209_1120 ();
 FILLER_ASAP7_75t_R FILLER_0_209_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_1128 ();
 DECAPx2_ASAP7_75t_R FILLER_0_209_1135 ();
 FILLER_ASAP7_75t_R FILLER_0_209_1141 ();
 FILLER_ASAP7_75t_R FILLER_0_209_1149 ();
 FILLER_ASAP7_75t_R FILLER_0_209_1157 ();
 DECAPx1_ASAP7_75t_R FILLER_0_209_1164 ();
 DECAPx6_ASAP7_75t_R FILLER_0_209_1174 ();
 FILLER_ASAP7_75t_R FILLER_0_209_1188 ();
 FILLER_ASAP7_75t_R FILLER_0_209_1195 ();
 DECAPx1_ASAP7_75t_R FILLER_0_209_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_1211 ();
 DECAPx2_ASAP7_75t_R FILLER_0_209_1218 ();
 FILLER_ASAP7_75t_R FILLER_0_209_1224 ();
 FILLER_ASAP7_75t_R FILLER_0_209_1233 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_1235 ();
 DECAPx1_ASAP7_75t_R FILLER_0_209_1242 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_1246 ();
 FILLER_ASAP7_75t_R FILLER_0_209_1253 ();
 FILLER_ASAP7_75t_R FILLER_0_209_1260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_209_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_0_209_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_0_209_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_0_209_1333 ();
 DECAPx10_ASAP7_75t_R FILLER_0_209_1355 ();
 DECAPx1_ASAP7_75t_R FILLER_0_209_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_210_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_210_9 ();
 DECAPx2_ASAP7_75t_R FILLER_0_210_29 ();
 FILLER_ASAP7_75t_R FILLER_0_210_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210_44 ();
 DECAPx2_ASAP7_75t_R FILLER_0_210_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210_63 ();
 FILLER_ASAP7_75t_R FILLER_0_210_69 ();
 FILLER_ASAP7_75t_R FILLER_0_210_77 ();
 DECAPx2_ASAP7_75t_R FILLER_0_210_84 ();
 DECAPx1_ASAP7_75t_R FILLER_0_210_96 ();
 FILLER_ASAP7_75t_R FILLER_0_210_110 ();
 FILLER_ASAP7_75t_R FILLER_0_210_122 ();
 DECAPx1_ASAP7_75t_R FILLER_0_210_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210_134 ();
 FILLER_ASAP7_75t_R FILLER_0_210_141 ();
 DECAPx6_ASAP7_75t_R FILLER_0_210_148 ();
 DECAPx4_ASAP7_75t_R FILLER_0_210_170 ();
 FILLER_ASAP7_75t_R FILLER_0_210_180 ();
 FILLER_ASAP7_75t_R FILLER_0_210_188 ();
 FILLER_ASAP7_75t_R FILLER_0_210_195 ();
 DECAPx10_ASAP7_75t_R FILLER_0_210_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210_224 ();
 FILLER_ASAP7_75t_R FILLER_0_210_235 ();
 DECAPx10_ASAP7_75t_R FILLER_0_210_244 ();
 DECAPx6_ASAP7_75t_R FILLER_0_210_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210_280 ();
 DECAPx1_ASAP7_75t_R FILLER_0_210_287 ();
 DECAPx1_ASAP7_75t_R FILLER_0_210_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210_301 ();
 DECAPx1_ASAP7_75t_R FILLER_0_210_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210_313 ();
 DECAPx1_ASAP7_75t_R FILLER_0_210_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210_321 ();
 FILLER_ASAP7_75t_R FILLER_0_210_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210_334 ();
 DECAPx1_ASAP7_75t_R FILLER_0_210_341 ();
 DECAPx1_ASAP7_75t_R FILLER_0_210_353 ();
 DECAPx6_ASAP7_75t_R FILLER_0_210_367 ();
 DECAPx2_ASAP7_75t_R FILLER_0_210_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210_387 ();
 DECAPx2_ASAP7_75t_R FILLER_0_210_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210_397 ();
 DECAPx1_ASAP7_75t_R FILLER_0_210_401 ();
 FILLER_ASAP7_75t_R FILLER_0_210_411 ();
 FILLER_ASAP7_75t_R FILLER_0_210_419 ();
 DECAPx2_ASAP7_75t_R FILLER_0_210_427 ();
 FILLER_ASAP7_75t_R FILLER_0_210_433 ();
 FILLER_ASAP7_75t_R FILLER_0_210_438 ();
 DECAPx6_ASAP7_75t_R FILLER_0_210_446 ();
 FILLER_ASAP7_75t_R FILLER_0_210_460 ();
 FILLER_ASAP7_75t_R FILLER_0_210_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210_466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_210_479 ();
 DECAPx4_ASAP7_75t_R FILLER_0_210_501 ();
 FILLER_ASAP7_75t_R FILLER_0_210_514 ();
 FILLER_ASAP7_75t_R FILLER_0_210_522 ();
 FILLER_ASAP7_75t_R FILLER_0_210_534 ();
 DECAPx2_ASAP7_75t_R FILLER_0_210_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210_554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_210_562 ();
 DECAPx6_ASAP7_75t_R FILLER_0_210_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210_598 ();
 DECAPx2_ASAP7_75t_R FILLER_0_210_611 ();
 FILLER_ASAP7_75t_R FILLER_0_210_625 ();
 DECAPx1_ASAP7_75t_R FILLER_0_210_630 ();
 DECAPx6_ASAP7_75t_R FILLER_0_210_646 ();
 FILLER_ASAP7_75t_R FILLER_0_210_660 ();
 FILLER_ASAP7_75t_R FILLER_0_210_670 ();
 DECAPx10_ASAP7_75t_R FILLER_0_210_678 ();
 FILLER_ASAP7_75t_R FILLER_0_210_700 ();
 FILLER_ASAP7_75t_R FILLER_0_210_708 ();
 DECAPx2_ASAP7_75t_R FILLER_0_210_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210_726 ();
 FILLER_ASAP7_75t_R FILLER_0_210_733 ();
 FILLER_ASAP7_75t_R FILLER_0_210_740 ();
 FILLER_ASAP7_75t_R FILLER_0_210_749 ();
 DECAPx1_ASAP7_75t_R FILLER_0_210_761 ();
 FILLER_ASAP7_75t_R FILLER_0_210_771 ();
 DECAPx1_ASAP7_75t_R FILLER_0_210_783 ();
 DECAPx1_ASAP7_75t_R FILLER_0_210_793 ();
 FILLER_ASAP7_75t_R FILLER_0_210_800 ();
 FILLER_ASAP7_75t_R FILLER_0_210_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210_814 ();
 DECAPx2_ASAP7_75t_R FILLER_0_210_835 ();
 DECAPx6_ASAP7_75t_R FILLER_0_210_851 ();
 DECAPx1_ASAP7_75t_R FILLER_0_210_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210_869 ();
 FILLER_ASAP7_75t_R FILLER_0_210_882 ();
 DECAPx4_ASAP7_75t_R FILLER_0_210_894 ();
 DECAPx1_ASAP7_75t_R FILLER_0_210_909 ();
 DECAPx6_ASAP7_75t_R FILLER_0_210_918 ();
 DECAPx2_ASAP7_75t_R FILLER_0_210_938 ();
 FILLER_ASAP7_75t_R FILLER_0_210_944 ();
 DECAPx10_ASAP7_75t_R FILLER_0_210_952 ();
 DECAPx6_ASAP7_75t_R FILLER_0_210_974 ();
 DECAPx1_ASAP7_75t_R FILLER_0_210_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210_992 ();
 FILLER_ASAP7_75t_R FILLER_0_210_998 ();
 DECAPx4_ASAP7_75t_R FILLER_0_210_1003 ();
 FILLER_ASAP7_75t_R FILLER_0_210_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210_1015 ();
 FILLER_ASAP7_75t_R FILLER_0_210_1026 ();
 FILLER_ASAP7_75t_R FILLER_0_210_1056 ();
 FILLER_ASAP7_75t_R FILLER_0_210_1064 ();
 FILLER_ASAP7_75t_R FILLER_0_210_1072 ();
 FILLER_ASAP7_75t_R FILLER_0_210_1080 ();
 DECAPx1_ASAP7_75t_R FILLER_0_210_1088 ();
 DECAPx1_ASAP7_75t_R FILLER_0_210_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210_1104 ();
 FILLER_ASAP7_75t_R FILLER_0_210_1111 ();
 FILLER_ASAP7_75t_R FILLER_0_210_1123 ();
 DECAPx6_ASAP7_75t_R FILLER_0_210_1131 ();
 DECAPx2_ASAP7_75t_R FILLER_0_210_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210_1151 ();
 DECAPx2_ASAP7_75t_R FILLER_0_210_1160 ();
 DECAPx2_ASAP7_75t_R FILLER_0_210_1176 ();
 FILLER_ASAP7_75t_R FILLER_0_210_1192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_210_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210_1218 ();
 FILLER_ASAP7_75t_R FILLER_0_210_1225 ();
 FILLER_ASAP7_75t_R FILLER_0_210_1233 ();
 FILLER_ASAP7_75t_R FILLER_0_210_1241 ();
 FILLER_ASAP7_75t_R FILLER_0_210_1253 ();
 FILLER_ASAP7_75t_R FILLER_0_210_1260 ();
 DECAPx2_ASAP7_75t_R FILLER_0_210_1265 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210_1271 ();
 DECAPx10_ASAP7_75t_R FILLER_0_210_1282 ();
 DECAPx1_ASAP7_75t_R FILLER_0_210_1326 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210_1330 ();
 DECAPx10_ASAP7_75t_R FILLER_0_210_1334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_210_1356 ();
 DECAPx1_ASAP7_75t_R FILLER_0_210_1378 ();
 DECAPx6_ASAP7_75t_R FILLER_0_211_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_16 ();
 DECAPx1_ASAP7_75t_R FILLER_0_211_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_26 ();
 FILLER_ASAP7_75t_R FILLER_0_211_32 ();
 DECAPx1_ASAP7_75t_R FILLER_0_211_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_44 ();
 DECAPx2_ASAP7_75t_R FILLER_0_211_52 ();
 DECAPx2_ASAP7_75t_R FILLER_0_211_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_70 ();
 FILLER_ASAP7_75t_R FILLER_0_211_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_85 ();
 FILLER_ASAP7_75t_R FILLER_0_211_91 ();
 FILLER_ASAP7_75t_R FILLER_0_211_100 ();
 FILLER_ASAP7_75t_R FILLER_0_211_112 ();
 DECAPx2_ASAP7_75t_R FILLER_0_211_124 ();
 FILLER_ASAP7_75t_R FILLER_0_211_130 ();
 FILLER_ASAP7_75t_R FILLER_0_211_138 ();
 DECAPx4_ASAP7_75t_R FILLER_0_211_146 ();
 FILLER_ASAP7_75t_R FILLER_0_211_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_158 ();
 DECAPx1_ASAP7_75t_R FILLER_0_211_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_175 ();
 FILLER_ASAP7_75t_R FILLER_0_211_182 ();
 DECAPx2_ASAP7_75t_R FILLER_0_211_190 ();
 FILLER_ASAP7_75t_R FILLER_0_211_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_198 ();
 DECAPx6_ASAP7_75t_R FILLER_0_211_211 ();
 FILLER_ASAP7_75t_R FILLER_0_211_225 ();
 FILLER_ASAP7_75t_R FILLER_0_211_242 ();
 DECAPx1_ASAP7_75t_R FILLER_0_211_247 ();
 DECAPx2_ASAP7_75t_R FILLER_0_211_257 ();
 FILLER_ASAP7_75t_R FILLER_0_211_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_265 ();
 DECAPx10_ASAP7_75t_R FILLER_0_211_272 ();
 DECAPx2_ASAP7_75t_R FILLER_0_211_297 ();
 DECAPx6_ASAP7_75t_R FILLER_0_211_309 ();
 DECAPx1_ASAP7_75t_R FILLER_0_211_323 ();
 FILLER_ASAP7_75t_R FILLER_0_211_337 ();
 FILLER_ASAP7_75t_R FILLER_0_211_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_347 ();
 DECAPx2_ASAP7_75t_R FILLER_0_211_354 ();
 DECAPx1_ASAP7_75t_R FILLER_0_211_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_370 ();
 FILLER_ASAP7_75t_R FILLER_0_211_377 ();
 DECAPx6_ASAP7_75t_R FILLER_0_211_385 ();
 DECAPx2_ASAP7_75t_R FILLER_0_211_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_405 ();
 FILLER_ASAP7_75t_R FILLER_0_211_414 ();
 DECAPx1_ASAP7_75t_R FILLER_0_211_422 ();
 DECAPx1_ASAP7_75t_R FILLER_0_211_432 ();
 DECAPx6_ASAP7_75t_R FILLER_0_211_444 ();
 DECAPx4_ASAP7_75t_R FILLER_0_211_470 ();
 FILLER_ASAP7_75t_R FILLER_0_211_480 ();
 FILLER_ASAP7_75t_R FILLER_0_211_494 ();
 DECAPx6_ASAP7_75t_R FILLER_0_211_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_531 ();
 DECAPx2_ASAP7_75t_R FILLER_0_211_544 ();
 FILLER_ASAP7_75t_R FILLER_0_211_550 ();
 DECAPx2_ASAP7_75t_R FILLER_0_211_559 ();
 FILLER_ASAP7_75t_R FILLER_0_211_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_567 ();
 FILLER_ASAP7_75t_R FILLER_0_211_588 ();
 DECAPx2_ASAP7_75t_R FILLER_0_211_611 ();
 FILLER_ASAP7_75t_R FILLER_0_211_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_619 ();
 FILLER_ASAP7_75t_R FILLER_0_211_628 ();
 DECAPx1_ASAP7_75t_R FILLER_0_211_636 ();
 DECAPx4_ASAP7_75t_R FILLER_0_211_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_662 ();
 FILLER_ASAP7_75t_R FILLER_0_211_671 ();
 DECAPx2_ASAP7_75t_R FILLER_0_211_676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_211_688 ();
 FILLER_ASAP7_75t_R FILLER_0_211_694 ();
 FILLER_ASAP7_75t_R FILLER_0_211_699 ();
 DECAPx10_ASAP7_75t_R FILLER_0_211_707 ();
 DECAPx6_ASAP7_75t_R FILLER_0_211_729 ();
 FILLER_ASAP7_75t_R FILLER_0_211_743 ();
 FILLER_ASAP7_75t_R FILLER_0_211_751 ();
 DECAPx2_ASAP7_75t_R FILLER_0_211_759 ();
 FILLER_ASAP7_75t_R FILLER_0_211_771 ();
 DECAPx1_ASAP7_75t_R FILLER_0_211_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_787 ();
 FILLER_ASAP7_75t_R FILLER_0_211_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_795 ();
 FILLER_ASAP7_75t_R FILLER_0_211_801 ();
 FILLER_ASAP7_75t_R FILLER_0_211_808 ();
 FILLER_ASAP7_75t_R FILLER_0_211_815 ();
 FILLER_ASAP7_75t_R FILLER_0_211_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_826 ();
 DECAPx4_ASAP7_75t_R FILLER_0_211_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_857 ();
 FILLER_ASAP7_75t_R FILLER_0_211_865 ();
 DECAPx1_ASAP7_75t_R FILLER_0_211_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_883 ();
 DECAPx1_ASAP7_75t_R FILLER_0_211_896 ();
 FILLER_ASAP7_75t_R FILLER_0_211_910 ();
 DECAPx2_ASAP7_75t_R FILLER_0_211_919 ();
 DECAPx2_ASAP7_75t_R FILLER_0_211_927 ();
 FILLER_ASAP7_75t_R FILLER_0_211_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_935 ();
 DECAPx1_ASAP7_75t_R FILLER_0_211_942 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_946 ();
 FILLER_ASAP7_75t_R FILLER_0_211_958 ();
 DECAPx2_ASAP7_75t_R FILLER_0_211_966 ();
 FILLER_ASAP7_75t_R FILLER_0_211_978 ();
 DECAPx2_ASAP7_75t_R FILLER_0_211_986 ();
 DECAPx6_ASAP7_75t_R FILLER_0_211_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_1018 ();
 FILLER_ASAP7_75t_R FILLER_0_211_1024 ();
 FILLER_ASAP7_75t_R FILLER_0_211_1054 ();
 FILLER_ASAP7_75t_R FILLER_0_211_1064 ();
 DECAPx2_ASAP7_75t_R FILLER_0_211_1071 ();
 DECAPx1_ASAP7_75t_R FILLER_0_211_1084 ();
 FILLER_ASAP7_75t_R FILLER_0_211_1100 ();
 FILLER_ASAP7_75t_R FILLER_0_211_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_1112 ();
 DECAPx2_ASAP7_75t_R FILLER_0_211_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_0_211_1137 ();
 DECAPx2_ASAP7_75t_R FILLER_0_211_1159 ();
 DECAPx6_ASAP7_75t_R FILLER_0_211_1171 ();
 FILLER_ASAP7_75t_R FILLER_0_211_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_211_1198 ();
 DECAPx4_ASAP7_75t_R FILLER_0_211_1220 ();
 FILLER_ASAP7_75t_R FILLER_0_211_1230 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_1232 ();
 DECAPx2_ASAP7_75t_R FILLER_0_211_1241 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_1247 ();
 FILLER_ASAP7_75t_R FILLER_0_211_1260 ();
 FILLER_ASAP7_75t_R FILLER_0_211_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_211_1277 ();
 DECAPx2_ASAP7_75t_R FILLER_0_211_1299 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_1305 ();
 DECAPx10_ASAP7_75t_R FILLER_0_211_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_0_211_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_0_211_1353 ();
 DECAPx2_ASAP7_75t_R FILLER_0_211_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211_1381 ();
 DECAPx6_ASAP7_75t_R FILLER_0_212_2 ();
 FILLER_ASAP7_75t_R FILLER_0_212_22 ();
 FILLER_ASAP7_75t_R FILLER_0_212_30 ();
 DECAPx2_ASAP7_75t_R FILLER_0_212_42 ();
 FILLER_ASAP7_75t_R FILLER_0_212_78 ();
 FILLER_ASAP7_75t_R FILLER_0_212_90 ();
 DECAPx1_ASAP7_75t_R FILLER_0_212_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_102 ();
 FILLER_ASAP7_75t_R FILLER_0_212_111 ();
 FILLER_ASAP7_75t_R FILLER_0_212_123 ();
 DECAPx2_ASAP7_75t_R FILLER_0_212_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_137 ();
 DECAPx2_ASAP7_75t_R FILLER_0_212_144 ();
 FILLER_ASAP7_75t_R FILLER_0_212_155 ();
 FILLER_ASAP7_75t_R FILLER_0_212_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_165 ();
 FILLER_ASAP7_75t_R FILLER_0_212_172 ();
 FILLER_ASAP7_75t_R FILLER_0_212_179 ();
 FILLER_ASAP7_75t_R FILLER_0_212_187 ();
 DECAPx10_ASAP7_75t_R FILLER_0_212_195 ();
 DECAPx2_ASAP7_75t_R FILLER_0_212_217 ();
 FILLER_ASAP7_75t_R FILLER_0_212_223 ();
 FILLER_ASAP7_75t_R FILLER_0_212_231 ();
 FILLER_ASAP7_75t_R FILLER_0_212_238 ();
 FILLER_ASAP7_75t_R FILLER_0_212_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_245 ();
 DECAPx2_ASAP7_75t_R FILLER_0_212_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_260 ();
 FILLER_ASAP7_75t_R FILLER_0_212_269 ();
 DECAPx2_ASAP7_75t_R FILLER_0_212_277 ();
 FILLER_ASAP7_75t_R FILLER_0_212_283 ();
 FILLER_ASAP7_75t_R FILLER_0_212_291 ();
 DECAPx1_ASAP7_75t_R FILLER_0_212_299 ();
 FILLER_ASAP7_75t_R FILLER_0_212_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_311 ();
 FILLER_ASAP7_75t_R FILLER_0_212_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_324 ();
 FILLER_ASAP7_75t_R FILLER_0_212_335 ();
 DECAPx4_ASAP7_75t_R FILLER_0_212_345 ();
 FILLER_ASAP7_75t_R FILLER_0_212_355 ();
 FILLER_ASAP7_75t_R FILLER_0_212_363 ();
 DECAPx1_ASAP7_75t_R FILLER_0_212_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_375 ();
 FILLER_ASAP7_75t_R FILLER_0_212_384 ();
 FILLER_ASAP7_75t_R FILLER_0_212_389 ();
 DECAPx4_ASAP7_75t_R FILLER_0_212_397 ();
 FILLER_ASAP7_75t_R FILLER_0_212_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_409 ();
 DECAPx2_ASAP7_75t_R FILLER_0_212_417 ();
 FILLER_ASAP7_75t_R FILLER_0_212_429 ();
 FILLER_ASAP7_75t_R FILLER_0_212_434 ();
 DECAPx6_ASAP7_75t_R FILLER_0_212_444 ();
 DECAPx1_ASAP7_75t_R FILLER_0_212_458 ();
 DECAPx1_ASAP7_75t_R FILLER_0_212_464 ();
 DECAPx2_ASAP7_75t_R FILLER_0_212_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_486 ();
 DECAPx1_ASAP7_75t_R FILLER_0_212_499 ();
 DECAPx2_ASAP7_75t_R FILLER_0_212_509 ();
 DECAPx6_ASAP7_75t_R FILLER_0_212_518 ();
 FILLER_ASAP7_75t_R FILLER_0_212_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_534 ();
 DECAPx4_ASAP7_75t_R FILLER_0_212_540 ();
 FILLER_ASAP7_75t_R FILLER_0_212_550 ();
 FILLER_ASAP7_75t_R FILLER_0_212_563 ();
 FILLER_ASAP7_75t_R FILLER_0_212_572 ();
 DECAPx2_ASAP7_75t_R FILLER_0_212_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_591 ();
 DECAPx2_ASAP7_75t_R FILLER_0_212_595 ();
 DECAPx4_ASAP7_75t_R FILLER_0_212_612 ();
 FILLER_ASAP7_75t_R FILLER_0_212_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_630 ();
 DECAPx2_ASAP7_75t_R FILLER_0_212_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_640 ();
 DECAPx6_ASAP7_75t_R FILLER_0_212_653 ();
 DECAPx2_ASAP7_75t_R FILLER_0_212_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_673 ();
 FILLER_ASAP7_75t_R FILLER_0_212_686 ();
 DECAPx1_ASAP7_75t_R FILLER_0_212_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_698 ();
 FILLER_ASAP7_75t_R FILLER_0_212_705 ();
 DECAPx1_ASAP7_75t_R FILLER_0_212_713 ();
 DECAPx10_ASAP7_75t_R FILLER_0_212_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_212_750 ();
 FILLER_ASAP7_75t_R FILLER_0_212_756 ();
 FILLER_ASAP7_75t_R FILLER_0_212_763 ();
 FILLER_ASAP7_75t_R FILLER_0_212_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_770 ();
 DECAPx2_ASAP7_75t_R FILLER_0_212_776 ();
 FILLER_ASAP7_75t_R FILLER_0_212_792 ();
 FILLER_ASAP7_75t_R FILLER_0_212_804 ();
 FILLER_ASAP7_75t_R FILLER_0_212_816 ();
 FILLER_ASAP7_75t_R FILLER_0_212_838 ();
 DECAPx2_ASAP7_75t_R FILLER_0_212_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_852 ();
 DECAPx2_ASAP7_75t_R FILLER_0_212_865 ();
 FILLER_ASAP7_75t_R FILLER_0_212_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_873 ();
 FILLER_ASAP7_75t_R FILLER_0_212_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_886 ();
 FILLER_ASAP7_75t_R FILLER_0_212_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_897 ();
 DECAPx2_ASAP7_75t_R FILLER_0_212_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_910 ();
 FILLER_ASAP7_75t_R FILLER_0_212_917 ();
 FILLER_ASAP7_75t_R FILLER_0_212_930 ();
 DECAPx1_ASAP7_75t_R FILLER_0_212_935 ();
 DECAPx1_ASAP7_75t_R FILLER_0_212_946 ();
 DECAPx10_ASAP7_75t_R FILLER_0_212_956 ();
 DECAPx6_ASAP7_75t_R FILLER_0_212_978 ();
 DECAPx2_ASAP7_75t_R FILLER_0_212_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_998 ();
 FILLER_ASAP7_75t_R FILLER_0_212_1020 ();
 FILLER_ASAP7_75t_R FILLER_0_212_1032 ();
 FILLER_ASAP7_75t_R FILLER_0_212_1039 ();
 FILLER_ASAP7_75t_R FILLER_0_212_1059 ();
 FILLER_ASAP7_75t_R FILLER_0_212_1067 ();
 FILLER_ASAP7_75t_R FILLER_0_212_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_1077 ();
 FILLER_ASAP7_75t_R FILLER_0_212_1084 ();
 FILLER_ASAP7_75t_R FILLER_0_212_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_1091 ();
 DECAPx10_ASAP7_75t_R FILLER_0_212_1098 ();
 DECAPx6_ASAP7_75t_R FILLER_0_212_1120 ();
 FILLER_ASAP7_75t_R FILLER_0_212_1134 ();
 FILLER_ASAP7_75t_R FILLER_0_212_1142 ();
 DECAPx4_ASAP7_75t_R FILLER_0_212_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_1161 ();
 FILLER_ASAP7_75t_R FILLER_0_212_1168 ();
 DECAPx2_ASAP7_75t_R FILLER_0_212_1176 ();
 DECAPx1_ASAP7_75t_R FILLER_0_212_1188 ();
 DECAPx4_ASAP7_75t_R FILLER_0_212_1198 ();
 DECAPx4_ASAP7_75t_R FILLER_0_212_1214 ();
 FILLER_ASAP7_75t_R FILLER_0_212_1230 ();
 DECAPx4_ASAP7_75t_R FILLER_0_212_1238 ();
 DECAPx2_ASAP7_75t_R FILLER_0_212_1258 ();
 FILLER_ASAP7_75t_R FILLER_0_212_1264 ();
 FILLER_ASAP7_75t_R FILLER_0_212_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_212_1277 ();
 DECAPx10_ASAP7_75t_R FILLER_0_212_1299 ();
 DECAPx10_ASAP7_75t_R FILLER_0_212_1321 ();
 DECAPx10_ASAP7_75t_R FILLER_0_212_1343 ();
 DECAPx6_ASAP7_75t_R FILLER_0_212_1365 ();
 FILLER_ASAP7_75t_R FILLER_0_212_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212_1381 ();
 DECAPx6_ASAP7_75t_R FILLER_0_213_2 ();
 FILLER_ASAP7_75t_R FILLER_0_213_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213_18 ();
 FILLER_ASAP7_75t_R FILLER_0_213_25 ();
 DECAPx1_ASAP7_75t_R FILLER_0_213_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_213_48 ();
 FILLER_ASAP7_75t_R FILLER_0_213_54 ();
 FILLER_ASAP7_75t_R FILLER_0_213_62 ();
 FILLER_ASAP7_75t_R FILLER_0_213_76 ();
 DECAPx1_ASAP7_75t_R FILLER_0_213_83 ();
 DECAPx2_ASAP7_75t_R FILLER_0_213_99 ();
 FILLER_ASAP7_75t_R FILLER_0_213_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213_112 ();
 FILLER_ASAP7_75t_R FILLER_0_213_123 ();
 FILLER_ASAP7_75t_R FILLER_0_213_130 ();
 DECAPx1_ASAP7_75t_R FILLER_0_213_144 ();
 FILLER_ASAP7_75t_R FILLER_0_213_159 ();
 FILLER_ASAP7_75t_R FILLER_0_213_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213_173 ();
 DECAPx2_ASAP7_75t_R FILLER_0_213_179 ();
 FILLER_ASAP7_75t_R FILLER_0_213_191 ();
 DECAPx10_ASAP7_75t_R FILLER_0_213_201 ();
 DECAPx4_ASAP7_75t_R FILLER_0_213_223 ();
 FILLER_ASAP7_75t_R FILLER_0_213_233 ();
 FILLER_ASAP7_75t_R FILLER_0_213_241 ();
 FILLER_ASAP7_75t_R FILLER_0_213_246 ();
 DECAPx1_ASAP7_75t_R FILLER_0_213_254 ();
 FILLER_ASAP7_75t_R FILLER_0_213_264 ();
 FILLER_ASAP7_75t_R FILLER_0_213_274 ();
 DECAPx2_ASAP7_75t_R FILLER_0_213_282 ();
 FILLER_ASAP7_75t_R FILLER_0_213_295 ();
 DECAPx10_ASAP7_75t_R FILLER_0_213_303 ();
 DECAPx2_ASAP7_75t_R FILLER_0_213_325 ();
 FILLER_ASAP7_75t_R FILLER_0_213_341 ();
 DECAPx1_ASAP7_75t_R FILLER_0_213_353 ();
 FILLER_ASAP7_75t_R FILLER_0_213_363 ();
 DECAPx6_ASAP7_75t_R FILLER_0_213_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213_387 ();
 FILLER_ASAP7_75t_R FILLER_0_213_396 ();
 DECAPx10_ASAP7_75t_R FILLER_0_213_401 ();
 DECAPx1_ASAP7_75t_R FILLER_0_213_423 ();
 FILLER_ASAP7_75t_R FILLER_0_213_433 ();
 FILLER_ASAP7_75t_R FILLER_0_213_441 ();
 DECAPx10_ASAP7_75t_R FILLER_0_213_446 ();
 DECAPx6_ASAP7_75t_R FILLER_0_213_468 ();
 FILLER_ASAP7_75t_R FILLER_0_213_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213_484 ();
 DECAPx2_ASAP7_75t_R FILLER_0_213_497 ();
 FILLER_ASAP7_75t_R FILLER_0_213_503 ();
 DECAPx10_ASAP7_75t_R FILLER_0_213_509 ();
 FILLER_ASAP7_75t_R FILLER_0_213_552 ();
 FILLER_ASAP7_75t_R FILLER_0_213_561 ();
 DECAPx2_ASAP7_75t_R FILLER_0_213_569 ();
 FILLER_ASAP7_75t_R FILLER_0_213_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213_577 ();
 DECAPx1_ASAP7_75t_R FILLER_0_213_585 ();
 DECAPx10_ASAP7_75t_R FILLER_0_213_597 ();
 DECAPx6_ASAP7_75t_R FILLER_0_213_619 ();
 DECAPx1_ASAP7_75t_R FILLER_0_213_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213_637 ();
 FILLER_ASAP7_75t_R FILLER_0_213_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213_652 ();
 DECAPx4_ASAP7_75t_R FILLER_0_213_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213_675 ();
 DECAPx1_ASAP7_75t_R FILLER_0_213_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213_686 ();
 DECAPx2_ASAP7_75t_R FILLER_0_213_694 ();
 FILLER_ASAP7_75t_R FILLER_0_213_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213_702 ();
 FILLER_ASAP7_75t_R FILLER_0_213_709 ();
 FILLER_ASAP7_75t_R FILLER_0_213_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213_719 ();
 DECAPx6_ASAP7_75t_R FILLER_0_213_726 ();
 DECAPx1_ASAP7_75t_R FILLER_0_213_740 ();
 DECAPx6_ASAP7_75t_R FILLER_0_213_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213_764 ();
 DECAPx2_ASAP7_75t_R FILLER_0_213_772 ();
 FILLER_ASAP7_75t_R FILLER_0_213_790 ();
 DECAPx1_ASAP7_75t_R FILLER_0_213_798 ();
 FILLER_ASAP7_75t_R FILLER_0_213_809 ();
 FILLER_ASAP7_75t_R FILLER_0_213_821 ();
 FILLER_ASAP7_75t_R FILLER_0_213_833 ();
 DECAPx1_ASAP7_75t_R FILLER_0_213_842 ();
 DECAPx1_ASAP7_75t_R FILLER_0_213_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213_860 ();
 FILLER_ASAP7_75t_R FILLER_0_213_867 ();
 DECAPx10_ASAP7_75t_R FILLER_0_213_875 ();
 DECAPx4_ASAP7_75t_R FILLER_0_213_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213_907 ();
 DECAPx4_ASAP7_75t_R FILLER_0_213_915 ();
 FILLER_ASAP7_75t_R FILLER_0_213_927 ();
 DECAPx6_ASAP7_75t_R FILLER_0_213_935 ();
 DECAPx2_ASAP7_75t_R FILLER_0_213_949 ();
 FILLER_ASAP7_75t_R FILLER_0_213_961 ();
 DECAPx6_ASAP7_75t_R FILLER_0_213_969 ();
 FILLER_ASAP7_75t_R FILLER_0_213_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213_985 ();
 FILLER_ASAP7_75t_R FILLER_0_213_1007 ();
 DECAPx2_ASAP7_75t_R FILLER_0_213_1015 ();
 FILLER_ASAP7_75t_R FILLER_0_213_1026 ();
 FILLER_ASAP7_75t_R FILLER_0_213_1038 ();
 FILLER_ASAP7_75t_R FILLER_0_213_1050 ();
 FILLER_ASAP7_75t_R FILLER_0_213_1062 ();
 FILLER_ASAP7_75t_R FILLER_0_213_1070 ();
 FILLER_ASAP7_75t_R FILLER_0_213_1083 ();
 FILLER_ASAP7_75t_R FILLER_0_213_1090 ();
 DECAPx2_ASAP7_75t_R FILLER_0_213_1097 ();
 FILLER_ASAP7_75t_R FILLER_0_213_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213_1105 ();
 DECAPx2_ASAP7_75t_R FILLER_0_213_1112 ();
 FILLER_ASAP7_75t_R FILLER_0_213_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213_1120 ();
 FILLER_ASAP7_75t_R FILLER_0_213_1127 ();
 FILLER_ASAP7_75t_R FILLER_0_213_1135 ();
 DECAPx1_ASAP7_75t_R FILLER_0_213_1142 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213_1146 ();
 DECAPx4_ASAP7_75t_R FILLER_0_213_1153 ();
 DECAPx2_ASAP7_75t_R FILLER_0_213_1171 ();
 FILLER_ASAP7_75t_R FILLER_0_213_1177 ();
 FILLER_ASAP7_75t_R FILLER_0_213_1185 ();
 DECAPx1_ASAP7_75t_R FILLER_0_213_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213_1194 ();
 DECAPx2_ASAP7_75t_R FILLER_0_213_1201 ();
 FILLER_ASAP7_75t_R FILLER_0_213_1207 ();
 DECAPx2_ASAP7_75t_R FILLER_0_213_1220 ();
 DECAPx2_ASAP7_75t_R FILLER_0_213_1232 ();
 FILLER_ASAP7_75t_R FILLER_0_213_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213_1240 ();
 FILLER_ASAP7_75t_R FILLER_0_213_1252 ();
 DECAPx2_ASAP7_75t_R FILLER_0_213_1260 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213_1266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_213_1273 ();
 DECAPx10_ASAP7_75t_R FILLER_0_213_1295 ();
 DECAPx10_ASAP7_75t_R FILLER_0_213_1317 ();
 DECAPx10_ASAP7_75t_R FILLER_0_213_1339 ();
 DECAPx6_ASAP7_75t_R FILLER_0_213_1361 ();
 DECAPx2_ASAP7_75t_R FILLER_0_213_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213_1381 ();
 DECAPx2_ASAP7_75t_R FILLER_0_214_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_8 ();
 FILLER_ASAP7_75t_R FILLER_0_214_15 ();
 FILLER_ASAP7_75t_R FILLER_0_214_23 ();
 FILLER_ASAP7_75t_R FILLER_0_214_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_33 ();
 DECAPx1_ASAP7_75t_R FILLER_0_214_54 ();
 DECAPx1_ASAP7_75t_R FILLER_0_214_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_68 ();
 FILLER_ASAP7_75t_R FILLER_0_214_79 ();
 FILLER_ASAP7_75t_R FILLER_0_214_91 ();
 FILLER_ASAP7_75t_R FILLER_0_214_103 ();
 FILLER_ASAP7_75t_R FILLER_0_214_110 ();
 FILLER_ASAP7_75t_R FILLER_0_214_122 ();
 FILLER_ASAP7_75t_R FILLER_0_214_129 ();
 FILLER_ASAP7_75t_R FILLER_0_214_134 ();
 DECAPx2_ASAP7_75t_R FILLER_0_214_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_160 ();
 DECAPx2_ASAP7_75t_R FILLER_0_214_171 ();
 FILLER_ASAP7_75t_R FILLER_0_214_188 ();
 DECAPx2_ASAP7_75t_R FILLER_0_214_195 ();
 DECAPx10_ASAP7_75t_R FILLER_0_214_211 ();
 FILLER_ASAP7_75t_R FILLER_0_214_233 ();
 FILLER_ASAP7_75t_R FILLER_0_214_241 ();
 DECAPx2_ASAP7_75t_R FILLER_0_214_249 ();
 FILLER_ASAP7_75t_R FILLER_0_214_261 ();
 DECAPx6_ASAP7_75t_R FILLER_0_214_271 ();
 FILLER_ASAP7_75t_R FILLER_0_214_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_287 ();
 DECAPx1_ASAP7_75t_R FILLER_0_214_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_298 ();
 FILLER_ASAP7_75t_R FILLER_0_214_319 ();
 DECAPx4_ASAP7_75t_R FILLER_0_214_343 ();
 FILLER_ASAP7_75t_R FILLER_0_214_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_361 ();
 FILLER_ASAP7_75t_R FILLER_0_214_368 ();
 DECAPx2_ASAP7_75t_R FILLER_0_214_376 ();
 FILLER_ASAP7_75t_R FILLER_0_214_382 ();
 FILLER_ASAP7_75t_R FILLER_0_214_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_214_399 ();
 DECAPx4_ASAP7_75t_R FILLER_0_214_421 ();
 FILLER_ASAP7_75t_R FILLER_0_214_439 ();
 DECAPx6_ASAP7_75t_R FILLER_0_214_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_214_464 ();
 DECAPx1_ASAP7_75t_R FILLER_0_214_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_490 ();
 DECAPx1_ASAP7_75t_R FILLER_0_214_512 ();
 DECAPx4_ASAP7_75t_R FILLER_0_214_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_532 ();
 DECAPx4_ASAP7_75t_R FILLER_0_214_536 ();
 FILLER_ASAP7_75t_R FILLER_0_214_549 ();
 FILLER_ASAP7_75t_R FILLER_0_214_561 ();
 DECAPx2_ASAP7_75t_R FILLER_0_214_571 ();
 FILLER_ASAP7_75t_R FILLER_0_214_588 ();
 DECAPx4_ASAP7_75t_R FILLER_0_214_596 ();
 FILLER_ASAP7_75t_R FILLER_0_214_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_608 ();
 FILLER_ASAP7_75t_R FILLER_0_214_617 ();
 FILLER_ASAP7_75t_R FILLER_0_214_625 ();
 FILLER_ASAP7_75t_R FILLER_0_214_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_641 ();
 FILLER_ASAP7_75t_R FILLER_0_214_653 ();
 FILLER_ASAP7_75t_R FILLER_0_214_676 ();
 DECAPx1_ASAP7_75t_R FILLER_0_214_689 ();
 DECAPx1_ASAP7_75t_R FILLER_0_214_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_703 ();
 FILLER_ASAP7_75t_R FILLER_0_214_710 ();
 DECAPx2_ASAP7_75t_R FILLER_0_214_715 ();
 FILLER_ASAP7_75t_R FILLER_0_214_724 ();
 DECAPx10_ASAP7_75t_R FILLER_0_214_732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_214_754 ();
 FILLER_ASAP7_75t_R FILLER_0_214_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_778 ();
 DECAPx4_ASAP7_75t_R FILLER_0_214_789 ();
 FILLER_ASAP7_75t_R FILLER_0_214_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_801 ();
 FILLER_ASAP7_75t_R FILLER_0_214_808 ();
 FILLER_ASAP7_75t_R FILLER_0_214_815 ();
 FILLER_ASAP7_75t_R FILLER_0_214_822 ();
 FILLER_ASAP7_75t_R FILLER_0_214_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_831 ();
 FILLER_ASAP7_75t_R FILLER_0_214_838 ();
 DECAPx1_ASAP7_75t_R FILLER_0_214_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_214_856 ();
 DECAPx6_ASAP7_75t_R FILLER_0_214_878 ();
 DECAPx1_ASAP7_75t_R FILLER_0_214_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_896 ();
 DECAPx4_ASAP7_75t_R FILLER_0_214_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_913 ();
 FILLER_ASAP7_75t_R FILLER_0_214_938 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_940 ();
 DECAPx2_ASAP7_75t_R FILLER_0_214_948 ();
 FILLER_ASAP7_75t_R FILLER_0_214_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_956 ();
 DECAPx2_ASAP7_75t_R FILLER_0_214_963 ();
 FILLER_ASAP7_75t_R FILLER_0_214_975 ();
 DECAPx1_ASAP7_75t_R FILLER_0_214_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_987 ();
 DECAPx4_ASAP7_75t_R FILLER_0_214_991 ();
 DECAPx6_ASAP7_75t_R FILLER_0_214_1004 ();
 DECAPx1_ASAP7_75t_R FILLER_0_214_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_1022 ();
 FILLER_ASAP7_75t_R FILLER_0_214_1033 ();
 FILLER_ASAP7_75t_R FILLER_0_214_1045 ();
 FILLER_ASAP7_75t_R FILLER_0_214_1057 ();
 FILLER_ASAP7_75t_R FILLER_0_214_1069 ();
 FILLER_ASAP7_75t_R FILLER_0_214_1077 ();
 FILLER_ASAP7_75t_R FILLER_0_214_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_1087 ();
 DECAPx2_ASAP7_75t_R FILLER_0_214_1094 ();
 FILLER_ASAP7_75t_R FILLER_0_214_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_1102 ();
 FILLER_ASAP7_75t_R FILLER_0_214_1114 ();
 FILLER_ASAP7_75t_R FILLER_0_214_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_1123 ();
 FILLER_ASAP7_75t_R FILLER_0_214_1130 ();
 FILLER_ASAP7_75t_R FILLER_0_214_1138 ();
 DECAPx4_ASAP7_75t_R FILLER_0_214_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_1156 ();
 DECAPx2_ASAP7_75t_R FILLER_0_214_1167 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_1173 ();
 FILLER_ASAP7_75t_R FILLER_0_214_1182 ();
 FILLER_ASAP7_75t_R FILLER_0_214_1190 ();
 FILLER_ASAP7_75t_R FILLER_0_214_1198 ();
 DECAPx1_ASAP7_75t_R FILLER_0_214_1206 ();
 DECAPx1_ASAP7_75t_R FILLER_0_214_1216 ();
 FILLER_ASAP7_75t_R FILLER_0_214_1228 ();
 FILLER_ASAP7_75t_R FILLER_0_214_1236 ();
 FILLER_ASAP7_75t_R FILLER_0_214_1243 ();
 FILLER_ASAP7_75t_R FILLER_0_214_1255 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214_1257 ();
 DECAPx10_ASAP7_75t_R FILLER_0_214_1268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_214_1290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_214_1312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_214_1334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_214_1356 ();
 DECAPx1_ASAP7_75t_R FILLER_0_214_1378 ();
 DECAPx2_ASAP7_75t_R FILLER_0_215_2 ();
 FILLER_ASAP7_75t_R FILLER_0_215_8 ();
 DECAPx2_ASAP7_75t_R FILLER_0_215_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_23 ();
 DECAPx2_ASAP7_75t_R FILLER_0_215_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_37 ();
 FILLER_ASAP7_75t_R FILLER_0_215_44 ();
 FILLER_ASAP7_75t_R FILLER_0_215_58 ();
 FILLER_ASAP7_75t_R FILLER_0_215_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_68 ();
 FILLER_ASAP7_75t_R FILLER_0_215_77 ();
 FILLER_ASAP7_75t_R FILLER_0_215_89 ();
 FILLER_ASAP7_75t_R FILLER_0_215_97 ();
 FILLER_ASAP7_75t_R FILLER_0_215_109 ();
 FILLER_ASAP7_75t_R FILLER_0_215_119 ();
 FILLER_ASAP7_75t_R FILLER_0_215_126 ();
 FILLER_ASAP7_75t_R FILLER_0_215_134 ();
 FILLER_ASAP7_75t_R FILLER_0_215_142 ();
 FILLER_ASAP7_75t_R FILLER_0_215_154 ();
 DECAPx2_ASAP7_75t_R FILLER_0_215_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_172 ();
 DECAPx6_ASAP7_75t_R FILLER_0_215_185 ();
 DECAPx1_ASAP7_75t_R FILLER_0_215_199 ();
 FILLER_ASAP7_75t_R FILLER_0_215_213 ();
 DECAPx1_ASAP7_75t_R FILLER_0_215_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_227 ();
 FILLER_ASAP7_75t_R FILLER_0_215_235 ();
 FILLER_ASAP7_75t_R FILLER_0_215_243 ();
 DECAPx1_ASAP7_75t_R FILLER_0_215_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_252 ();
 DECAPx10_ASAP7_75t_R FILLER_0_215_261 ();
 DECAPx2_ASAP7_75t_R FILLER_0_215_283 ();
 FILLER_ASAP7_75t_R FILLER_0_215_295 ();
 DECAPx10_ASAP7_75t_R FILLER_0_215_300 ();
 DECAPx2_ASAP7_75t_R FILLER_0_215_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_328 ();
 FILLER_ASAP7_75t_R FILLER_0_215_339 ();
 FILLER_ASAP7_75t_R FILLER_0_215_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_346 ();
 FILLER_ASAP7_75t_R FILLER_0_215_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_355 ();
 FILLER_ASAP7_75t_R FILLER_0_215_362 ();
 DECAPx2_ASAP7_75t_R FILLER_0_215_371 ();
 DECAPx2_ASAP7_75t_R FILLER_0_215_388 ();
 FILLER_ASAP7_75t_R FILLER_0_215_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_396 ();
 FILLER_ASAP7_75t_R FILLER_0_215_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_410 ();
 FILLER_ASAP7_75t_R FILLER_0_215_418 ();
 FILLER_ASAP7_75t_R FILLER_0_215_426 ();
 FILLER_ASAP7_75t_R FILLER_0_215_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_433 ();
 DECAPx6_ASAP7_75t_R FILLER_0_215_440 ();
 FILLER_ASAP7_75t_R FILLER_0_215_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_456 ();
 DECAPx1_ASAP7_75t_R FILLER_0_215_467 ();
 DECAPx4_ASAP7_75t_R FILLER_0_215_481 ();
 FILLER_ASAP7_75t_R FILLER_0_215_499 ();
 DECAPx4_ASAP7_75t_R FILLER_0_215_504 ();
 FILLER_ASAP7_75t_R FILLER_0_215_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_516 ();
 FILLER_ASAP7_75t_R FILLER_0_215_525 ();
 DECAPx4_ASAP7_75t_R FILLER_0_215_533 ();
 FILLER_ASAP7_75t_R FILLER_0_215_543 ();
 FILLER_ASAP7_75t_R FILLER_0_215_566 ();
 DECAPx2_ASAP7_75t_R FILLER_0_215_589 ();
 DECAPx4_ASAP7_75t_R FILLER_0_215_607 ();
 FILLER_ASAP7_75t_R FILLER_0_215_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_215_626 ();
 DECAPx2_ASAP7_75t_R FILLER_0_215_648 ();
 FILLER_ASAP7_75t_R FILLER_0_215_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_656 ();
 DECAPx6_ASAP7_75t_R FILLER_0_215_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_674 ();
 FILLER_ASAP7_75t_R FILLER_0_215_687 ();
 DECAPx2_ASAP7_75t_R FILLER_0_215_699 ();
 FILLER_ASAP7_75t_R FILLER_0_215_711 ();
 DECAPx1_ASAP7_75t_R FILLER_0_215_716 ();
 FILLER_ASAP7_75t_R FILLER_0_215_726 ();
 FILLER_ASAP7_75t_R FILLER_0_215_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_736 ();
 FILLER_ASAP7_75t_R FILLER_0_215_743 ();
 DECAPx2_ASAP7_75t_R FILLER_0_215_751 ();
 FILLER_ASAP7_75t_R FILLER_0_215_757 ();
 DECAPx2_ASAP7_75t_R FILLER_0_215_766 ();
 FILLER_ASAP7_75t_R FILLER_0_215_784 ();
 DECAPx1_ASAP7_75t_R FILLER_0_215_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_797 ();
 DECAPx2_ASAP7_75t_R FILLER_0_215_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_811 ();
 FILLER_ASAP7_75t_R FILLER_0_215_818 ();
 FILLER_ASAP7_75t_R FILLER_0_215_826 ();
 FILLER_ASAP7_75t_R FILLER_0_215_834 ();
 FILLER_ASAP7_75t_R FILLER_0_215_842 ();
 FILLER_ASAP7_75t_R FILLER_0_215_855 ();
 FILLER_ASAP7_75t_R FILLER_0_215_863 ();
 FILLER_ASAP7_75t_R FILLER_0_215_871 ();
 DECAPx1_ASAP7_75t_R FILLER_0_215_879 ();
 FILLER_ASAP7_75t_R FILLER_0_215_889 ();
 DECAPx10_ASAP7_75t_R FILLER_0_215_903 ();
 FILLER_ASAP7_75t_R FILLER_0_215_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_929 ();
 FILLER_ASAP7_75t_R FILLER_0_215_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_938 ();
 FILLER_ASAP7_75t_R FILLER_0_215_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_947 ();
 FILLER_ASAP7_75t_R FILLER_0_215_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_956 ();
 FILLER_ASAP7_75t_R FILLER_0_215_963 ();
 FILLER_ASAP7_75t_R FILLER_0_215_971 ();
 DECAPx1_ASAP7_75t_R FILLER_0_215_979 ();
 DECAPx10_ASAP7_75t_R FILLER_0_215_989 ();
 DECAPx2_ASAP7_75t_R FILLER_0_215_1011 ();
 FILLER_ASAP7_75t_R FILLER_0_215_1027 ();
 FILLER_ASAP7_75t_R FILLER_0_215_1047 ();
 DECAPx1_ASAP7_75t_R FILLER_0_215_1055 ();
 FILLER_ASAP7_75t_R FILLER_0_215_1070 ();
 DECAPx2_ASAP7_75t_R FILLER_0_215_1082 ();
 DECAPx4_ASAP7_75t_R FILLER_0_215_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_1109 ();
 FILLER_ASAP7_75t_R FILLER_0_215_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_1118 ();
 FILLER_ASAP7_75t_R FILLER_0_215_1122 ();
 FILLER_ASAP7_75t_R FILLER_0_215_1130 ();
 DECAPx4_ASAP7_75t_R FILLER_0_215_1139 ();
 DECAPx1_ASAP7_75t_R FILLER_0_215_1159 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_1163 ();
 FILLER_ASAP7_75t_R FILLER_0_215_1174 ();
 FILLER_ASAP7_75t_R FILLER_0_215_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_215_1194 ();
 FILLER_ASAP7_75t_R FILLER_0_215_1202 ();
 DECAPx1_ASAP7_75t_R FILLER_0_215_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_1214 ();
 FILLER_ASAP7_75t_R FILLER_0_215_1225 ();
 FILLER_ASAP7_75t_R FILLER_0_215_1237 ();
 FILLER_ASAP7_75t_R FILLER_0_215_1242 ();
 FILLER_ASAP7_75t_R FILLER_0_215_1252 ();
 DECAPx10_ASAP7_75t_R FILLER_0_215_1259 ();
 DECAPx10_ASAP7_75t_R FILLER_0_215_1281 ();
 DECAPx10_ASAP7_75t_R FILLER_0_215_1303 ();
 DECAPx10_ASAP7_75t_R FILLER_0_215_1325 ();
 DECAPx10_ASAP7_75t_R FILLER_0_215_1347 ();
 DECAPx4_ASAP7_75t_R FILLER_0_215_1369 ();
 FILLER_ASAP7_75t_R FILLER_0_215_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_216_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_4 ();
 FILLER_ASAP7_75t_R FILLER_0_216_11 ();
 DECAPx1_ASAP7_75t_R FILLER_0_216_23 ();
 FILLER_ASAP7_75t_R FILLER_0_216_35 ();
 FILLER_ASAP7_75t_R FILLER_0_216_47 ();
 DECAPx2_ASAP7_75t_R FILLER_0_216_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_65 ();
 FILLER_ASAP7_75t_R FILLER_0_216_72 ();
 DECAPx1_ASAP7_75t_R FILLER_0_216_84 ();
 DECAPx1_ASAP7_75t_R FILLER_0_216_98 ();
 FILLER_ASAP7_75t_R FILLER_0_216_112 ();
 FILLER_ASAP7_75t_R FILLER_0_216_126 ();
 FILLER_ASAP7_75t_R FILLER_0_216_133 ();
 FILLER_ASAP7_75t_R FILLER_0_216_147 ();
 FILLER_ASAP7_75t_R FILLER_0_216_154 ();
 FILLER_ASAP7_75t_R FILLER_0_216_164 ();
 DECAPx6_ASAP7_75t_R FILLER_0_216_174 ();
 DECAPx2_ASAP7_75t_R FILLER_0_216_188 ();
 FILLER_ASAP7_75t_R FILLER_0_216_214 ();
 DECAPx6_ASAP7_75t_R FILLER_0_216_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_240 ();
 DECAPx1_ASAP7_75t_R FILLER_0_216_247 ();
 DECAPx1_ASAP7_75t_R FILLER_0_216_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_258 ();
 FILLER_ASAP7_75t_R FILLER_0_216_269 ();
 FILLER_ASAP7_75t_R FILLER_0_216_277 ();
 FILLER_ASAP7_75t_R FILLER_0_216_285 ();
 FILLER_ASAP7_75t_R FILLER_0_216_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_297 ();
 FILLER_ASAP7_75t_R FILLER_0_216_304 ();
 FILLER_ASAP7_75t_R FILLER_0_216_312 ();
 DECAPx6_ASAP7_75t_R FILLER_0_216_320 ();
 FILLER_ASAP7_75t_R FILLER_0_216_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_336 ();
 DECAPx4_ASAP7_75t_R FILLER_0_216_341 ();
 FILLER_ASAP7_75t_R FILLER_0_216_351 ();
 FILLER_ASAP7_75t_R FILLER_0_216_358 ();
 FILLER_ASAP7_75t_R FILLER_0_216_366 ();
 DECAPx1_ASAP7_75t_R FILLER_0_216_374 ();
 DECAPx2_ASAP7_75t_R FILLER_0_216_381 ();
 DECAPx2_ASAP7_75t_R FILLER_0_216_393 ();
 DECAPx2_ASAP7_75t_R FILLER_0_216_405 ();
 DECAPx2_ASAP7_75t_R FILLER_0_216_419 ();
 FILLER_ASAP7_75t_R FILLER_0_216_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_427 ();
 DECAPx1_ASAP7_75t_R FILLER_0_216_436 ();
 DECAPx6_ASAP7_75t_R FILLER_0_216_443 ();
 DECAPx1_ASAP7_75t_R FILLER_0_216_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_461 ();
 DECAPx2_ASAP7_75t_R FILLER_0_216_464 ();
 DECAPx2_ASAP7_75t_R FILLER_0_216_478 ();
 FILLER_ASAP7_75t_R FILLER_0_216_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_486 ();
 DECAPx6_ASAP7_75t_R FILLER_0_216_499 ();
 DECAPx1_ASAP7_75t_R FILLER_0_216_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_517 ();
 DECAPx2_ASAP7_75t_R FILLER_0_216_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_532 ();
 FILLER_ASAP7_75t_R FILLER_0_216_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_546 ();
 DECAPx6_ASAP7_75t_R FILLER_0_216_550 ();
 FILLER_ASAP7_75t_R FILLER_0_216_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_566 ();
 FILLER_ASAP7_75t_R FILLER_0_216_573 ();
 DECAPx1_ASAP7_75t_R FILLER_0_216_578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_216_603 ();
 FILLER_ASAP7_75t_R FILLER_0_216_617 ();
 DECAPx1_ASAP7_75t_R FILLER_0_216_630 ();
 DECAPx1_ASAP7_75t_R FILLER_0_216_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_216_650 ();
 DECAPx1_ASAP7_75t_R FILLER_0_216_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_676 ();
 DECAPx1_ASAP7_75t_R FILLER_0_216_689 ();
 DECAPx2_ASAP7_75t_R FILLER_0_216_714 ();
 FILLER_ASAP7_75t_R FILLER_0_216_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_216_736 ();
 DECAPx1_ASAP7_75t_R FILLER_0_216_748 ();
 FILLER_ASAP7_75t_R FILLER_0_216_759 ();
 FILLER_ASAP7_75t_R FILLER_0_216_766 ();
 DECAPx4_ASAP7_75t_R FILLER_0_216_774 ();
 DECAPx4_ASAP7_75t_R FILLER_0_216_787 ();
 FILLER_ASAP7_75t_R FILLER_0_216_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_799 ();
 FILLER_ASAP7_75t_R FILLER_0_216_806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_216_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_828 ();
 FILLER_ASAP7_75t_R FILLER_0_216_835 ();
 DECAPx2_ASAP7_75t_R FILLER_0_216_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_849 ();
 DECAPx2_ASAP7_75t_R FILLER_0_216_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_862 ();
 FILLER_ASAP7_75t_R FILLER_0_216_869 ();
 FILLER_ASAP7_75t_R FILLER_0_216_881 ();
 DECAPx1_ASAP7_75t_R FILLER_0_216_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_893 ();
 DECAPx2_ASAP7_75t_R FILLER_0_216_902 ();
 FILLER_ASAP7_75t_R FILLER_0_216_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_910 ();
 FILLER_ASAP7_75t_R FILLER_0_216_917 ();
 FILLER_ASAP7_75t_R FILLER_0_216_929 ();
 FILLER_ASAP7_75t_R FILLER_0_216_941 ();
 FILLER_ASAP7_75t_R FILLER_0_216_949 ();
 FILLER_ASAP7_75t_R FILLER_0_216_957 ();
 FILLER_ASAP7_75t_R FILLER_0_216_965 ();
 FILLER_ASAP7_75t_R FILLER_0_216_973 ();
 FILLER_ASAP7_75t_R FILLER_0_216_981 ();
 FILLER_ASAP7_75t_R FILLER_0_216_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_991 ();
 DECAPx6_ASAP7_75t_R FILLER_0_216_1013 ();
 FILLER_ASAP7_75t_R FILLER_0_216_1065 ();
 DECAPx1_ASAP7_75t_R FILLER_0_216_1073 ();
 FILLER_ASAP7_75t_R FILLER_0_216_1085 ();
 FILLER_ASAP7_75t_R FILLER_0_216_1093 ();
 FILLER_ASAP7_75t_R FILLER_0_216_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_1103 ();
 DECAPx2_ASAP7_75t_R FILLER_0_216_1110 ();
 FILLER_ASAP7_75t_R FILLER_0_216_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_1118 ();
 FILLER_ASAP7_75t_R FILLER_0_216_1122 ();
 FILLER_ASAP7_75t_R FILLER_0_216_1129 ();
 FILLER_ASAP7_75t_R FILLER_0_216_1137 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_1139 ();
 FILLER_ASAP7_75t_R FILLER_0_216_1143 ();
 FILLER_ASAP7_75t_R FILLER_0_216_1151 ();
 DECAPx2_ASAP7_75t_R FILLER_0_216_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_1169 ();
 FILLER_ASAP7_75t_R FILLER_0_216_1180 ();
 FILLER_ASAP7_75t_R FILLER_0_216_1192 ();
 FILLER_ASAP7_75t_R FILLER_0_216_1200 ();
 FILLER_ASAP7_75t_R FILLER_0_216_1207 ();
 DECAPx1_ASAP7_75t_R FILLER_0_216_1219 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_1223 ();
 FILLER_ASAP7_75t_R FILLER_0_216_1235 ();
 FILLER_ASAP7_75t_R FILLER_0_216_1243 ();
 FILLER_ASAP7_75t_R FILLER_0_216_1251 ();
 DECAPx10_ASAP7_75t_R FILLER_0_216_1259 ();
 DECAPx10_ASAP7_75t_R FILLER_0_216_1281 ();
 DECAPx10_ASAP7_75t_R FILLER_0_216_1303 ();
 DECAPx10_ASAP7_75t_R FILLER_0_216_1325 ();
 DECAPx10_ASAP7_75t_R FILLER_0_216_1347 ();
 DECAPx4_ASAP7_75t_R FILLER_0_216_1369 ();
 FILLER_ASAP7_75t_R FILLER_0_216_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216_1381 ();
 FILLER_ASAP7_75t_R FILLER_0_217_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_4 ();
 FILLER_ASAP7_75t_R FILLER_0_217_21 ();
 FILLER_ASAP7_75t_R FILLER_0_217_33 ();
 FILLER_ASAP7_75t_R FILLER_0_217_41 ();
 FILLER_ASAP7_75t_R FILLER_0_217_53 ();
 DECAPx2_ASAP7_75t_R FILLER_0_217_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_68 ();
 FILLER_ASAP7_75t_R FILLER_0_217_75 ();
 FILLER_ASAP7_75t_R FILLER_0_217_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_89 ();
 FILLER_ASAP7_75t_R FILLER_0_217_100 ();
 FILLER_ASAP7_75t_R FILLER_0_217_112 ();
 FILLER_ASAP7_75t_R FILLER_0_217_124 ();
 DECAPx2_ASAP7_75t_R FILLER_0_217_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_140 ();
 FILLER_ASAP7_75t_R FILLER_0_217_147 ();
 DECAPx1_ASAP7_75t_R FILLER_0_217_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_160 ();
 DECAPx2_ASAP7_75t_R FILLER_0_217_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_172 ();
 FILLER_ASAP7_75t_R FILLER_0_217_203 ();
 DECAPx1_ASAP7_75t_R FILLER_0_217_215 ();
 FILLER_ASAP7_75t_R FILLER_0_217_224 ();
 DECAPx6_ASAP7_75t_R FILLER_0_217_231 ();
 FILLER_ASAP7_75t_R FILLER_0_217_245 ();
 FILLER_ASAP7_75t_R FILLER_0_217_251 ();
 DECAPx2_ASAP7_75t_R FILLER_0_217_261 ();
 FILLER_ASAP7_75t_R FILLER_0_217_267 ();
 DECAPx2_ASAP7_75t_R FILLER_0_217_275 ();
 DECAPx4_ASAP7_75t_R FILLER_0_217_284 ();
 FILLER_ASAP7_75t_R FILLER_0_217_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_296 ();
 DECAPx6_ASAP7_75t_R FILLER_0_217_300 ();
 FILLER_ASAP7_75t_R FILLER_0_217_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_316 ();
 FILLER_ASAP7_75t_R FILLER_0_217_323 ();
 DECAPx4_ASAP7_75t_R FILLER_0_217_335 ();
 FILLER_ASAP7_75t_R FILLER_0_217_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_347 ();
 DECAPx2_ASAP7_75t_R FILLER_0_217_353 ();
 FILLER_ASAP7_75t_R FILLER_0_217_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_361 ();
 FILLER_ASAP7_75t_R FILLER_0_217_366 ();
 FILLER_ASAP7_75t_R FILLER_0_217_374 ();
 DECAPx4_ASAP7_75t_R FILLER_0_217_382 ();
 FILLER_ASAP7_75t_R FILLER_0_217_392 ();
 FILLER_ASAP7_75t_R FILLER_0_217_400 ();
 FILLER_ASAP7_75t_R FILLER_0_217_408 ();
 DECAPx2_ASAP7_75t_R FILLER_0_217_413 ();
 FILLER_ASAP7_75t_R FILLER_0_217_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_421 ();
 FILLER_ASAP7_75t_R FILLER_0_217_428 ();
 DECAPx1_ASAP7_75t_R FILLER_0_217_436 ();
 DECAPx6_ASAP7_75t_R FILLER_0_217_446 ();
 DECAPx2_ASAP7_75t_R FILLER_0_217_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_466 ();
 FILLER_ASAP7_75t_R FILLER_0_217_475 ();
 FILLER_ASAP7_75t_R FILLER_0_217_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_485 ();
 DECAPx6_ASAP7_75t_R FILLER_0_217_498 ();
 DECAPx1_ASAP7_75t_R FILLER_0_217_512 ();
 DECAPx6_ASAP7_75t_R FILLER_0_217_522 ();
 FILLER_ASAP7_75t_R FILLER_0_217_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_538 ();
 DECAPx4_ASAP7_75t_R FILLER_0_217_545 ();
 FILLER_ASAP7_75t_R FILLER_0_217_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_217_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_583 ();
 DECAPx4_ASAP7_75t_R FILLER_0_217_587 ();
 FILLER_ASAP7_75t_R FILLER_0_217_609 ();
 DECAPx2_ASAP7_75t_R FILLER_0_217_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_629 ();
 FILLER_ASAP7_75t_R FILLER_0_217_651 ();
 DECAPx6_ASAP7_75t_R FILLER_0_217_674 ();
 DECAPx2_ASAP7_75t_R FILLER_0_217_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_694 ();
 DECAPx10_ASAP7_75t_R FILLER_0_217_698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_217_720 ();
 FILLER_ASAP7_75t_R FILLER_0_217_748 ();
 DECAPx2_ASAP7_75t_R FILLER_0_217_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_762 ();
 DECAPx2_ASAP7_75t_R FILLER_0_217_766 ();
 FILLER_ASAP7_75t_R FILLER_0_217_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_780 ();
 FILLER_ASAP7_75t_R FILLER_0_217_784 ();
 DECAPx2_ASAP7_75t_R FILLER_0_217_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_802 ();
 FILLER_ASAP7_75t_R FILLER_0_217_811 ();
 DECAPx4_ASAP7_75t_R FILLER_0_217_819 ();
 FILLER_ASAP7_75t_R FILLER_0_217_829 ();
 DECAPx4_ASAP7_75t_R FILLER_0_217_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_847 ();
 DECAPx6_ASAP7_75t_R FILLER_0_217_854 ();
 DECAPx1_ASAP7_75t_R FILLER_0_217_868 ();
 FILLER_ASAP7_75t_R FILLER_0_217_878 ();
 DECAPx6_ASAP7_75t_R FILLER_0_217_886 ();
 FILLER_ASAP7_75t_R FILLER_0_217_900 ();
 DECAPx1_ASAP7_75t_R FILLER_0_217_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_912 ();
 DECAPx2_ASAP7_75t_R FILLER_0_217_919 ();
 DECAPx6_ASAP7_75t_R FILLER_0_217_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_941 ();
 FILLER_ASAP7_75t_R FILLER_0_217_948 ();
 DECAPx4_ASAP7_75t_R FILLER_0_217_956 ();
 DECAPx10_ASAP7_75t_R FILLER_0_217_972 ();
 DECAPx4_ASAP7_75t_R FILLER_0_217_997 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_1007 ();
 DECAPx4_ASAP7_75t_R FILLER_0_217_1011 ();
 FILLER_ASAP7_75t_R FILLER_0_217_1021 ();
 FILLER_ASAP7_75t_R FILLER_0_217_1026 ();
 FILLER_ASAP7_75t_R FILLER_0_217_1039 ();
 DECAPx2_ASAP7_75t_R FILLER_0_217_1051 ();
 FILLER_ASAP7_75t_R FILLER_0_217_1065 ();
 DECAPx1_ASAP7_75t_R FILLER_0_217_1073 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_1077 ();
 DECAPx2_ASAP7_75t_R FILLER_0_217_1090 ();
 DECAPx2_ASAP7_75t_R FILLER_0_217_1102 ();
 FILLER_ASAP7_75t_R FILLER_0_217_1115 ();
 DECAPx1_ASAP7_75t_R FILLER_0_217_1123 ();
 DECAPx2_ASAP7_75t_R FILLER_0_217_1131 ();
 FILLER_ASAP7_75t_R FILLER_0_217_1143 ();
 DECAPx1_ASAP7_75t_R FILLER_0_217_1151 ();
 FILLER_ASAP7_75t_R FILLER_0_217_1158 ();
 FILLER_ASAP7_75t_R FILLER_0_217_1170 ();
 FILLER_ASAP7_75t_R FILLER_0_217_1182 ();
 FILLER_ASAP7_75t_R FILLER_0_217_1194 ();
 FILLER_ASAP7_75t_R FILLER_0_217_1202 ();
 FILLER_ASAP7_75t_R FILLER_0_217_1214 ();
 FILLER_ASAP7_75t_R FILLER_0_217_1228 ();
 FILLER_ASAP7_75t_R FILLER_0_217_1235 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_1237 ();
 DECAPx10_ASAP7_75t_R FILLER_0_217_1243 ();
 DECAPx10_ASAP7_75t_R FILLER_0_217_1265 ();
 DECAPx10_ASAP7_75t_R FILLER_0_217_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_0_217_1309 ();
 DECAPx10_ASAP7_75t_R FILLER_0_217_1331 ();
 DECAPx10_ASAP7_75t_R FILLER_0_217_1353 ();
 DECAPx2_ASAP7_75t_R FILLER_0_217_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217_1381 ();
 DECAPx6_ASAP7_75t_R FILLER_0_218_2 ();
 FILLER_ASAP7_75t_R FILLER_0_218_16 ();
 FILLER_ASAP7_75t_R FILLER_0_218_23 ();
 DECAPx1_ASAP7_75t_R FILLER_0_218_35 ();
 FILLER_ASAP7_75t_R FILLER_0_218_45 ();
 FILLER_ASAP7_75t_R FILLER_0_218_53 ();
 FILLER_ASAP7_75t_R FILLER_0_218_62 ();
 FILLER_ASAP7_75t_R FILLER_0_218_71 ();
 FILLER_ASAP7_75t_R FILLER_0_218_83 ();
 FILLER_ASAP7_75t_R FILLER_0_218_95 ();
 FILLER_ASAP7_75t_R FILLER_0_218_107 ();
 FILLER_ASAP7_75t_R FILLER_0_218_119 ();
 FILLER_ASAP7_75t_R FILLER_0_218_131 ();
 FILLER_ASAP7_75t_R FILLER_0_218_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_145 ();
 FILLER_ASAP7_75t_R FILLER_0_218_156 ();
 FILLER_ASAP7_75t_R FILLER_0_218_164 ();
 DECAPx1_ASAP7_75t_R FILLER_0_218_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_175 ();
 DECAPx1_ASAP7_75t_R FILLER_0_218_184 ();
 FILLER_ASAP7_75t_R FILLER_0_218_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_218_221 ();
 DECAPx2_ASAP7_75t_R FILLER_0_218_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_249 ();
 FILLER_ASAP7_75t_R FILLER_0_218_256 ();
 FILLER_ASAP7_75t_R FILLER_0_218_261 ();
 FILLER_ASAP7_75t_R FILLER_0_218_269 ();
 DECAPx2_ASAP7_75t_R FILLER_0_218_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_285 ();
 DECAPx2_ASAP7_75t_R FILLER_0_218_294 ();
 FILLER_ASAP7_75t_R FILLER_0_218_300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_218_305 ();
 DECAPx10_ASAP7_75t_R FILLER_0_218_327 ();
 DECAPx10_ASAP7_75t_R FILLER_0_218_349 ();
 DECAPx2_ASAP7_75t_R FILLER_0_218_371 ();
 FILLER_ASAP7_75t_R FILLER_0_218_377 ();
 DECAPx1_ASAP7_75t_R FILLER_0_218_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_391 ();
 DECAPx6_ASAP7_75t_R FILLER_0_218_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_409 ();
 FILLER_ASAP7_75t_R FILLER_0_218_422 ();
 FILLER_ASAP7_75t_R FILLER_0_218_430 ();
 FILLER_ASAP7_75t_R FILLER_0_218_435 ();
 DECAPx6_ASAP7_75t_R FILLER_0_218_440 ();
 FILLER_ASAP7_75t_R FILLER_0_218_460 ();
 DECAPx2_ASAP7_75t_R FILLER_0_218_464 ();
 FILLER_ASAP7_75t_R FILLER_0_218_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_472 ();
 FILLER_ASAP7_75t_R FILLER_0_218_485 ();
 DECAPx2_ASAP7_75t_R FILLER_0_218_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_505 ();
 DECAPx10_ASAP7_75t_R FILLER_0_218_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_538 ();
 FILLER_ASAP7_75t_R FILLER_0_218_545 ();
 DECAPx2_ASAP7_75t_R FILLER_0_218_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_556 ();
 FILLER_ASAP7_75t_R FILLER_0_218_563 ();
 DECAPx10_ASAP7_75t_R FILLER_0_218_568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_218_590 ();
 DECAPx2_ASAP7_75t_R FILLER_0_218_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_618 ();
 DECAPx2_ASAP7_75t_R FILLER_0_218_626 ();
 DECAPx6_ASAP7_75t_R FILLER_0_218_635 ();
 FILLER_ASAP7_75t_R FILLER_0_218_655 ();
 DECAPx10_ASAP7_75t_R FILLER_0_218_660 ();
 DECAPx1_ASAP7_75t_R FILLER_0_218_682 ();
 DECAPx10_ASAP7_75t_R FILLER_0_218_707 ();
 DECAPx6_ASAP7_75t_R FILLER_0_218_729 ();
 DECAPx2_ASAP7_75t_R FILLER_0_218_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_769 ();
 FILLER_ASAP7_75t_R FILLER_0_218_780 ();
 FILLER_ASAP7_75t_R FILLER_0_218_788 ();
 DECAPx4_ASAP7_75t_R FILLER_0_218_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_218_817 ();
 FILLER_ASAP7_75t_R FILLER_0_218_831 ();
 DECAPx1_ASAP7_75t_R FILLER_0_218_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_843 ();
 FILLER_ASAP7_75t_R FILLER_0_218_850 ();
 DECAPx6_ASAP7_75t_R FILLER_0_218_859 ();
 DECAPx2_ASAP7_75t_R FILLER_0_218_873 ();
 FILLER_ASAP7_75t_R FILLER_0_218_885 ();
 FILLER_ASAP7_75t_R FILLER_0_218_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_895 ();
 FILLER_ASAP7_75t_R FILLER_0_218_902 ();
 DECAPx4_ASAP7_75t_R FILLER_0_218_910 ();
 FILLER_ASAP7_75t_R FILLER_0_218_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_922 ();
 FILLER_ASAP7_75t_R FILLER_0_218_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_931 ();
 DECAPx10_ASAP7_75t_R FILLER_0_218_938 ();
 FILLER_ASAP7_75t_R FILLER_0_218_966 ();
 DECAPx1_ASAP7_75t_R FILLER_0_218_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_978 ();
 DECAPx1_ASAP7_75t_R FILLER_0_218_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_1005 ();
 FILLER_ASAP7_75t_R FILLER_0_218_1028 ();
 FILLER_ASAP7_75t_R FILLER_0_218_1040 ();
 FILLER_ASAP7_75t_R FILLER_0_218_1052 ();
 FILLER_ASAP7_75t_R FILLER_0_218_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_1059 ();
 DECAPx2_ASAP7_75t_R FILLER_0_218_1090 ();
 FILLER_ASAP7_75t_R FILLER_0_218_1096 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_1098 ();
 FILLER_ASAP7_75t_R FILLER_0_218_1102 ();
 FILLER_ASAP7_75t_R FILLER_0_218_1110 ();
 FILLER_ASAP7_75t_R FILLER_0_218_1118 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_1120 ();
 DECAPx2_ASAP7_75t_R FILLER_0_218_1127 ();
 FILLER_ASAP7_75t_R FILLER_0_218_1133 ();
 FILLER_ASAP7_75t_R FILLER_0_218_1147 ();
 DECAPx4_ASAP7_75t_R FILLER_0_218_1152 ();
 FILLER_ASAP7_75t_R FILLER_0_218_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_1164 ();
 FILLER_ASAP7_75t_R FILLER_0_218_1183 ();
 DECAPx4_ASAP7_75t_R FILLER_0_218_1195 ();
 FILLER_ASAP7_75t_R FILLER_0_218_1205 ();
 FILLER_ASAP7_75t_R FILLER_0_218_1212 ();
 FILLER_ASAP7_75t_R FILLER_0_218_1220 ();
 FILLER_ASAP7_75t_R FILLER_0_218_1227 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_1229 ();
 DECAPx10_ASAP7_75t_R FILLER_0_218_1233 ();
 DECAPx10_ASAP7_75t_R FILLER_0_218_1255 ();
 DECAPx10_ASAP7_75t_R FILLER_0_218_1277 ();
 DECAPx10_ASAP7_75t_R FILLER_0_218_1299 ();
 DECAPx10_ASAP7_75t_R FILLER_0_218_1321 ();
 DECAPx10_ASAP7_75t_R FILLER_0_218_1343 ();
 DECAPx6_ASAP7_75t_R FILLER_0_218_1365 ();
 FILLER_ASAP7_75t_R FILLER_0_218_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218_1381 ();
 DECAPx4_ASAP7_75t_R FILLER_0_219_2 ();
 FILLER_ASAP7_75t_R FILLER_0_219_17 ();
 FILLER_ASAP7_75t_R FILLER_0_219_24 ();
 DECAPx1_ASAP7_75t_R FILLER_0_219_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_40 ();
 FILLER_ASAP7_75t_R FILLER_0_219_47 ();
 FILLER_ASAP7_75t_R FILLER_0_219_55 ();
 FILLER_ASAP7_75t_R FILLER_0_219_65 ();
 FILLER_ASAP7_75t_R FILLER_0_219_77 ();
 FILLER_ASAP7_75t_R FILLER_0_219_89 ();
 FILLER_ASAP7_75t_R FILLER_0_219_101 ();
 FILLER_ASAP7_75t_R FILLER_0_219_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_123 ();
 FILLER_ASAP7_75t_R FILLER_0_219_130 ();
 FILLER_ASAP7_75t_R FILLER_0_219_142 ();
 FILLER_ASAP7_75t_R FILLER_0_219_152 ();
 FILLER_ASAP7_75t_R FILLER_0_219_159 ();
 FILLER_ASAP7_75t_R FILLER_0_219_167 ();
 FILLER_ASAP7_75t_R FILLER_0_219_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_177 ();
 FILLER_ASAP7_75t_R FILLER_0_219_184 ();
 FILLER_ASAP7_75t_R FILLER_0_219_192 ();
 FILLER_ASAP7_75t_R FILLER_0_219_202 ();
 DECAPx6_ASAP7_75t_R FILLER_0_219_214 ();
 DECAPx1_ASAP7_75t_R FILLER_0_219_228 ();
 DECAPx1_ASAP7_75t_R FILLER_0_219_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_242 ();
 DECAPx10_ASAP7_75t_R FILLER_0_219_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_271 ();
 DECAPx4_ASAP7_75t_R FILLER_0_219_278 ();
 DECAPx2_ASAP7_75t_R FILLER_0_219_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_297 ();
 FILLER_ASAP7_75t_R FILLER_0_219_304 ();
 FILLER_ASAP7_75t_R FILLER_0_219_312 ();
 DECAPx4_ASAP7_75t_R FILLER_0_219_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_329 ();
 FILLER_ASAP7_75t_R FILLER_0_219_358 ();
 FILLER_ASAP7_75t_R FILLER_0_219_366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_219_376 ();
 FILLER_ASAP7_75t_R FILLER_0_219_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_384 ();
 DECAPx2_ASAP7_75t_R FILLER_0_219_392 ();
 FILLER_ASAP7_75t_R FILLER_0_219_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_400 ();
 FILLER_ASAP7_75t_R FILLER_0_219_425 ();
 FILLER_ASAP7_75t_R FILLER_0_219_435 ();
 DECAPx1_ASAP7_75t_R FILLER_0_219_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_447 ();
 FILLER_ASAP7_75t_R FILLER_0_219_454 ();
 DECAPx2_ASAP7_75t_R FILLER_0_219_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_484 ();
 FILLER_ASAP7_75t_R FILLER_0_219_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_492 ();
 FILLER_ASAP7_75t_R FILLER_0_219_504 ();
 DECAPx10_ASAP7_75t_R FILLER_0_219_514 ();
 FILLER_ASAP7_75t_R FILLER_0_219_536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_219_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_554 ();
 DECAPx2_ASAP7_75t_R FILLER_0_219_561 ();
 DECAPx2_ASAP7_75t_R FILLER_0_219_575 ();
 DECAPx2_ASAP7_75t_R FILLER_0_219_589 ();
 FILLER_ASAP7_75t_R FILLER_0_219_607 ();
 DECAPx6_ASAP7_75t_R FILLER_0_219_621 ();
 DECAPx1_ASAP7_75t_R FILLER_0_219_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_639 ();
 FILLER_ASAP7_75t_R FILLER_0_219_643 ();
 DECAPx4_ASAP7_75t_R FILLER_0_219_653 ();
 FILLER_ASAP7_75t_R FILLER_0_219_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_686 ();
 FILLER_ASAP7_75t_R FILLER_0_219_693 ();
 DECAPx4_ASAP7_75t_R FILLER_0_219_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_708 ();
 FILLER_ASAP7_75t_R FILLER_0_219_712 ();
 DECAPx6_ASAP7_75t_R FILLER_0_219_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_734 ();
 FILLER_ASAP7_75t_R FILLER_0_219_745 ();
 DECAPx10_ASAP7_75t_R FILLER_0_219_753 ();
 DECAPx4_ASAP7_75t_R FILLER_0_219_775 ();
 DECAPx4_ASAP7_75t_R FILLER_0_219_792 ();
 DECAPx1_ASAP7_75t_R FILLER_0_219_822 ();
 DECAPx2_ASAP7_75t_R FILLER_0_219_846 ();
 DECAPx2_ASAP7_75t_R FILLER_0_219_858 ();
 FILLER_ASAP7_75t_R FILLER_0_219_864 ();
 FILLER_ASAP7_75t_R FILLER_0_219_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_874 ();
 DECAPx1_ASAP7_75t_R FILLER_0_219_878 ();
 DECAPx4_ASAP7_75t_R FILLER_0_219_892 ();
 FILLER_ASAP7_75t_R FILLER_0_219_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_904 ();
 DECAPx1_ASAP7_75t_R FILLER_0_219_911 ();
 FILLER_ASAP7_75t_R FILLER_0_219_923 ();
 DECAPx4_ASAP7_75t_R FILLER_0_219_927 ();
 DECAPx2_ASAP7_75t_R FILLER_0_219_940 ();
 FILLER_ASAP7_75t_R FILLER_0_219_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_954 ();
 DECAPx1_ASAP7_75t_R FILLER_0_219_961 ();
 DECAPx2_ASAP7_75t_R FILLER_0_219_973 ();
 FILLER_ASAP7_75t_R FILLER_0_219_979 ();
 DECAPx4_ASAP7_75t_R FILLER_0_219_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_994 ();
 FILLER_ASAP7_75t_R FILLER_0_219_998 ();
 FILLER_ASAP7_75t_R FILLER_0_219_1018 ();
 FILLER_ASAP7_75t_R FILLER_0_219_1025 ();
 FILLER_ASAP7_75t_R FILLER_0_219_1037 ();
 FILLER_ASAP7_75t_R FILLER_0_219_1047 ();
 DECAPx4_ASAP7_75t_R FILLER_0_219_1057 ();
 FILLER_ASAP7_75t_R FILLER_0_219_1067 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_1069 ();
 FILLER_ASAP7_75t_R FILLER_0_219_1073 ();
 FILLER_ASAP7_75t_R FILLER_0_219_1081 ();
 FILLER_ASAP7_75t_R FILLER_0_219_1089 ();
 DECAPx10_ASAP7_75t_R FILLER_0_219_1097 ();
 DECAPx6_ASAP7_75t_R FILLER_0_219_1119 ();
 DECAPx1_ASAP7_75t_R FILLER_0_219_1133 ();
 DECAPx4_ASAP7_75t_R FILLER_0_219_1158 ();
 FILLER_ASAP7_75t_R FILLER_0_219_1173 ();
 DECAPx10_ASAP7_75t_R FILLER_0_219_1183 ();
 DECAPx4_ASAP7_75t_R FILLER_0_219_1205 ();
 FILLER_ASAP7_75t_R FILLER_0_219_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_1217 ();
 DECAPx6_ASAP7_75t_R FILLER_0_219_1221 ();
 DECAPx1_ASAP7_75t_R FILLER_0_219_1235 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_1239 ();
 DECAPx6_ASAP7_75t_R FILLER_0_219_1246 ();
 FILLER_ASAP7_75t_R FILLER_0_219_1266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_219_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_0_219_1301 ();
 DECAPx10_ASAP7_75t_R FILLER_0_219_1323 ();
 DECAPx10_ASAP7_75t_R FILLER_0_219_1345 ();
 DECAPx6_ASAP7_75t_R FILLER_0_219_1367 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219_1381 ();
 DECAPx4_ASAP7_75t_R FILLER_0_220_2 ();
 FILLER_ASAP7_75t_R FILLER_0_220_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_14 ();
 DECAPx1_ASAP7_75t_R FILLER_0_220_21 ();
 FILLER_ASAP7_75t_R FILLER_0_220_31 ();
 FILLER_ASAP7_75t_R FILLER_0_220_39 ();
 DECAPx2_ASAP7_75t_R FILLER_0_220_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_55 ();
 FILLER_ASAP7_75t_R FILLER_0_220_63 ();
 FILLER_ASAP7_75t_R FILLER_0_220_71 ();
 FILLER_ASAP7_75t_R FILLER_0_220_83 ();
 FILLER_ASAP7_75t_R FILLER_0_220_95 ();
 FILLER_ASAP7_75t_R FILLER_0_220_107 ();
 FILLER_ASAP7_75t_R FILLER_0_220_119 ();
 FILLER_ASAP7_75t_R FILLER_0_220_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_133 ();
 DECAPx1_ASAP7_75t_R FILLER_0_220_144 ();
 FILLER_ASAP7_75t_R FILLER_0_220_154 ();
 FILLER_ASAP7_75t_R FILLER_0_220_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_169 ();
 FILLER_ASAP7_75t_R FILLER_0_220_176 ();
 FILLER_ASAP7_75t_R FILLER_0_220_184 ();
 FILLER_ASAP7_75t_R FILLER_0_220_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_194 ();
 DECAPx2_ASAP7_75t_R FILLER_0_220_201 ();
 FILLER_ASAP7_75t_R FILLER_0_220_207 ();
 DECAPx6_ASAP7_75t_R FILLER_0_220_216 ();
 DECAPx2_ASAP7_75t_R FILLER_0_220_230 ();
 DECAPx1_ASAP7_75t_R FILLER_0_220_239 ();
 FILLER_ASAP7_75t_R FILLER_0_220_250 ();
 DECAPx1_ASAP7_75t_R FILLER_0_220_258 ();
 FILLER_ASAP7_75t_R FILLER_0_220_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_270 ();
 FILLER_ASAP7_75t_R FILLER_0_220_277 ();
 FILLER_ASAP7_75t_R FILLER_0_220_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_301 ();
 FILLER_ASAP7_75t_R FILLER_0_220_309 ();
 DECAPx2_ASAP7_75t_R FILLER_0_220_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_323 ();
 DECAPx2_ASAP7_75t_R FILLER_0_220_334 ();
 FILLER_ASAP7_75t_R FILLER_0_220_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_342 ();
 FILLER_ASAP7_75t_R FILLER_0_220_349 ();
 FILLER_ASAP7_75t_R FILLER_0_220_357 ();
 DECAPx2_ASAP7_75t_R FILLER_0_220_366 ();
 FILLER_ASAP7_75t_R FILLER_0_220_372 ();
 FILLER_ASAP7_75t_R FILLER_0_220_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_382 ();
 FILLER_ASAP7_75t_R FILLER_0_220_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_391 ();
 FILLER_ASAP7_75t_R FILLER_0_220_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_400 ();
 DECAPx6_ASAP7_75t_R FILLER_0_220_407 ();
 FILLER_ASAP7_75t_R FILLER_0_220_421 ();
 DECAPx6_ASAP7_75t_R FILLER_0_220_429 ();
 DECAPx1_ASAP7_75t_R FILLER_0_220_443 ();
 DECAPx1_ASAP7_75t_R FILLER_0_220_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_461 ();
 FILLER_ASAP7_75t_R FILLER_0_220_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_466 ();
 DECAPx4_ASAP7_75t_R FILLER_0_220_488 ();
 FILLER_ASAP7_75t_R FILLER_0_220_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_500 ();
 FILLER_ASAP7_75t_R FILLER_0_220_504 ();
 FILLER_ASAP7_75t_R FILLER_0_220_512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_220_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_544 ();
 FILLER_ASAP7_75t_R FILLER_0_220_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_555 ();
 FILLER_ASAP7_75t_R FILLER_0_220_562 ();
 DECAPx2_ASAP7_75t_R FILLER_0_220_572 ();
 FILLER_ASAP7_75t_R FILLER_0_220_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_580 ();
 DECAPx2_ASAP7_75t_R FILLER_0_220_602 ();
 DECAPx2_ASAP7_75t_R FILLER_0_220_620 ();
 FILLER_ASAP7_75t_R FILLER_0_220_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_628 ();
 DECAPx4_ASAP7_75t_R FILLER_0_220_634 ();
 DECAPx4_ASAP7_75t_R FILLER_0_220_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_665 ();
 FILLER_ASAP7_75t_R FILLER_0_220_672 ();
 DECAPx6_ASAP7_75t_R FILLER_0_220_677 ();
 FILLER_ASAP7_75t_R FILLER_0_220_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_693 ();
 DECAPx2_ASAP7_75t_R FILLER_0_220_704 ();
 DECAPx6_ASAP7_75t_R FILLER_0_220_716 ();
 FILLER_ASAP7_75t_R FILLER_0_220_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_220_753 ();
 DECAPx2_ASAP7_75t_R FILLER_0_220_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_781 ();
 FILLER_ASAP7_75t_R FILLER_0_220_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_790 ();
 DECAPx6_ASAP7_75t_R FILLER_0_220_797 ();
 DECAPx1_ASAP7_75t_R FILLER_0_220_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_815 ();
 DECAPx2_ASAP7_75t_R FILLER_0_220_822 ();
 FILLER_ASAP7_75t_R FILLER_0_220_828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_220_840 ();
 DECAPx2_ASAP7_75t_R FILLER_0_220_862 ();
 FILLER_ASAP7_75t_R FILLER_0_220_868 ();
 DECAPx6_ASAP7_75t_R FILLER_0_220_875 ();
 DECAPx1_ASAP7_75t_R FILLER_0_220_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_893 ();
 DECAPx1_ASAP7_75t_R FILLER_0_220_900 ();
 DECAPx1_ASAP7_75t_R FILLER_0_220_910 ();
 DECAPx2_ASAP7_75t_R FILLER_0_220_925 ();
 FILLER_ASAP7_75t_R FILLER_0_220_937 ();
 FILLER_ASAP7_75t_R FILLER_0_220_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_952 ();
 DECAPx6_ASAP7_75t_R FILLER_0_220_974 ();
 FILLER_ASAP7_75t_R FILLER_0_220_988 ();
 FILLER_ASAP7_75t_R FILLER_0_220_996 ();
 FILLER_ASAP7_75t_R FILLER_0_220_1001 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_1003 ();
 FILLER_ASAP7_75t_R FILLER_0_220_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_1012 ();
 FILLER_ASAP7_75t_R FILLER_0_220_1019 ();
 FILLER_ASAP7_75t_R FILLER_0_220_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_1029 ();
 DECAPx1_ASAP7_75t_R FILLER_0_220_1036 ();
 DECAPx2_ASAP7_75t_R FILLER_0_220_1048 ();
 DECAPx2_ASAP7_75t_R FILLER_0_220_1075 ();
 FILLER_ASAP7_75t_R FILLER_0_220_1081 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_1083 ();
 DECAPx10_ASAP7_75t_R FILLER_0_220_1096 ();
 FILLER_ASAP7_75t_R FILLER_0_220_1118 ();
 FILLER_ASAP7_75t_R FILLER_0_220_1142 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_1144 ();
 FILLER_ASAP7_75t_R FILLER_0_220_1149 ();
 DECAPx1_ASAP7_75t_R FILLER_0_220_1156 ();
 FILLER_ASAP7_75t_R FILLER_0_220_1170 ();
 FILLER_ASAP7_75t_R FILLER_0_220_1182 ();
 FILLER_ASAP7_75t_R FILLER_0_220_1190 ();
 DECAPx4_ASAP7_75t_R FILLER_0_220_1198 ();
 FILLER_ASAP7_75t_R FILLER_0_220_1208 ();
 FILLER_ASAP7_75t_R FILLER_0_220_1216 ();
 FILLER_ASAP7_75t_R FILLER_0_220_1224 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_1226 ();
 DECAPx1_ASAP7_75t_R FILLER_0_220_1233 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_1237 ();
 DECAPx2_ASAP7_75t_R FILLER_0_220_1244 ();
 FILLER_ASAP7_75t_R FILLER_0_220_1250 ();
 FILLER_ASAP7_75t_R FILLER_0_220_1263 ();
 FILLER_ASAP7_75t_R FILLER_0_220_1271 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220_1273 ();
 DECAPx4_ASAP7_75t_R FILLER_0_220_1280 ();
 DECAPx4_ASAP7_75t_R FILLER_0_220_1296 ();
 DECAPx10_ASAP7_75t_R FILLER_0_220_1312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_220_1334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_220_1356 ();
 DECAPx1_ASAP7_75t_R FILLER_0_220_1378 ();
 DECAPx1_ASAP7_75t_R FILLER_0_221_2 ();
 FILLER_ASAP7_75t_R FILLER_0_221_12 ();
 DECAPx2_ASAP7_75t_R FILLER_0_221_24 ();
 DECAPx2_ASAP7_75t_R FILLER_0_221_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_56 ();
 DECAPx2_ASAP7_75t_R FILLER_0_221_67 ();
 FILLER_ASAP7_75t_R FILLER_0_221_83 ();
 FILLER_ASAP7_75t_R FILLER_0_221_95 ();
 FILLER_ASAP7_75t_R FILLER_0_221_107 ();
 FILLER_ASAP7_75t_R FILLER_0_221_119 ();
 DECAPx2_ASAP7_75t_R FILLER_0_221_131 ();
 DECAPx1_ASAP7_75t_R FILLER_0_221_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_151 ();
 FILLER_ASAP7_75t_R FILLER_0_221_158 ();
 FILLER_ASAP7_75t_R FILLER_0_221_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_168 ();
 DECAPx1_ASAP7_75t_R FILLER_0_221_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_179 ();
 FILLER_ASAP7_75t_R FILLER_0_221_188 ();
 DECAPx6_ASAP7_75t_R FILLER_0_221_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_207 ();
 DECAPx10_ASAP7_75t_R FILLER_0_221_213 ();
 DECAPx2_ASAP7_75t_R FILLER_0_221_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_241 ();
 FILLER_ASAP7_75t_R FILLER_0_221_250 ();
 DECAPx1_ASAP7_75t_R FILLER_0_221_258 ();
 FILLER_ASAP7_75t_R FILLER_0_221_265 ();
 FILLER_ASAP7_75t_R FILLER_0_221_273 ();
 FILLER_ASAP7_75t_R FILLER_0_221_282 ();
 DECAPx1_ASAP7_75t_R FILLER_0_221_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_294 ();
 DECAPx2_ASAP7_75t_R FILLER_0_221_301 ();
 FILLER_ASAP7_75t_R FILLER_0_221_307 ();
 DECAPx10_ASAP7_75t_R FILLER_0_221_317 ();
 FILLER_ASAP7_75t_R FILLER_0_221_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_341 ();
 DECAPx2_ASAP7_75t_R FILLER_0_221_348 ();
 FILLER_ASAP7_75t_R FILLER_0_221_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_362 ();
 DECAPx2_ASAP7_75t_R FILLER_0_221_369 ();
 FILLER_ASAP7_75t_R FILLER_0_221_375 ();
 FILLER_ASAP7_75t_R FILLER_0_221_383 ();
 FILLER_ASAP7_75t_R FILLER_0_221_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_390 ();
 FILLER_ASAP7_75t_R FILLER_0_221_397 ();
 DECAPx10_ASAP7_75t_R FILLER_0_221_405 ();
 FILLER_ASAP7_75t_R FILLER_0_221_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_429 ();
 FILLER_ASAP7_75t_R FILLER_0_221_433 ();
 DECAPx4_ASAP7_75t_R FILLER_0_221_441 ();
 FILLER_ASAP7_75t_R FILLER_0_221_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_453 ();
 FILLER_ASAP7_75t_R FILLER_0_221_457 ();
 FILLER_ASAP7_75t_R FILLER_0_221_462 ();
 DECAPx2_ASAP7_75t_R FILLER_0_221_470 ();
 FILLER_ASAP7_75t_R FILLER_0_221_488 ();
 FILLER_ASAP7_75t_R FILLER_0_221_495 ();
 DECAPx2_ASAP7_75t_R FILLER_0_221_509 ();
 FILLER_ASAP7_75t_R FILLER_0_221_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_517 ();
 DECAPx2_ASAP7_75t_R FILLER_0_221_539 ();
 DECAPx4_ASAP7_75t_R FILLER_0_221_551 ();
 FILLER_ASAP7_75t_R FILLER_0_221_561 ();
 DECAPx10_ASAP7_75t_R FILLER_0_221_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_595 ();
 FILLER_ASAP7_75t_R FILLER_0_221_599 ();
 FILLER_ASAP7_75t_R FILLER_0_221_613 ();
 DECAPx10_ASAP7_75t_R FILLER_0_221_621 ();
 DECAPx2_ASAP7_75t_R FILLER_0_221_643 ();
 FILLER_ASAP7_75t_R FILLER_0_221_649 ();
 DECAPx10_ASAP7_75t_R FILLER_0_221_654 ();
 DECAPx4_ASAP7_75t_R FILLER_0_221_676 ();
 DECAPx4_ASAP7_75t_R FILLER_0_221_690 ();
 FILLER_ASAP7_75t_R FILLER_0_221_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_702 ();
 FILLER_ASAP7_75t_R FILLER_0_221_723 ();
 FILLER_ASAP7_75t_R FILLER_0_221_731 ();
 FILLER_ASAP7_75t_R FILLER_0_221_739 ();
 DECAPx1_ASAP7_75t_R FILLER_0_221_747 ();
 FILLER_ASAP7_75t_R FILLER_0_221_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_759 ();
 DECAPx1_ASAP7_75t_R FILLER_0_221_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_770 ();
 DECAPx1_ASAP7_75t_R FILLER_0_221_777 ();
 DECAPx1_ASAP7_75t_R FILLER_0_221_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_791 ();
 FILLER_ASAP7_75t_R FILLER_0_221_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_800 ();
 DECAPx1_ASAP7_75t_R FILLER_0_221_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_812 ();
 DECAPx2_ASAP7_75t_R FILLER_0_221_819 ();
 FILLER_ASAP7_75t_R FILLER_0_221_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_827 ();
 FILLER_ASAP7_75t_R FILLER_0_221_838 ();
 FILLER_ASAP7_75t_R FILLER_0_221_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_848 ();
 FILLER_ASAP7_75t_R FILLER_0_221_855 ();
 FILLER_ASAP7_75t_R FILLER_0_221_863 ();
 FILLER_ASAP7_75t_R FILLER_0_221_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_873 ();
 FILLER_ASAP7_75t_R FILLER_0_221_880 ();
 FILLER_ASAP7_75t_R FILLER_0_221_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_891 ();
 FILLER_ASAP7_75t_R FILLER_0_221_898 ();
 DECAPx6_ASAP7_75t_R FILLER_0_221_906 ();
 DECAPx1_ASAP7_75t_R FILLER_0_221_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_924 ();
 DECAPx10_ASAP7_75t_R FILLER_0_221_927 ();
 DECAPx1_ASAP7_75t_R FILLER_0_221_949 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_953 ();
 FILLER_ASAP7_75t_R FILLER_0_221_957 ();
 DECAPx10_ASAP7_75t_R FILLER_0_221_965 ();
 FILLER_ASAP7_75t_R FILLER_0_221_993 ();
 DECAPx1_ASAP7_75t_R FILLER_0_221_998 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_1002 ();
 DECAPx10_ASAP7_75t_R FILLER_0_221_1009 ();
 DECAPx2_ASAP7_75t_R FILLER_0_221_1031 ();
 DECAPx1_ASAP7_75t_R FILLER_0_221_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_1045 ();
 FILLER_ASAP7_75t_R FILLER_0_221_1052 ();
 FILLER_ASAP7_75t_R FILLER_0_221_1057 ();
 DECAPx2_ASAP7_75t_R FILLER_0_221_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_1068 ();
 FILLER_ASAP7_75t_R FILLER_0_221_1072 ();
 DECAPx4_ASAP7_75t_R FILLER_0_221_1084 ();
 FILLER_ASAP7_75t_R FILLER_0_221_1094 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_1096 ();
 FILLER_ASAP7_75t_R FILLER_0_221_1119 ();
 FILLER_ASAP7_75t_R FILLER_0_221_1142 ();
 DECAPx1_ASAP7_75t_R FILLER_0_221_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_1158 ();
 FILLER_ASAP7_75t_R FILLER_0_221_1169 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_1171 ();
 FILLER_ASAP7_75t_R FILLER_0_221_1210 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_1212 ();
 DECAPx1_ASAP7_75t_R FILLER_0_221_1225 ();
 FILLER_ASAP7_75t_R FILLER_0_221_1241 ();
 DECAPx4_ASAP7_75t_R FILLER_0_221_1246 ();
 FILLER_ASAP7_75t_R FILLER_0_221_1268 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_1270 ();
 DECAPx1_ASAP7_75t_R FILLER_0_221_1279 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_1283 ();
 DECAPx4_ASAP7_75t_R FILLER_0_221_1296 ();
 DECAPx1_ASAP7_75t_R FILLER_0_221_1316 ();
 FILLER_ASAP7_75t_R FILLER_0_221_1330 ();
 DECAPx2_ASAP7_75t_R FILLER_0_221_1337 ();
 FILLER_ASAP7_75t_R FILLER_0_221_1343 ();
 DECAPx2_ASAP7_75t_R FILLER_0_221_1351 ();
 FILLER_ASAP7_75t_R FILLER_0_221_1357 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_1359 ();
 DECAPx6_ASAP7_75t_R FILLER_0_221_1363 ();
 DECAPx1_ASAP7_75t_R FILLER_0_221_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221_1381 ();
 DECAPx4_ASAP7_75t_R FILLER_0_222_2 ();
 FILLER_ASAP7_75t_R FILLER_0_222_20 ();
 FILLER_ASAP7_75t_R FILLER_0_222_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_27 ();
 DECAPx1_ASAP7_75t_R FILLER_0_222_48 ();
 FILLER_ASAP7_75t_R FILLER_0_222_63 ();
 FILLER_ASAP7_75t_R FILLER_0_222_71 ();
 FILLER_ASAP7_75t_R FILLER_0_222_83 ();
 FILLER_ASAP7_75t_R FILLER_0_222_95 ();
 FILLER_ASAP7_75t_R FILLER_0_222_107 ();
 FILLER_ASAP7_75t_R FILLER_0_222_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_121 ();
 DECAPx2_ASAP7_75t_R FILLER_0_222_132 ();
 DECAPx2_ASAP7_75t_R FILLER_0_222_144 ();
 FILLER_ASAP7_75t_R FILLER_0_222_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_163 ();
 FILLER_ASAP7_75t_R FILLER_0_222_170 ();
 FILLER_ASAP7_75t_R FILLER_0_222_178 ();
 DECAPx6_ASAP7_75t_R FILLER_0_222_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_200 ();
 FILLER_ASAP7_75t_R FILLER_0_222_211 ();
 FILLER_ASAP7_75t_R FILLER_0_222_223 ();
 DECAPx10_ASAP7_75t_R FILLER_0_222_228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_222_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_272 ();
 DECAPx1_ASAP7_75t_R FILLER_0_222_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_283 ();
 DECAPx2_ASAP7_75t_R FILLER_0_222_290 ();
 FILLER_ASAP7_75t_R FILLER_0_222_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_298 ();
 FILLER_ASAP7_75t_R FILLER_0_222_305 ();
 FILLER_ASAP7_75t_R FILLER_0_222_313 ();
 DECAPx4_ASAP7_75t_R FILLER_0_222_335 ();
 FILLER_ASAP7_75t_R FILLER_0_222_351 ();
 DECAPx4_ASAP7_75t_R FILLER_0_222_361 ();
 FILLER_ASAP7_75t_R FILLER_0_222_371 ();
 DECAPx1_ASAP7_75t_R FILLER_0_222_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_385 ();
 DECAPx6_ASAP7_75t_R FILLER_0_222_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_403 ();
 FILLER_ASAP7_75t_R FILLER_0_222_410 ();
 DECAPx2_ASAP7_75t_R FILLER_0_222_415 ();
 FILLER_ASAP7_75t_R FILLER_0_222_427 ();
 FILLER_ASAP7_75t_R FILLER_0_222_437 ();
 DECAPx6_ASAP7_75t_R FILLER_0_222_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_222_456 ();
 FILLER_ASAP7_75t_R FILLER_0_222_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_466 ();
 DECAPx4_ASAP7_75t_R FILLER_0_222_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_498 ();
 DECAPx4_ASAP7_75t_R FILLER_0_222_511 ();
 FILLER_ASAP7_75t_R FILLER_0_222_527 ();
 DECAPx10_ASAP7_75t_R FILLER_0_222_532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_222_554 ();
 DECAPx2_ASAP7_75t_R FILLER_0_222_576 ();
 FILLER_ASAP7_75t_R FILLER_0_222_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_584 ();
 FILLER_ASAP7_75t_R FILLER_0_222_597 ();
 DECAPx2_ASAP7_75t_R FILLER_0_222_610 ();
 DECAPx2_ASAP7_75t_R FILLER_0_222_637 ();
 FILLER_ASAP7_75t_R FILLER_0_222_643 ();
 FILLER_ASAP7_75t_R FILLER_0_222_655 ();
 FILLER_ASAP7_75t_R FILLER_0_222_678 ();
 FILLER_ASAP7_75t_R FILLER_0_222_692 ();
 DECAPx10_ASAP7_75t_R FILLER_0_222_700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_222_722 ();
 DECAPx2_ASAP7_75t_R FILLER_0_222_744 ();
 FILLER_ASAP7_75t_R FILLER_0_222_750 ();
 DECAPx2_ASAP7_75t_R FILLER_0_222_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_222_771 ();
 DECAPx1_ASAP7_75t_R FILLER_0_222_793 ();
 FILLER_ASAP7_75t_R FILLER_0_222_803 ();
 DECAPx2_ASAP7_75t_R FILLER_0_222_812 ();
 FILLER_ASAP7_75t_R FILLER_0_222_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_827 ();
 DECAPx2_ASAP7_75t_R FILLER_0_222_848 ();
 FILLER_ASAP7_75t_R FILLER_0_222_854 ();
 FILLER_ASAP7_75t_R FILLER_0_222_867 ();
 FILLER_ASAP7_75t_R FILLER_0_222_875 ();
 DECAPx10_ASAP7_75t_R FILLER_0_222_883 ();
 DECAPx4_ASAP7_75t_R FILLER_0_222_905 ();
 FILLER_ASAP7_75t_R FILLER_0_222_915 ();
 DECAPx2_ASAP7_75t_R FILLER_0_222_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_929 ();
 DECAPx2_ASAP7_75t_R FILLER_0_222_942 ();
 FILLER_ASAP7_75t_R FILLER_0_222_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_950 ();
 FILLER_ASAP7_75t_R FILLER_0_222_954 ();
 FILLER_ASAP7_75t_R FILLER_0_222_967 ();
 DECAPx6_ASAP7_75t_R FILLER_0_222_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_989 ();
 DECAPx4_ASAP7_75t_R FILLER_0_222_996 ();
 DECAPx2_ASAP7_75t_R FILLER_0_222_1012 ();
 FILLER_ASAP7_75t_R FILLER_0_222_1024 ();
 FILLER_ASAP7_75t_R FILLER_0_222_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_1031 ();
 FILLER_ASAP7_75t_R FILLER_0_222_1042 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_1044 ();
 DECAPx4_ASAP7_75t_R FILLER_0_222_1051 ();
 FILLER_ASAP7_75t_R FILLER_0_222_1061 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_1063 ();
 FILLER_ASAP7_75t_R FILLER_0_222_1070 ();
 DECAPx4_ASAP7_75t_R FILLER_0_222_1078 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_1088 ();
 FILLER_ASAP7_75t_R FILLER_0_222_1110 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_1112 ();
 FILLER_ASAP7_75t_R FILLER_0_222_1116 ();
 FILLER_ASAP7_75t_R FILLER_0_222_1136 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_1138 ();
 FILLER_ASAP7_75t_R FILLER_0_222_1144 ();
 FILLER_ASAP7_75t_R FILLER_0_222_1156 ();
 FILLER_ASAP7_75t_R FILLER_0_222_1168 ();
 FILLER_ASAP7_75t_R FILLER_0_222_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_1179 ();
 FILLER_ASAP7_75t_R FILLER_0_222_1198 ();
 DECAPx1_ASAP7_75t_R FILLER_0_222_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_1210 ();
 FILLER_ASAP7_75t_R FILLER_0_222_1222 ();
 FILLER_ASAP7_75t_R FILLER_0_222_1230 ();
 DECAPx4_ASAP7_75t_R FILLER_0_222_1238 ();
 FILLER_ASAP7_75t_R FILLER_0_222_1248 ();
 FILLER_ASAP7_75t_R FILLER_0_222_1256 ();
 DECAPx4_ASAP7_75t_R FILLER_0_222_1264 ();
 DECAPx1_ASAP7_75t_R FILLER_0_222_1280 ();
 FILLER_ASAP7_75t_R FILLER_0_222_1289 ();
 FILLER_ASAP7_75t_R FILLER_0_222_1321 ();
 DECAPx4_ASAP7_75t_R FILLER_0_222_1335 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_1345 ();
 FILLER_ASAP7_75t_R FILLER_0_222_1353 ();
 FILLER_ASAP7_75t_R FILLER_0_222_1361 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222_1363 ();
 FILLER_ASAP7_75t_R FILLER_0_222_1371 ();
 DECAPx1_ASAP7_75t_R FILLER_0_222_1378 ();
 DECAPx4_ASAP7_75t_R FILLER_0_223_2 ();
 FILLER_ASAP7_75t_R FILLER_0_223_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_14 ();
 DECAPx4_ASAP7_75t_R FILLER_0_223_23 ();
 FILLER_ASAP7_75t_R FILLER_0_223_43 ();
 FILLER_ASAP7_75t_R FILLER_0_223_50 ();
 FILLER_ASAP7_75t_R FILLER_0_223_58 ();
 FILLER_ASAP7_75t_R FILLER_0_223_66 ();
 FILLER_ASAP7_75t_R FILLER_0_223_78 ();
 FILLER_ASAP7_75t_R FILLER_0_223_90 ();
 FILLER_ASAP7_75t_R FILLER_0_223_102 ();
 DECAPx2_ASAP7_75t_R FILLER_0_223_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_120 ();
 FILLER_ASAP7_75t_R FILLER_0_223_127 ();
 FILLER_ASAP7_75t_R FILLER_0_223_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_137 ();
 FILLER_ASAP7_75t_R FILLER_0_223_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_146 ();
 FILLER_ASAP7_75t_R FILLER_0_223_153 ();
 FILLER_ASAP7_75t_R FILLER_0_223_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_162 ();
 FILLER_ASAP7_75t_R FILLER_0_223_169 ();
 FILLER_ASAP7_75t_R FILLER_0_223_181 ();
 FILLER_ASAP7_75t_R FILLER_0_223_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_192 ();
 FILLER_ASAP7_75t_R FILLER_0_223_203 ();
 FILLER_ASAP7_75t_R FILLER_0_223_215 ();
 DECAPx6_ASAP7_75t_R FILLER_0_223_227 ();
 DECAPx2_ASAP7_75t_R FILLER_0_223_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_247 ();
 DECAPx6_ASAP7_75t_R FILLER_0_223_251 ();
 DECAPx6_ASAP7_75t_R FILLER_0_223_271 ();
 DECAPx1_ASAP7_75t_R FILLER_0_223_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_289 ();
 FILLER_ASAP7_75t_R FILLER_0_223_296 ();
 FILLER_ASAP7_75t_R FILLER_0_223_306 ();
 FILLER_ASAP7_75t_R FILLER_0_223_314 ();
 FILLER_ASAP7_75t_R FILLER_0_223_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_324 ();
 FILLER_ASAP7_75t_R FILLER_0_223_328 ();
 DECAPx6_ASAP7_75t_R FILLER_0_223_358 ();
 DECAPx1_ASAP7_75t_R FILLER_0_223_378 ();
 DECAPx4_ASAP7_75t_R FILLER_0_223_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_400 ();
 FILLER_ASAP7_75t_R FILLER_0_223_404 ();
 DECAPx1_ASAP7_75t_R FILLER_0_223_412 ();
 FILLER_ASAP7_75t_R FILLER_0_223_426 ();
 FILLER_ASAP7_75t_R FILLER_0_223_431 ();
 FILLER_ASAP7_75t_R FILLER_0_223_436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_223_444 ();
 FILLER_ASAP7_75t_R FILLER_0_223_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_468 ();
 DECAPx2_ASAP7_75t_R FILLER_0_223_472 ();
 DECAPx10_ASAP7_75t_R FILLER_0_223_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_512 ();
 DECAPx6_ASAP7_75t_R FILLER_0_223_525 ();
 FILLER_ASAP7_75t_R FILLER_0_223_547 ();
 DECAPx4_ASAP7_75t_R FILLER_0_223_555 ();
 FILLER_ASAP7_75t_R FILLER_0_223_565 ();
 FILLER_ASAP7_75t_R FILLER_0_223_588 ();
 DECAPx2_ASAP7_75t_R FILLER_0_223_596 ();
 FILLER_ASAP7_75t_R FILLER_0_223_602 ();
 DECAPx2_ASAP7_75t_R FILLER_0_223_608 ();
 FILLER_ASAP7_75t_R FILLER_0_223_614 ();
 DECAPx4_ASAP7_75t_R FILLER_0_223_622 ();
 FILLER_ASAP7_75t_R FILLER_0_223_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_634 ();
 FILLER_ASAP7_75t_R FILLER_0_223_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_640 ();
 FILLER_ASAP7_75t_R FILLER_0_223_661 ();
 DECAPx1_ASAP7_75t_R FILLER_0_223_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_673 ();
 DECAPx2_ASAP7_75t_R FILLER_0_223_686 ();
 FILLER_ASAP7_75t_R FILLER_0_223_692 ();
 DECAPx1_ASAP7_75t_R FILLER_0_223_702 ();
 FILLER_ASAP7_75t_R FILLER_0_223_718 ();
 FILLER_ASAP7_75t_R FILLER_0_223_731 ();
 DECAPx4_ASAP7_75t_R FILLER_0_223_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_754 ();
 DECAPx2_ASAP7_75t_R FILLER_0_223_766 ();
 FILLER_ASAP7_75t_R FILLER_0_223_772 ();
 DECAPx4_ASAP7_75t_R FILLER_0_223_780 ();
 FILLER_ASAP7_75t_R FILLER_0_223_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_792 ();
 FILLER_ASAP7_75t_R FILLER_0_223_798 ();
 DECAPx1_ASAP7_75t_R FILLER_0_223_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_815 ();
 DECAPx2_ASAP7_75t_R FILLER_0_223_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_223_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_842 ();
 DECAPx2_ASAP7_75t_R FILLER_0_223_849 ();
 DECAPx6_ASAP7_75t_R FILLER_0_223_861 ();
 DECAPx1_ASAP7_75t_R FILLER_0_223_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_879 ();
 FILLER_ASAP7_75t_R FILLER_0_223_886 ();
 FILLER_ASAP7_75t_R FILLER_0_223_894 ();
 DECAPx4_ASAP7_75t_R FILLER_0_223_899 ();
 FILLER_ASAP7_75t_R FILLER_0_223_912 ();
 FILLER_ASAP7_75t_R FILLER_0_223_917 ();
 FILLER_ASAP7_75t_R FILLER_0_223_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_924 ();
 DECAPx1_ASAP7_75t_R FILLER_0_223_927 ();
 DECAPx10_ASAP7_75t_R FILLER_0_223_952 ();
 FILLER_ASAP7_75t_R FILLER_0_223_974 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_976 ();
 DECAPx10_ASAP7_75t_R FILLER_0_223_987 ();
 DECAPx10_ASAP7_75t_R FILLER_0_223_1009 ();
 DECAPx4_ASAP7_75t_R FILLER_0_223_1031 ();
 FILLER_ASAP7_75t_R FILLER_0_223_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_1043 ();
 DECAPx1_ASAP7_75t_R FILLER_0_223_1047 ();
 DECAPx4_ASAP7_75t_R FILLER_0_223_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_1067 ();
 DECAPx4_ASAP7_75t_R FILLER_0_223_1071 ();
 FILLER_ASAP7_75t_R FILLER_0_223_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_1086 ();
 FILLER_ASAP7_75t_R FILLER_0_223_1093 ();
 FILLER_ASAP7_75t_R FILLER_0_223_1098 ();
 DECAPx6_ASAP7_75t_R FILLER_0_223_1103 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_1117 ();
 DECAPx2_ASAP7_75t_R FILLER_0_223_1128 ();
 DECAPx1_ASAP7_75t_R FILLER_0_223_1140 ();
 FILLER_ASAP7_75t_R FILLER_0_223_1152 ();
 DECAPx2_ASAP7_75t_R FILLER_0_223_1172 ();
 FILLER_ASAP7_75t_R FILLER_0_223_1178 ();
 DECAPx1_ASAP7_75t_R FILLER_0_223_1190 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_1194 ();
 FILLER_ASAP7_75t_R FILLER_0_223_1205 ();
 FILLER_ASAP7_75t_R FILLER_0_223_1225 ();
 FILLER_ASAP7_75t_R FILLER_0_223_1233 ();
 DECAPx2_ASAP7_75t_R FILLER_0_223_1241 ();
 FILLER_ASAP7_75t_R FILLER_0_223_1253 ();
 FILLER_ASAP7_75t_R FILLER_0_223_1260 ();
 DECAPx1_ASAP7_75t_R FILLER_0_223_1267 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_1271 ();
 FILLER_ASAP7_75t_R FILLER_0_223_1278 ();
 FILLER_ASAP7_75t_R FILLER_0_223_1286 ();
 DECAPx2_ASAP7_75t_R FILLER_0_223_1295 ();
 FILLER_ASAP7_75t_R FILLER_0_223_1306 ();
 DECAPx2_ASAP7_75t_R FILLER_0_223_1318 ();
 FILLER_ASAP7_75t_R FILLER_0_223_1324 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_1326 ();
 FILLER_ASAP7_75t_R FILLER_0_223_1335 ();
 DECAPx1_ASAP7_75t_R FILLER_0_223_1343 ();
 DECAPx1_ASAP7_75t_R FILLER_0_223_1357 ();
 DECAPx4_ASAP7_75t_R FILLER_0_223_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223_1381 ();
 DECAPx4_ASAP7_75t_R FILLER_0_224_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224_12 ();
 FILLER_ASAP7_75t_R FILLER_0_224_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224_21 ();
 FILLER_ASAP7_75t_R FILLER_0_224_28 ();
 FILLER_ASAP7_75t_R FILLER_0_224_36 ();
 FILLER_ASAP7_75t_R FILLER_0_224_44 ();
 FILLER_ASAP7_75t_R FILLER_0_224_52 ();
 FILLER_ASAP7_75t_R FILLER_0_224_60 ();
 FILLER_ASAP7_75t_R FILLER_0_224_68 ();
 FILLER_ASAP7_75t_R FILLER_0_224_76 ();
 DECAPx1_ASAP7_75t_R FILLER_0_224_86 ();
 FILLER_ASAP7_75t_R FILLER_0_224_96 ();
 DECAPx2_ASAP7_75t_R FILLER_0_224_108 ();
 FILLER_ASAP7_75t_R FILLER_0_224_120 ();
 DECAPx1_ASAP7_75t_R FILLER_0_224_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224_132 ();
 FILLER_ASAP7_75t_R FILLER_0_224_140 ();
 FILLER_ASAP7_75t_R FILLER_0_224_148 ();
 FILLER_ASAP7_75t_R FILLER_0_224_155 ();
 FILLER_ASAP7_75t_R FILLER_0_224_162 ();
 DECAPx1_ASAP7_75t_R FILLER_0_224_167 ();
 DECAPx2_ASAP7_75t_R FILLER_0_224_179 ();
 FILLER_ASAP7_75t_R FILLER_0_224_185 ();
 DECAPx4_ASAP7_75t_R FILLER_0_224_193 ();
 DECAPx2_ASAP7_75t_R FILLER_0_224_213 ();
 FILLER_ASAP7_75t_R FILLER_0_224_225 ();
 DECAPx6_ASAP7_75t_R FILLER_0_224_230 ();
 DECAPx2_ASAP7_75t_R FILLER_0_224_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224_250 ();
 DECAPx1_ASAP7_75t_R FILLER_0_224_261 ();
 FILLER_ASAP7_75t_R FILLER_0_224_273 ();
 FILLER_ASAP7_75t_R FILLER_0_224_283 ();
 FILLER_ASAP7_75t_R FILLER_0_224_293 ();
 DECAPx10_ASAP7_75t_R FILLER_0_224_301 ();
 DECAPx4_ASAP7_75t_R FILLER_0_224_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224_333 ();
 DECAPx2_ASAP7_75t_R FILLER_0_224_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224_345 ();
 FILLER_ASAP7_75t_R FILLER_0_224_352 ();
 FILLER_ASAP7_75t_R FILLER_0_224_376 ();
 DECAPx2_ASAP7_75t_R FILLER_0_224_386 ();
 DECAPx4_ASAP7_75t_R FILLER_0_224_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224_408 ();
 DECAPx10_ASAP7_75t_R FILLER_0_224_412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_224_434 ();
 DECAPx2_ASAP7_75t_R FILLER_0_224_456 ();
 DECAPx2_ASAP7_75t_R FILLER_0_224_464 ();
 FILLER_ASAP7_75t_R FILLER_0_224_478 ();
 FILLER_ASAP7_75t_R FILLER_0_224_492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_224_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224_515 ();
 DECAPx4_ASAP7_75t_R FILLER_0_224_537 ();
 FILLER_ASAP7_75t_R FILLER_0_224_559 ();
 FILLER_ASAP7_75t_R FILLER_0_224_573 ();
 DECAPx2_ASAP7_75t_R FILLER_0_224_578 ();
 FILLER_ASAP7_75t_R FILLER_0_224_584 ();
 DECAPx10_ASAP7_75t_R FILLER_0_224_607 ();
 DECAPx4_ASAP7_75t_R FILLER_0_224_629 ();
 FILLER_ASAP7_75t_R FILLER_0_224_647 ();
 DECAPx2_ASAP7_75t_R FILLER_0_224_652 ();
 DECAPx2_ASAP7_75t_R FILLER_0_224_670 ();
 DECAPx1_ASAP7_75t_R FILLER_0_224_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224_683 ();
 DECAPx2_ASAP7_75t_R FILLER_0_224_696 ();
 FILLER_ASAP7_75t_R FILLER_0_224_702 ();
 DECAPx4_ASAP7_75t_R FILLER_0_224_716 ();
 DECAPx4_ASAP7_75t_R FILLER_0_224_737 ();
 FILLER_ASAP7_75t_R FILLER_0_224_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224_749 ();
 DECAPx4_ASAP7_75t_R FILLER_0_224_760 ();
 FILLER_ASAP7_75t_R FILLER_0_224_770 ();
 FILLER_ASAP7_75t_R FILLER_0_224_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224_777 ();
 DECAPx6_ASAP7_75t_R FILLER_0_224_784 ();
 DECAPx1_ASAP7_75t_R FILLER_0_224_798 ();
 DECAPx2_ASAP7_75t_R FILLER_0_224_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224_814 ();
 DECAPx6_ASAP7_75t_R FILLER_0_224_821 ();
 FILLER_ASAP7_75t_R FILLER_0_224_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224_837 ();
 DECAPx1_ASAP7_75t_R FILLER_0_224_844 ();
 DECAPx1_ASAP7_75t_R FILLER_0_224_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224_858 ();
 DECAPx10_ASAP7_75t_R FILLER_0_224_865 ();
 DECAPx2_ASAP7_75t_R FILLER_0_224_887 ();
 FILLER_ASAP7_75t_R FILLER_0_224_893 ();
 FILLER_ASAP7_75t_R FILLER_0_224_901 ();
 FILLER_ASAP7_75t_R FILLER_0_224_909 ();
 FILLER_ASAP7_75t_R FILLER_0_224_917 ();
 DECAPx10_ASAP7_75t_R FILLER_0_224_925 ();
 FILLER_ASAP7_75t_R FILLER_0_224_947 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224_949 ();
 DECAPx6_ASAP7_75t_R FILLER_0_224_953 ();
 FILLER_ASAP7_75t_R FILLER_0_224_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224_969 ();
 FILLER_ASAP7_75t_R FILLER_0_224_973 ();
 DECAPx6_ASAP7_75t_R FILLER_0_224_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224_995 ();
 FILLER_ASAP7_75t_R FILLER_0_224_999 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224_1001 ();
 DECAPx1_ASAP7_75t_R FILLER_0_224_1008 ();
 DECAPx2_ASAP7_75t_R FILLER_0_224_1018 ();
 FILLER_ASAP7_75t_R FILLER_0_224_1024 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224_1026 ();
 FILLER_ASAP7_75t_R FILLER_0_224_1030 ();
 FILLER_ASAP7_75t_R FILLER_0_224_1038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_224_1046 ();
 DECAPx2_ASAP7_75t_R FILLER_0_224_1068 ();
 FILLER_ASAP7_75t_R FILLER_0_224_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_224_1082 ();
 DECAPx6_ASAP7_75t_R FILLER_0_224_1104 ();
 DECAPx1_ASAP7_75t_R FILLER_0_224_1118 ();
 FILLER_ASAP7_75t_R FILLER_0_224_1125 ();
 FILLER_ASAP7_75t_R FILLER_0_224_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224_1167 ();
 FILLER_ASAP7_75t_R FILLER_0_224_1175 ();
 FILLER_ASAP7_75t_R FILLER_0_224_1183 ();
 FILLER_ASAP7_75t_R FILLER_0_224_1191 ();
 FILLER_ASAP7_75t_R FILLER_0_224_1198 ();
 FILLER_ASAP7_75t_R FILLER_0_224_1210 ();
 DECAPx2_ASAP7_75t_R FILLER_0_224_1223 ();
 FILLER_ASAP7_75t_R FILLER_0_224_1236 ();
 DECAPx1_ASAP7_75t_R FILLER_0_224_1244 ();
 FILLER_ASAP7_75t_R FILLER_0_224_1254 ();
 DECAPx4_ASAP7_75t_R FILLER_0_224_1259 ();
 FILLER_ASAP7_75t_R FILLER_0_224_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224_1271 ();
 FILLER_ASAP7_75t_R FILLER_0_224_1278 ();
 DECAPx1_ASAP7_75t_R FILLER_0_224_1286 ();
 FILLER_ASAP7_75t_R FILLER_0_224_1297 ();
 DECAPx2_ASAP7_75t_R FILLER_0_224_1305 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224_1311 ();
 FILLER_ASAP7_75t_R FILLER_0_224_1324 ();
 FILLER_ASAP7_75t_R FILLER_0_224_1333 ();
 FILLER_ASAP7_75t_R FILLER_0_224_1355 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_224_1364 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224_1366 ();
 DECAPx1_ASAP7_75t_R FILLER_0_224_1378 ();
 DECAPx2_ASAP7_75t_R FILLER_0_225_2 ();
 FILLER_ASAP7_75t_R FILLER_0_225_8 ();
 FILLER_ASAP7_75t_R FILLER_0_225_16 ();
 FILLER_ASAP7_75t_R FILLER_0_225_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_26 ();
 FILLER_ASAP7_75t_R FILLER_0_225_37 ();
 FILLER_ASAP7_75t_R FILLER_0_225_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_49 ();
 FILLER_ASAP7_75t_R FILLER_0_225_62 ();
 DECAPx2_ASAP7_75t_R FILLER_0_225_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_77 ();
 DECAPx2_ASAP7_75t_R FILLER_0_225_88 ();
 FILLER_ASAP7_75t_R FILLER_0_225_104 ();
 FILLER_ASAP7_75t_R FILLER_0_225_116 ();
 FILLER_ASAP7_75t_R FILLER_0_225_124 ();
 FILLER_ASAP7_75t_R FILLER_0_225_133 ();
 FILLER_ASAP7_75t_R FILLER_0_225_142 ();
 DECAPx2_ASAP7_75t_R FILLER_0_225_149 ();
 DECAPx4_ASAP7_75t_R FILLER_0_225_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_172 ();
 DECAPx4_ASAP7_75t_R FILLER_0_225_181 ();
 FILLER_ASAP7_75t_R FILLER_0_225_191 ();
 FILLER_ASAP7_75t_R FILLER_0_225_203 ();
 FILLER_ASAP7_75t_R FILLER_0_225_215 ();
 FILLER_ASAP7_75t_R FILLER_0_225_225 ();
 DECAPx4_ASAP7_75t_R FILLER_0_225_233 ();
 DECAPx2_ASAP7_75t_R FILLER_0_225_253 ();
 FILLER_ASAP7_75t_R FILLER_0_225_265 ();
 DECAPx4_ASAP7_75t_R FILLER_0_225_270 ();
 FILLER_ASAP7_75t_R FILLER_0_225_286 ();
 DECAPx10_ASAP7_75t_R FILLER_0_225_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_316 ();
 DECAPx4_ASAP7_75t_R FILLER_0_225_339 ();
 FILLER_ASAP7_75t_R FILLER_0_225_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_357 ();
 FILLER_ASAP7_75t_R FILLER_0_225_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_366 ();
 FILLER_ASAP7_75t_R FILLER_0_225_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_375 ();
 FILLER_ASAP7_75t_R FILLER_0_225_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_384 ();
 FILLER_ASAP7_75t_R FILLER_0_225_391 ();
 DECAPx4_ASAP7_75t_R FILLER_0_225_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_406 ();
 FILLER_ASAP7_75t_R FILLER_0_225_413 ();
 DECAPx10_ASAP7_75t_R FILLER_0_225_425 ();
 FILLER_ASAP7_75t_R FILLER_0_225_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_449 ();
 DECAPx4_ASAP7_75t_R FILLER_0_225_471 ();
 DECAPx4_ASAP7_75t_R FILLER_0_225_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_503 ();
 DECAPx2_ASAP7_75t_R FILLER_0_225_508 ();
 FILLER_ASAP7_75t_R FILLER_0_225_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_516 ();
 FILLER_ASAP7_75t_R FILLER_0_225_525 ();
 DECAPx4_ASAP7_75t_R FILLER_0_225_530 ();
 FILLER_ASAP7_75t_R FILLER_0_225_546 ();
 DECAPx4_ASAP7_75t_R FILLER_0_225_560 ();
 FILLER_ASAP7_75t_R FILLER_0_225_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_583 ();
 FILLER_ASAP7_75t_R FILLER_0_225_587 ();
 FILLER_ASAP7_75t_R FILLER_0_225_594 ();
 FILLER_ASAP7_75t_R FILLER_0_225_602 ();
 DECAPx2_ASAP7_75t_R FILLER_0_225_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_618 ();
 DECAPx6_ASAP7_75t_R FILLER_0_225_627 ();
 FILLER_ASAP7_75t_R FILLER_0_225_641 ();
 FILLER_ASAP7_75t_R FILLER_0_225_651 ();
 DECAPx2_ASAP7_75t_R FILLER_0_225_656 ();
 FILLER_ASAP7_75t_R FILLER_0_225_662 ();
 FILLER_ASAP7_75t_R FILLER_0_225_685 ();
 FILLER_ASAP7_75t_R FILLER_0_225_693 ();
 DECAPx1_ASAP7_75t_R FILLER_0_225_703 ();
 DECAPx6_ASAP7_75t_R FILLER_0_225_728 ();
 DECAPx1_ASAP7_75t_R FILLER_0_225_742 ();
 DECAPx1_ASAP7_75t_R FILLER_0_225_766 ();
 DECAPx1_ASAP7_75t_R FILLER_0_225_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_780 ();
 DECAPx6_ASAP7_75t_R FILLER_0_225_787 ();
 FILLER_ASAP7_75t_R FILLER_0_225_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_803 ();
 DECAPx2_ASAP7_75t_R FILLER_0_225_810 ();
 FILLER_ASAP7_75t_R FILLER_0_225_822 ();
 DECAPx10_ASAP7_75t_R FILLER_0_225_830 ();
 FILLER_ASAP7_75t_R FILLER_0_225_852 ();
 FILLER_ASAP7_75t_R FILLER_0_225_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_859 ();
 DECAPx10_ASAP7_75t_R FILLER_0_225_870 ();
 FILLER_ASAP7_75t_R FILLER_0_225_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_894 ();
 DECAPx6_ASAP7_75t_R FILLER_0_225_905 ();
 DECAPx2_ASAP7_75t_R FILLER_0_225_919 ();
 DECAPx6_ASAP7_75t_R FILLER_0_225_927 ();
 DECAPx2_ASAP7_75t_R FILLER_0_225_941 ();
 DECAPx6_ASAP7_75t_R FILLER_0_225_953 ();
 DECAPx1_ASAP7_75t_R FILLER_0_225_967 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_971 ();
 DECAPx1_ASAP7_75t_R FILLER_0_225_982 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_986 ();
 FILLER_ASAP7_75t_R FILLER_0_225_997 ();
 FILLER_ASAP7_75t_R FILLER_0_225_1009 ();
 FILLER_ASAP7_75t_R FILLER_0_225_1017 ();
 DECAPx4_ASAP7_75t_R FILLER_0_225_1025 ();
 DECAPx2_ASAP7_75t_R FILLER_0_225_1041 ();
 FILLER_ASAP7_75t_R FILLER_0_225_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_1049 ();
 DECAPx6_ASAP7_75t_R FILLER_0_225_1061 ();
 FILLER_ASAP7_75t_R FILLER_0_225_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_1077 ();
 DECAPx4_ASAP7_75t_R FILLER_0_225_1084 ();
 DECAPx6_ASAP7_75t_R FILLER_0_225_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_1115 ();
 FILLER_ASAP7_75t_R FILLER_0_225_1120 ();
 DECAPx1_ASAP7_75t_R FILLER_0_225_1132 ();
 FILLER_ASAP7_75t_R FILLER_0_225_1144 ();
 DECAPx1_ASAP7_75t_R FILLER_0_225_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_1164 ();
 FILLER_ASAP7_75t_R FILLER_0_225_1175 ();
 FILLER_ASAP7_75t_R FILLER_0_225_1187 ();
 FILLER_ASAP7_75t_R FILLER_0_225_1199 ();
 FILLER_ASAP7_75t_R FILLER_0_225_1211 ();
 FILLER_ASAP7_75t_R FILLER_0_225_1223 ();
 FILLER_ASAP7_75t_R FILLER_0_225_1231 ();
 FILLER_ASAP7_75t_R FILLER_0_225_1239 ();
 FILLER_ASAP7_75t_R FILLER_0_225_1247 ();
 DECAPx1_ASAP7_75t_R FILLER_0_225_1252 ();
 FILLER_ASAP7_75t_R FILLER_0_225_1266 ();
 FILLER_ASAP7_75t_R FILLER_0_225_1276 ();
 DECAPx6_ASAP7_75t_R FILLER_0_225_1286 ();
 FILLER_ASAP7_75t_R FILLER_0_225_1300 ();
 DECAPx1_ASAP7_75t_R FILLER_0_225_1308 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225_1312 ();
 FILLER_ASAP7_75t_R FILLER_0_225_1319 ();
 FILLER_ASAP7_75t_R FILLER_0_225_1341 ();
 FILLER_ASAP7_75t_R FILLER_0_225_1353 ();
 DECAPx1_ASAP7_75t_R FILLER_0_225_1358 ();
 FILLER_ASAP7_75t_R FILLER_0_225_1368 ();
 DECAPx2_ASAP7_75t_R FILLER_0_225_1376 ();
 DECAPx4_ASAP7_75t_R FILLER_0_226_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_12 ();
 DECAPx1_ASAP7_75t_R FILLER_0_226_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_27 ();
 FILLER_ASAP7_75t_R FILLER_0_226_31 ();
 FILLER_ASAP7_75t_R FILLER_0_226_53 ();
 DECAPx1_ASAP7_75t_R FILLER_0_226_61 ();
 DECAPx2_ASAP7_75t_R FILLER_0_226_71 ();
 FILLER_ASAP7_75t_R FILLER_0_226_87 ();
 FILLER_ASAP7_75t_R FILLER_0_226_99 ();
 FILLER_ASAP7_75t_R FILLER_0_226_111 ();
 FILLER_ASAP7_75t_R FILLER_0_226_123 ();
 FILLER_ASAP7_75t_R FILLER_0_226_132 ();
 FILLER_ASAP7_75t_R FILLER_0_226_140 ();
 DECAPx1_ASAP7_75t_R FILLER_0_226_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_157 ();
 DECAPx4_ASAP7_75t_R FILLER_0_226_164 ();
 FILLER_ASAP7_75t_R FILLER_0_226_174 ();
 FILLER_ASAP7_75t_R FILLER_0_226_182 ();
 DECAPx2_ASAP7_75t_R FILLER_0_226_190 ();
 FILLER_ASAP7_75t_R FILLER_0_226_202 ();
 FILLER_ASAP7_75t_R FILLER_0_226_214 ();
 FILLER_ASAP7_75t_R FILLER_0_226_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_223 ();
 DECAPx4_ASAP7_75t_R FILLER_0_226_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_244 ();
 FILLER_ASAP7_75t_R FILLER_0_226_253 ();
 DECAPx1_ASAP7_75t_R FILLER_0_226_258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_226_273 ();
 DECAPx6_ASAP7_75t_R FILLER_0_226_295 ();
 DECAPx1_ASAP7_75t_R FILLER_0_226_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_313 ();
 DECAPx6_ASAP7_75t_R FILLER_0_226_319 ();
 DECAPx2_ASAP7_75t_R FILLER_0_226_333 ();
 FILLER_ASAP7_75t_R FILLER_0_226_343 ();
 FILLER_ASAP7_75t_R FILLER_0_226_351 ();
 FILLER_ASAP7_75t_R FILLER_0_226_358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_226_370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_226_392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_226_414 ();
 DECAPx2_ASAP7_75t_R FILLER_0_226_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_442 ();
 FILLER_ASAP7_75t_R FILLER_0_226_446 ();
 DECAPx2_ASAP7_75t_R FILLER_0_226_454 ();
 FILLER_ASAP7_75t_R FILLER_0_226_460 ();
 DECAPx1_ASAP7_75t_R FILLER_0_226_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_226_472 ();
 DECAPx1_ASAP7_75t_R FILLER_0_226_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_498 ();
 DECAPx4_ASAP7_75t_R FILLER_0_226_520 ();
 FILLER_ASAP7_75t_R FILLER_0_226_530 ();
 FILLER_ASAP7_75t_R FILLER_0_226_544 ();
 FILLER_ASAP7_75t_R FILLER_0_226_558 ();
 DECAPx10_ASAP7_75t_R FILLER_0_226_570 ();
 DECAPx4_ASAP7_75t_R FILLER_0_226_592 ();
 DECAPx4_ASAP7_75t_R FILLER_0_226_608 ();
 FILLER_ASAP7_75t_R FILLER_0_226_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_620 ();
 DECAPx6_ASAP7_75t_R FILLER_0_226_629 ();
 FILLER_ASAP7_75t_R FILLER_0_226_643 ();
 FILLER_ASAP7_75t_R FILLER_0_226_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_655 ();
 DECAPx1_ASAP7_75t_R FILLER_0_226_668 ();
 FILLER_ASAP7_75t_R FILLER_0_226_682 ();
 FILLER_ASAP7_75t_R FILLER_0_226_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_696 ();
 FILLER_ASAP7_75t_R FILLER_0_226_701 ();
 FILLER_ASAP7_75t_R FILLER_0_226_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_226_712 ();
 DECAPx6_ASAP7_75t_R FILLER_0_226_734 ();
 DECAPx4_ASAP7_75t_R FILLER_0_226_753 ();
 FILLER_ASAP7_75t_R FILLER_0_226_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_765 ();
 FILLER_ASAP7_75t_R FILLER_0_226_777 ();
 DECAPx2_ASAP7_75t_R FILLER_0_226_785 ();
 FILLER_ASAP7_75t_R FILLER_0_226_798 ();
 FILLER_ASAP7_75t_R FILLER_0_226_810 ();
 DECAPx1_ASAP7_75t_R FILLER_0_226_822 ();
 DECAPx2_ASAP7_75t_R FILLER_0_226_832 ();
 FILLER_ASAP7_75t_R FILLER_0_226_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_840 ();
 FILLER_ASAP7_75t_R FILLER_0_226_851 ();
 FILLER_ASAP7_75t_R FILLER_0_226_859 ();
 DECAPx10_ASAP7_75t_R FILLER_0_226_864 ();
 DECAPx1_ASAP7_75t_R FILLER_0_226_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_890 ();
 DECAPx2_ASAP7_75t_R FILLER_0_226_897 ();
 FILLER_ASAP7_75t_R FILLER_0_226_903 ();
 DECAPx6_ASAP7_75t_R FILLER_0_226_909 ();
 DECAPx1_ASAP7_75t_R FILLER_0_226_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_927 ();
 DECAPx2_ASAP7_75t_R FILLER_0_226_938 ();
 FILLER_ASAP7_75t_R FILLER_0_226_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_946 ();
 DECAPx6_ASAP7_75t_R FILLER_0_226_955 ();
 FILLER_ASAP7_75t_R FILLER_0_226_969 ();
 FILLER_ASAP7_75t_R FILLER_0_226_977 ();
 DECAPx10_ASAP7_75t_R FILLER_0_226_985 ();
 FILLER_ASAP7_75t_R FILLER_0_226_1007 ();
 DECAPx1_ASAP7_75t_R FILLER_0_226_1015 ();
 FILLER_ASAP7_75t_R FILLER_0_226_1029 ();
 FILLER_ASAP7_75t_R FILLER_0_226_1037 ();
 DECAPx1_ASAP7_75t_R FILLER_0_226_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_1049 ();
 DECAPx2_ASAP7_75t_R FILLER_0_226_1056 ();
 FILLER_ASAP7_75t_R FILLER_0_226_1062 ();
 FILLER_ASAP7_75t_R FILLER_0_226_1075 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_1077 ();
 DECAPx1_ASAP7_75t_R FILLER_0_226_1084 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_1088 ();
 FILLER_ASAP7_75t_R FILLER_0_226_1095 ();
 DECAPx4_ASAP7_75t_R FILLER_0_226_1103 ();
 FILLER_ASAP7_75t_R FILLER_0_226_1113 ();
 FILLER_ASAP7_75t_R FILLER_0_226_1125 ();
 DECAPx2_ASAP7_75t_R FILLER_0_226_1133 ();
 DECAPx2_ASAP7_75t_R FILLER_0_226_1151 ();
 FILLER_ASAP7_75t_R FILLER_0_226_1157 ();
 FILLER_ASAP7_75t_R FILLER_0_226_1169 ();
 DECAPx2_ASAP7_75t_R FILLER_0_226_1177 ();
 FILLER_ASAP7_75t_R FILLER_0_226_1183 ();
 FILLER_ASAP7_75t_R FILLER_0_226_1195 ();
 FILLER_ASAP7_75t_R FILLER_0_226_1207 ();
 FILLER_ASAP7_75t_R FILLER_0_226_1219 ();
 FILLER_ASAP7_75t_R FILLER_0_226_1229 ();
 FILLER_ASAP7_75t_R FILLER_0_226_1238 ();
 DECAPx4_ASAP7_75t_R FILLER_0_226_1246 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_1256 ();
 FILLER_ASAP7_75t_R FILLER_0_226_1262 ();
 DECAPx1_ASAP7_75t_R FILLER_0_226_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_1274 ();
 DECAPx2_ASAP7_75t_R FILLER_0_226_1281 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_1287 ();
 FILLER_ASAP7_75t_R FILLER_0_226_1295 ();
 DECAPx6_ASAP7_75t_R FILLER_0_226_1303 ();
 DECAPx1_ASAP7_75t_R FILLER_0_226_1317 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_1321 ();
 DECAPx2_ASAP7_75t_R FILLER_0_226_1329 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226_1335 ();
 DECAPx1_ASAP7_75t_R FILLER_0_226_1346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_226_1356 ();
 DECAPx1_ASAP7_75t_R FILLER_0_226_1378 ();
 DECAPx4_ASAP7_75t_R FILLER_0_227_2 ();
 FILLER_ASAP7_75t_R FILLER_0_227_12 ();
 DECAPx2_ASAP7_75t_R FILLER_0_227_20 ();
 FILLER_ASAP7_75t_R FILLER_0_227_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_28 ();
 DECAPx4_ASAP7_75t_R FILLER_0_227_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_49 ();
 FILLER_ASAP7_75t_R FILLER_0_227_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_58 ();
 FILLER_ASAP7_75t_R FILLER_0_227_64 ();
 FILLER_ASAP7_75t_R FILLER_0_227_72 ();
 FILLER_ASAP7_75t_R FILLER_0_227_84 ();
 FILLER_ASAP7_75t_R FILLER_0_227_96 ();
 FILLER_ASAP7_75t_R FILLER_0_227_112 ();
 DECAPx1_ASAP7_75t_R FILLER_0_227_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_128 ();
 FILLER_ASAP7_75t_R FILLER_0_227_144 ();
 DECAPx1_ASAP7_75t_R FILLER_0_227_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_156 ();
 FILLER_ASAP7_75t_R FILLER_0_227_168 ();
 DECAPx1_ASAP7_75t_R FILLER_0_227_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_184 ();
 FILLER_ASAP7_75t_R FILLER_0_227_191 ();
 DECAPx2_ASAP7_75t_R FILLER_0_227_204 ();
 FILLER_ASAP7_75t_R FILLER_0_227_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_227_223 ();
 DECAPx6_ASAP7_75t_R FILLER_0_227_245 ();
 DECAPx6_ASAP7_75t_R FILLER_0_227_280 ();
 FILLER_ASAP7_75t_R FILLER_0_227_297 ();
 DECAPx1_ASAP7_75t_R FILLER_0_227_309 ();
 DECAPx2_ASAP7_75t_R FILLER_0_227_323 ();
 FILLER_ASAP7_75t_R FILLER_0_227_339 ();
 DECAPx2_ASAP7_75t_R FILLER_0_227_351 ();
 FILLER_ASAP7_75t_R FILLER_0_227_357 ();
 FILLER_ASAP7_75t_R FILLER_0_227_369 ();
 FILLER_ASAP7_75t_R FILLER_0_227_378 ();
 FILLER_ASAP7_75t_R FILLER_0_227_386 ();
 DECAPx10_ASAP7_75t_R FILLER_0_227_393 ();
 DECAPx2_ASAP7_75t_R FILLER_0_227_415 ();
 FILLER_ASAP7_75t_R FILLER_0_227_421 ();
 DECAPx2_ASAP7_75t_R FILLER_0_227_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_439 ();
 DECAPx2_ASAP7_75t_R FILLER_0_227_451 ();
 DECAPx1_ASAP7_75t_R FILLER_0_227_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_464 ();
 DECAPx6_ASAP7_75t_R FILLER_0_227_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_485 ();
 DECAPx4_ASAP7_75t_R FILLER_0_227_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_517 ();
 DECAPx2_ASAP7_75t_R FILLER_0_227_521 ();
 FILLER_ASAP7_75t_R FILLER_0_227_532 ();
 FILLER_ASAP7_75t_R FILLER_0_227_540 ();
 DECAPx1_ASAP7_75t_R FILLER_0_227_548 ();
 FILLER_ASAP7_75t_R FILLER_0_227_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_227_573 ();
 DECAPx2_ASAP7_75t_R FILLER_0_227_595 ();
 FILLER_ASAP7_75t_R FILLER_0_227_609 ();
 FILLER_ASAP7_75t_R FILLER_0_227_619 ();
 DECAPx2_ASAP7_75t_R FILLER_0_227_629 ();
 FILLER_ASAP7_75t_R FILLER_0_227_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_637 ();
 FILLER_ASAP7_75t_R FILLER_0_227_641 ();
 DECAPx10_ASAP7_75t_R FILLER_0_227_651 ();
 DECAPx4_ASAP7_75t_R FILLER_0_227_673 ();
 FILLER_ASAP7_75t_R FILLER_0_227_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_685 ();
 FILLER_ASAP7_75t_R FILLER_0_227_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_694 ();
 DECAPx4_ASAP7_75t_R FILLER_0_227_716 ();
 FILLER_ASAP7_75t_R FILLER_0_227_732 ();
 FILLER_ASAP7_75t_R FILLER_0_227_744 ();
 FILLER_ASAP7_75t_R FILLER_0_227_767 ();
 FILLER_ASAP7_75t_R FILLER_0_227_772 ();
 DECAPx2_ASAP7_75t_R FILLER_0_227_780 ();
 FILLER_ASAP7_75t_R FILLER_0_227_786 ();
 DECAPx6_ASAP7_75t_R FILLER_0_227_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_814 ();
 DECAPx4_ASAP7_75t_R FILLER_0_227_820 ();
 FILLER_ASAP7_75t_R FILLER_0_227_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_832 ();
 FILLER_ASAP7_75t_R FILLER_0_227_839 ();
 FILLER_ASAP7_75t_R FILLER_0_227_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_853 ();
 DECAPx6_ASAP7_75t_R FILLER_0_227_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_874 ();
 DECAPx2_ASAP7_75t_R FILLER_0_227_885 ();
 FILLER_ASAP7_75t_R FILLER_0_227_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_893 ();
 DECAPx4_ASAP7_75t_R FILLER_0_227_897 ();
 DECAPx1_ASAP7_75t_R FILLER_0_227_913 ();
 FILLER_ASAP7_75t_R FILLER_0_227_923 ();
 FILLER_ASAP7_75t_R FILLER_0_227_927 ();
 DECAPx2_ASAP7_75t_R FILLER_0_227_940 ();
 FILLER_ASAP7_75t_R FILLER_0_227_949 ();
 DECAPx6_ASAP7_75t_R FILLER_0_227_957 ();
 DECAPx2_ASAP7_75t_R FILLER_0_227_974 ();
 DECAPx4_ASAP7_75t_R FILLER_0_227_986 ();
 FILLER_ASAP7_75t_R FILLER_0_227_996 ();
 DECAPx1_ASAP7_75t_R FILLER_0_227_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_1008 ();
 DECAPx1_ASAP7_75t_R FILLER_0_227_1029 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_1033 ();
 DECAPx1_ASAP7_75t_R FILLER_0_227_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_1044 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1051 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1059 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1067 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1075 ();
 DECAPx2_ASAP7_75t_R FILLER_0_227_1083 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1089 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1097 ();
 DECAPx10_ASAP7_75t_R FILLER_0_227_1105 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_1129 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1136 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1141 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_1148 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1154 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1166 ();
 DECAPx2_ASAP7_75t_R FILLER_0_227_1174 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1180 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1188 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1200 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1207 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1219 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1227 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1235 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1243 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_1245 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1251 ();
 DECAPx6_ASAP7_75t_R FILLER_0_227_1263 ();
 DECAPx1_ASAP7_75t_R FILLER_0_227_1277 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1288 ();
 DECAPx2_ASAP7_75t_R FILLER_0_227_1301 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1307 ();
 DECAPx6_ASAP7_75t_R FILLER_0_227_1319 ();
 DECAPx2_ASAP7_75t_R FILLER_0_227_1333 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_1339 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1348 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1356 ();
 FILLER_ASAP7_75t_R FILLER_0_227_1369 ();
 DECAPx1_ASAP7_75t_R FILLER_0_227_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227_1381 ();
 DECAPx2_ASAP7_75t_R FILLER_0_228_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_228_8 ();
 FILLER_ASAP7_75t_R FILLER_0_228_15 ();
 DECAPx1_ASAP7_75t_R FILLER_0_228_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_228_27 ();
 DECAPx2_ASAP7_75t_R FILLER_0_228_34 ();
 FILLER_ASAP7_75t_R FILLER_0_228_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_228_42 ();
 FILLER_ASAP7_75t_R FILLER_0_228_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_228_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_228_63 ();
 FILLER_ASAP7_75t_R FILLER_0_228_69 ();
 FILLER_ASAP7_75t_R FILLER_0_228_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_228_93 ();
 FILLER_ASAP7_75t_R FILLER_0_228_102 ();
 FILLER_ASAP7_75t_R FILLER_0_228_114 ();
 DECAPx2_ASAP7_75t_R FILLER_0_228_128 ();
 FILLER_ASAP7_75t_R FILLER_0_228_141 ();
 FILLER_ASAP7_75t_R FILLER_0_228_148 ();
 FILLER_ASAP7_75t_R FILLER_0_228_156 ();
 FILLER_ASAP7_75t_R FILLER_0_228_164 ();
 FILLER_ASAP7_75t_R FILLER_0_228_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_228_174 ();
 FILLER_ASAP7_75t_R FILLER_0_228_183 ();
 DECAPx6_ASAP7_75t_R FILLER_0_228_191 ();
 DECAPx1_ASAP7_75t_R FILLER_0_228_205 ();
 DECAPx10_ASAP7_75t_R FILLER_0_228_215 ();
 DECAPx6_ASAP7_75t_R FILLER_0_228_237 ();
 DECAPx1_ASAP7_75t_R FILLER_0_228_251 ();
 FILLER_ASAP7_75t_R FILLER_0_228_258 ();
 FILLER_ASAP7_75t_R FILLER_0_228_266 ();
 DECAPx4_ASAP7_75t_R FILLER_0_228_274 ();
 FILLER_ASAP7_75t_R FILLER_0_228_284 ();
 DECAPx4_ASAP7_75t_R FILLER_0_228_292 ();
 FILLER_ASAP7_75t_R FILLER_0_228_312 ();
 FILLER_ASAP7_75t_R FILLER_0_228_319 ();
 DECAPx2_ASAP7_75t_R FILLER_0_228_331 ();
 DECAPx1_ASAP7_75t_R FILLER_0_228_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_228_351 ();
 FILLER_ASAP7_75t_R FILLER_0_228_362 ();
 DECAPx1_ASAP7_75t_R FILLER_0_228_374 ();
 FILLER_ASAP7_75t_R FILLER_0_228_388 ();
 DECAPx1_ASAP7_75t_R FILLER_0_228_400 ();
 FILLER_ASAP7_75t_R FILLER_0_228_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_228_409 ();
 DECAPx1_ASAP7_75t_R FILLER_0_228_416 ();
 DECAPx1_ASAP7_75t_R FILLER_0_228_440 ();
 DECAPx1_ASAP7_75t_R FILLER_0_228_450 ();
 FILLER_ASAP7_75t_R FILLER_0_228_460 ();
 FILLER_ASAP7_75t_R FILLER_0_228_464 ();
 DECAPx4_ASAP7_75t_R FILLER_0_228_472 ();
 FILLER_ASAP7_75t_R FILLER_0_228_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_228_484 ();
 FILLER_ASAP7_75t_R FILLER_0_228_493 ();
 DECAPx2_ASAP7_75t_R FILLER_0_228_498 ();
 FILLER_ASAP7_75t_R FILLER_0_228_510 ();
 DECAPx6_ASAP7_75t_R FILLER_0_228_515 ();
 DECAPx1_ASAP7_75t_R FILLER_0_228_529 ();
 FILLER_ASAP7_75t_R FILLER_0_228_544 ();
 FILLER_ASAP7_75t_R FILLER_0_228_549 ();
 DECAPx2_ASAP7_75t_R FILLER_0_228_559 ();
 FILLER_ASAP7_75t_R FILLER_0_228_565 ();
 DECAPx10_ASAP7_75t_R FILLER_0_228_575 ();
 FILLER_ASAP7_75t_R FILLER_0_228_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_228_599 ();
 DECAPx1_ASAP7_75t_R FILLER_0_228_606 ();
 DECAPx1_ASAP7_75t_R FILLER_0_228_617 ();
 DECAPx4_ASAP7_75t_R FILLER_0_228_629 ();
 FILLER_ASAP7_75t_R FILLER_0_228_639 ();
 DECAPx10_ASAP7_75t_R FILLER_0_228_649 ();
 DECAPx2_ASAP7_75t_R FILLER_0_228_671 ();
 FILLER_ASAP7_75t_R FILLER_0_228_677 ();
 FILLER_ASAP7_75t_R FILLER_0_228_687 ();
 FILLER_ASAP7_75t_R FILLER_0_228_695 ();
 FILLER_ASAP7_75t_R FILLER_0_228_703 ();
 DECAPx1_ASAP7_75t_R FILLER_0_228_708 ();
 FILLER_ASAP7_75t_R FILLER_0_228_720 ();
 DECAPx2_ASAP7_75t_R FILLER_0_228_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_228_742 ();
 FILLER_ASAP7_75t_R FILLER_0_228_754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_228_759 ();
 DECAPx4_ASAP7_75t_R FILLER_0_228_781 ();
 FILLER_ASAP7_75t_R FILLER_0_228_803 ();
 DECAPx10_ASAP7_75t_R FILLER_0_228_825 ();
 DECAPx6_ASAP7_75t_R FILLER_0_228_847 ();
 FILLER_ASAP7_75t_R FILLER_0_228_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_228_869 ();
 FILLER_ASAP7_75t_R FILLER_0_228_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_228_882 ();
 FILLER_ASAP7_75t_R FILLER_0_228_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_228_888 ();
 DECAPx4_ASAP7_75t_R FILLER_0_228_896 ();
 FILLER_ASAP7_75t_R FILLER_0_228_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_228_908 ();
 FILLER_ASAP7_75t_R FILLER_0_228_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_228_917 ();
 FILLER_ASAP7_75t_R FILLER_0_228_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_228_936 ();
 DECAPx1_ASAP7_75t_R FILLER_0_228_940 ();
 FILLER_ASAP7_75t_R FILLER_0_228_950 ();
 DECAPx4_ASAP7_75t_R FILLER_0_228_958 ();
 FILLER_ASAP7_75t_R FILLER_0_228_968 ();
 DECAPx4_ASAP7_75t_R FILLER_0_228_981 ();
 FILLER_ASAP7_75t_R FILLER_0_228_997 ();
 FILLER_ASAP7_75t_R FILLER_0_228_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_228_1011 ();
 FILLER_ASAP7_75t_R FILLER_0_228_1018 ();
 DECAPx4_ASAP7_75t_R FILLER_0_228_1026 ();
 FILLER_ASAP7_75t_R FILLER_0_228_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_228_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_228_1066 ();
 DECAPx2_ASAP7_75t_R FILLER_0_228_1073 ();
 DECAPx4_ASAP7_75t_R FILLER_0_228_1085 ();
 FILLER_ASAP7_75t_R FILLER_0_228_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_0_228_1103 ();
 FILLER_ASAP7_75t_R FILLER_0_228_1125 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_228_1127 ();
 DECAPx2_ASAP7_75t_R FILLER_0_228_1131 ();
 FILLER_ASAP7_75t_R FILLER_0_228_1143 ();
 FILLER_ASAP7_75t_R FILLER_0_228_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_228_1153 ();
 FILLER_ASAP7_75t_R FILLER_0_228_1162 ();
 FILLER_ASAP7_75t_R FILLER_0_228_1170 ();
 FILLER_ASAP7_75t_R FILLER_0_228_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_228_1180 ();
 FILLER_ASAP7_75t_R FILLER_0_228_1187 ();
 FILLER_ASAP7_75t_R FILLER_0_228_1195 ();
 FILLER_ASAP7_75t_R FILLER_0_228_1200 ();
 FILLER_ASAP7_75t_R FILLER_0_228_1212 ();
 FILLER_ASAP7_75t_R FILLER_0_228_1220 ();
 FILLER_ASAP7_75t_R FILLER_0_228_1228 ();
 FILLER_ASAP7_75t_R FILLER_0_228_1236 ();
 FILLER_ASAP7_75t_R FILLER_0_228_1243 ();
 FILLER_ASAP7_75t_R FILLER_0_228_1255 ();
 DECAPx10_ASAP7_75t_R FILLER_0_228_1262 ();
 DECAPx2_ASAP7_75t_R FILLER_0_228_1284 ();
 FILLER_ASAP7_75t_R FILLER_0_228_1290 ();
 FILLER_ASAP7_75t_R FILLER_0_228_1297 ();
 DECAPx2_ASAP7_75t_R FILLER_0_228_1305 ();
 FILLER_ASAP7_75t_R FILLER_0_228_1311 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_228_1313 ();
 FILLER_ASAP7_75t_R FILLER_0_228_1326 ();
 DECAPx2_ASAP7_75t_R FILLER_0_228_1338 ();
 DECAPx2_ASAP7_75t_R FILLER_0_228_1355 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_228_1361 ();
 DECAPx6_ASAP7_75t_R FILLER_0_228_1368 ();
 DECAPx1_ASAP7_75t_R FILLER_0_229_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229_6 ();
 FILLER_ASAP7_75t_R FILLER_0_229_17 ();
 DECAPx1_ASAP7_75t_R FILLER_0_229_24 ();
 FILLER_ASAP7_75t_R FILLER_0_229_34 ();
 DECAPx4_ASAP7_75t_R FILLER_0_229_42 ();
 FILLER_ASAP7_75t_R FILLER_0_229_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229_54 ();
 DECAPx2_ASAP7_75t_R FILLER_0_229_61 ();
 FILLER_ASAP7_75t_R FILLER_0_229_67 ();
 FILLER_ASAP7_75t_R FILLER_0_229_75 ();
 FILLER_ASAP7_75t_R FILLER_0_229_83 ();
 FILLER_ASAP7_75t_R FILLER_0_229_91 ();
 FILLER_ASAP7_75t_R FILLER_0_229_103 ();
 FILLER_ASAP7_75t_R FILLER_0_229_115 ();
 FILLER_ASAP7_75t_R FILLER_0_229_127 ();
 DECAPx2_ASAP7_75t_R FILLER_0_229_135 ();
 FILLER_ASAP7_75t_R FILLER_0_229_141 ();
 FILLER_ASAP7_75t_R FILLER_0_229_149 ();
 DECAPx4_ASAP7_75t_R FILLER_0_229_154 ();
 FILLER_ASAP7_75t_R FILLER_0_229_164 ();
 FILLER_ASAP7_75t_R FILLER_0_229_172 ();
 FILLER_ASAP7_75t_R FILLER_0_229_192 ();
 FILLER_ASAP7_75t_R FILLER_0_229_199 ();
 DECAPx4_ASAP7_75t_R FILLER_0_229_204 ();
 FILLER_ASAP7_75t_R FILLER_0_229_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229_216 ();
 FILLER_ASAP7_75t_R FILLER_0_229_239 ();
 FILLER_ASAP7_75t_R FILLER_0_229_271 ();
 DECAPx2_ASAP7_75t_R FILLER_0_229_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229_285 ();
 DECAPx2_ASAP7_75t_R FILLER_0_229_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229_298 ();
 FILLER_ASAP7_75t_R FILLER_0_229_304 ();
 DECAPx2_ASAP7_75t_R FILLER_0_229_316 ();
 FILLER_ASAP7_75t_R FILLER_0_229_332 ();
 DECAPx1_ASAP7_75t_R FILLER_0_229_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229_348 ();
 DECAPx2_ASAP7_75t_R FILLER_0_229_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229_360 ();
 FILLER_ASAP7_75t_R FILLER_0_229_381 ();
 FILLER_ASAP7_75t_R FILLER_0_229_403 ();
 DECAPx6_ASAP7_75t_R FILLER_0_229_411 ();
 FILLER_ASAP7_75t_R FILLER_0_229_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229_427 ();
 DECAPx6_ASAP7_75t_R FILLER_0_229_434 ();
 DECAPx2_ASAP7_75t_R FILLER_0_229_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229_454 ();
 DECAPx4_ASAP7_75t_R FILLER_0_229_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229_471 ();
 DECAPx6_ASAP7_75t_R FILLER_0_229_482 ();
 DECAPx2_ASAP7_75t_R FILLER_0_229_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229_502 ();
 FILLER_ASAP7_75t_R FILLER_0_229_514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_229_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229_532 ();
 DECAPx1_ASAP7_75t_R FILLER_0_229_541 ();
 FILLER_ASAP7_75t_R FILLER_0_229_567 ();
 FILLER_ASAP7_75t_R FILLER_0_229_577 ();
 DECAPx2_ASAP7_75t_R FILLER_0_229_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229_597 ();
 FILLER_ASAP7_75t_R FILLER_0_229_610 ();
 FILLER_ASAP7_75t_R FILLER_0_229_619 ();
 DECAPx4_ASAP7_75t_R FILLER_0_229_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229_639 ();
 FILLER_ASAP7_75t_R FILLER_0_229_646 ();
 DECAPx10_ASAP7_75t_R FILLER_0_229_651 ();
 DECAPx2_ASAP7_75t_R FILLER_0_229_673 ();
 DECAPx10_ASAP7_75t_R FILLER_0_229_685 ();
 DECAPx6_ASAP7_75t_R FILLER_0_229_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229_721 ();
 DECAPx1_ASAP7_75t_R FILLER_0_229_732 ();
 DECAPx6_ASAP7_75t_R FILLER_0_229_742 ();
 DECAPx6_ASAP7_75t_R FILLER_0_229_768 ();
 DECAPx6_ASAP7_75t_R FILLER_0_229_794 ();
 FILLER_ASAP7_75t_R FILLER_0_229_808 ();
 DECAPx6_ASAP7_75t_R FILLER_0_229_820 ();
 DECAPx2_ASAP7_75t_R FILLER_0_229_834 ();
 DECAPx10_ASAP7_75t_R FILLER_0_229_843 ();
 FILLER_ASAP7_75t_R FILLER_0_229_885 ();
 FILLER_ASAP7_75t_R FILLER_0_229_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229_895 ();
 DECAPx4_ASAP7_75t_R FILLER_0_229_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229_912 ();
 DECAPx2_ASAP7_75t_R FILLER_0_229_919 ();
 FILLER_ASAP7_75t_R FILLER_0_229_927 ();
 DECAPx4_ASAP7_75t_R FILLER_0_229_935 ();
 FILLER_ASAP7_75t_R FILLER_0_229_945 ();
 DECAPx2_ASAP7_75t_R FILLER_0_229_950 ();
 FILLER_ASAP7_75t_R FILLER_0_229_956 ();
 DECAPx4_ASAP7_75t_R FILLER_0_229_965 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229_975 ();
 FILLER_ASAP7_75t_R FILLER_0_229_983 ();
 FILLER_ASAP7_75t_R FILLER_0_229_990 ();
 FILLER_ASAP7_75t_R FILLER_0_229_998 ();
 FILLER_ASAP7_75t_R FILLER_0_229_1006 ();
 DECAPx4_ASAP7_75t_R FILLER_0_229_1013 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229_1023 ();
 DECAPx1_ASAP7_75t_R FILLER_0_229_1030 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229_1034 ();
 DECAPx1_ASAP7_75t_R FILLER_0_229_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229_1045 ();
 FILLER_ASAP7_75t_R FILLER_0_229_1052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_229_1061 ();
 DECAPx1_ASAP7_75t_R FILLER_0_229_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229_1087 ();
 FILLER_ASAP7_75t_R FILLER_0_229_1094 ();
 DECAPx6_ASAP7_75t_R FILLER_0_229_1116 ();
 DECAPx1_ASAP7_75t_R FILLER_0_229_1130 ();
 DECAPx6_ASAP7_75t_R FILLER_0_229_1145 ();
 DECAPx1_ASAP7_75t_R FILLER_0_229_1169 ();
 DECAPx1_ASAP7_75t_R FILLER_0_229_1184 ();
 FILLER_ASAP7_75t_R FILLER_0_229_1198 ();
 DECAPx4_ASAP7_75t_R FILLER_0_229_1211 ();
 DECAPx2_ASAP7_75t_R FILLER_0_229_1231 ();
 FILLER_ASAP7_75t_R FILLER_0_229_1237 ();
 DECAPx1_ASAP7_75t_R FILLER_0_229_1245 ();
 DECAPx6_ASAP7_75t_R FILLER_0_229_1259 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229_1273 ();
 FILLER_ASAP7_75t_R FILLER_0_229_1281 ();
 FILLER_ASAP7_75t_R FILLER_0_229_1289 ();
 FILLER_ASAP7_75t_R FILLER_0_229_1301 ();
 DECAPx4_ASAP7_75t_R FILLER_0_229_1308 ();
 FILLER_ASAP7_75t_R FILLER_0_229_1318 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229_1320 ();
 DECAPx1_ASAP7_75t_R FILLER_0_229_1328 ();
 DECAPx1_ASAP7_75t_R FILLER_0_229_1338 ();
 FILLER_ASAP7_75t_R FILLER_0_229_1348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_229_1356 ();
 DECAPx1_ASAP7_75t_R FILLER_0_229_1378 ();
 DECAPx2_ASAP7_75t_R FILLER_0_230_2 ();
 FILLER_ASAP7_75t_R FILLER_0_230_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_10 ();
 DECAPx2_ASAP7_75t_R FILLER_0_230_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_27 ();
 FILLER_ASAP7_75t_R FILLER_0_230_34 ();
 DECAPx4_ASAP7_75t_R FILLER_0_230_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_52 ();
 FILLER_ASAP7_75t_R FILLER_0_230_59 ();
 DECAPx1_ASAP7_75t_R FILLER_0_230_67 ();
 FILLER_ASAP7_75t_R FILLER_0_230_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_93 ();
 FILLER_ASAP7_75t_R FILLER_0_230_97 ();
 FILLER_ASAP7_75t_R FILLER_0_230_109 ();
 FILLER_ASAP7_75t_R FILLER_0_230_122 ();
 DECAPx2_ASAP7_75t_R FILLER_0_230_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_136 ();
 FILLER_ASAP7_75t_R FILLER_0_230_144 ();
 DECAPx10_ASAP7_75t_R FILLER_0_230_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_173 ();
 FILLER_ASAP7_75t_R FILLER_0_230_181 ();
 FILLER_ASAP7_75t_R FILLER_0_230_195 ();
 FILLER_ASAP7_75t_R FILLER_0_230_203 ();
 DECAPx2_ASAP7_75t_R FILLER_0_230_211 ();
 FILLER_ASAP7_75t_R FILLER_0_230_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_219 ();
 DECAPx4_ASAP7_75t_R FILLER_0_230_223 ();
 FILLER_ASAP7_75t_R FILLER_0_230_245 ();
 DECAPx2_ASAP7_75t_R FILLER_0_230_267 ();
 DECAPx1_ASAP7_75t_R FILLER_0_230_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_285 ();
 DECAPx2_ASAP7_75t_R FILLER_0_230_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_298 ();
 FILLER_ASAP7_75t_R FILLER_0_230_309 ();
 FILLER_ASAP7_75t_R FILLER_0_230_329 ();
 FILLER_ASAP7_75t_R FILLER_0_230_337 ();
 FILLER_ASAP7_75t_R FILLER_0_230_359 ();
 DECAPx2_ASAP7_75t_R FILLER_0_230_371 ();
 FILLER_ASAP7_75t_R FILLER_0_230_377 ();
 FILLER_ASAP7_75t_R FILLER_0_230_389 ();
 FILLER_ASAP7_75t_R FILLER_0_230_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_399 ();
 DECAPx6_ASAP7_75t_R FILLER_0_230_411 ();
 DECAPx1_ASAP7_75t_R FILLER_0_230_436 ();
 FILLER_ASAP7_75t_R FILLER_0_230_460 ();
 DECAPx4_ASAP7_75t_R FILLER_0_230_464 ();
 FILLER_ASAP7_75t_R FILLER_0_230_474 ();
 DECAPx6_ASAP7_75t_R FILLER_0_230_482 ();
 DECAPx2_ASAP7_75t_R FILLER_0_230_496 ();
 DECAPx1_ASAP7_75t_R FILLER_0_230_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_230_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_531 ();
 FILLER_ASAP7_75t_R FILLER_0_230_540 ();
 DECAPx2_ASAP7_75t_R FILLER_0_230_548 ();
 FILLER_ASAP7_75t_R FILLER_0_230_564 ();
 DECAPx6_ASAP7_75t_R FILLER_0_230_572 ();
 DECAPx10_ASAP7_75t_R FILLER_0_230_592 ();
 DECAPx1_ASAP7_75t_R FILLER_0_230_614 ();
 DECAPx4_ASAP7_75t_R FILLER_0_230_625 ();
 FILLER_ASAP7_75t_R FILLER_0_230_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_637 ();
 DECAPx2_ASAP7_75t_R FILLER_0_230_649 ();
 DECAPx1_ASAP7_75t_R FILLER_0_230_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_667 ();
 DECAPx6_ASAP7_75t_R FILLER_0_230_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_692 ();
 DECAPx10_ASAP7_75t_R FILLER_0_230_701 ();
 FILLER_ASAP7_75t_R FILLER_0_230_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_725 ();
 DECAPx10_ASAP7_75t_R FILLER_0_230_732 ();
 DECAPx4_ASAP7_75t_R FILLER_0_230_754 ();
 FILLER_ASAP7_75t_R FILLER_0_230_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_230_775 ();
 DECAPx10_ASAP7_75t_R FILLER_0_230_797 ();
 DECAPx4_ASAP7_75t_R FILLER_0_230_819 ();
 FILLER_ASAP7_75t_R FILLER_0_230_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_831 ();
 FILLER_ASAP7_75t_R FILLER_0_230_838 ();
 FILLER_ASAP7_75t_R FILLER_0_230_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_847 ();
 DECAPx6_ASAP7_75t_R FILLER_0_230_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_868 ();
 DECAPx4_ASAP7_75t_R FILLER_0_230_875 ();
 FILLER_ASAP7_75t_R FILLER_0_230_885 ();
 FILLER_ASAP7_75t_R FILLER_0_230_893 ();
 DECAPx2_ASAP7_75t_R FILLER_0_230_902 ();
 DECAPx2_ASAP7_75t_R FILLER_0_230_914 ();
 DECAPx6_ASAP7_75t_R FILLER_0_230_923 ();
 FILLER_ASAP7_75t_R FILLER_0_230_937 ();
 DECAPx2_ASAP7_75t_R FILLER_0_230_944 ();
 FILLER_ASAP7_75t_R FILLER_0_230_961 ();
 DECAPx1_ASAP7_75t_R FILLER_0_230_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_973 ();
 DECAPx1_ASAP7_75t_R FILLER_0_230_984 ();
 FILLER_ASAP7_75t_R FILLER_0_230_998 ();
 DECAPx2_ASAP7_75t_R FILLER_0_230_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_1012 ();
 FILLER_ASAP7_75t_R FILLER_0_230_1019 ();
 DECAPx2_ASAP7_75t_R FILLER_0_230_1027 ();
 FILLER_ASAP7_75t_R FILLER_0_230_1033 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_1035 ();
 FILLER_ASAP7_75t_R FILLER_0_230_1060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_230_1068 ();
 DECAPx1_ASAP7_75t_R FILLER_0_230_1100 ();
 DECAPx6_ASAP7_75t_R FILLER_0_230_1114 ();
 DECAPx2_ASAP7_75t_R FILLER_0_230_1128 ();
 FILLER_ASAP7_75t_R FILLER_0_230_1140 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_1142 ();
 DECAPx6_ASAP7_75t_R FILLER_0_230_1149 ();
 FILLER_ASAP7_75t_R FILLER_0_230_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_1165 ();
 DECAPx2_ASAP7_75t_R FILLER_0_230_1172 ();
 FILLER_ASAP7_75t_R FILLER_0_230_1178 ();
 DECAPx4_ASAP7_75t_R FILLER_0_230_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_230_1196 ();
 FILLER_ASAP7_75t_R FILLER_0_230_1205 ();
 DECAPx6_ASAP7_75t_R FILLER_0_230_1212 ();
 DECAPx1_ASAP7_75t_R FILLER_0_230_1226 ();
 FILLER_ASAP7_75t_R FILLER_0_230_1236 ();
 FILLER_ASAP7_75t_R FILLER_0_230_1244 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_1246 ();
 FILLER_ASAP7_75t_R FILLER_0_230_1252 ();
 FILLER_ASAP7_75t_R FILLER_0_230_1260 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_1262 ();
 FILLER_ASAP7_75t_R FILLER_0_230_1270 ();
 DECAPx2_ASAP7_75t_R FILLER_0_230_1283 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_1289 ();
 FILLER_ASAP7_75t_R FILLER_0_230_1297 ();
 FILLER_ASAP7_75t_R FILLER_0_230_1305 ();
 DECAPx6_ASAP7_75t_R FILLER_0_230_1313 ();
 DECAPx4_ASAP7_75t_R FILLER_0_230_1333 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_1343 ();
 DECAPx2_ASAP7_75t_R FILLER_0_230_1350 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230_1356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_230_1360 ();
 DECAPx2_ASAP7_75t_R FILLER_0_231_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_8 ();
 FILLER_ASAP7_75t_R FILLER_0_231_21 ();
 FILLER_ASAP7_75t_R FILLER_0_231_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_231_36 ();
 FILLER_ASAP7_75t_R FILLER_0_231_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_52 ();
 DECAPx1_ASAP7_75t_R FILLER_0_231_59 ();
 FILLER_ASAP7_75t_R FILLER_0_231_69 ();
 FILLER_ASAP7_75t_R FILLER_0_231_77 ();
 DECAPx1_ASAP7_75t_R FILLER_0_231_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_93 ();
 FILLER_ASAP7_75t_R FILLER_0_231_104 ();
 FILLER_ASAP7_75t_R FILLER_0_231_112 ();
 FILLER_ASAP7_75t_R FILLER_0_231_120 ();
 DECAPx2_ASAP7_75t_R FILLER_0_231_127 ();
 DECAPx4_ASAP7_75t_R FILLER_0_231_141 ();
 FILLER_ASAP7_75t_R FILLER_0_231_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_153 ();
 FILLER_ASAP7_75t_R FILLER_0_231_160 ();
 DECAPx2_ASAP7_75t_R FILLER_0_231_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_178 ();
 FILLER_ASAP7_75t_R FILLER_0_231_185 ();
 FILLER_ASAP7_75t_R FILLER_0_231_203 ();
 DECAPx2_ASAP7_75t_R FILLER_0_231_211 ();
 FILLER_ASAP7_75t_R FILLER_0_231_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_219 ();
 FILLER_ASAP7_75t_R FILLER_0_231_241 ();
 FILLER_ASAP7_75t_R FILLER_0_231_261 ();
 DECAPx1_ASAP7_75t_R FILLER_0_231_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_275 ();
 FILLER_ASAP7_75t_R FILLER_0_231_282 ();
 DECAPx4_ASAP7_75t_R FILLER_0_231_290 ();
 FILLER_ASAP7_75t_R FILLER_0_231_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_302 ();
 FILLER_ASAP7_75t_R FILLER_0_231_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_312 ();
 FILLER_ASAP7_75t_R FILLER_0_231_323 ();
 FILLER_ASAP7_75t_R FILLER_0_231_349 ();
 DECAPx2_ASAP7_75t_R FILLER_0_231_361 ();
 DECAPx2_ASAP7_75t_R FILLER_0_231_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_383 ();
 DECAPx2_ASAP7_75t_R FILLER_0_231_394 ();
 FILLER_ASAP7_75t_R FILLER_0_231_408 ();
 DECAPx2_ASAP7_75t_R FILLER_0_231_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_421 ();
 FILLER_ASAP7_75t_R FILLER_0_231_430 ();
 FILLER_ASAP7_75t_R FILLER_0_231_437 ();
 FILLER_ASAP7_75t_R FILLER_0_231_445 ();
 DECAPx2_ASAP7_75t_R FILLER_0_231_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_231_468 ();
 DECAPx4_ASAP7_75t_R FILLER_0_231_490 ();
 FILLER_ASAP7_75t_R FILLER_0_231_500 ();
 DECAPx2_ASAP7_75t_R FILLER_0_231_505 ();
 FILLER_ASAP7_75t_R FILLER_0_231_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_513 ();
 DECAPx6_ASAP7_75t_R FILLER_0_231_526 ();
 FILLER_ASAP7_75t_R FILLER_0_231_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_542 ();
 FILLER_ASAP7_75t_R FILLER_0_231_553 ();
 DECAPx2_ASAP7_75t_R FILLER_0_231_561 ();
 FILLER_ASAP7_75t_R FILLER_0_231_567 ();
 DECAPx4_ASAP7_75t_R FILLER_0_231_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_590 ();
 DECAPx4_ASAP7_75t_R FILLER_0_231_597 ();
 FILLER_ASAP7_75t_R FILLER_0_231_617 ();
 DECAPx2_ASAP7_75t_R FILLER_0_231_626 ();
 FILLER_ASAP7_75t_R FILLER_0_231_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_634 ();
 DECAPx1_ASAP7_75t_R FILLER_0_231_645 ();
 DECAPx2_ASAP7_75t_R FILLER_0_231_660 ();
 DECAPx1_ASAP7_75t_R FILLER_0_231_676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_231_688 ();
 DECAPx1_ASAP7_75t_R FILLER_0_231_700 ();
 DECAPx4_ASAP7_75t_R FILLER_0_231_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_720 ();
 FILLER_ASAP7_75t_R FILLER_0_231_727 ();
 DECAPx10_ASAP7_75t_R FILLER_0_231_737 ();
 FILLER_ASAP7_75t_R FILLER_0_231_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_761 ();
 FILLER_ASAP7_75t_R FILLER_0_231_765 ();
 FILLER_ASAP7_75t_R FILLER_0_231_778 ();
 DECAPx2_ASAP7_75t_R FILLER_0_231_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_792 ();
 DECAPx6_ASAP7_75t_R FILLER_0_231_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_817 ();
 FILLER_ASAP7_75t_R FILLER_0_231_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_830 ();
 FILLER_ASAP7_75t_R FILLER_0_231_837 ();
 DECAPx1_ASAP7_75t_R FILLER_0_231_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_849 ();
 FILLER_ASAP7_75t_R FILLER_0_231_856 ();
 DECAPx6_ASAP7_75t_R FILLER_0_231_861 ();
 DECAPx1_ASAP7_75t_R FILLER_0_231_875 ();
 DECAPx4_ASAP7_75t_R FILLER_0_231_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_895 ();
 FILLER_ASAP7_75t_R FILLER_0_231_906 ();
 FILLER_ASAP7_75t_R FILLER_0_231_914 ();
 FILLER_ASAP7_75t_R FILLER_0_231_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_924 ();
 FILLER_ASAP7_75t_R FILLER_0_231_927 ();
 DECAPx4_ASAP7_75t_R FILLER_0_231_936 ();
 FILLER_ASAP7_75t_R FILLER_0_231_946 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_948 ();
 DECAPx2_ASAP7_75t_R FILLER_0_231_955 ();
 FILLER_ASAP7_75t_R FILLER_0_231_961 ();
 DECAPx2_ASAP7_75t_R FILLER_0_231_983 ();
 FILLER_ASAP7_75t_R FILLER_0_231_989 ();
 FILLER_ASAP7_75t_R FILLER_0_231_1003 ();
 FILLER_ASAP7_75t_R FILLER_0_231_1011 ();
 FILLER_ASAP7_75t_R FILLER_0_231_1019 ();
 FILLER_ASAP7_75t_R FILLER_0_231_1027 ();
 FILLER_ASAP7_75t_R FILLER_0_231_1035 ();
 DECAPx4_ASAP7_75t_R FILLER_0_231_1043 ();
 FILLER_ASAP7_75t_R FILLER_0_231_1053 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_1055 ();
 DECAPx2_ASAP7_75t_R FILLER_0_231_1062 ();
 FILLER_ASAP7_75t_R FILLER_0_231_1068 ();
 FILLER_ASAP7_75t_R FILLER_0_231_1076 ();
 DECAPx1_ASAP7_75t_R FILLER_0_231_1085 ();
 FILLER_ASAP7_75t_R FILLER_0_231_1095 ();
 DECAPx4_ASAP7_75t_R FILLER_0_231_1117 ();
 FILLER_ASAP7_75t_R FILLER_0_231_1127 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_1129 ();
 FILLER_ASAP7_75t_R FILLER_0_231_1140 ();
 DECAPx4_ASAP7_75t_R FILLER_0_231_1152 ();
 DECAPx2_ASAP7_75t_R FILLER_0_231_1170 ();
 FILLER_ASAP7_75t_R FILLER_0_231_1176 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_1178 ();
 FILLER_ASAP7_75t_R FILLER_0_231_1182 ();
 DECAPx2_ASAP7_75t_R FILLER_0_231_1194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_231_1208 ();
 DECAPx2_ASAP7_75t_R FILLER_0_231_1230 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_1236 ();
 DECAPx2_ASAP7_75t_R FILLER_0_231_1247 ();
 FILLER_ASAP7_75t_R FILLER_0_231_1253 ();
 DECAPx10_ASAP7_75t_R FILLER_0_231_1263 ();
 DECAPx1_ASAP7_75t_R FILLER_0_231_1285 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_1289 ();
 DECAPx2_ASAP7_75t_R FILLER_0_231_1302 ();
 DECAPx4_ASAP7_75t_R FILLER_0_231_1316 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_1326 ();
 DECAPx1_ASAP7_75t_R FILLER_0_231_1334 ();
 DECAPx2_ASAP7_75t_R FILLER_0_231_1341 ();
 FILLER_ASAP7_75t_R FILLER_0_231_1353 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231_1355 ();
 FILLER_ASAP7_75t_R FILLER_0_231_1362 ();
 DECAPx4_ASAP7_75t_R FILLER_0_231_1370 ();
 FILLER_ASAP7_75t_R FILLER_0_231_1380 ();
 DECAPx2_ASAP7_75t_R FILLER_0_232_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_8 ();
 DECAPx4_ASAP7_75t_R FILLER_0_232_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_27 ();
 FILLER_ASAP7_75t_R FILLER_0_232_38 ();
 DECAPx6_ASAP7_75t_R FILLER_0_232_46 ();
 FILLER_ASAP7_75t_R FILLER_0_232_60 ();
 DECAPx2_ASAP7_75t_R FILLER_0_232_68 ();
 FILLER_ASAP7_75t_R FILLER_0_232_74 ();
 DECAPx2_ASAP7_75t_R FILLER_0_232_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_92 ();
 DECAPx1_ASAP7_75t_R FILLER_0_232_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_103 ();
 FILLER_ASAP7_75t_R FILLER_0_232_110 ();
 FILLER_ASAP7_75t_R FILLER_0_232_118 ();
 DECAPx2_ASAP7_75t_R FILLER_0_232_125 ();
 FILLER_ASAP7_75t_R FILLER_0_232_131 ();
 FILLER_ASAP7_75t_R FILLER_0_232_139 ();
 FILLER_ASAP7_75t_R FILLER_0_232_147 ();
 FILLER_ASAP7_75t_R FILLER_0_232_160 ();
 DECAPx4_ASAP7_75t_R FILLER_0_232_168 ();
 FILLER_ASAP7_75t_R FILLER_0_232_178 ();
 DECAPx6_ASAP7_75t_R FILLER_0_232_186 ();
 DECAPx6_ASAP7_75t_R FILLER_0_232_206 ();
 FILLER_ASAP7_75t_R FILLER_0_232_220 ();
 DECAPx6_ASAP7_75t_R FILLER_0_232_225 ();
 FILLER_ASAP7_75t_R FILLER_0_232_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_241 ();
 FILLER_ASAP7_75t_R FILLER_0_232_254 ();
 DECAPx2_ASAP7_75t_R FILLER_0_232_274 ();
 FILLER_ASAP7_75t_R FILLER_0_232_290 ();
 FILLER_ASAP7_75t_R FILLER_0_232_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_300 ();
 DECAPx2_ASAP7_75t_R FILLER_0_232_307 ();
 DECAPx1_ASAP7_75t_R FILLER_0_232_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_323 ();
 FILLER_ASAP7_75t_R FILLER_0_232_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_332 ();
 DECAPx1_ASAP7_75t_R FILLER_0_232_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_343 ();
 FILLER_ASAP7_75t_R FILLER_0_232_350 ();
 DECAPx6_ASAP7_75t_R FILLER_0_232_366 ();
 FILLER_ASAP7_75t_R FILLER_0_232_380 ();
 DECAPx4_ASAP7_75t_R FILLER_0_232_392 ();
 FILLER_ASAP7_75t_R FILLER_0_232_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_414 ();
 DECAPx1_ASAP7_75t_R FILLER_0_232_421 ();
 DECAPx1_ASAP7_75t_R FILLER_0_232_432 ();
 DECAPx1_ASAP7_75t_R FILLER_0_232_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_446 ();
 DECAPx2_ASAP7_75t_R FILLER_0_232_453 ();
 FILLER_ASAP7_75t_R FILLER_0_232_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_461 ();
 FILLER_ASAP7_75t_R FILLER_0_232_464 ();
 FILLER_ASAP7_75t_R FILLER_0_232_472 ();
 FILLER_ASAP7_75t_R FILLER_0_232_480 ();
 DECAPx4_ASAP7_75t_R FILLER_0_232_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_498 ();
 DECAPx2_ASAP7_75t_R FILLER_0_232_519 ();
 FILLER_ASAP7_75t_R FILLER_0_232_525 ();
 FILLER_ASAP7_75t_R FILLER_0_232_537 ();
 DECAPx4_ASAP7_75t_R FILLER_0_232_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_559 ();
 DECAPx1_ASAP7_75t_R FILLER_0_232_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_570 ();
 DECAPx4_ASAP7_75t_R FILLER_0_232_579 ();
 FILLER_ASAP7_75t_R FILLER_0_232_589 ();
 DECAPx1_ASAP7_75t_R FILLER_0_232_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_601 ();
 FILLER_ASAP7_75t_R FILLER_0_232_612 ();
 FILLER_ASAP7_75t_R FILLER_0_232_624 ();
 FILLER_ASAP7_75t_R FILLER_0_232_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_635 ();
 DECAPx1_ASAP7_75t_R FILLER_0_232_647 ();
 FILLER_ASAP7_75t_R FILLER_0_232_657 ();
 FILLER_ASAP7_75t_R FILLER_0_232_665 ();
 FILLER_ASAP7_75t_R FILLER_0_232_678 ();
 DECAPx1_ASAP7_75t_R FILLER_0_232_686 ();
 FILLER_ASAP7_75t_R FILLER_0_232_694 ();
 FILLER_ASAP7_75t_R FILLER_0_232_699 ();
 DECAPx4_ASAP7_75t_R FILLER_0_232_707 ();
 DECAPx10_ASAP7_75t_R FILLER_0_232_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_751 ();
 DECAPx1_ASAP7_75t_R FILLER_0_232_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_768 ();
 FILLER_ASAP7_75t_R FILLER_0_232_772 ();
 FILLER_ASAP7_75t_R FILLER_0_232_796 ();
 DECAPx2_ASAP7_75t_R FILLER_0_232_819 ();
 FILLER_ASAP7_75t_R FILLER_0_232_825 ();
 DECAPx4_ASAP7_75t_R FILLER_0_232_830 ();
 DECAPx1_ASAP7_75t_R FILLER_0_232_846 ();
 DECAPx4_ASAP7_75t_R FILLER_0_232_861 ();
 DECAPx1_ASAP7_75t_R FILLER_0_232_874 ();
 FILLER_ASAP7_75t_R FILLER_0_232_884 ();
 FILLER_ASAP7_75t_R FILLER_0_232_892 ();
 DECAPx2_ASAP7_75t_R FILLER_0_232_900 ();
 FILLER_ASAP7_75t_R FILLER_0_232_906 ();
 FILLER_ASAP7_75t_R FILLER_0_232_928 ();
 DECAPx4_ASAP7_75t_R FILLER_0_232_941 ();
 FILLER_ASAP7_75t_R FILLER_0_232_951 ();
 DECAPx4_ASAP7_75t_R FILLER_0_232_959 ();
 FILLER_ASAP7_75t_R FILLER_0_232_979 ();
 DECAPx1_ASAP7_75t_R FILLER_0_232_986 ();
 FILLER_ASAP7_75t_R FILLER_0_232_997 ();
 DECAPx2_ASAP7_75t_R FILLER_0_232_1005 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_1011 ();
 FILLER_ASAP7_75t_R FILLER_0_232_1022 ();
 DECAPx1_ASAP7_75t_R FILLER_0_232_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_1031 ();
 FILLER_ASAP7_75t_R FILLER_0_232_1038 ();
 DECAPx1_ASAP7_75t_R FILLER_0_232_1046 ();
 DECAPx2_ASAP7_75t_R FILLER_0_232_1056 ();
 FILLER_ASAP7_75t_R FILLER_0_232_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_1064 ();
 DECAPx2_ASAP7_75t_R FILLER_0_232_1070 ();
 FILLER_ASAP7_75t_R FILLER_0_232_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_1078 ();
 DECAPx2_ASAP7_75t_R FILLER_0_232_1089 ();
 FILLER_ASAP7_75t_R FILLER_0_232_1095 ();
 DECAPx2_ASAP7_75t_R FILLER_0_232_1103 ();
 FILLER_ASAP7_75t_R FILLER_0_232_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_1111 ();
 FILLER_ASAP7_75t_R FILLER_0_232_1118 ();
 DECAPx1_ASAP7_75t_R FILLER_0_232_1130 ();
 FILLER_ASAP7_75t_R FILLER_0_232_1144 ();
 FILLER_ASAP7_75t_R FILLER_0_232_1152 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_1154 ();
 DECAPx4_ASAP7_75t_R FILLER_0_232_1175 ();
 DECAPx2_ASAP7_75t_R FILLER_0_232_1191 ();
 DECAPx1_ASAP7_75t_R FILLER_0_232_1205 ();
 FILLER_ASAP7_75t_R FILLER_0_232_1221 ();
 DECAPx2_ASAP7_75t_R FILLER_0_232_1229 ();
 DECAPx2_ASAP7_75t_R FILLER_0_232_1243 ();
 FILLER_ASAP7_75t_R FILLER_0_232_1249 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_1251 ();
 FILLER_ASAP7_75t_R FILLER_0_232_1258 ();
 FILLER_ASAP7_75t_R FILLER_0_232_1266 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_1268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_232_1275 ();
 FILLER_ASAP7_75t_R FILLER_0_232_1289 ();
 FILLER_ASAP7_75t_R FILLER_0_232_1297 ();
 DECAPx2_ASAP7_75t_R FILLER_0_232_1305 ();
 FILLER_ASAP7_75t_R FILLER_0_232_1311 ();
 FILLER_ASAP7_75t_R FILLER_0_232_1320 ();
 FILLER_ASAP7_75t_R FILLER_0_232_1329 ();
 FILLER_ASAP7_75t_R FILLER_0_232_1341 ();
 DECAPx6_ASAP7_75t_R FILLER_0_232_1349 ();
 FILLER_ASAP7_75t_R FILLER_0_232_1363 ();
 DECAPx4_ASAP7_75t_R FILLER_0_232_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232_1381 ();
 DECAPx4_ASAP7_75t_R FILLER_0_233_2 ();
 FILLER_ASAP7_75t_R FILLER_0_233_18 ();
 DECAPx4_ASAP7_75t_R FILLER_0_233_28 ();
 FILLER_ASAP7_75t_R FILLER_0_233_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_40 ();
 DECAPx10_ASAP7_75t_R FILLER_0_233_47 ();
 DECAPx6_ASAP7_75t_R FILLER_0_233_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_83 ();
 FILLER_ASAP7_75t_R FILLER_0_233_89 ();
 FILLER_ASAP7_75t_R FILLER_0_233_96 ();
 FILLER_ASAP7_75t_R FILLER_0_233_108 ();
 DECAPx2_ASAP7_75t_R FILLER_0_233_120 ();
 FILLER_ASAP7_75t_R FILLER_0_233_133 ();
 DECAPx10_ASAP7_75t_R FILLER_0_233_147 ();
 DECAPx4_ASAP7_75t_R FILLER_0_233_169 ();
 FILLER_ASAP7_75t_R FILLER_0_233_179 ();
 FILLER_ASAP7_75t_R FILLER_0_233_187 ();
 DECAPx4_ASAP7_75t_R FILLER_0_233_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_205 ();
 FILLER_ASAP7_75t_R FILLER_0_233_212 ();
 DECAPx6_ASAP7_75t_R FILLER_0_233_220 ();
 DECAPx1_ASAP7_75t_R FILLER_0_233_262 ();
 FILLER_ASAP7_75t_R FILLER_0_233_272 ();
 DECAPx2_ASAP7_75t_R FILLER_0_233_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_300 ();
 FILLER_ASAP7_75t_R FILLER_0_233_311 ();
 FILLER_ASAP7_75t_R FILLER_0_233_317 ();
 FILLER_ASAP7_75t_R FILLER_0_233_326 ();
 DECAPx1_ASAP7_75t_R FILLER_0_233_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_344 ();
 FILLER_ASAP7_75t_R FILLER_0_233_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_353 ();
 DECAPx2_ASAP7_75t_R FILLER_0_233_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_372 ();
 FILLER_ASAP7_75t_R FILLER_0_233_383 ();
 DECAPx4_ASAP7_75t_R FILLER_0_233_395 ();
 FILLER_ASAP7_75t_R FILLER_0_233_405 ();
 FILLER_ASAP7_75t_R FILLER_0_233_427 ();
 DECAPx2_ASAP7_75t_R FILLER_0_233_441 ();
 DECAPx1_ASAP7_75t_R FILLER_0_233_453 ();
 DECAPx2_ASAP7_75t_R FILLER_0_233_463 ();
 DECAPx2_ASAP7_75t_R FILLER_0_233_475 ();
 FILLER_ASAP7_75t_R FILLER_0_233_481 ();
 FILLER_ASAP7_75t_R FILLER_0_233_489 ();
 DECAPx2_ASAP7_75t_R FILLER_0_233_497 ();
 FILLER_ASAP7_75t_R FILLER_0_233_503 ();
 DECAPx1_ASAP7_75t_R FILLER_0_233_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_519 ();
 DECAPx2_ASAP7_75t_R FILLER_0_233_532 ();
 DECAPx1_ASAP7_75t_R FILLER_0_233_558 ();
 FILLER_ASAP7_75t_R FILLER_0_233_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_570 ();
 DECAPx2_ASAP7_75t_R FILLER_0_233_577 ();
 FILLER_ASAP7_75t_R FILLER_0_233_583 ();
 FILLER_ASAP7_75t_R FILLER_0_233_591 ();
 DECAPx2_ASAP7_75t_R FILLER_0_233_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_607 ();
 FILLER_ASAP7_75t_R FILLER_0_233_616 ();
 DECAPx10_ASAP7_75t_R FILLER_0_233_628 ();
 DECAPx10_ASAP7_75t_R FILLER_0_233_650 ();
 DECAPx2_ASAP7_75t_R FILLER_0_233_672 ();
 FILLER_ASAP7_75t_R FILLER_0_233_678 ();
 DECAPx6_ASAP7_75t_R FILLER_0_233_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_700 ();
 FILLER_ASAP7_75t_R FILLER_0_233_713 ();
 FILLER_ASAP7_75t_R FILLER_0_233_727 ();
 FILLER_ASAP7_75t_R FILLER_0_233_740 ();
 FILLER_ASAP7_75t_R FILLER_0_233_754 ();
 DECAPx6_ASAP7_75t_R FILLER_0_233_762 ();
 DECAPx6_ASAP7_75t_R FILLER_0_233_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_793 ();
 FILLER_ASAP7_75t_R FILLER_0_233_804 ();
 DECAPx4_ASAP7_75t_R FILLER_0_233_816 ();
 DECAPx4_ASAP7_75t_R FILLER_0_233_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_842 ();
 DECAPx6_ASAP7_75t_R FILLER_0_233_846 ();
 DECAPx1_ASAP7_75t_R FILLER_0_233_860 ();
 FILLER_ASAP7_75t_R FILLER_0_233_870 ();
 FILLER_ASAP7_75t_R FILLER_0_233_878 ();
 DECAPx4_ASAP7_75t_R FILLER_0_233_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_896 ();
 DECAPx4_ASAP7_75t_R FILLER_0_233_903 ();
 FILLER_ASAP7_75t_R FILLER_0_233_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_915 ();
 FILLER_ASAP7_75t_R FILLER_0_233_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_924 ();
 DECAPx2_ASAP7_75t_R FILLER_0_233_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_933 ();
 FILLER_ASAP7_75t_R FILLER_0_233_944 ();
 FILLER_ASAP7_75t_R FILLER_0_233_952 ();
 DECAPx1_ASAP7_75t_R FILLER_0_233_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_966 ();
 FILLER_ASAP7_75t_R FILLER_0_233_972 ();
 DECAPx2_ASAP7_75t_R FILLER_0_233_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_998 ();
 FILLER_ASAP7_75t_R FILLER_0_233_1007 ();
 DECAPx6_ASAP7_75t_R FILLER_0_233_1014 ();
 DECAPx6_ASAP7_75t_R FILLER_0_233_1034 ();
 FILLER_ASAP7_75t_R FILLER_0_233_1054 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_1056 ();
 DECAPx10_ASAP7_75t_R FILLER_0_233_1064 ();
 DECAPx2_ASAP7_75t_R FILLER_0_233_1108 ();
 FILLER_ASAP7_75t_R FILLER_0_233_1114 ();
 FILLER_ASAP7_75t_R FILLER_0_233_1126 ();
 FILLER_ASAP7_75t_R FILLER_0_233_1138 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_1140 ();
 FILLER_ASAP7_75t_R FILLER_0_233_1151 ();
 DECAPx10_ASAP7_75t_R FILLER_0_233_1158 ();
 DECAPx2_ASAP7_75t_R FILLER_0_233_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_233_1197 ();
 DECAPx2_ASAP7_75t_R FILLER_0_233_1211 ();
 FILLER_ASAP7_75t_R FILLER_0_233_1217 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_1219 ();
 FILLER_ASAP7_75t_R FILLER_0_233_1229 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_1231 ();
 DECAPx1_ASAP7_75t_R FILLER_0_233_1252 ();
 DECAPx1_ASAP7_75t_R FILLER_0_233_1263 ();
 DECAPx1_ASAP7_75t_R FILLER_0_233_1277 ();
 DECAPx1_ASAP7_75t_R FILLER_0_233_1287 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_1291 ();
 FILLER_ASAP7_75t_R FILLER_0_233_1297 ();
 FILLER_ASAP7_75t_R FILLER_0_233_1310 ();
 DECAPx6_ASAP7_75t_R FILLER_0_233_1317 ();
 FILLER_ASAP7_75t_R FILLER_0_233_1351 ();
 FILLER_ASAP7_75t_R FILLER_0_233_1359 ();
 DECAPx6_ASAP7_75t_R FILLER_0_233_1367 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233_1381 ();
 DECAPx2_ASAP7_75t_R FILLER_0_234_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_8 ();
 DECAPx1_ASAP7_75t_R FILLER_0_234_15 ();
 DECAPx1_ASAP7_75t_R FILLER_0_234_25 ();
 FILLER_ASAP7_75t_R FILLER_0_234_35 ();
 DECAPx1_ASAP7_75t_R FILLER_0_234_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_47 ();
 FILLER_ASAP7_75t_R FILLER_0_234_55 ();
 DECAPx1_ASAP7_75t_R FILLER_0_234_63 ();
 DECAPx1_ASAP7_75t_R FILLER_0_234_73 ();
 FILLER_ASAP7_75t_R FILLER_0_234_83 ();
 FILLER_ASAP7_75t_R FILLER_0_234_91 ();
 FILLER_ASAP7_75t_R FILLER_0_234_103 ();
 FILLER_ASAP7_75t_R FILLER_0_234_115 ();
 FILLER_ASAP7_75t_R FILLER_0_234_128 ();
 FILLER_ASAP7_75t_R FILLER_0_234_136 ();
 DECAPx4_ASAP7_75t_R FILLER_0_234_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_153 ();
 FILLER_ASAP7_75t_R FILLER_0_234_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_170 ();
 FILLER_ASAP7_75t_R FILLER_0_234_181 ();
 DECAPx1_ASAP7_75t_R FILLER_0_234_189 ();
 FILLER_ASAP7_75t_R FILLER_0_234_203 ();
 DECAPx6_ASAP7_75t_R FILLER_0_234_211 ();
 FILLER_ASAP7_75t_R FILLER_0_234_230 ();
 FILLER_ASAP7_75t_R FILLER_0_234_242 ();
 FILLER_ASAP7_75t_R FILLER_0_234_254 ();
 FILLER_ASAP7_75t_R FILLER_0_234_274 ();
 FILLER_ASAP7_75t_R FILLER_0_234_284 ();
 FILLER_ASAP7_75t_R FILLER_0_234_292 ();
 DECAPx2_ASAP7_75t_R FILLER_0_234_300 ();
 DECAPx2_ASAP7_75t_R FILLER_0_234_311 ();
 DECAPx1_ASAP7_75t_R FILLER_0_234_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_327 ();
 DECAPx2_ASAP7_75t_R FILLER_0_234_338 ();
 FILLER_ASAP7_75t_R FILLER_0_234_344 ();
 DECAPx2_ASAP7_75t_R FILLER_0_234_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_362 ();
 DECAPx1_ASAP7_75t_R FILLER_0_234_383 ();
 FILLER_ASAP7_75t_R FILLER_0_234_397 ();
 DECAPx6_ASAP7_75t_R FILLER_0_234_404 ();
 DECAPx4_ASAP7_75t_R FILLER_0_234_424 ();
 FILLER_ASAP7_75t_R FILLER_0_234_434 ();
 FILLER_ASAP7_75t_R FILLER_0_234_442 ();
 DECAPx1_ASAP7_75t_R FILLER_0_234_450 ();
 FILLER_ASAP7_75t_R FILLER_0_234_460 ();
 FILLER_ASAP7_75t_R FILLER_0_234_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_466 ();
 FILLER_ASAP7_75t_R FILLER_0_234_473 ();
 DECAPx6_ASAP7_75t_R FILLER_0_234_485 ();
 DECAPx10_ASAP7_75t_R FILLER_0_234_505 ();
 DECAPx6_ASAP7_75t_R FILLER_0_234_527 ();
 FILLER_ASAP7_75t_R FILLER_0_234_541 ();
 FILLER_ASAP7_75t_R FILLER_0_234_553 ();
 DECAPx2_ASAP7_75t_R FILLER_0_234_563 ();
 DECAPx4_ASAP7_75t_R FILLER_0_234_575 ();
 FILLER_ASAP7_75t_R FILLER_0_234_585 ();
 DECAPx6_ASAP7_75t_R FILLER_0_234_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_611 ();
 DECAPx6_ASAP7_75t_R FILLER_0_234_620 ();
 FILLER_ASAP7_75t_R FILLER_0_234_646 ();
 FILLER_ASAP7_75t_R FILLER_0_234_656 ();
 FILLER_ASAP7_75t_R FILLER_0_234_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_668 ();
 DECAPx6_ASAP7_75t_R FILLER_0_234_672 ();
 FILLER_ASAP7_75t_R FILLER_0_234_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_234_699 ();
 DECAPx2_ASAP7_75t_R FILLER_0_234_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_727 ();
 DECAPx2_ASAP7_75t_R FILLER_0_234_739 ();
 DECAPx10_ASAP7_75t_R FILLER_0_234_757 ();
 DECAPx6_ASAP7_75t_R FILLER_0_234_779 ();
 DECAPx2_ASAP7_75t_R FILLER_0_234_793 ();
 DECAPx6_ASAP7_75t_R FILLER_0_234_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_816 ();
 DECAPx4_ASAP7_75t_R FILLER_0_234_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_837 ();
 DECAPx6_ASAP7_75t_R FILLER_0_234_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_872 ();
 FILLER_ASAP7_75t_R FILLER_0_234_879 ();
 DECAPx6_ASAP7_75t_R FILLER_0_234_887 ();
 FILLER_ASAP7_75t_R FILLER_0_234_911 ();
 DECAPx2_ASAP7_75t_R FILLER_0_234_921 ();
 DECAPx10_ASAP7_75t_R FILLER_0_234_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_955 ();
 DECAPx4_ASAP7_75t_R FILLER_0_234_962 ();
 FILLER_ASAP7_75t_R FILLER_0_234_972 ();
 DECAPx2_ASAP7_75t_R FILLER_0_234_984 ();
 FILLER_ASAP7_75t_R FILLER_0_234_990 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_992 ();
 FILLER_ASAP7_75t_R FILLER_0_234_998 ();
 FILLER_ASAP7_75t_R FILLER_0_234_1006 ();
 FILLER_ASAP7_75t_R FILLER_0_234_1018 ();
 FILLER_ASAP7_75t_R FILLER_0_234_1026 ();
 FILLER_ASAP7_75t_R FILLER_0_234_1034 ();
 DECAPx2_ASAP7_75t_R FILLER_0_234_1044 ();
 DECAPx4_ASAP7_75t_R FILLER_0_234_1056 ();
 FILLER_ASAP7_75t_R FILLER_0_234_1066 ();
 DECAPx2_ASAP7_75t_R FILLER_0_234_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_1080 ();
 FILLER_ASAP7_75t_R FILLER_0_234_1091 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_1093 ();
 FILLER_ASAP7_75t_R FILLER_0_234_1100 ();
 DECAPx2_ASAP7_75t_R FILLER_0_234_1107 ();
 DECAPx1_ASAP7_75t_R FILLER_0_234_1123 ();
 FILLER_ASAP7_75t_R FILLER_0_234_1137 ();
 FILLER_ASAP7_75t_R FILLER_0_234_1151 ();
 FILLER_ASAP7_75t_R FILLER_0_234_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_1163 ();
 DECAPx4_ASAP7_75t_R FILLER_0_234_1178 ();
 FILLER_ASAP7_75t_R FILLER_0_234_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_1190 ();
 FILLER_ASAP7_75t_R FILLER_0_234_1201 ();
 FILLER_ASAP7_75t_R FILLER_0_234_1213 ();
 FILLER_ASAP7_75t_R FILLER_0_234_1221 ();
 FILLER_ASAP7_75t_R FILLER_0_234_1229 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_1231 ();
 DECAPx2_ASAP7_75t_R FILLER_0_234_1239 ();
 FILLER_ASAP7_75t_R FILLER_0_234_1245 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_1247 ();
 FILLER_ASAP7_75t_R FILLER_0_234_1258 ();
 DECAPx1_ASAP7_75t_R FILLER_0_234_1265 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_1269 ();
 FILLER_ASAP7_75t_R FILLER_0_234_1276 ();
 FILLER_ASAP7_75t_R FILLER_0_234_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_1290 ();
 FILLER_ASAP7_75t_R FILLER_0_234_1294 ();
 FILLER_ASAP7_75t_R FILLER_0_234_1302 ();
 DECAPx1_ASAP7_75t_R FILLER_0_234_1312 ();
 DECAPx1_ASAP7_75t_R FILLER_0_234_1326 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_1330 ();
 DECAPx6_ASAP7_75t_R FILLER_0_234_1337 ();
 FILLER_ASAP7_75t_R FILLER_0_234_1351 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_1353 ();
 FILLER_ASAP7_75t_R FILLER_0_234_1360 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_1362 ();
 DECAPx2_ASAP7_75t_R FILLER_0_234_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_234_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234_1381 ();
 DECAPx6_ASAP7_75t_R FILLER_0_235_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_235_16 ();
 FILLER_ASAP7_75t_R FILLER_0_235_23 ();
 FILLER_ASAP7_75t_R FILLER_0_235_35 ();
 DECAPx1_ASAP7_75t_R FILLER_0_235_43 ();
 DECAPx2_ASAP7_75t_R FILLER_0_235_54 ();
 DECAPx1_ASAP7_75t_R FILLER_0_235_67 ();
 FILLER_ASAP7_75t_R FILLER_0_235_91 ();
 FILLER_ASAP7_75t_R FILLER_0_235_98 ();
 DECAPx1_ASAP7_75t_R FILLER_0_235_106 ();
 FILLER_ASAP7_75t_R FILLER_0_235_116 ();
 FILLER_ASAP7_75t_R FILLER_0_235_124 ();
 FILLER_ASAP7_75t_R FILLER_0_235_132 ();
 DECAPx6_ASAP7_75t_R FILLER_0_235_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_235_155 ();
 FILLER_ASAP7_75t_R FILLER_0_235_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_235_168 ();
 DECAPx4_ASAP7_75t_R FILLER_0_235_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_235_199 ();
 DECAPx1_ASAP7_75t_R FILLER_0_235_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_235_216 ();
 FILLER_ASAP7_75t_R FILLER_0_235_239 ();
 FILLER_ASAP7_75t_R FILLER_0_235_269 ();
 DECAPx2_ASAP7_75t_R FILLER_0_235_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_235_287 ();
 DECAPx2_ASAP7_75t_R FILLER_0_235_294 ();
 FILLER_ASAP7_75t_R FILLER_0_235_306 ();
 FILLER_ASAP7_75t_R FILLER_0_235_324 ();
 DECAPx2_ASAP7_75t_R FILLER_0_235_332 ();
 FILLER_ASAP7_75t_R FILLER_0_235_338 ();
 FILLER_ASAP7_75t_R FILLER_0_235_345 ();
 FILLER_ASAP7_75t_R FILLER_0_235_357 ();
 DECAPx2_ASAP7_75t_R FILLER_0_235_369 ();
 DECAPx2_ASAP7_75t_R FILLER_0_235_383 ();
 DECAPx2_ASAP7_75t_R FILLER_0_235_409 ();
 FILLER_ASAP7_75t_R FILLER_0_235_415 ();
 DECAPx10_ASAP7_75t_R FILLER_0_235_427 ();
 FILLER_ASAP7_75t_R FILLER_0_235_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_235_451 ();
 DECAPx4_ASAP7_75t_R FILLER_0_235_458 ();
 FILLER_ASAP7_75t_R FILLER_0_235_468 ();
 FILLER_ASAP7_75t_R FILLER_0_235_476 ();
 DECAPx4_ASAP7_75t_R FILLER_0_235_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_235_499 ();
 DECAPx2_ASAP7_75t_R FILLER_0_235_506 ();
 FILLER_ASAP7_75t_R FILLER_0_235_512 ();
 DECAPx2_ASAP7_75t_R FILLER_0_235_526 ();
 FILLER_ASAP7_75t_R FILLER_0_235_532 ();
 DECAPx1_ASAP7_75t_R FILLER_0_235_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_235_549 ();
 DECAPx1_ASAP7_75t_R FILLER_0_235_556 ();
 FILLER_ASAP7_75t_R FILLER_0_235_580 ();
 FILLER_ASAP7_75t_R FILLER_0_235_592 ();
 DECAPx2_ASAP7_75t_R FILLER_0_235_600 ();
 DECAPx6_ASAP7_75t_R FILLER_0_235_622 ();
 DECAPx1_ASAP7_75t_R FILLER_0_235_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_235_640 ();
 FILLER_ASAP7_75t_R FILLER_0_235_647 ();
 DECAPx2_ASAP7_75t_R FILLER_0_235_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_235_666 ();
 FILLER_ASAP7_75t_R FILLER_0_235_673 ();
 DECAPx6_ASAP7_75t_R FILLER_0_235_681 ();
 FILLER_ASAP7_75t_R FILLER_0_235_695 ();
 DECAPx2_ASAP7_75t_R FILLER_0_235_705 ();
 FILLER_ASAP7_75t_R FILLER_0_235_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_235_713 ();
 DECAPx6_ASAP7_75t_R FILLER_0_235_724 ();
 DECAPx6_ASAP7_75t_R FILLER_0_235_748 ();
 DECAPx1_ASAP7_75t_R FILLER_0_235_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_235_766 ();
 FILLER_ASAP7_75t_R FILLER_0_235_779 ();
 DECAPx10_ASAP7_75t_R FILLER_0_235_793 ();
 FILLER_ASAP7_75t_R FILLER_0_235_815 ();
 FILLER_ASAP7_75t_R FILLER_0_235_837 ();
 DECAPx6_ASAP7_75t_R FILLER_0_235_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_235_860 ();
 FILLER_ASAP7_75t_R FILLER_0_235_867 ();
 FILLER_ASAP7_75t_R FILLER_0_235_875 ();
 FILLER_ASAP7_75t_R FILLER_0_235_883 ();
 DECAPx1_ASAP7_75t_R FILLER_0_235_891 ();
 DECAPx4_ASAP7_75t_R FILLER_0_235_915 ();
 DECAPx6_ASAP7_75t_R FILLER_0_235_927 ();
 DECAPx2_ASAP7_75t_R FILLER_0_235_941 ();
 DECAPx2_ASAP7_75t_R FILLER_0_235_953 ();
 FILLER_ASAP7_75t_R FILLER_0_235_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_235_961 ();
 FILLER_ASAP7_75t_R FILLER_0_235_977 ();
 DECAPx2_ASAP7_75t_R FILLER_0_235_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_235_992 ();
 DECAPx1_ASAP7_75t_R FILLER_0_235_1003 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_235_1007 ();
 FILLER_ASAP7_75t_R FILLER_0_235_1018 ();
 FILLER_ASAP7_75t_R FILLER_0_235_1032 ();
 FILLER_ASAP7_75t_R FILLER_0_235_1044 ();
 FILLER_ASAP7_75t_R FILLER_0_235_1052 ();
 DECAPx2_ASAP7_75t_R FILLER_0_235_1060 ();
 DECAPx2_ASAP7_75t_R FILLER_0_235_1074 ();
 FILLER_ASAP7_75t_R FILLER_0_235_1080 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_235_1082 ();
 FILLER_ASAP7_75t_R FILLER_0_235_1089 ();
 FILLER_ASAP7_75t_R FILLER_0_235_1097 ();
 DECAPx6_ASAP7_75t_R FILLER_0_235_1109 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_235_1123 ();
 DECAPx6_ASAP7_75t_R FILLER_0_235_1134 ();
 FILLER_ASAP7_75t_R FILLER_0_235_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_235_1150 ();
 FILLER_ASAP7_75t_R FILLER_0_235_1161 ();
 DECAPx2_ASAP7_75t_R FILLER_0_235_1169 ();
 FILLER_ASAP7_75t_R FILLER_0_235_1181 ();
 FILLER_ASAP7_75t_R FILLER_0_235_1201 ();
 FILLER_ASAP7_75t_R FILLER_0_235_1213 ();
 FILLER_ASAP7_75t_R FILLER_0_235_1223 ();
 FILLER_ASAP7_75t_R FILLER_0_235_1230 ();
 FILLER_ASAP7_75t_R FILLER_0_235_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_235_1240 ();
 FILLER_ASAP7_75t_R FILLER_0_235_1251 ();
 FILLER_ASAP7_75t_R FILLER_0_235_1271 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_235_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_0_235_1286 ();
 FILLER_ASAP7_75t_R FILLER_0_235_1292 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_235_1294 ();
 FILLER_ASAP7_75t_R FILLER_0_235_1301 ();
 FILLER_ASAP7_75t_R FILLER_0_235_1310 ();
 DECAPx2_ASAP7_75t_R FILLER_0_235_1319 ();
 DECAPx2_ASAP7_75t_R FILLER_0_235_1328 ();
 FILLER_ASAP7_75t_R FILLER_0_235_1340 ();
 DECAPx2_ASAP7_75t_R FILLER_0_235_1345 ();
 FILLER_ASAP7_75t_R FILLER_0_235_1351 ();
 FILLER_ASAP7_75t_R FILLER_0_235_1359 ();
 DECAPx6_ASAP7_75t_R FILLER_0_235_1364 ();
 DECAPx1_ASAP7_75t_R FILLER_0_235_1378 ();
 DECAPx2_ASAP7_75t_R FILLER_0_236_2 ();
 FILLER_ASAP7_75t_R FILLER_0_236_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_10 ();
 FILLER_ASAP7_75t_R FILLER_0_236_17 ();
 DECAPx4_ASAP7_75t_R FILLER_0_236_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_35 ();
 DECAPx6_ASAP7_75t_R FILLER_0_236_42 ();
 DECAPx2_ASAP7_75t_R FILLER_0_236_56 ();
 FILLER_ASAP7_75t_R FILLER_0_236_68 ();
 FILLER_ASAP7_75t_R FILLER_0_236_76 ();
 DECAPx2_ASAP7_75t_R FILLER_0_236_85 ();
 FILLER_ASAP7_75t_R FILLER_0_236_91 ();
 DECAPx2_ASAP7_75t_R FILLER_0_236_105 ();
 FILLER_ASAP7_75t_R FILLER_0_236_121 ();
 FILLER_ASAP7_75t_R FILLER_0_236_129 ();
 FILLER_ASAP7_75t_R FILLER_0_236_136 ();
 DECAPx6_ASAP7_75t_R FILLER_0_236_141 ();
 DECAPx1_ASAP7_75t_R FILLER_0_236_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_159 ();
 DECAPx1_ASAP7_75t_R FILLER_0_236_166 ();
 FILLER_ASAP7_75t_R FILLER_0_236_180 ();
 FILLER_ASAP7_75t_R FILLER_0_236_190 ();
 FILLER_ASAP7_75t_R FILLER_0_236_198 ();
 DECAPx6_ASAP7_75t_R FILLER_0_236_205 ();
 DECAPx2_ASAP7_75t_R FILLER_0_236_219 ();
 FILLER_ASAP7_75t_R FILLER_0_236_230 ();
 FILLER_ASAP7_75t_R FILLER_0_236_238 ();
 DECAPx1_ASAP7_75t_R FILLER_0_236_250 ();
 DECAPx1_ASAP7_75t_R FILLER_0_236_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_276 ();
 FILLER_ASAP7_75t_R FILLER_0_236_287 ();
 FILLER_ASAP7_75t_R FILLER_0_236_295 ();
 DECAPx2_ASAP7_75t_R FILLER_0_236_303 ();
 FILLER_ASAP7_75t_R FILLER_0_236_309 ();
 DECAPx2_ASAP7_75t_R FILLER_0_236_322 ();
 FILLER_ASAP7_75t_R FILLER_0_236_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_330 ();
 DECAPx2_ASAP7_75t_R FILLER_0_236_341 ();
 FILLER_ASAP7_75t_R FILLER_0_236_355 ();
 DECAPx2_ASAP7_75t_R FILLER_0_236_364 ();
 FILLER_ASAP7_75t_R FILLER_0_236_390 ();
 DECAPx4_ASAP7_75t_R FILLER_0_236_402 ();
 FILLER_ASAP7_75t_R FILLER_0_236_412 ();
 FILLER_ASAP7_75t_R FILLER_0_236_424 ();
 FILLER_ASAP7_75t_R FILLER_0_236_436 ();
 DECAPx2_ASAP7_75t_R FILLER_0_236_444 ();
 FILLER_ASAP7_75t_R FILLER_0_236_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_452 ();
 FILLER_ASAP7_75t_R FILLER_0_236_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_461 ();
 DECAPx6_ASAP7_75t_R FILLER_0_236_464 ();
 FILLER_ASAP7_75t_R FILLER_0_236_478 ();
 DECAPx6_ASAP7_75t_R FILLER_0_236_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_236_506 ();
 DECAPx10_ASAP7_75t_R FILLER_0_236_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_550 ();
 DECAPx1_ASAP7_75t_R FILLER_0_236_561 ();
 DECAPx2_ASAP7_75t_R FILLER_0_236_576 ();
 FILLER_ASAP7_75t_R FILLER_0_236_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_584 ();
 DECAPx2_ASAP7_75t_R FILLER_0_236_593 ();
 FILLER_ASAP7_75t_R FILLER_0_236_599 ();
 FILLER_ASAP7_75t_R FILLER_0_236_609 ();
 DECAPx2_ASAP7_75t_R FILLER_0_236_619 ();
 FILLER_ASAP7_75t_R FILLER_0_236_625 ();
 DECAPx2_ASAP7_75t_R FILLER_0_236_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_645 ();
 DECAPx1_ASAP7_75t_R FILLER_0_236_649 ();
 DECAPx1_ASAP7_75t_R FILLER_0_236_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_665 ();
 FILLER_ASAP7_75t_R FILLER_0_236_674 ();
 FILLER_ASAP7_75t_R FILLER_0_236_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_688 ();
 FILLER_ASAP7_75t_R FILLER_0_236_701 ();
 DECAPx2_ASAP7_75t_R FILLER_0_236_709 ();
 FILLER_ASAP7_75t_R FILLER_0_236_735 ();
 FILLER_ASAP7_75t_R FILLER_0_236_745 ();
 DECAPx4_ASAP7_75t_R FILLER_0_236_753 ();
 FILLER_ASAP7_75t_R FILLER_0_236_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_765 ();
 FILLER_ASAP7_75t_R FILLER_0_236_778 ();
 FILLER_ASAP7_75t_R FILLER_0_236_801 ();
 FILLER_ASAP7_75t_R FILLER_0_236_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_826 ();
 FILLER_ASAP7_75t_R FILLER_0_236_832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_236_839 ();
 DECAPx1_ASAP7_75t_R FILLER_0_236_861 ();
 DECAPx4_ASAP7_75t_R FILLER_0_236_871 ();
 FILLER_ASAP7_75t_R FILLER_0_236_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_883 ();
 FILLER_ASAP7_75t_R FILLER_0_236_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_896 ();
 DECAPx4_ASAP7_75t_R FILLER_0_236_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_914 ();
 DECAPx6_ASAP7_75t_R FILLER_0_236_923 ();
 FILLER_ASAP7_75t_R FILLER_0_236_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_945 ();
 DECAPx6_ASAP7_75t_R FILLER_0_236_956 ();
 FILLER_ASAP7_75t_R FILLER_0_236_970 ();
 DECAPx4_ASAP7_75t_R FILLER_0_236_978 ();
 FILLER_ASAP7_75t_R FILLER_0_236_996 ();
 DECAPx1_ASAP7_75t_R FILLER_0_236_1006 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_1010 ();
 FILLER_ASAP7_75t_R FILLER_0_236_1022 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_1024 ();
 FILLER_ASAP7_75t_R FILLER_0_236_1035 ();
 FILLER_ASAP7_75t_R FILLER_0_236_1043 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_1045 ();
 DECAPx6_ASAP7_75t_R FILLER_0_236_1052 ();
 DECAPx2_ASAP7_75t_R FILLER_0_236_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_1072 ();
 FILLER_ASAP7_75t_R FILLER_0_236_1093 ();
 FILLER_ASAP7_75t_R FILLER_0_236_1101 ();
 DECAPx4_ASAP7_75t_R FILLER_0_236_1109 ();
 DECAPx1_ASAP7_75t_R FILLER_0_236_1123 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_1127 ();
 FILLER_ASAP7_75t_R FILLER_0_236_1138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_236_1145 ();
 FILLER_ASAP7_75t_R FILLER_0_236_1161 ();
 FILLER_ASAP7_75t_R FILLER_0_236_1171 ();
 DECAPx2_ASAP7_75t_R FILLER_0_236_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_1184 ();
 FILLER_ASAP7_75t_R FILLER_0_236_1193 ();
 FILLER_ASAP7_75t_R FILLER_0_236_1215 ();
 FILLER_ASAP7_75t_R FILLER_0_236_1223 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_1225 ();
 FILLER_ASAP7_75t_R FILLER_0_236_1232 ();
 DECAPx1_ASAP7_75t_R FILLER_0_236_1239 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_1243 ();
 FILLER_ASAP7_75t_R FILLER_0_236_1251 ();
 FILLER_ASAP7_75t_R FILLER_0_236_1263 ();
 FILLER_ASAP7_75t_R FILLER_0_236_1270 ();
 DECAPx4_ASAP7_75t_R FILLER_0_236_1283 ();
 FILLER_ASAP7_75t_R FILLER_0_236_1293 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_1295 ();
 FILLER_ASAP7_75t_R FILLER_0_236_1303 ();
 DECAPx4_ASAP7_75t_R FILLER_0_236_1311 ();
 FILLER_ASAP7_75t_R FILLER_0_236_1321 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236_1323 ();
 FILLER_ASAP7_75t_R FILLER_0_236_1330 ();
 FILLER_ASAP7_75t_R FILLER_0_236_1338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_236_1346 ();
 DECAPx2_ASAP7_75t_R FILLER_0_236_1374 ();
 FILLER_ASAP7_75t_R FILLER_0_236_1380 ();
 DECAPx4_ASAP7_75t_R FILLER_0_237_2 ();
 FILLER_ASAP7_75t_R FILLER_0_237_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_14 ();
 FILLER_ASAP7_75t_R FILLER_0_237_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_23 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_30 ();
 DECAPx10_ASAP7_75t_R FILLER_0_237_42 ();
 DECAPx1_ASAP7_75t_R FILLER_0_237_64 ();
 FILLER_ASAP7_75t_R FILLER_0_237_73 ();
 FILLER_ASAP7_75t_R FILLER_0_237_80 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_92 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_114 ();
 FILLER_ASAP7_75t_R FILLER_0_237_121 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_129 ();
 FILLER_ASAP7_75t_R FILLER_0_237_141 ();
 FILLER_ASAP7_75t_R FILLER_0_237_149 ();
 FILLER_ASAP7_75t_R FILLER_0_237_157 ();
 DECAPx6_ASAP7_75t_R FILLER_0_237_165 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_179 ();
 FILLER_ASAP7_75t_R FILLER_0_237_201 ();
 DECAPx6_ASAP7_75t_R FILLER_0_237_209 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_229 ();
 FILLER_ASAP7_75t_R FILLER_0_237_233 ();
 FILLER_ASAP7_75t_R FILLER_0_237_241 ();
 FILLER_ASAP7_75t_R FILLER_0_237_249 ();
 FILLER_ASAP7_75t_R FILLER_0_237_261 ();
 FILLER_ASAP7_75t_R FILLER_0_237_271 ();
 FILLER_ASAP7_75t_R FILLER_0_237_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_281 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_296 ();
 FILLER_ASAP7_75t_R FILLER_0_237_305 ();
 DECAPx1_ASAP7_75t_R FILLER_0_237_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_316 ();
 FILLER_ASAP7_75t_R FILLER_0_237_324 ();
 FILLER_ASAP7_75t_R FILLER_0_237_332 ();
 DECAPx1_ASAP7_75t_R FILLER_0_237_344 ();
 FILLER_ASAP7_75t_R FILLER_0_237_353 ();
 FILLER_ASAP7_75t_R FILLER_0_237_361 ();
 FILLER_ASAP7_75t_R FILLER_0_237_391 ();
 FILLER_ASAP7_75t_R FILLER_0_237_399 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_414 ();
 FILLER_ASAP7_75t_R FILLER_0_237_421 ();
 FILLER_ASAP7_75t_R FILLER_0_237_429 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_442 ();
 FILLER_ASAP7_75t_R FILLER_0_237_448 ();
 DECAPx1_ASAP7_75t_R FILLER_0_237_456 ();
 FILLER_ASAP7_75t_R FILLER_0_237_467 ();
 FILLER_ASAP7_75t_R FILLER_0_237_475 ();
 FILLER_ASAP7_75t_R FILLER_0_237_483 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_491 ();
 DECAPx6_ASAP7_75t_R FILLER_0_237_503 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_523 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_541 ();
 FILLER_ASAP7_75t_R FILLER_0_237_553 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_558 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_564 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_581 ();
 FILLER_ASAP7_75t_R FILLER_0_237_592 ();
 DECAPx10_ASAP7_75t_R FILLER_0_237_605 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_627 ();
 FILLER_ASAP7_75t_R FILLER_0_237_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_635 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_648 ();
 FILLER_ASAP7_75t_R FILLER_0_237_654 ();
 FILLER_ASAP7_75t_R FILLER_0_237_664 ();
 FILLER_ASAP7_75t_R FILLER_0_237_669 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_682 ();
 DECAPx1_ASAP7_75t_R FILLER_0_237_698 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_716 ();
 FILLER_ASAP7_75t_R FILLER_0_237_725 ();
 FILLER_ASAP7_75t_R FILLER_0_237_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_735 ();
 DECAPx4_ASAP7_75t_R FILLER_0_237_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_758 ();
 DECAPx6_ASAP7_75t_R FILLER_0_237_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_781 ();
 DECAPx4_ASAP7_75t_R FILLER_0_237_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_795 ();
 FILLER_ASAP7_75t_R FILLER_0_237_804 ();
 DECAPx4_ASAP7_75t_R FILLER_0_237_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_819 ();
 FILLER_ASAP7_75t_R FILLER_0_237_826 ();
 FILLER_ASAP7_75t_R FILLER_0_237_833 ();
 DECAPx6_ASAP7_75t_R FILLER_0_237_845 ();
 DECAPx1_ASAP7_75t_R FILLER_0_237_859 ();
 DECAPx4_ASAP7_75t_R FILLER_0_237_871 ();
 FILLER_ASAP7_75t_R FILLER_0_237_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_883 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_889 ();
 FILLER_ASAP7_75t_R FILLER_0_237_895 ();
 DECAPx1_ASAP7_75t_R FILLER_0_237_907 ();
 FILLER_ASAP7_75t_R FILLER_0_237_923 ();
 FILLER_ASAP7_75t_R FILLER_0_237_927 ();
 FILLER_ASAP7_75t_R FILLER_0_237_939 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_941 ();
 FILLER_ASAP7_75t_R FILLER_0_237_947 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_955 ();
 FILLER_ASAP7_75t_R FILLER_0_237_967 ();
 FILLER_ASAP7_75t_R FILLER_0_237_980 ();
 FILLER_ASAP7_75t_R FILLER_0_237_987 ();
 FILLER_ASAP7_75t_R FILLER_0_237_999 ();
 FILLER_ASAP7_75t_R FILLER_0_237_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_0_237_1018 ();
 FILLER_ASAP7_75t_R FILLER_0_237_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_1042 ();
 DECAPx10_ASAP7_75t_R FILLER_0_237_1049 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_1077 ();
 DECAPx1_ASAP7_75t_R FILLER_0_237_1084 ();
 DECAPx6_ASAP7_75t_R FILLER_0_237_1094 ();
 DECAPx1_ASAP7_75t_R FILLER_0_237_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_1112 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_1120 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_1126 ();
 DECAPx1_ASAP7_75t_R FILLER_0_237_1137 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_1141 ();
 DECAPx1_ASAP7_75t_R FILLER_0_237_1152 ();
 FILLER_ASAP7_75t_R FILLER_0_237_1174 ();
 FILLER_ASAP7_75t_R FILLER_0_237_1182 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_1190 ();
 FILLER_ASAP7_75t_R FILLER_0_237_1206 ();
 FILLER_ASAP7_75t_R FILLER_0_237_1214 ();
 FILLER_ASAP7_75t_R FILLER_0_237_1221 ();
 FILLER_ASAP7_75t_R FILLER_0_237_1226 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_1228 ();
 FILLER_ASAP7_75t_R FILLER_0_237_1235 ();
 FILLER_ASAP7_75t_R FILLER_0_237_1243 ();
 FILLER_ASAP7_75t_R FILLER_0_237_1253 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_1261 ();
 FILLER_ASAP7_75t_R FILLER_0_237_1267 ();
 FILLER_ASAP7_75t_R FILLER_0_237_1276 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_1284 ();
 FILLER_ASAP7_75t_R FILLER_0_237_1290 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_237_1299 ();
 DECAPx4_ASAP7_75t_R FILLER_0_237_1321 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_1331 ();
 DECAPx6_ASAP7_75t_R FILLER_0_237_1338 ();
 DECAPx1_ASAP7_75t_R FILLER_0_237_1352 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237_1356 ();
 FILLER_ASAP7_75t_R FILLER_0_237_1363 ();
 DECAPx2_ASAP7_75t_R FILLER_0_237_1376 ();
 DECAPx4_ASAP7_75t_R FILLER_0_238_2 ();
 FILLER_ASAP7_75t_R FILLER_0_238_12 ();
 FILLER_ASAP7_75t_R FILLER_0_238_20 ();
 DECAPx4_ASAP7_75t_R FILLER_0_238_32 ();
 FILLER_ASAP7_75t_R FILLER_0_238_48 ();
 FILLER_ASAP7_75t_R FILLER_0_238_56 ();
 FILLER_ASAP7_75t_R FILLER_0_238_64 ();
 DECAPx2_ASAP7_75t_R FILLER_0_238_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_83 ();
 FILLER_ASAP7_75t_R FILLER_0_238_89 ();
 FILLER_ASAP7_75t_R FILLER_0_238_101 ();
 FILLER_ASAP7_75t_R FILLER_0_238_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_115 ();
 FILLER_ASAP7_75t_R FILLER_0_238_122 ();
 DECAPx1_ASAP7_75t_R FILLER_0_238_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_134 ();
 FILLER_ASAP7_75t_R FILLER_0_238_143 ();
 DECAPx2_ASAP7_75t_R FILLER_0_238_148 ();
 DECAPx2_ASAP7_75t_R FILLER_0_238_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_238_191 ();
 DECAPx6_ASAP7_75t_R FILLER_0_238_213 ();
 DECAPx2_ASAP7_75t_R FILLER_0_238_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_233 ();
 FILLER_ASAP7_75t_R FILLER_0_238_244 ();
 FILLER_ASAP7_75t_R FILLER_0_238_256 ();
 FILLER_ASAP7_75t_R FILLER_0_238_268 ();
 FILLER_ASAP7_75t_R FILLER_0_238_278 ();
 FILLER_ASAP7_75t_R FILLER_0_238_286 ();
 FILLER_ASAP7_75t_R FILLER_0_238_294 ();
 DECAPx2_ASAP7_75t_R FILLER_0_238_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_307 ();
 DECAPx4_ASAP7_75t_R FILLER_0_238_314 ();
 FILLER_ASAP7_75t_R FILLER_0_238_330 ();
 DECAPx4_ASAP7_75t_R FILLER_0_238_339 ();
 FILLER_ASAP7_75t_R FILLER_0_238_349 ();
 FILLER_ASAP7_75t_R FILLER_0_238_354 ();
 FILLER_ASAP7_75t_R FILLER_0_238_362 ();
 DECAPx10_ASAP7_75t_R FILLER_0_238_369 ();
 DECAPx10_ASAP7_75t_R FILLER_0_238_391 ();
 FILLER_ASAP7_75t_R FILLER_0_238_413 ();
 FILLER_ASAP7_75t_R FILLER_0_238_421 ();
 DECAPx2_ASAP7_75t_R FILLER_0_238_430 ();
 FILLER_ASAP7_75t_R FILLER_0_238_436 ();
 DECAPx1_ASAP7_75t_R FILLER_0_238_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_238_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_461 ();
 DECAPx1_ASAP7_75t_R FILLER_0_238_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_468 ();
 DECAPx4_ASAP7_75t_R FILLER_0_238_475 ();
 FILLER_ASAP7_75t_R FILLER_0_238_491 ();
 FILLER_ASAP7_75t_R FILLER_0_238_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_502 ();
 FILLER_ASAP7_75t_R FILLER_0_238_513 ();
 FILLER_ASAP7_75t_R FILLER_0_238_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_535 ();
 DECAPx1_ASAP7_75t_R FILLER_0_238_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_548 ();
 DECAPx10_ASAP7_75t_R FILLER_0_238_560 ();
 DECAPx1_ASAP7_75t_R FILLER_0_238_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_238_592 ();
 DECAPx10_ASAP7_75t_R FILLER_0_238_614 ();
 DECAPx1_ASAP7_75t_R FILLER_0_238_636 ();
 DECAPx2_ASAP7_75t_R FILLER_0_238_646 ();
 FILLER_ASAP7_75t_R FILLER_0_238_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_238_661 ();
 FILLER_ASAP7_75t_R FILLER_0_238_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_677 ();
 DECAPx10_ASAP7_75t_R FILLER_0_238_688 ();
 DECAPx2_ASAP7_75t_R FILLER_0_238_710 ();
 DECAPx1_ASAP7_75t_R FILLER_0_238_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_726 ();
 FILLER_ASAP7_75t_R FILLER_0_238_739 ();
 FILLER_ASAP7_75t_R FILLER_0_238_749 ();
 DECAPx1_ASAP7_75t_R FILLER_0_238_759 ();
 FILLER_ASAP7_75t_R FILLER_0_238_766 ();
 FILLER_ASAP7_75t_R FILLER_0_238_776 ();
 DECAPx1_ASAP7_75t_R FILLER_0_238_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_790 ();
 FILLER_ASAP7_75t_R FILLER_0_238_801 ();
 DECAPx1_ASAP7_75t_R FILLER_0_238_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_817 ();
 DECAPx1_ASAP7_75t_R FILLER_0_238_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_832 ();
 FILLER_ASAP7_75t_R FILLER_0_238_839 ();
 DECAPx1_ASAP7_75t_R FILLER_0_238_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_855 ();
 FILLER_ASAP7_75t_R FILLER_0_238_868 ();
 FILLER_ASAP7_75t_R FILLER_0_238_880 ();
 DECAPx4_ASAP7_75t_R FILLER_0_238_892 ();
 FILLER_ASAP7_75t_R FILLER_0_238_912 ();
 FILLER_ASAP7_75t_R FILLER_0_238_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_922 ();
 DECAPx4_ASAP7_75t_R FILLER_0_238_929 ();
 FILLER_ASAP7_75t_R FILLER_0_238_945 ();
 DECAPx1_ASAP7_75t_R FILLER_0_238_953 ();
 FILLER_ASAP7_75t_R FILLER_0_238_962 ();
 DECAPx1_ASAP7_75t_R FILLER_0_238_970 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_974 ();
 FILLER_ASAP7_75t_R FILLER_0_238_985 ();
 FILLER_ASAP7_75t_R FILLER_0_238_997 ();
 FILLER_ASAP7_75t_R FILLER_0_238_1005 ();
 DECAPx2_ASAP7_75t_R FILLER_0_238_1013 ();
 DECAPx2_ASAP7_75t_R FILLER_0_238_1027 ();
 FILLER_ASAP7_75t_R FILLER_0_238_1033 ();
 DECAPx1_ASAP7_75t_R FILLER_0_238_1045 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_1049 ();
 FILLER_ASAP7_75t_R FILLER_0_238_1060 ();
 FILLER_ASAP7_75t_R FILLER_0_238_1069 ();
 DECAPx1_ASAP7_75t_R FILLER_0_238_1077 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_1081 ();
 DECAPx2_ASAP7_75t_R FILLER_0_238_1088 ();
 FILLER_ASAP7_75t_R FILLER_0_238_1094 ();
 DECAPx2_ASAP7_75t_R FILLER_0_238_1102 ();
 FILLER_ASAP7_75t_R FILLER_0_238_1108 ();
 DECAPx1_ASAP7_75t_R FILLER_0_238_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_1134 ();
 FILLER_ASAP7_75t_R FILLER_0_238_1139 ();
 DECAPx2_ASAP7_75t_R FILLER_0_238_1146 ();
 FILLER_ASAP7_75t_R FILLER_0_238_1152 ();
 FILLER_ASAP7_75t_R FILLER_0_238_1164 ();
 FILLER_ASAP7_75t_R FILLER_0_238_1172 ();
 FILLER_ASAP7_75t_R FILLER_0_238_1180 ();
 FILLER_ASAP7_75t_R FILLER_0_238_1188 ();
 FILLER_ASAP7_75t_R FILLER_0_238_1196 ();
 FILLER_ASAP7_75t_R FILLER_0_238_1204 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_1206 ();
 DECAPx6_ASAP7_75t_R FILLER_0_238_1214 ();
 DECAPx1_ASAP7_75t_R FILLER_0_238_1228 ();
 FILLER_ASAP7_75t_R FILLER_0_238_1238 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_1240 ();
 FILLER_ASAP7_75t_R FILLER_0_238_1247 ();
 DECAPx1_ASAP7_75t_R FILLER_0_238_1257 ();
 DECAPx2_ASAP7_75t_R FILLER_0_238_1271 ();
 FILLER_ASAP7_75t_R FILLER_0_238_1277 ();
 DECAPx2_ASAP7_75t_R FILLER_0_238_1285 ();
 FILLER_ASAP7_75t_R FILLER_0_238_1291 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_1293 ();
 FILLER_ASAP7_75t_R FILLER_0_238_1300 ();
 DECAPx4_ASAP7_75t_R FILLER_0_238_1307 ();
 FILLER_ASAP7_75t_R FILLER_0_238_1317 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238_1319 ();
 DECAPx1_ASAP7_75t_R FILLER_0_238_1328 ();
 FILLER_ASAP7_75t_R FILLER_0_238_1338 ();
 DECAPx6_ASAP7_75t_R FILLER_0_238_1346 ();
 DECAPx1_ASAP7_75t_R FILLER_0_238_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_238_1376 ();
 FILLER_ASAP7_75t_R FILLER_0_239_2 ();
 FILLER_ASAP7_75t_R FILLER_0_239_20 ();
 FILLER_ASAP7_75t_R FILLER_0_239_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_29 ();
 FILLER_ASAP7_75t_R FILLER_0_239_40 ();
 FILLER_ASAP7_75t_R FILLER_0_239_48 ();
 DECAPx1_ASAP7_75t_R FILLER_0_239_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_60 ();
 FILLER_ASAP7_75t_R FILLER_0_239_64 ();
 DECAPx1_ASAP7_75t_R FILLER_0_239_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_75 ();
 DECAPx2_ASAP7_75t_R FILLER_0_239_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_102 ();
 FILLER_ASAP7_75t_R FILLER_0_239_113 ();
 FILLER_ASAP7_75t_R FILLER_0_239_125 ();
 FILLER_ASAP7_75t_R FILLER_0_239_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_132 ();
 FILLER_ASAP7_75t_R FILLER_0_239_140 ();
 FILLER_ASAP7_75t_R FILLER_0_239_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_150 ();
 FILLER_ASAP7_75t_R FILLER_0_239_159 ();
 FILLER_ASAP7_75t_R FILLER_0_239_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_169 ();
 FILLER_ASAP7_75t_R FILLER_0_239_177 ();
 DECAPx10_ASAP7_75t_R FILLER_0_239_185 ();
 DECAPx10_ASAP7_75t_R FILLER_0_239_215 ();
 DECAPx4_ASAP7_75t_R FILLER_0_239_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_247 ();
 DECAPx1_ASAP7_75t_R FILLER_0_239_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_274 ();
 FILLER_ASAP7_75t_R FILLER_0_239_281 ();
 FILLER_ASAP7_75t_R FILLER_0_239_289 ();
 FILLER_ASAP7_75t_R FILLER_0_239_295 ();
 FILLER_ASAP7_75t_R FILLER_0_239_303 ();
 DECAPx6_ASAP7_75t_R FILLER_0_239_311 ();
 DECAPx2_ASAP7_75t_R FILLER_0_239_325 ();
 DECAPx2_ASAP7_75t_R FILLER_0_239_337 ();
 FILLER_ASAP7_75t_R FILLER_0_239_343 ();
 DECAPx2_ASAP7_75t_R FILLER_0_239_351 ();
 DECAPx2_ASAP7_75t_R FILLER_0_239_363 ();
 FILLER_ASAP7_75t_R FILLER_0_239_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_371 ();
 FILLER_ASAP7_75t_R FILLER_0_239_378 ();
 DECAPx2_ASAP7_75t_R FILLER_0_239_388 ();
 FILLER_ASAP7_75t_R FILLER_0_239_394 ();
 FILLER_ASAP7_75t_R FILLER_0_239_402 ();
 FILLER_ASAP7_75t_R FILLER_0_239_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_412 ();
 DECAPx4_ASAP7_75t_R FILLER_0_239_416 ();
 DECAPx2_ASAP7_75t_R FILLER_0_239_432 ();
 FILLER_ASAP7_75t_R FILLER_0_239_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_440 ();
 DECAPx4_ASAP7_75t_R FILLER_0_239_449 ();
 DECAPx10_ASAP7_75t_R FILLER_0_239_466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_239_488 ();
 DECAPx1_ASAP7_75t_R FILLER_0_239_510 ();
 DECAPx2_ASAP7_75t_R FILLER_0_239_534 ();
 FILLER_ASAP7_75t_R FILLER_0_239_540 ();
 FILLER_ASAP7_75t_R FILLER_0_239_550 ();
 FILLER_ASAP7_75t_R FILLER_0_239_556 ();
 FILLER_ASAP7_75t_R FILLER_0_239_561 ();
 DECAPx1_ASAP7_75t_R FILLER_0_239_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_579 ();
 DECAPx4_ASAP7_75t_R FILLER_0_239_588 ();
 FILLER_ASAP7_75t_R FILLER_0_239_598 ();
 FILLER_ASAP7_75t_R FILLER_0_239_612 ();
 DECAPx2_ASAP7_75t_R FILLER_0_239_617 ();
 FILLER_ASAP7_75t_R FILLER_0_239_623 ();
 FILLER_ASAP7_75t_R FILLER_0_239_633 ();
 DECAPx2_ASAP7_75t_R FILLER_0_239_645 ();
 FILLER_ASAP7_75t_R FILLER_0_239_651 ();
 DECAPx4_ASAP7_75t_R FILLER_0_239_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_673 ();
 DECAPx1_ASAP7_75t_R FILLER_0_239_685 ();
 DECAPx6_ASAP7_75t_R FILLER_0_239_700 ();
 FILLER_ASAP7_75t_R FILLER_0_239_714 ();
 DECAPx4_ASAP7_75t_R FILLER_0_239_728 ();
 FILLER_ASAP7_75t_R FILLER_0_239_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_740 ();
 DECAPx2_ASAP7_75t_R FILLER_0_239_753 ();
 FILLER_ASAP7_75t_R FILLER_0_239_759 ();
 DECAPx2_ASAP7_75t_R FILLER_0_239_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_777 ();
 FILLER_ASAP7_75t_R FILLER_0_239_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_788 ();
 FILLER_ASAP7_75t_R FILLER_0_239_800 ();
 DECAPx6_ASAP7_75t_R FILLER_0_239_813 ();
 FILLER_ASAP7_75t_R FILLER_0_239_827 ();
 FILLER_ASAP7_75t_R FILLER_0_239_839 ();
 DECAPx4_ASAP7_75t_R FILLER_0_239_851 ();
 FILLER_ASAP7_75t_R FILLER_0_239_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_863 ();
 FILLER_ASAP7_75t_R FILLER_0_239_880 ();
 FILLER_ASAP7_75t_R FILLER_0_239_902 ();
 FILLER_ASAP7_75t_R FILLER_0_239_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_913 ();
 DECAPx1_ASAP7_75t_R FILLER_0_239_921 ();
 DECAPx6_ASAP7_75t_R FILLER_0_239_927 ();
 DECAPx1_ASAP7_75t_R FILLER_0_239_941 ();
 DECAPx1_ASAP7_75t_R FILLER_0_239_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_959 ();
 FILLER_ASAP7_75t_R FILLER_0_239_970 ();
 DECAPx4_ASAP7_75t_R FILLER_0_239_982 ();
 FILLER_ASAP7_75t_R FILLER_0_239_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_994 ();
 DECAPx1_ASAP7_75t_R FILLER_0_239_1000 ();
 DECAPx1_ASAP7_75t_R FILLER_0_239_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_1018 ();
 FILLER_ASAP7_75t_R FILLER_0_239_1025 ();
 DECAPx2_ASAP7_75t_R FILLER_0_239_1033 ();
 FILLER_ASAP7_75t_R FILLER_0_239_1039 ();
 DECAPx1_ASAP7_75t_R FILLER_0_239_1047 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_1051 ();
 DECAPx1_ASAP7_75t_R FILLER_0_239_1058 ();
 DECAPx1_ASAP7_75t_R FILLER_0_239_1068 ();
 DECAPx1_ASAP7_75t_R FILLER_0_239_1092 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_1096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_239_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_1130 ();
 DECAPx10_ASAP7_75t_R FILLER_0_239_1141 ();
 DECAPx10_ASAP7_75t_R FILLER_0_239_1163 ();
 DECAPx6_ASAP7_75t_R FILLER_0_239_1185 ();
 FILLER_ASAP7_75t_R FILLER_0_239_1199 ();
 FILLER_ASAP7_75t_R FILLER_0_239_1207 ();
 FILLER_ASAP7_75t_R FILLER_0_239_1215 ();
 FILLER_ASAP7_75t_R FILLER_0_239_1223 ();
 FILLER_ASAP7_75t_R FILLER_0_239_1231 ();
 FILLER_ASAP7_75t_R FILLER_0_239_1239 ();
 FILLER_ASAP7_75t_R FILLER_0_239_1247 ();
 FILLER_ASAP7_75t_R FILLER_0_239_1254 ();
 DECAPx4_ASAP7_75t_R FILLER_0_239_1278 ();
 FILLER_ASAP7_75t_R FILLER_0_239_1294 ();
 FILLER_ASAP7_75t_R FILLER_0_239_1307 ();
 FILLER_ASAP7_75t_R FILLER_0_239_1316 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_1318 ();
 DECAPx1_ASAP7_75t_R FILLER_0_239_1325 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_1329 ();
 FILLER_ASAP7_75t_R FILLER_0_239_1342 ();
 FILLER_ASAP7_75t_R FILLER_0_239_1350 ();
 DECAPx1_ASAP7_75t_R FILLER_0_239_1358 ();
 FILLER_ASAP7_75t_R FILLER_0_239_1370 ();
 DECAPx1_ASAP7_75t_R FILLER_0_239_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239_1381 ();
 DECAPx6_ASAP7_75t_R FILLER_0_240_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_240_16 ();
 DECAPx6_ASAP7_75t_R FILLER_0_240_28 ();
 DECAPx1_ASAP7_75t_R FILLER_0_240_42 ();
 DECAPx2_ASAP7_75t_R FILLER_0_240_52 ();
 FILLER_ASAP7_75t_R FILLER_0_240_58 ();
 DECAPx2_ASAP7_75t_R FILLER_0_240_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_78 ();
 FILLER_ASAP7_75t_R FILLER_0_240_82 ();
 FILLER_ASAP7_75t_R FILLER_0_240_94 ();
 FILLER_ASAP7_75t_R FILLER_0_240_114 ();
 DECAPx1_ASAP7_75t_R FILLER_0_240_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_126 ();
 FILLER_ASAP7_75t_R FILLER_0_240_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_135 ();
 FILLER_ASAP7_75t_R FILLER_0_240_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_158 ();
 DECAPx2_ASAP7_75t_R FILLER_0_240_165 ();
 FILLER_ASAP7_75t_R FILLER_0_240_177 ();
 FILLER_ASAP7_75t_R FILLER_0_240_185 ();
 DECAPx4_ASAP7_75t_R FILLER_0_240_193 ();
 FILLER_ASAP7_75t_R FILLER_0_240_203 ();
 DECAPx10_ASAP7_75t_R FILLER_0_240_217 ();
 DECAPx1_ASAP7_75t_R FILLER_0_240_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_243 ();
 FILLER_ASAP7_75t_R FILLER_0_240_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_254 ();
 DECAPx1_ASAP7_75t_R FILLER_0_240_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_271 ();
 FILLER_ASAP7_75t_R FILLER_0_240_282 ();
 FILLER_ASAP7_75t_R FILLER_0_240_295 ();
 FILLER_ASAP7_75t_R FILLER_0_240_303 ();
 DECAPx6_ASAP7_75t_R FILLER_0_240_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_324 ();
 FILLER_ASAP7_75t_R FILLER_0_240_331 ();
 DECAPx1_ASAP7_75t_R FILLER_0_240_339 ();
 DECAPx1_ASAP7_75t_R FILLER_0_240_353 ();
 DECAPx1_ASAP7_75t_R FILLER_0_240_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_367 ();
 FILLER_ASAP7_75t_R FILLER_0_240_374 ();
 DECAPx2_ASAP7_75t_R FILLER_0_240_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_385 ();
 FILLER_ASAP7_75t_R FILLER_0_240_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_391 ();
 FILLER_ASAP7_75t_R FILLER_0_240_398 ();
 DECAPx2_ASAP7_75t_R FILLER_0_240_406 ();
 FILLER_ASAP7_75t_R FILLER_0_240_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_422 ();
 FILLER_ASAP7_75t_R FILLER_0_240_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_431 ();
 FILLER_ASAP7_75t_R FILLER_0_240_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_439 ();
 DECAPx6_ASAP7_75t_R FILLER_0_240_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_461 ();
 DECAPx2_ASAP7_75t_R FILLER_0_240_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_470 ();
 FILLER_ASAP7_75t_R FILLER_0_240_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_479 ();
 FILLER_ASAP7_75t_R FILLER_0_240_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_490 ();
 FILLER_ASAP7_75t_R FILLER_0_240_497 ();
 DECAPx6_ASAP7_75t_R FILLER_0_240_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_523 ();
 DECAPx2_ASAP7_75t_R FILLER_0_240_534 ();
 FILLER_ASAP7_75t_R FILLER_0_240_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_542 ();
 FILLER_ASAP7_75t_R FILLER_0_240_551 ();
 DECAPx2_ASAP7_75t_R FILLER_0_240_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_567 ();
 DECAPx2_ASAP7_75t_R FILLER_0_240_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_580 ();
 DECAPx10_ASAP7_75t_R FILLER_0_240_589 ();
 FILLER_ASAP7_75t_R FILLER_0_240_611 ();
 FILLER_ASAP7_75t_R FILLER_0_240_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_627 ();
 DECAPx1_ASAP7_75t_R FILLER_0_240_634 ();
 FILLER_ASAP7_75t_R FILLER_0_240_649 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_651 ();
 DECAPx2_ASAP7_75t_R FILLER_0_240_662 ();
 FILLER_ASAP7_75t_R FILLER_0_240_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_680 ();
 FILLER_ASAP7_75t_R FILLER_0_240_684 ();
 DECAPx1_ASAP7_75t_R FILLER_0_240_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_698 ();
 DECAPx6_ASAP7_75t_R FILLER_0_240_705 ();
 DECAPx1_ASAP7_75t_R FILLER_0_240_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_723 ();
 DECAPx2_ASAP7_75t_R FILLER_0_240_734 ();
 DECAPx4_ASAP7_75t_R FILLER_0_240_750 ();
 FILLER_ASAP7_75t_R FILLER_0_240_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_762 ();
 FILLER_ASAP7_75t_R FILLER_0_240_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_777 ();
 FILLER_ASAP7_75t_R FILLER_0_240_784 ();
 FILLER_ASAP7_75t_R FILLER_0_240_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_795 ();
 FILLER_ASAP7_75t_R FILLER_0_240_801 ();
 FILLER_ASAP7_75t_R FILLER_0_240_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_826 ();
 FILLER_ASAP7_75t_R FILLER_0_240_837 ();
 DECAPx2_ASAP7_75t_R FILLER_0_240_849 ();
 FILLER_ASAP7_75t_R FILLER_0_240_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_857 ();
 DECAPx6_ASAP7_75t_R FILLER_0_240_868 ();
 FILLER_ASAP7_75t_R FILLER_0_240_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_884 ();
 DECAPx1_ASAP7_75t_R FILLER_0_240_897 ();
 FILLER_ASAP7_75t_R FILLER_0_240_911 ();
 DECAPx1_ASAP7_75t_R FILLER_0_240_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_922 ();
 FILLER_ASAP7_75t_R FILLER_0_240_929 ();
 DECAPx4_ASAP7_75t_R FILLER_0_240_937 ();
 FILLER_ASAP7_75t_R FILLER_0_240_947 ();
 FILLER_ASAP7_75t_R FILLER_0_240_961 ();
 DECAPx6_ASAP7_75t_R FILLER_0_240_969 ();
 DECAPx2_ASAP7_75t_R FILLER_0_240_983 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_989 ();
 DECAPx1_ASAP7_75t_R FILLER_0_240_1000 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_1004 ();
 DECAPx2_ASAP7_75t_R FILLER_0_240_1015 ();
 FILLER_ASAP7_75t_R FILLER_0_240_1021 ();
 FILLER_ASAP7_75t_R FILLER_0_240_1043 ();
 DECAPx10_ASAP7_75t_R FILLER_0_240_1051 ();
 DECAPx4_ASAP7_75t_R FILLER_0_240_1073 ();
 DECAPx2_ASAP7_75t_R FILLER_0_240_1089 ();
 DECAPx2_ASAP7_75t_R FILLER_0_240_1101 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_1107 ();
 FILLER_ASAP7_75t_R FILLER_0_240_1120 ();
 FILLER_ASAP7_75t_R FILLER_0_240_1132 ();
 DECAPx4_ASAP7_75t_R FILLER_0_240_1144 ();
 DECAPx6_ASAP7_75t_R FILLER_0_240_1157 ();
 DECAPx1_ASAP7_75t_R FILLER_0_240_1171 ();
 DECAPx6_ASAP7_75t_R FILLER_0_240_1185 ();
 DECAPx6_ASAP7_75t_R FILLER_0_240_1219 ();
 DECAPx2_ASAP7_75t_R FILLER_0_240_1233 ();
 FILLER_ASAP7_75t_R FILLER_0_240_1249 ();
 FILLER_ASAP7_75t_R FILLER_0_240_1257 ();
 FILLER_ASAP7_75t_R FILLER_0_240_1269 ();
 FILLER_ASAP7_75t_R FILLER_0_240_1277 ();
 FILLER_ASAP7_75t_R FILLER_0_240_1285 ();
 FILLER_ASAP7_75t_R FILLER_0_240_1293 ();
 FILLER_ASAP7_75t_R FILLER_0_240_1301 ();
 DECAPx1_ASAP7_75t_R FILLER_0_240_1309 ();
 FILLER_ASAP7_75t_R FILLER_0_240_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_0_240_1332 ();
 DECAPx6_ASAP7_75t_R FILLER_0_240_1354 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240_1368 ();
 FILLER_ASAP7_75t_R FILLER_0_240_1375 ();
 FILLER_ASAP7_75t_R FILLER_0_240_1380 ();
 DECAPx2_ASAP7_75t_R FILLER_0_241_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_8 ();
 DECAPx1_ASAP7_75t_R FILLER_0_241_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_19 ();
 DECAPx4_ASAP7_75t_R FILLER_0_241_26 ();
 DECAPx2_ASAP7_75t_R FILLER_0_241_42 ();
 DECAPx4_ASAP7_75t_R FILLER_0_241_54 ();
 FILLER_ASAP7_75t_R FILLER_0_241_64 ();
 FILLER_ASAP7_75t_R FILLER_0_241_72 ();
 FILLER_ASAP7_75t_R FILLER_0_241_84 ();
 FILLER_ASAP7_75t_R FILLER_0_241_96 ();
 FILLER_ASAP7_75t_R FILLER_0_241_108 ();
 FILLER_ASAP7_75t_R FILLER_0_241_116 ();
 DECAPx1_ASAP7_75t_R FILLER_0_241_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_127 ();
 FILLER_ASAP7_75t_R FILLER_0_241_134 ();
 DECAPx2_ASAP7_75t_R FILLER_0_241_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_147 ();
 DECAPx6_ASAP7_75t_R FILLER_0_241_156 ();
 DECAPx2_ASAP7_75t_R FILLER_0_241_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_176 ();
 FILLER_ASAP7_75t_R FILLER_0_241_183 ();
 DECAPx10_ASAP7_75t_R FILLER_0_241_195 ();
 DECAPx10_ASAP7_75t_R FILLER_0_241_217 ();
 DECAPx2_ASAP7_75t_R FILLER_0_241_239 ();
 FILLER_ASAP7_75t_R FILLER_0_241_245 ();
 FILLER_ASAP7_75t_R FILLER_0_241_253 ();
 FILLER_ASAP7_75t_R FILLER_0_241_266 ();
 DECAPx1_ASAP7_75t_R FILLER_0_241_274 ();
 DECAPx2_ASAP7_75t_R FILLER_0_241_284 ();
 DECAPx1_ASAP7_75t_R FILLER_0_241_297 ();
 FILLER_ASAP7_75t_R FILLER_0_241_307 ();
 DECAPx10_ASAP7_75t_R FILLER_0_241_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_336 ();
 DECAPx4_ASAP7_75t_R FILLER_0_241_343 ();
 FILLER_ASAP7_75t_R FILLER_0_241_353 ();
 FILLER_ASAP7_75t_R FILLER_0_241_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_363 ();
 FILLER_ASAP7_75t_R FILLER_0_241_370 ();
 FILLER_ASAP7_75t_R FILLER_0_241_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_381 ();
 DECAPx4_ASAP7_75t_R FILLER_0_241_388 ();
 DECAPx1_ASAP7_75t_R FILLER_0_241_408 ();
 DECAPx4_ASAP7_75t_R FILLER_0_241_420 ();
 FILLER_ASAP7_75t_R FILLER_0_241_436 ();
 DECAPx2_ASAP7_75t_R FILLER_0_241_449 ();
 FILLER_ASAP7_75t_R FILLER_0_241_455 ();
 FILLER_ASAP7_75t_R FILLER_0_241_463 ();
 FILLER_ASAP7_75t_R FILLER_0_241_471 ();
 FILLER_ASAP7_75t_R FILLER_0_241_484 ();
 DECAPx4_ASAP7_75t_R FILLER_0_241_492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_241_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_241_530 ();
 DECAPx4_ASAP7_75t_R FILLER_0_241_552 ();
 FILLER_ASAP7_75t_R FILLER_0_241_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_564 ();
 FILLER_ASAP7_75t_R FILLER_0_241_577 ();
 FILLER_ASAP7_75t_R FILLER_0_241_585 ();
 FILLER_ASAP7_75t_R FILLER_0_241_593 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_595 ();
 FILLER_ASAP7_75t_R FILLER_0_241_608 ();
 FILLER_ASAP7_75t_R FILLER_0_241_622 ();
 DECAPx4_ASAP7_75t_R FILLER_0_241_630 ();
 FILLER_ASAP7_75t_R FILLER_0_241_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_642 ();
 DECAPx6_ASAP7_75t_R FILLER_0_241_655 ();
 DECAPx2_ASAP7_75t_R FILLER_0_241_679 ();
 FILLER_ASAP7_75t_R FILLER_0_241_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_687 ();
 FILLER_ASAP7_75t_R FILLER_0_241_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_693 ();
 DECAPx2_ASAP7_75t_R FILLER_0_241_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_705 ();
 FILLER_ASAP7_75t_R FILLER_0_241_716 ();
 DECAPx2_ASAP7_75t_R FILLER_0_241_724 ();
 FILLER_ASAP7_75t_R FILLER_0_241_730 ();
 DECAPx1_ASAP7_75t_R FILLER_0_241_744 ();
 DECAPx6_ASAP7_75t_R FILLER_0_241_758 ();
 DECAPx1_ASAP7_75t_R FILLER_0_241_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_776 ();
 DECAPx4_ASAP7_75t_R FILLER_0_241_785 ();
 DECAPx2_ASAP7_75t_R FILLER_0_241_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_804 ();
 DECAPx10_ASAP7_75t_R FILLER_0_241_808 ();
 DECAPx2_ASAP7_75t_R FILLER_0_241_830 ();
 FILLER_ASAP7_75t_R FILLER_0_241_840 ();
 FILLER_ASAP7_75t_R FILLER_0_241_852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_241_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_882 ();
 FILLER_ASAP7_75t_R FILLER_0_241_895 ();
 FILLER_ASAP7_75t_R FILLER_0_241_904 ();
 FILLER_ASAP7_75t_R FILLER_0_241_916 ();
 FILLER_ASAP7_75t_R FILLER_0_241_923 ();
 FILLER_ASAP7_75t_R FILLER_0_241_927 ();
 FILLER_ASAP7_75t_R FILLER_0_241_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_938 ();
 FILLER_ASAP7_75t_R FILLER_0_241_945 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_947 ();
 DECAPx2_ASAP7_75t_R FILLER_0_241_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_960 ();
 FILLER_ASAP7_75t_R FILLER_0_241_968 ();
 DECAPx1_ASAP7_75t_R FILLER_0_241_978 ();
 FILLER_ASAP7_75t_R FILLER_0_241_1002 ();
 FILLER_ASAP7_75t_R FILLER_0_241_1014 ();
 FILLER_ASAP7_75t_R FILLER_0_241_1022 ();
 FILLER_ASAP7_75t_R FILLER_0_241_1030 ();
 DECAPx2_ASAP7_75t_R FILLER_0_241_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_1043 ();
 DECAPx2_ASAP7_75t_R FILLER_0_241_1050 ();
 FILLER_ASAP7_75t_R FILLER_0_241_1062 ();
 DECAPx1_ASAP7_75t_R FILLER_0_241_1069 ();
 FILLER_ASAP7_75t_R FILLER_0_241_1079 ();
 DECAPx10_ASAP7_75t_R FILLER_0_241_1091 ();
 DECAPx1_ASAP7_75t_R FILLER_0_241_1113 ();
 FILLER_ASAP7_75t_R FILLER_0_241_1127 ();
 FILLER_ASAP7_75t_R FILLER_0_241_1134 ();
 DECAPx2_ASAP7_75t_R FILLER_0_241_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_1152 ();
 FILLER_ASAP7_75t_R FILLER_0_241_1161 ();
 FILLER_ASAP7_75t_R FILLER_0_241_1169 ();
 FILLER_ASAP7_75t_R FILLER_0_241_1176 ();
 FILLER_ASAP7_75t_R FILLER_0_241_1184 ();
 DECAPx4_ASAP7_75t_R FILLER_0_241_1191 ();
 DECAPx10_ASAP7_75t_R FILLER_0_241_1211 ();
 DECAPx1_ASAP7_75t_R FILLER_0_241_1233 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_1237 ();
 DECAPx2_ASAP7_75t_R FILLER_0_241_1248 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_1254 ();
 FILLER_ASAP7_75t_R FILLER_0_241_1260 ();
 FILLER_ASAP7_75t_R FILLER_0_241_1272 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_1274 ();
 FILLER_ASAP7_75t_R FILLER_0_241_1285 ();
 DECAPx2_ASAP7_75t_R FILLER_0_241_1293 ();
 FILLER_ASAP7_75t_R FILLER_0_241_1299 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_1301 ();
 FILLER_ASAP7_75t_R FILLER_0_241_1310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_241_1317 ();
 DECAPx2_ASAP7_75t_R FILLER_0_241_1339 ();
 FILLER_ASAP7_75t_R FILLER_0_241_1345 ();
 DECAPx2_ASAP7_75t_R FILLER_0_241_1353 ();
 FILLER_ASAP7_75t_R FILLER_0_241_1359 ();
 DECAPx2_ASAP7_75t_R FILLER_0_241_1367 ();
 FILLER_ASAP7_75t_R FILLER_0_241_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241_1381 ();
 DECAPx2_ASAP7_75t_R FILLER_0_242_2 ();
 FILLER_ASAP7_75t_R FILLER_0_242_8 ();
 DECAPx2_ASAP7_75t_R FILLER_0_242_18 ();
 FILLER_ASAP7_75t_R FILLER_0_242_24 ();
 DECAPx4_ASAP7_75t_R FILLER_0_242_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_42 ();
 DECAPx2_ASAP7_75t_R FILLER_0_242_49 ();
 FILLER_ASAP7_75t_R FILLER_0_242_55 ();
 DECAPx4_ASAP7_75t_R FILLER_0_242_63 ();
 FILLER_ASAP7_75t_R FILLER_0_242_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_81 ();
 FILLER_ASAP7_75t_R FILLER_0_242_88 ();
 FILLER_ASAP7_75t_R FILLER_0_242_100 ();
 FILLER_ASAP7_75t_R FILLER_0_242_108 ();
 DECAPx6_ASAP7_75t_R FILLER_0_242_115 ();
 DECAPx2_ASAP7_75t_R FILLER_0_242_129 ();
 DECAPx1_ASAP7_75t_R FILLER_0_242_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_145 ();
 DECAPx6_ASAP7_75t_R FILLER_0_242_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_166 ();
 FILLER_ASAP7_75t_R FILLER_0_242_173 ();
 FILLER_ASAP7_75t_R FILLER_0_242_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_183 ();
 DECAPx2_ASAP7_75t_R FILLER_0_242_190 ();
 DECAPx1_ASAP7_75t_R FILLER_0_242_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_206 ();
 DECAPx4_ASAP7_75t_R FILLER_0_242_228 ();
 FILLER_ASAP7_75t_R FILLER_0_242_243 ();
 DECAPx2_ASAP7_75t_R FILLER_0_242_261 ();
 DECAPx1_ASAP7_75t_R FILLER_0_242_277 ();
 DECAPx2_ASAP7_75t_R FILLER_0_242_290 ();
 FILLER_ASAP7_75t_R FILLER_0_242_306 ();
 DECAPx2_ASAP7_75t_R FILLER_0_242_314 ();
 FILLER_ASAP7_75t_R FILLER_0_242_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_322 ();
 DECAPx6_ASAP7_75t_R FILLER_0_242_329 ();
 DECAPx2_ASAP7_75t_R FILLER_0_242_343 ();
 FILLER_ASAP7_75t_R FILLER_0_242_355 ();
 DECAPx2_ASAP7_75t_R FILLER_0_242_363 ();
 FILLER_ASAP7_75t_R FILLER_0_242_369 ();
 DECAPx10_ASAP7_75t_R FILLER_0_242_377 ();
 DECAPx6_ASAP7_75t_R FILLER_0_242_399 ();
 FILLER_ASAP7_75t_R FILLER_0_242_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_415 ();
 DECAPx4_ASAP7_75t_R FILLER_0_242_422 ();
 FILLER_ASAP7_75t_R FILLER_0_242_432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_242_440 ();
 DECAPx1_ASAP7_75t_R FILLER_0_242_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_468 ();
 FILLER_ASAP7_75t_R FILLER_0_242_475 ();
 FILLER_ASAP7_75t_R FILLER_0_242_483 ();
 DECAPx10_ASAP7_75t_R FILLER_0_242_493 ();
 DECAPx1_ASAP7_75t_R FILLER_0_242_515 ();
 FILLER_ASAP7_75t_R FILLER_0_242_523 ();
 FILLER_ASAP7_75t_R FILLER_0_242_531 ();
 DECAPx2_ASAP7_75t_R FILLER_0_242_539 ();
 DECAPx10_ASAP7_75t_R FILLER_0_242_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_573 ();
 DECAPx4_ASAP7_75t_R FILLER_0_242_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_595 ();
 DECAPx4_ASAP7_75t_R FILLER_0_242_607 ();
 FILLER_ASAP7_75t_R FILLER_0_242_617 ();
 DECAPx10_ASAP7_75t_R FILLER_0_242_624 ();
 DECAPx10_ASAP7_75t_R FILLER_0_242_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_668 ();
 FILLER_ASAP7_75t_R FILLER_0_242_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_676 ();
 DECAPx4_ASAP7_75t_R FILLER_0_242_687 ();
 FILLER_ASAP7_75t_R FILLER_0_242_703 ();
 FILLER_ASAP7_75t_R FILLER_0_242_713 ();
 DECAPx4_ASAP7_75t_R FILLER_0_242_723 ();
 FILLER_ASAP7_75t_R FILLER_0_242_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_735 ();
 DECAPx4_ASAP7_75t_R FILLER_0_242_742 ();
 FILLER_ASAP7_75t_R FILLER_0_242_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_754 ();
 FILLER_ASAP7_75t_R FILLER_0_242_767 ();
 FILLER_ASAP7_75t_R FILLER_0_242_775 ();
 DECAPx2_ASAP7_75t_R FILLER_0_242_781 ();
 FILLER_ASAP7_75t_R FILLER_0_242_787 ();
 DECAPx10_ASAP7_75t_R FILLER_0_242_809 ();
 DECAPx4_ASAP7_75t_R FILLER_0_242_836 ();
 FILLER_ASAP7_75t_R FILLER_0_242_846 ();
 FILLER_ASAP7_75t_R FILLER_0_242_858 ();
 DECAPx1_ASAP7_75t_R FILLER_0_242_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_874 ();
 DECAPx2_ASAP7_75t_R FILLER_0_242_885 ();
 FILLER_ASAP7_75t_R FILLER_0_242_891 ();
 DECAPx2_ASAP7_75t_R FILLER_0_242_899 ();
 FILLER_ASAP7_75t_R FILLER_0_242_905 ();
 DECAPx4_ASAP7_75t_R FILLER_0_242_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_923 ();
 FILLER_ASAP7_75t_R FILLER_0_242_930 ();
 FILLER_ASAP7_75t_R FILLER_0_242_938 ();
 DECAPx2_ASAP7_75t_R FILLER_0_242_943 ();
 DECAPx1_ASAP7_75t_R FILLER_0_242_954 ();
 FILLER_ASAP7_75t_R FILLER_0_242_968 ();
 DECAPx1_ASAP7_75t_R FILLER_0_242_975 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_979 ();
 FILLER_ASAP7_75t_R FILLER_0_242_986 ();
 FILLER_ASAP7_75t_R FILLER_0_242_994 ();
 FILLER_ASAP7_75t_R FILLER_0_242_1002 ();
 DECAPx1_ASAP7_75t_R FILLER_0_242_1014 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_1018 ();
 FILLER_ASAP7_75t_R FILLER_0_242_1029 ();
 FILLER_ASAP7_75t_R FILLER_0_242_1037 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_1039 ();
 FILLER_ASAP7_75t_R FILLER_0_242_1051 ();
 DECAPx1_ASAP7_75t_R FILLER_0_242_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_1067 ();
 FILLER_ASAP7_75t_R FILLER_0_242_1076 ();
 DECAPx2_ASAP7_75t_R FILLER_0_242_1083 ();
 FILLER_ASAP7_75t_R FILLER_0_242_1089 ();
 DECAPx1_ASAP7_75t_R FILLER_0_242_1111 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_1115 ();
 DECAPx2_ASAP7_75t_R FILLER_0_242_1121 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_1127 ();
 FILLER_ASAP7_75t_R FILLER_0_242_1133 ();
 FILLER_ASAP7_75t_R FILLER_0_242_1145 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_1147 ();
 FILLER_ASAP7_75t_R FILLER_0_242_1154 ();
 FILLER_ASAP7_75t_R FILLER_0_242_1163 ();
 FILLER_ASAP7_75t_R FILLER_0_242_1171 ();
 FILLER_ASAP7_75t_R FILLER_0_242_1180 ();
 FILLER_ASAP7_75t_R FILLER_0_242_1188 ();
 FILLER_ASAP7_75t_R FILLER_0_242_1196 ();
 FILLER_ASAP7_75t_R FILLER_0_242_1204 ();
 FILLER_ASAP7_75t_R FILLER_0_242_1212 ();
 DECAPx1_ASAP7_75t_R FILLER_0_242_1220 ();
 DECAPx2_ASAP7_75t_R FILLER_0_242_1230 ();
 FILLER_ASAP7_75t_R FILLER_0_242_1236 ();
 FILLER_ASAP7_75t_R FILLER_0_242_1243 ();
 DECAPx2_ASAP7_75t_R FILLER_0_242_1251 ();
 FILLER_ASAP7_75t_R FILLER_0_242_1257 ();
 DECAPx4_ASAP7_75t_R FILLER_0_242_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_1279 ();
 FILLER_ASAP7_75t_R FILLER_0_242_1285 ();
 DECAPx1_ASAP7_75t_R FILLER_0_242_1297 ();
 DECAPx2_ASAP7_75t_R FILLER_0_242_1313 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_1319 ();
 FILLER_ASAP7_75t_R FILLER_0_242_1327 ();
 FILLER_ASAP7_75t_R FILLER_0_242_1335 ();
 FILLER_ASAP7_75t_R FILLER_0_242_1343 ();
 DECAPx2_ASAP7_75t_R FILLER_0_242_1351 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_242_1364 ();
 DECAPx1_ASAP7_75t_R FILLER_0_242_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242_1381 ();
 DECAPx2_ASAP7_75t_R FILLER_0_243_2 ();
 FILLER_ASAP7_75t_R FILLER_0_243_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_10 ();
 DECAPx4_ASAP7_75t_R FILLER_0_243_17 ();
 FILLER_ASAP7_75t_R FILLER_0_243_35 ();
 FILLER_ASAP7_75t_R FILLER_0_243_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_45 ();
 FILLER_ASAP7_75t_R FILLER_0_243_58 ();
 DECAPx2_ASAP7_75t_R FILLER_0_243_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_73 ();
 FILLER_ASAP7_75t_R FILLER_0_243_80 ();
 FILLER_ASAP7_75t_R FILLER_0_243_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_90 ();
 DECAPx1_ASAP7_75t_R FILLER_0_243_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_103 ();
 DECAPx2_ASAP7_75t_R FILLER_0_243_114 ();
 FILLER_ASAP7_75t_R FILLER_0_243_120 ();
 DECAPx1_ASAP7_75t_R FILLER_0_243_128 ();
 FILLER_ASAP7_75t_R FILLER_0_243_138 ();
 FILLER_ASAP7_75t_R FILLER_0_243_146 ();
 DECAPx4_ASAP7_75t_R FILLER_0_243_154 ();
 FILLER_ASAP7_75t_R FILLER_0_243_170 ();
 DECAPx2_ASAP7_75t_R FILLER_0_243_178 ();
 FILLER_ASAP7_75t_R FILLER_0_243_190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_243_198 ();
 DECAPx2_ASAP7_75t_R FILLER_0_243_220 ();
 FILLER_ASAP7_75t_R FILLER_0_243_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_231 ();
 FILLER_ASAP7_75t_R FILLER_0_243_237 ();
 FILLER_ASAP7_75t_R FILLER_0_243_245 ();
 FILLER_ASAP7_75t_R FILLER_0_243_253 ();
 FILLER_ASAP7_75t_R FILLER_0_243_265 ();
 FILLER_ASAP7_75t_R FILLER_0_243_270 ();
 FILLER_ASAP7_75t_R FILLER_0_243_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_284 ();
 DECAPx2_ASAP7_75t_R FILLER_0_243_291 ();
 FILLER_ASAP7_75t_R FILLER_0_243_303 ();
 DECAPx1_ASAP7_75t_R FILLER_0_243_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_317 ();
 DECAPx2_ASAP7_75t_R FILLER_0_243_324 ();
 FILLER_ASAP7_75t_R FILLER_0_243_330 ();
 DECAPx4_ASAP7_75t_R FILLER_0_243_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_350 ();
 DECAPx6_ASAP7_75t_R FILLER_0_243_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_371 ();
 DECAPx2_ASAP7_75t_R FILLER_0_243_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_384 ();
 DECAPx10_ASAP7_75t_R FILLER_0_243_391 ();
 FILLER_ASAP7_75t_R FILLER_0_243_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_415 ();
 DECAPx2_ASAP7_75t_R FILLER_0_243_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_428 ();
 FILLER_ASAP7_75t_R FILLER_0_243_435 ();
 DECAPx2_ASAP7_75t_R FILLER_0_243_444 ();
 FILLER_ASAP7_75t_R FILLER_0_243_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_452 ();
 FILLER_ASAP7_75t_R FILLER_0_243_459 ();
 DECAPx2_ASAP7_75t_R FILLER_0_243_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_473 ();
 DECAPx10_ASAP7_75t_R FILLER_0_243_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_506 ();
 DECAPx1_ASAP7_75t_R FILLER_0_243_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_517 ();
 FILLER_ASAP7_75t_R FILLER_0_243_524 ();
 FILLER_ASAP7_75t_R FILLER_0_243_532 ();
 FILLER_ASAP7_75t_R FILLER_0_243_542 ();
 FILLER_ASAP7_75t_R FILLER_0_243_552 ();
 FILLER_ASAP7_75t_R FILLER_0_243_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_559 ();
 DECAPx10_ASAP7_75t_R FILLER_0_243_571 ();
 DECAPx4_ASAP7_75t_R FILLER_0_243_593 ();
 FILLER_ASAP7_75t_R FILLER_0_243_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_605 ();
 FILLER_ASAP7_75t_R FILLER_0_243_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_619 ();
 FILLER_ASAP7_75t_R FILLER_0_243_632 ();
 FILLER_ASAP7_75t_R FILLER_0_243_645 ();
 DECAPx2_ASAP7_75t_R FILLER_0_243_658 ();
 FILLER_ASAP7_75t_R FILLER_0_243_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_666 ();
 FILLER_ASAP7_75t_R FILLER_0_243_675 ();
 FILLER_ASAP7_75t_R FILLER_0_243_687 ();
 FILLER_ASAP7_75t_R FILLER_0_243_701 ();
 DECAPx1_ASAP7_75t_R FILLER_0_243_713 ();
 DECAPx1_ASAP7_75t_R FILLER_0_243_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_731 ();
 DECAPx4_ASAP7_75t_R FILLER_0_243_744 ();
 FILLER_ASAP7_75t_R FILLER_0_243_754 ();
 DECAPx6_ASAP7_75t_R FILLER_0_243_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_776 ();
 DECAPx4_ASAP7_75t_R FILLER_0_243_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_793 ();
 DECAPx2_ASAP7_75t_R FILLER_0_243_802 ();
 FILLER_ASAP7_75t_R FILLER_0_243_816 ();
 DECAPx2_ASAP7_75t_R FILLER_0_243_838 ();
 FILLER_ASAP7_75t_R FILLER_0_243_844 ();
 DECAPx2_ASAP7_75t_R FILLER_0_243_852 ();
 DECAPx2_ASAP7_75t_R FILLER_0_243_868 ();
 DECAPx1_ASAP7_75t_R FILLER_0_243_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_884 ();
 DECAPx1_ASAP7_75t_R FILLER_0_243_905 ();
 FILLER_ASAP7_75t_R FILLER_0_243_915 ();
 FILLER_ASAP7_75t_R FILLER_0_243_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_924 ();
 DECAPx2_ASAP7_75t_R FILLER_0_243_927 ();
 FILLER_ASAP7_75t_R FILLER_0_243_933 ();
 DECAPx2_ASAP7_75t_R FILLER_0_243_941 ();
 DECAPx1_ASAP7_75t_R FILLER_0_243_953 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_957 ();
 FILLER_ASAP7_75t_R FILLER_0_243_968 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_970 ();
 FILLER_ASAP7_75t_R FILLER_0_243_981 ();
 FILLER_ASAP7_75t_R FILLER_0_243_993 ();
 FILLER_ASAP7_75t_R FILLER_0_243_1005 ();
 FILLER_ASAP7_75t_R FILLER_0_243_1017 ();
 FILLER_ASAP7_75t_R FILLER_0_243_1027 ();
 FILLER_ASAP7_75t_R FILLER_0_243_1035 ();
 FILLER_ASAP7_75t_R FILLER_0_243_1042 ();
 FILLER_ASAP7_75t_R FILLER_0_243_1064 ();
 FILLER_ASAP7_75t_R FILLER_0_243_1076 ();
 FILLER_ASAP7_75t_R FILLER_0_243_1081 ();
 FILLER_ASAP7_75t_R FILLER_0_243_1086 ();
 FILLER_ASAP7_75t_R FILLER_0_243_1095 ();
 DECAPx4_ASAP7_75t_R FILLER_0_243_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_1118 ();
 FILLER_ASAP7_75t_R FILLER_0_243_1123 ();
 DECAPx2_ASAP7_75t_R FILLER_0_243_1135 ();
 DECAPx1_ASAP7_75t_R FILLER_0_243_1151 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_1155 ();
 FILLER_ASAP7_75t_R FILLER_0_243_1161 ();
 FILLER_ASAP7_75t_R FILLER_0_243_1173 ();
 DECAPx1_ASAP7_75t_R FILLER_0_243_1181 ();
 FILLER_ASAP7_75t_R FILLER_0_243_1195 ();
 FILLER_ASAP7_75t_R FILLER_0_243_1203 ();
 DECAPx2_ASAP7_75t_R FILLER_0_243_1211 ();
 FILLER_ASAP7_75t_R FILLER_0_243_1224 ();
 DECAPx1_ASAP7_75t_R FILLER_0_243_1236 ();
 FILLER_ASAP7_75t_R FILLER_0_243_1250 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_1252 ();
 DECAPx2_ASAP7_75t_R FILLER_0_243_1258 ();
 FILLER_ASAP7_75t_R FILLER_0_243_1267 ();
 DECAPx2_ASAP7_75t_R FILLER_0_243_1272 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_1278 ();
 DECAPx2_ASAP7_75t_R FILLER_0_243_1299 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_1305 ();
 DECAPx4_ASAP7_75t_R FILLER_0_243_1312 ();
 FILLER_ASAP7_75t_R FILLER_0_243_1328 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243_1330 ();
 FILLER_ASAP7_75t_R FILLER_0_243_1338 ();
 FILLER_ASAP7_75t_R FILLER_0_243_1352 ();
 DECAPx10_ASAP7_75t_R FILLER_0_243_1360 ();
 DECAPx2_ASAP7_75t_R FILLER_0_244_2 ();
 FILLER_ASAP7_75t_R FILLER_0_244_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_10 ();
 DECAPx4_ASAP7_75t_R FILLER_0_244_17 ();
 DECAPx1_ASAP7_75t_R FILLER_0_244_33 ();
 FILLER_ASAP7_75t_R FILLER_0_244_43 ();
 FILLER_ASAP7_75t_R FILLER_0_244_51 ();
 FILLER_ASAP7_75t_R FILLER_0_244_59 ();
 FILLER_ASAP7_75t_R FILLER_0_244_67 ();
 FILLER_ASAP7_75t_R FILLER_0_244_75 ();
 DECAPx2_ASAP7_75t_R FILLER_0_244_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_90 ();
 DECAPx2_ASAP7_75t_R FILLER_0_244_101 ();
 FILLER_ASAP7_75t_R FILLER_0_244_113 ();
 FILLER_ASAP7_75t_R FILLER_0_244_121 ();
 DECAPx2_ASAP7_75t_R FILLER_0_244_129 ();
 DECAPx4_ASAP7_75t_R FILLER_0_244_141 ();
 DECAPx2_ASAP7_75t_R FILLER_0_244_157 ();
 FILLER_ASAP7_75t_R FILLER_0_244_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_165 ();
 DECAPx10_ASAP7_75t_R FILLER_0_244_172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_244_194 ();
 DECAPx6_ASAP7_75t_R FILLER_0_244_216 ();
 DECAPx2_ASAP7_75t_R FILLER_0_244_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_236 ();
 FILLER_ASAP7_75t_R FILLER_0_244_242 ();
 FILLER_ASAP7_75t_R FILLER_0_244_254 ();
 FILLER_ASAP7_75t_R FILLER_0_244_266 ();
 FILLER_ASAP7_75t_R FILLER_0_244_278 ();
 FILLER_ASAP7_75t_R FILLER_0_244_288 ();
 FILLER_ASAP7_75t_R FILLER_0_244_295 ();
 FILLER_ASAP7_75t_R FILLER_0_244_307 ();
 FILLER_ASAP7_75t_R FILLER_0_244_314 ();
 FILLER_ASAP7_75t_R FILLER_0_244_324 ();
 FILLER_ASAP7_75t_R FILLER_0_244_336 ();
 FILLER_ASAP7_75t_R FILLER_0_244_344 ();
 DECAPx1_ASAP7_75t_R FILLER_0_244_351 ();
 DECAPx2_ASAP7_75t_R FILLER_0_244_361 ();
 FILLER_ASAP7_75t_R FILLER_0_244_367 ();
 DECAPx2_ASAP7_75t_R FILLER_0_244_375 ();
 FILLER_ASAP7_75t_R FILLER_0_244_381 ();
 FILLER_ASAP7_75t_R FILLER_0_244_391 ();
 FILLER_ASAP7_75t_R FILLER_0_244_404 ();
 DECAPx1_ASAP7_75t_R FILLER_0_244_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_416 ();
 FILLER_ASAP7_75t_R FILLER_0_244_425 ();
 DECAPx10_ASAP7_75t_R FILLER_0_244_437 ();
 FILLER_ASAP7_75t_R FILLER_0_244_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_461 ();
 DECAPx1_ASAP7_75t_R FILLER_0_244_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_468 ();
 FILLER_ASAP7_75t_R FILLER_0_244_481 ();
 FILLER_ASAP7_75t_R FILLER_0_244_489 ();
 DECAPx2_ASAP7_75t_R FILLER_0_244_502 ();
 FILLER_ASAP7_75t_R FILLER_0_244_508 ();
 DECAPx2_ASAP7_75t_R FILLER_0_244_520 ();
 FILLER_ASAP7_75t_R FILLER_0_244_534 ();
 FILLER_ASAP7_75t_R FILLER_0_244_540 ();
 DECAPx1_ASAP7_75t_R FILLER_0_244_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_554 ();
 FILLER_ASAP7_75t_R FILLER_0_244_567 ();
 FILLER_ASAP7_75t_R FILLER_0_244_572 ();
 FILLER_ASAP7_75t_R FILLER_0_244_584 ();
 FILLER_ASAP7_75t_R FILLER_0_244_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_596 ();
 DECAPx4_ASAP7_75t_R FILLER_0_244_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_619 ();
 DECAPx2_ASAP7_75t_R FILLER_0_244_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_638 ();
 DECAPx1_ASAP7_75t_R FILLER_0_244_650 ();
 FILLER_ASAP7_75t_R FILLER_0_244_665 ();
 FILLER_ASAP7_75t_R FILLER_0_244_670 ();
 DECAPx4_ASAP7_75t_R FILLER_0_244_680 ();
 FILLER_ASAP7_75t_R FILLER_0_244_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_692 ();
 DECAPx2_ASAP7_75t_R FILLER_0_244_713 ();
 DECAPx2_ASAP7_75t_R FILLER_0_244_727 ();
 DECAPx2_ASAP7_75t_R FILLER_0_244_745 ();
 FILLER_ASAP7_75t_R FILLER_0_244_751 ();
 DECAPx4_ASAP7_75t_R FILLER_0_244_764 ();
 DECAPx4_ASAP7_75t_R FILLER_0_244_784 ();
 FILLER_ASAP7_75t_R FILLER_0_244_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_796 ();
 FILLER_ASAP7_75t_R FILLER_0_244_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_805 ();
 DECAPx1_ASAP7_75t_R FILLER_0_244_814 ();
 FILLER_ASAP7_75t_R FILLER_0_244_828 ();
 FILLER_ASAP7_75t_R FILLER_0_244_836 ();
 FILLER_ASAP7_75t_R FILLER_0_244_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_845 ();
 FILLER_ASAP7_75t_R FILLER_0_244_858 ();
 FILLER_ASAP7_75t_R FILLER_0_244_870 ();
 DECAPx2_ASAP7_75t_R FILLER_0_244_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_888 ();
 DECAPx4_ASAP7_75t_R FILLER_0_244_899 ();
 FILLER_ASAP7_75t_R FILLER_0_244_909 ();
 FILLER_ASAP7_75t_R FILLER_0_244_917 ();
 FILLER_ASAP7_75t_R FILLER_0_244_925 ();
 DECAPx2_ASAP7_75t_R FILLER_0_244_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_939 ();
 DECAPx6_ASAP7_75t_R FILLER_0_244_948 ();
 FILLER_ASAP7_75t_R FILLER_0_244_967 ();
 DECAPx6_ASAP7_75t_R FILLER_0_244_979 ();
 DECAPx2_ASAP7_75t_R FILLER_0_244_993 ();
 FILLER_ASAP7_75t_R FILLER_0_244_1002 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_1004 ();
 FILLER_ASAP7_75t_R FILLER_0_244_1015 ();
 FILLER_ASAP7_75t_R FILLER_0_244_1023 ();
 FILLER_ASAP7_75t_R FILLER_0_244_1035 ();
 DECAPx6_ASAP7_75t_R FILLER_0_244_1043 ();
 FILLER_ASAP7_75t_R FILLER_0_244_1063 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_1065 ();
 FILLER_ASAP7_75t_R FILLER_0_244_1076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_244_1084 ();
 DECAPx4_ASAP7_75t_R FILLER_0_244_1106 ();
 DECAPx2_ASAP7_75t_R FILLER_0_244_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_1132 ();
 DECAPx1_ASAP7_75t_R FILLER_0_244_1151 ();
 DECAPx1_ASAP7_75t_R FILLER_0_244_1161 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_1165 ();
 DECAPx1_ASAP7_75t_R FILLER_0_244_1174 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_1178 ();
 FILLER_ASAP7_75t_R FILLER_0_244_1189 ();
 FILLER_ASAP7_75t_R FILLER_0_244_1201 ();
 FILLER_ASAP7_75t_R FILLER_0_244_1209 ();
 FILLER_ASAP7_75t_R FILLER_0_244_1217 ();
 FILLER_ASAP7_75t_R FILLER_0_244_1225 ();
 DECAPx1_ASAP7_75t_R FILLER_0_244_1233 ();
 FILLER_ASAP7_75t_R FILLER_0_244_1242 ();
 DECAPx4_ASAP7_75t_R FILLER_0_244_1248 ();
 FILLER_ASAP7_75t_R FILLER_0_244_1268 ();
 DECAPx1_ASAP7_75t_R FILLER_0_244_1276 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_1280 ();
 FILLER_ASAP7_75t_R FILLER_0_244_1291 ();
 FILLER_ASAP7_75t_R FILLER_0_244_1300 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_1302 ();
 FILLER_ASAP7_75t_R FILLER_0_244_1309 ();
 DECAPx1_ASAP7_75t_R FILLER_0_244_1314 ();
 DECAPx6_ASAP7_75t_R FILLER_0_244_1330 ();
 FILLER_ASAP7_75t_R FILLER_0_244_1344 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_1346 ();
 DECAPx6_ASAP7_75t_R FILLER_0_244_1353 ();
 FILLER_ASAP7_75t_R FILLER_0_244_1367 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244_1369 ();
 FILLER_ASAP7_75t_R FILLER_0_244_1380 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_2 ();
 FILLER_ASAP7_75t_R FILLER_0_245_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_10 ();
 DECAPx6_ASAP7_75t_R FILLER_0_245_17 ();
 FILLER_ASAP7_75t_R FILLER_0_245_36 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_41 ();
 FILLER_ASAP7_75t_R FILLER_0_245_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_49 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_56 ();
 FILLER_ASAP7_75t_R FILLER_0_245_62 ();
 FILLER_ASAP7_75t_R FILLER_0_245_71 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_83 ();
 FILLER_ASAP7_75t_R FILLER_0_245_89 ();
 FILLER_ASAP7_75t_R FILLER_0_245_101 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_109 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_127 ();
 FILLER_ASAP7_75t_R FILLER_0_245_134 ();
 DECAPx6_ASAP7_75t_R FILLER_0_245_142 ();
 DECAPx1_ASAP7_75t_R FILLER_0_245_156 ();
 FILLER_ASAP7_75t_R FILLER_0_245_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_245_180 ();
 DECAPx6_ASAP7_75t_R FILLER_0_245_202 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_222 ();
 FILLER_ASAP7_75t_R FILLER_0_245_228 ();
 FILLER_ASAP7_75t_R FILLER_0_245_235 ();
 FILLER_ASAP7_75t_R FILLER_0_245_242 ();
 FILLER_ASAP7_75t_R FILLER_0_245_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_252 ();
 FILLER_ASAP7_75t_R FILLER_0_245_271 ();
 FILLER_ASAP7_75t_R FILLER_0_245_283 ();
 FILLER_ASAP7_75t_R FILLER_0_245_291 ();
 FILLER_ASAP7_75t_R FILLER_0_245_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_301 ();
 FILLER_ASAP7_75t_R FILLER_0_245_312 ();
 FILLER_ASAP7_75t_R FILLER_0_245_321 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_329 ();
 FILLER_ASAP7_75t_R FILLER_0_245_341 ();
 FILLER_ASAP7_75t_R FILLER_0_245_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_351 ();
 FILLER_ASAP7_75t_R FILLER_0_245_358 ();
 FILLER_ASAP7_75t_R FILLER_0_245_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_368 ();
 FILLER_ASAP7_75t_R FILLER_0_245_379 ();
 DECAPx6_ASAP7_75t_R FILLER_0_245_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_400 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_407 ();
 FILLER_ASAP7_75t_R FILLER_0_245_413 ();
 FILLER_ASAP7_75t_R FILLER_0_245_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_423 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_430 ();
 FILLER_ASAP7_75t_R FILLER_0_245_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_450 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_467 ();
 FILLER_ASAP7_75t_R FILLER_0_245_473 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_484 ();
 FILLER_ASAP7_75t_R FILLER_0_245_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_493 ();
 DECAPx10_ASAP7_75t_R FILLER_0_245_505 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_527 ();
 FILLER_ASAP7_75t_R FILLER_0_245_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_535 ();
 FILLER_ASAP7_75t_R FILLER_0_245_541 ();
 DECAPx6_ASAP7_75t_R FILLER_0_245_549 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_563 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_569 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_578 ();
 FILLER_ASAP7_75t_R FILLER_0_245_590 ();
 FILLER_ASAP7_75t_R FILLER_0_245_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_245_612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_245_634 ();
 DECAPx6_ASAP7_75t_R FILLER_0_245_656 ();
 FILLER_ASAP7_75t_R FILLER_0_245_670 ();
 FILLER_ASAP7_75t_R FILLER_0_245_680 ();
 DECAPx6_ASAP7_75t_R FILLER_0_245_690 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_704 ();
 FILLER_ASAP7_75t_R FILLER_0_245_715 ();
 FILLER_ASAP7_75t_R FILLER_0_245_723 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_728 ();
 DECAPx6_ASAP7_75t_R FILLER_0_245_742 ();
 DECAPx6_ASAP7_75t_R FILLER_0_245_762 ();
 FILLER_ASAP7_75t_R FILLER_0_245_776 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_784 ();
 FILLER_ASAP7_75t_R FILLER_0_245_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_792 ();
 FILLER_ASAP7_75t_R FILLER_0_245_801 ();
 FILLER_ASAP7_75t_R FILLER_0_245_809 ();
 FILLER_ASAP7_75t_R FILLER_0_245_815 ();
 FILLER_ASAP7_75t_R FILLER_0_245_821 ();
 FILLER_ASAP7_75t_R FILLER_0_245_833 ();
 FILLER_ASAP7_75t_R FILLER_0_245_845 ();
 DECAPx1_ASAP7_75t_R FILLER_0_245_857 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_877 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_894 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_903 ();
 FILLER_ASAP7_75t_R FILLER_0_245_915 ();
 FILLER_ASAP7_75t_R FILLER_0_245_923 ();
 DECAPx1_ASAP7_75t_R FILLER_0_245_927 ();
 DECAPx6_ASAP7_75t_R FILLER_0_245_938 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_952 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_958 ();
 DECAPx10_ASAP7_75t_R FILLER_0_245_964 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_986 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_992 ();
 FILLER_ASAP7_75t_R FILLER_0_245_999 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_1017 ();
 FILLER_ASAP7_75t_R FILLER_0_245_1028 ();
 FILLER_ASAP7_75t_R FILLER_0_245_1036 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_1043 ();
 FILLER_ASAP7_75t_R FILLER_0_245_1049 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_1051 ();
 DECAPx6_ASAP7_75t_R FILLER_0_245_1062 ();
 FILLER_ASAP7_75t_R FILLER_0_245_1082 ();
 FILLER_ASAP7_75t_R FILLER_0_245_1089 ();
 DECAPx6_ASAP7_75t_R FILLER_0_245_1094 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_1108 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_1114 ();
 FILLER_ASAP7_75t_R FILLER_0_245_1119 ();
 FILLER_ASAP7_75t_R FILLER_0_245_1126 ();
 FILLER_ASAP7_75t_R FILLER_0_245_1138 ();
 FILLER_ASAP7_75t_R FILLER_0_245_1150 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_1162 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_1168 ();
 FILLER_ASAP7_75t_R FILLER_0_245_1193 ();
 FILLER_ASAP7_75t_R FILLER_0_245_1207 ();
 FILLER_ASAP7_75t_R FILLER_0_245_1215 ();
 FILLER_ASAP7_75t_R FILLER_0_245_1223 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_1230 ();
 FILLER_ASAP7_75t_R FILLER_0_245_1236 ();
 FILLER_ASAP7_75t_R FILLER_0_245_1258 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_1270 ();
 FILLER_ASAP7_75t_R FILLER_0_245_1276 ();
 DECAPx1_ASAP7_75t_R FILLER_0_245_1283 ();
 DECAPx1_ASAP7_75t_R FILLER_0_245_1297 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245_1301 ();
 DECAPx10_ASAP7_75t_R FILLER_0_245_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_245_1336 ();
 DECAPx1_ASAP7_75t_R FILLER_0_245_1364 ();
 DECAPx2_ASAP7_75t_R FILLER_0_245_1374 ();
 FILLER_ASAP7_75t_R FILLER_0_245_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_246_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_24 ();
 FILLER_ASAP7_75t_R FILLER_0_246_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_246_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_50 ();
 DECAPx2_ASAP7_75t_R FILLER_0_246_57 ();
 DECAPx2_ASAP7_75t_R FILLER_0_246_83 ();
 FILLER_ASAP7_75t_R FILLER_0_246_94 ();
 FILLER_ASAP7_75t_R FILLER_0_246_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_103 ();
 FILLER_ASAP7_75t_R FILLER_0_246_114 ();
 FILLER_ASAP7_75t_R FILLER_0_246_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_123 ();
 DECAPx10_ASAP7_75t_R FILLER_0_246_130 ();
 DECAPx6_ASAP7_75t_R FILLER_0_246_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_166 ();
 DECAPx10_ASAP7_75t_R FILLER_0_246_172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_246_194 ();
 DECAPx2_ASAP7_75t_R FILLER_0_246_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_222 ();
 FILLER_ASAP7_75t_R FILLER_0_246_228 ();
 FILLER_ASAP7_75t_R FILLER_0_246_235 ();
 FILLER_ASAP7_75t_R FILLER_0_246_247 ();
 FILLER_ASAP7_75t_R FILLER_0_246_259 ();
 FILLER_ASAP7_75t_R FILLER_0_246_271 ();
 FILLER_ASAP7_75t_R FILLER_0_246_283 ();
 FILLER_ASAP7_75t_R FILLER_0_246_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_295 ();
 FILLER_ASAP7_75t_R FILLER_0_246_302 ();
 FILLER_ASAP7_75t_R FILLER_0_246_310 ();
 FILLER_ASAP7_75t_R FILLER_0_246_318 ();
 FILLER_ASAP7_75t_R FILLER_0_246_330 ();
 DECAPx6_ASAP7_75t_R FILLER_0_246_337 ();
 FILLER_ASAP7_75t_R FILLER_0_246_351 ();
 DECAPx4_ASAP7_75t_R FILLER_0_246_364 ();
 FILLER_ASAP7_75t_R FILLER_0_246_374 ();
 DECAPx6_ASAP7_75t_R FILLER_0_246_383 ();
 DECAPx1_ASAP7_75t_R FILLER_0_246_397 ();
 DECAPx6_ASAP7_75t_R FILLER_0_246_408 ();
 FILLER_ASAP7_75t_R FILLER_0_246_422 ();
 FILLER_ASAP7_75t_R FILLER_0_246_434 ();
 DECAPx6_ASAP7_75t_R FILLER_0_246_441 ();
 DECAPx2_ASAP7_75t_R FILLER_0_246_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_461 ();
 DECAPx1_ASAP7_75t_R FILLER_0_246_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_246_477 ();
 DECAPx10_ASAP7_75t_R FILLER_0_246_499 ();
 DECAPx10_ASAP7_75t_R FILLER_0_246_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_543 ();
 DECAPx6_ASAP7_75t_R FILLER_0_246_550 ();
 DECAPx2_ASAP7_75t_R FILLER_0_246_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_570 ();
 DECAPx2_ASAP7_75t_R FILLER_0_246_577 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_583 ();
 FILLER_ASAP7_75t_R FILLER_0_246_590 ();
 DECAPx4_ASAP7_75t_R FILLER_0_246_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_613 ();
 FILLER_ASAP7_75t_R FILLER_0_246_625 ();
 DECAPx1_ASAP7_75t_R FILLER_0_246_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_637 ();
 DECAPx6_ASAP7_75t_R FILLER_0_246_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_660 ();
 DECAPx2_ASAP7_75t_R FILLER_0_246_666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_246_680 ();
 FILLER_ASAP7_75t_R FILLER_0_246_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_704 ();
 FILLER_ASAP7_75t_R FILLER_0_246_708 ();
 FILLER_ASAP7_75t_R FILLER_0_246_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_718 ();
 DECAPx2_ASAP7_75t_R FILLER_0_246_724 ();
 FILLER_ASAP7_75t_R FILLER_0_246_730 ();
 FILLER_ASAP7_75t_R FILLER_0_246_738 ();
 FILLER_ASAP7_75t_R FILLER_0_246_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_246_759 ();
 DECAPx4_ASAP7_75t_R FILLER_0_246_781 ();
 FILLER_ASAP7_75t_R FILLER_0_246_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_793 ();
 DECAPx10_ASAP7_75t_R FILLER_0_246_798 ();
 FILLER_ASAP7_75t_R FILLER_0_246_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_822 ();
 DECAPx10_ASAP7_75t_R FILLER_0_246_831 ();
 FILLER_ASAP7_75t_R FILLER_0_246_853 ();
 FILLER_ASAP7_75t_R FILLER_0_246_865 ();
 FILLER_ASAP7_75t_R FILLER_0_246_875 ();
 DECAPx4_ASAP7_75t_R FILLER_0_246_883 ();
 FILLER_ASAP7_75t_R FILLER_0_246_903 ();
 FILLER_ASAP7_75t_R FILLER_0_246_915 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_917 ();
 DECAPx6_ASAP7_75t_R FILLER_0_246_923 ();
 DECAPx1_ASAP7_75t_R FILLER_0_246_937 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_941 ();
 DECAPx2_ASAP7_75t_R FILLER_0_246_949 ();
 FILLER_ASAP7_75t_R FILLER_0_246_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_957 ();
 FILLER_ASAP7_75t_R FILLER_0_246_963 ();
 DECAPx2_ASAP7_75t_R FILLER_0_246_985 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1001 ();
 DECAPx1_ASAP7_75t_R FILLER_0_246_1013 ();
 DECAPx1_ASAP7_75t_R FILLER_0_246_1023 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1034 ();
 DECAPx2_ASAP7_75t_R FILLER_0_246_1041 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1053 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1061 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1068 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_1070 ();
 DECAPx1_ASAP7_75t_R FILLER_0_246_1091 ();
 DECAPx2_ASAP7_75t_R FILLER_0_246_1105 ();
 DECAPx2_ASAP7_75t_R FILLER_0_246_1116 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1122 ();
 DECAPx1_ASAP7_75t_R FILLER_0_246_1134 ();
 DECAPx1_ASAP7_75t_R FILLER_0_246_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_1152 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1163 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1175 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1187 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1194 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1208 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1220 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1227 ();
 DECAPx2_ASAP7_75t_R FILLER_0_246_1234 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1246 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1254 ();
 DECAPx6_ASAP7_75t_R FILLER_0_246_1262 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1276 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_1278 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1299 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1307 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1315 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1321 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246_1323 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1330 ();
 DECAPx4_ASAP7_75t_R FILLER_0_246_1337 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1347 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1355 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1363 ();
 FILLER_ASAP7_75t_R FILLER_0_246_1371 ();
 DECAPx2_ASAP7_75t_R FILLER_0_246_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_247_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_247_24 ();
 FILLER_ASAP7_75t_R FILLER_0_247_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_38 ();
 FILLER_ASAP7_75t_R FILLER_0_247_45 ();
 DECAPx1_ASAP7_75t_R FILLER_0_247_50 ();
 DECAPx6_ASAP7_75t_R FILLER_0_247_60 ();
 FILLER_ASAP7_75t_R FILLER_0_247_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_76 ();
 DECAPx1_ASAP7_75t_R FILLER_0_247_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_87 ();
 FILLER_ASAP7_75t_R FILLER_0_247_93 ();
 DECAPx1_ASAP7_75t_R FILLER_0_247_105 ();
 DECAPx1_ASAP7_75t_R FILLER_0_247_115 ();
 DECAPx4_ASAP7_75t_R FILLER_0_247_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_132 ();
 FILLER_ASAP7_75t_R FILLER_0_247_139 ();
 FILLER_ASAP7_75t_R FILLER_0_247_144 ();
 DECAPx2_ASAP7_75t_R FILLER_0_247_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_158 ();
 DECAPx2_ASAP7_75t_R FILLER_0_247_165 ();
 DECAPx6_ASAP7_75t_R FILLER_0_247_174 ();
 DECAPx2_ASAP7_75t_R FILLER_0_247_188 ();
 DECAPx2_ASAP7_75t_R FILLER_0_247_216 ();
 FILLER_ASAP7_75t_R FILLER_0_247_227 ();
 FILLER_ASAP7_75t_R FILLER_0_247_235 ();
 FILLER_ASAP7_75t_R FILLER_0_247_247 ();
 FILLER_ASAP7_75t_R FILLER_0_247_259 ();
 FILLER_ASAP7_75t_R FILLER_0_247_279 ();
 FILLER_ASAP7_75t_R FILLER_0_247_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_293 ();
 FILLER_ASAP7_75t_R FILLER_0_247_297 ();
 FILLER_ASAP7_75t_R FILLER_0_247_309 ();
 FILLER_ASAP7_75t_R FILLER_0_247_317 ();
 FILLER_ASAP7_75t_R FILLER_0_247_327 ();
 FILLER_ASAP7_75t_R FILLER_0_247_335 ();
 DECAPx2_ASAP7_75t_R FILLER_0_247_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_347 ();
 DECAPx4_ASAP7_75t_R FILLER_0_247_354 ();
 DECAPx2_ASAP7_75t_R FILLER_0_247_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_378 ();
 DECAPx2_ASAP7_75t_R FILLER_0_247_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_397 ();
 FILLER_ASAP7_75t_R FILLER_0_247_418 ();
 FILLER_ASAP7_75t_R FILLER_0_247_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_430 ();
 DECAPx2_ASAP7_75t_R FILLER_0_247_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_443 ();
 DECAPx2_ASAP7_75t_R FILLER_0_247_450 ();
 DECAPx1_ASAP7_75t_R FILLER_0_247_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_466 ();
 FILLER_ASAP7_75t_R FILLER_0_247_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_489 ();
 FILLER_ASAP7_75t_R FILLER_0_247_493 ();
 DECAPx1_ASAP7_75t_R FILLER_0_247_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_511 ();
 DECAPx1_ASAP7_75t_R FILLER_0_247_518 ();
 DECAPx6_ASAP7_75t_R FILLER_0_247_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_557 ();
 DECAPx6_ASAP7_75t_R FILLER_0_247_579 ();
 DECAPx2_ASAP7_75t_R FILLER_0_247_593 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_599 ();
 DECAPx1_ASAP7_75t_R FILLER_0_247_610 ();
 FILLER_ASAP7_75t_R FILLER_0_247_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_627 ();
 FILLER_ASAP7_75t_R FILLER_0_247_638 ();
 DECAPx6_ASAP7_75t_R FILLER_0_247_648 ();
 DECAPx2_ASAP7_75t_R FILLER_0_247_662 ();
 DECAPx1_ASAP7_75t_R FILLER_0_247_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_680 ();
 DECAPx1_ASAP7_75t_R FILLER_0_247_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_693 ();
 DECAPx10_ASAP7_75t_R FILLER_0_247_702 ();
 DECAPx4_ASAP7_75t_R FILLER_0_247_724 ();
 FILLER_ASAP7_75t_R FILLER_0_247_734 ();
 DECAPx10_ASAP7_75t_R FILLER_0_247_742 ();
 DECAPx6_ASAP7_75t_R FILLER_0_247_764 ();
 DECAPx2_ASAP7_75t_R FILLER_0_247_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_792 ();
 FILLER_ASAP7_75t_R FILLER_0_247_801 ();
 DECAPx10_ASAP7_75t_R FILLER_0_247_811 ();
 FILLER_ASAP7_75t_R FILLER_0_247_833 ();
 DECAPx2_ASAP7_75t_R FILLER_0_247_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_851 ();
 DECAPx2_ASAP7_75t_R FILLER_0_247_858 ();
 FILLER_ASAP7_75t_R FILLER_0_247_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_866 ();
 DECAPx1_ASAP7_75t_R FILLER_0_247_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_879 ();
 FILLER_ASAP7_75t_R FILLER_0_247_886 ();
 DECAPx6_ASAP7_75t_R FILLER_0_247_894 ();
 FILLER_ASAP7_75t_R FILLER_0_247_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_910 ();
 FILLER_ASAP7_75t_R FILLER_0_247_923 ();
 DECAPx4_ASAP7_75t_R FILLER_0_247_927 ();
 FILLER_ASAP7_75t_R FILLER_0_247_937 ();
 FILLER_ASAP7_75t_R FILLER_0_247_951 ();
 FILLER_ASAP7_75t_R FILLER_0_247_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_961 ();
 DECAPx1_ASAP7_75t_R FILLER_0_247_970 ();
 FILLER_ASAP7_75t_R FILLER_0_247_980 ();
 FILLER_ASAP7_75t_R FILLER_0_247_988 ();
 DECAPx2_ASAP7_75t_R FILLER_0_247_998 ();
 DECAPx2_ASAP7_75t_R FILLER_0_247_1008 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1024 ();
 DECAPx4_ASAP7_75t_R FILLER_0_247_1034 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1044 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1049 ();
 DECAPx1_ASAP7_75t_R FILLER_0_247_1062 ();
 DECAPx1_ASAP7_75t_R FILLER_0_247_1078 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1088 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1096 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1104 ();
 DECAPx1_ASAP7_75t_R FILLER_0_247_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_1120 ();
 DECAPx2_ASAP7_75t_R FILLER_0_247_1131 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1147 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1159 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1171 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1183 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1195 ();
 DECAPx1_ASAP7_75t_R FILLER_0_247_1207 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1221 ();
 DECAPx1_ASAP7_75t_R FILLER_0_247_1233 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_1237 ();
 DECAPx2_ASAP7_75t_R FILLER_0_247_1244 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1250 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1260 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1272 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1281 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1293 ();
 DECAPx2_ASAP7_75t_R FILLER_0_247_1301 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1307 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_1309 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1318 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1326 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247_1328 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1335 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1343 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1351 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1359 ();
 DECAPx6_ASAP7_75t_R FILLER_0_247_1366 ();
 FILLER_ASAP7_75t_R FILLER_0_247_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_248_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_24 ();
 FILLER_ASAP7_75t_R FILLER_0_248_36 ();
 DECAPx6_ASAP7_75t_R FILLER_0_248_44 ();
 FILLER_ASAP7_75t_R FILLER_0_248_58 ();
 FILLER_ASAP7_75t_R FILLER_0_248_66 ();
 DECAPx6_ASAP7_75t_R FILLER_0_248_78 ();
 FILLER_ASAP7_75t_R FILLER_0_248_92 ();
 DECAPx6_ASAP7_75t_R FILLER_0_248_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_118 ();
 DECAPx1_ASAP7_75t_R FILLER_0_248_129 ();
 FILLER_ASAP7_75t_R FILLER_0_248_139 ();
 FILLER_ASAP7_75t_R FILLER_0_248_147 ();
 DECAPx1_ASAP7_75t_R FILLER_0_248_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_159 ();
 FILLER_ASAP7_75t_R FILLER_0_248_163 ();
 DECAPx10_ASAP7_75t_R FILLER_0_248_171 ();
 DECAPx6_ASAP7_75t_R FILLER_0_248_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_207 ();
 FILLER_ASAP7_75t_R FILLER_0_248_213 ();
 DECAPx2_ASAP7_75t_R FILLER_0_248_225 ();
 FILLER_ASAP7_75t_R FILLER_0_248_231 ();
 FILLER_ASAP7_75t_R FILLER_0_248_241 ();
 FILLER_ASAP7_75t_R FILLER_0_248_253 ();
 FILLER_ASAP7_75t_R FILLER_0_248_265 ();
 FILLER_ASAP7_75t_R FILLER_0_248_277 ();
 FILLER_ASAP7_75t_R FILLER_0_248_289 ();
 DECAPx1_ASAP7_75t_R FILLER_0_248_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_301 ();
 FILLER_ASAP7_75t_R FILLER_0_248_312 ();
 FILLER_ASAP7_75t_R FILLER_0_248_319 ();
 DECAPx1_ASAP7_75t_R FILLER_0_248_329 ();
 DECAPx2_ASAP7_75t_R FILLER_0_248_338 ();
 DECAPx1_ASAP7_75t_R FILLER_0_248_355 ();
 FILLER_ASAP7_75t_R FILLER_0_248_366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_248_374 ();
 FILLER_ASAP7_75t_R FILLER_0_248_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_398 ();
 FILLER_ASAP7_75t_R FILLER_0_248_419 ();
 FILLER_ASAP7_75t_R FILLER_0_248_428 ();
 DECAPx1_ASAP7_75t_R FILLER_0_248_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_440 ();
 FILLER_ASAP7_75t_R FILLER_0_248_447 ();
 DECAPx2_ASAP7_75t_R FILLER_0_248_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_461 ();
 DECAPx2_ASAP7_75t_R FILLER_0_248_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_470 ();
 FILLER_ASAP7_75t_R FILLER_0_248_477 ();
 FILLER_ASAP7_75t_R FILLER_0_248_485 ();
 DECAPx2_ASAP7_75t_R FILLER_0_248_497 ();
 FILLER_ASAP7_75t_R FILLER_0_248_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_517 ();
 DECAPx1_ASAP7_75t_R FILLER_0_248_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_528 ();
 DECAPx6_ASAP7_75t_R FILLER_0_248_539 ();
 DECAPx2_ASAP7_75t_R FILLER_0_248_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_559 ();
 FILLER_ASAP7_75t_R FILLER_0_248_563 ();
 DECAPx10_ASAP7_75t_R FILLER_0_248_570 ();
 DECAPx1_ASAP7_75t_R FILLER_0_248_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_596 ();
 DECAPx6_ASAP7_75t_R FILLER_0_248_607 ();
 DECAPx1_ASAP7_75t_R FILLER_0_248_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_625 ();
 DECAPx2_ASAP7_75t_R FILLER_0_248_632 ();
 DECAPx1_ASAP7_75t_R FILLER_0_248_646 ();
 DECAPx2_ASAP7_75t_R FILLER_0_248_658 ();
 DECAPx2_ASAP7_75t_R FILLER_0_248_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_680 ();
 FILLER_ASAP7_75t_R FILLER_0_248_691 ();
 FILLER_ASAP7_75t_R FILLER_0_248_701 ();
 DECAPx2_ASAP7_75t_R FILLER_0_248_707 ();
 FILLER_ASAP7_75t_R FILLER_0_248_713 ();
 DECAPx6_ASAP7_75t_R FILLER_0_248_721 ();
 FILLER_ASAP7_75t_R FILLER_0_248_735 ();
 DECAPx1_ASAP7_75t_R FILLER_0_248_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_752 ();
 FILLER_ASAP7_75t_R FILLER_0_248_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_763 ();
 FILLER_ASAP7_75t_R FILLER_0_248_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_774 ();
 FILLER_ASAP7_75t_R FILLER_0_248_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_780 ();
 FILLER_ASAP7_75t_R FILLER_0_248_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_791 ();
 FILLER_ASAP7_75t_R FILLER_0_248_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_802 ();
 FILLER_ASAP7_75t_R FILLER_0_248_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_811 ();
 FILLER_ASAP7_75t_R FILLER_0_248_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_817 ();
 FILLER_ASAP7_75t_R FILLER_0_248_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_828 ();
 DECAPx1_ASAP7_75t_R FILLER_0_248_849 ();
 FILLER_ASAP7_75t_R FILLER_0_248_864 ();
 DECAPx1_ASAP7_75t_R FILLER_0_248_872 ();
 FILLER_ASAP7_75t_R FILLER_0_248_883 ();
 FILLER_ASAP7_75t_R FILLER_0_248_891 ();
 DECAPx2_ASAP7_75t_R FILLER_0_248_901 ();
 FILLER_ASAP7_75t_R FILLER_0_248_907 ();
 FILLER_ASAP7_75t_R FILLER_0_248_921 ();
 FILLER_ASAP7_75t_R FILLER_0_248_931 ();
 DECAPx2_ASAP7_75t_R FILLER_0_248_940 ();
 FILLER_ASAP7_75t_R FILLER_0_248_946 ();
 FILLER_ASAP7_75t_R FILLER_0_248_954 ();
 FILLER_ASAP7_75t_R FILLER_0_248_966 ();
 FILLER_ASAP7_75t_R FILLER_0_248_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_978 ();
 FILLER_ASAP7_75t_R FILLER_0_248_989 ();
 FILLER_ASAP7_75t_R FILLER_0_248_1001 ();
 DECAPx1_ASAP7_75t_R FILLER_0_248_1013 ();
 FILLER_ASAP7_75t_R FILLER_0_248_1023 ();
 DECAPx1_ASAP7_75t_R FILLER_0_248_1037 ();
 FILLER_ASAP7_75t_R FILLER_0_248_1049 ();
 DECAPx1_ASAP7_75t_R FILLER_0_248_1057 ();
 DECAPx6_ASAP7_75t_R FILLER_0_248_1066 ();
 FILLER_ASAP7_75t_R FILLER_0_248_1086 ();
 FILLER_ASAP7_75t_R FILLER_0_248_1094 ();
 DECAPx6_ASAP7_75t_R FILLER_0_248_1102 ();
 DECAPx2_ASAP7_75t_R FILLER_0_248_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_1122 ();
 DECAPx2_ASAP7_75t_R FILLER_0_248_1133 ();
 DECAPx1_ASAP7_75t_R FILLER_0_248_1149 ();
 FILLER_ASAP7_75t_R FILLER_0_248_1163 ();
 FILLER_ASAP7_75t_R FILLER_0_248_1175 ();
 FILLER_ASAP7_75t_R FILLER_0_248_1187 ();
 FILLER_ASAP7_75t_R FILLER_0_248_1199 ();
 FILLER_ASAP7_75t_R FILLER_0_248_1207 ();
 FILLER_ASAP7_75t_R FILLER_0_248_1214 ();
 DECAPx1_ASAP7_75t_R FILLER_0_248_1226 ();
 FILLER_ASAP7_75t_R FILLER_0_248_1240 ();
 FILLER_ASAP7_75t_R FILLER_0_248_1250 ();
 FILLER_ASAP7_75t_R FILLER_0_248_1258 ();
 FILLER_ASAP7_75t_R FILLER_0_248_1270 ();
 DECAPx1_ASAP7_75t_R FILLER_0_248_1277 ();
 DECAPx1_ASAP7_75t_R FILLER_0_248_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_1292 ();
 FILLER_ASAP7_75t_R FILLER_0_248_1296 ();
 FILLER_ASAP7_75t_R FILLER_0_248_1308 ();
 FILLER_ASAP7_75t_R FILLER_0_248_1320 ();
 DECAPx10_ASAP7_75t_R FILLER_0_248_1330 ();
 DECAPx10_ASAP7_75t_R FILLER_0_248_1352 ();
 DECAPx2_ASAP7_75t_R FILLER_0_248_1374 ();
 FILLER_ASAP7_75t_R FILLER_0_248_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_249_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_249_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_249_46 ();
 DECAPx6_ASAP7_75t_R FILLER_0_249_68 ();
 DECAPx2_ASAP7_75t_R FILLER_0_249_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_88 ();
 FILLER_ASAP7_75t_R FILLER_0_249_99 ();
 DECAPx10_ASAP7_75t_R FILLER_0_249_107 ();
 DECAPx2_ASAP7_75t_R FILLER_0_249_129 ();
 DECAPx2_ASAP7_75t_R FILLER_0_249_138 ();
 FILLER_ASAP7_75t_R FILLER_0_249_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_249_157 ();
 DECAPx10_ASAP7_75t_R FILLER_0_249_179 ();
 DECAPx4_ASAP7_75t_R FILLER_0_249_201 ();
 FILLER_ASAP7_75t_R FILLER_0_249_211 ();
 DECAPx1_ASAP7_75t_R FILLER_0_249_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_220 ();
 FILLER_ASAP7_75t_R FILLER_0_249_226 ();
 FILLER_ASAP7_75t_R FILLER_0_249_236 ();
 FILLER_ASAP7_75t_R FILLER_0_249_248 ();
 FILLER_ASAP7_75t_R FILLER_0_249_260 ();
 FILLER_ASAP7_75t_R FILLER_0_249_272 ();
 FILLER_ASAP7_75t_R FILLER_0_249_284 ();
 FILLER_ASAP7_75t_R FILLER_0_249_296 ();
 FILLER_ASAP7_75t_R FILLER_0_249_306 ();
 DECAPx2_ASAP7_75t_R FILLER_0_249_315 ();
 FILLER_ASAP7_75t_R FILLER_0_249_327 ();
 FILLER_ASAP7_75t_R FILLER_0_249_335 ();
 DECAPx1_ASAP7_75t_R FILLER_0_249_353 ();
 DECAPx6_ASAP7_75t_R FILLER_0_249_363 ();
 DECAPx1_ASAP7_75t_R FILLER_0_249_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_381 ();
 FILLER_ASAP7_75t_R FILLER_0_249_389 ();
 DECAPx2_ASAP7_75t_R FILLER_0_249_397 ();
 FILLER_ASAP7_75t_R FILLER_0_249_403 ();
 FILLER_ASAP7_75t_R FILLER_0_249_411 ();
 DECAPx4_ASAP7_75t_R FILLER_0_249_425 ();
 FILLER_ASAP7_75t_R FILLER_0_249_435 ();
 DECAPx1_ASAP7_75t_R FILLER_0_249_443 ();
 DECAPx1_ASAP7_75t_R FILLER_0_249_454 ();
 FILLER_ASAP7_75t_R FILLER_0_249_463 ();
 FILLER_ASAP7_75t_R FILLER_0_249_471 ();
 DECAPx2_ASAP7_75t_R FILLER_0_249_479 ();
 DECAPx1_ASAP7_75t_R FILLER_0_249_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_500 ();
 DECAPx4_ASAP7_75t_R FILLER_0_249_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_523 ();
 DECAPx6_ASAP7_75t_R FILLER_0_249_527 ();
 FILLER_ASAP7_75t_R FILLER_0_249_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_543 ();
 FILLER_ASAP7_75t_R FILLER_0_249_552 ();
 FILLER_ASAP7_75t_R FILLER_0_249_564 ();
 DECAPx2_ASAP7_75t_R FILLER_0_249_576 ();
 FILLER_ASAP7_75t_R FILLER_0_249_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_584 ();
 FILLER_ASAP7_75t_R FILLER_0_249_593 ();
 DECAPx10_ASAP7_75t_R FILLER_0_249_601 ();
 FILLER_ASAP7_75t_R FILLER_0_249_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_625 ();
 FILLER_ASAP7_75t_R FILLER_0_249_636 ();
 FILLER_ASAP7_75t_R FILLER_0_249_646 ();
 DECAPx4_ASAP7_75t_R FILLER_0_249_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_666 ();
 DECAPx2_ASAP7_75t_R FILLER_0_249_675 ();
 FILLER_ASAP7_75t_R FILLER_0_249_689 ();
 FILLER_ASAP7_75t_R FILLER_0_249_699 ();
 FILLER_ASAP7_75t_R FILLER_0_249_709 ();
 FILLER_ASAP7_75t_R FILLER_0_249_721 ();
 FILLER_ASAP7_75t_R FILLER_0_249_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_731 ();
 FILLER_ASAP7_75t_R FILLER_0_249_743 ();
 DECAPx1_ASAP7_75t_R FILLER_0_249_750 ();
 FILLER_ASAP7_75t_R FILLER_0_249_760 ();
 FILLER_ASAP7_75t_R FILLER_0_249_768 ();
 DECAPx1_ASAP7_75t_R FILLER_0_249_776 ();
 DECAPx1_ASAP7_75t_R FILLER_0_249_790 ();
 DECAPx1_ASAP7_75t_R FILLER_0_249_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_804 ();
 FILLER_ASAP7_75t_R FILLER_0_249_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_813 ();
 DECAPx1_ASAP7_75t_R FILLER_0_249_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_826 ();
 FILLER_ASAP7_75t_R FILLER_0_249_835 ();
 FILLER_ASAP7_75t_R FILLER_0_249_840 ();
 DECAPx6_ASAP7_75t_R FILLER_0_249_845 ();
 DECAPx2_ASAP7_75t_R FILLER_0_249_865 ();
 FILLER_ASAP7_75t_R FILLER_0_249_871 ();
 FILLER_ASAP7_75t_R FILLER_0_249_883 ();
 FILLER_ASAP7_75t_R FILLER_0_249_895 ();
 DECAPx2_ASAP7_75t_R FILLER_0_249_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_909 ();
 DECAPx1_ASAP7_75t_R FILLER_0_249_921 ();
 FILLER_ASAP7_75t_R FILLER_0_249_927 ();
 FILLER_ASAP7_75t_R FILLER_0_249_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_936 ();
 FILLER_ASAP7_75t_R FILLER_0_249_952 ();
 FILLER_ASAP7_75t_R FILLER_0_249_964 ();
 FILLER_ASAP7_75t_R FILLER_0_249_972 ();
 FILLER_ASAP7_75t_R FILLER_0_249_994 ();
 FILLER_ASAP7_75t_R FILLER_0_249_1002 ();
 DECAPx1_ASAP7_75t_R FILLER_0_249_1009 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_1013 ();
 FILLER_ASAP7_75t_R FILLER_0_249_1020 ();
 DECAPx1_ASAP7_75t_R FILLER_0_249_1028 ();
 DECAPx1_ASAP7_75t_R FILLER_0_249_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_1042 ();
 DECAPx10_ASAP7_75t_R FILLER_0_249_1049 ();
 FILLER_ASAP7_75t_R FILLER_0_249_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_1073 ();
 DECAPx10_ASAP7_75t_R FILLER_0_249_1080 ();
 DECAPx2_ASAP7_75t_R FILLER_0_249_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_1108 ();
 DECAPx4_ASAP7_75t_R FILLER_0_249_1121 ();
 FILLER_ASAP7_75t_R FILLER_0_249_1137 ();
 DECAPx2_ASAP7_75t_R FILLER_0_249_1149 ();
 FILLER_ASAP7_75t_R FILLER_0_249_1165 ();
 FILLER_ASAP7_75t_R FILLER_0_249_1177 ();
 FILLER_ASAP7_75t_R FILLER_0_249_1189 ();
 FILLER_ASAP7_75t_R FILLER_0_249_1203 ();
 FILLER_ASAP7_75t_R FILLER_0_249_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_1210 ();
 DECAPx1_ASAP7_75t_R FILLER_0_249_1219 ();
 DECAPx2_ASAP7_75t_R FILLER_0_249_1229 ();
 DECAPx2_ASAP7_75t_R FILLER_0_249_1243 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_1249 ();
 FILLER_ASAP7_75t_R FILLER_0_249_1260 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_1262 ();
 FILLER_ASAP7_75t_R FILLER_0_249_1273 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_1275 ();
 DECAPx6_ASAP7_75t_R FILLER_0_249_1286 ();
 DECAPx2_ASAP7_75t_R FILLER_0_249_1300 ();
 DECAPx1_ASAP7_75t_R FILLER_0_249_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_0_249_1325 ();
 DECAPx2_ASAP7_75t_R FILLER_0_249_1347 ();
 FILLER_ASAP7_75t_R FILLER_0_249_1353 ();
 DECAPx2_ASAP7_75t_R FILLER_0_249_1363 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_1369 ();
 FILLER_ASAP7_75t_R FILLER_0_249_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_250_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_250_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_250_46 ();
 DECAPx6_ASAP7_75t_R FILLER_0_250_68 ();
 DECAPx2_ASAP7_75t_R FILLER_0_250_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_88 ();
 DECAPx10_ASAP7_75t_R FILLER_0_250_99 ();
 DECAPx10_ASAP7_75t_R FILLER_0_250_121 ();
 DECAPx10_ASAP7_75t_R FILLER_0_250_143 ();
 DECAPx10_ASAP7_75t_R FILLER_0_250_165 ();
 DECAPx10_ASAP7_75t_R FILLER_0_250_187 ();
 DECAPx4_ASAP7_75t_R FILLER_0_250_209 ();
 FILLER_ASAP7_75t_R FILLER_0_250_219 ();
 FILLER_ASAP7_75t_R FILLER_0_250_226 ();
 FILLER_ASAP7_75t_R FILLER_0_250_234 ();
 FILLER_ASAP7_75t_R FILLER_0_250_246 ();
 FILLER_ASAP7_75t_R FILLER_0_250_258 ();
 FILLER_ASAP7_75t_R FILLER_0_250_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_272 ();
 FILLER_ASAP7_75t_R FILLER_0_250_295 ();
 FILLER_ASAP7_75t_R FILLER_0_250_302 ();
 FILLER_ASAP7_75t_R FILLER_0_250_314 ();
 FILLER_ASAP7_75t_R FILLER_0_250_326 ();
 DECAPx2_ASAP7_75t_R FILLER_0_250_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_344 ();
 DECAPx1_ASAP7_75t_R FILLER_0_250_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_359 ();
 FILLER_ASAP7_75t_R FILLER_0_250_366 ();
 DECAPx1_ASAP7_75t_R FILLER_0_250_376 ();
 FILLER_ASAP7_75t_R FILLER_0_250_386 ();
 DECAPx2_ASAP7_75t_R FILLER_0_250_398 ();
 FILLER_ASAP7_75t_R FILLER_0_250_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_406 ();
 DECAPx1_ASAP7_75t_R FILLER_0_250_417 ();
 DECAPx10_ASAP7_75t_R FILLER_0_250_427 ();
 DECAPx4_ASAP7_75t_R FILLER_0_250_449 ();
 FILLER_ASAP7_75t_R FILLER_0_250_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_461 ();
 FILLER_ASAP7_75t_R FILLER_0_250_464 ();
 FILLER_ASAP7_75t_R FILLER_0_250_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_474 ();
 DECAPx4_ASAP7_75t_R FILLER_0_250_481 ();
 DECAPx6_ASAP7_75t_R FILLER_0_250_497 ();
 FILLER_ASAP7_75t_R FILLER_0_250_511 ();
 DECAPx6_ASAP7_75t_R FILLER_0_250_516 ();
 DECAPx2_ASAP7_75t_R FILLER_0_250_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_536 ();
 FILLER_ASAP7_75t_R FILLER_0_250_543 ();
 FILLER_ASAP7_75t_R FILLER_0_250_551 ();
 FILLER_ASAP7_75t_R FILLER_0_250_561 ();
 DECAPx1_ASAP7_75t_R FILLER_0_250_571 ();
 FILLER_ASAP7_75t_R FILLER_0_250_583 ();
 FILLER_ASAP7_75t_R FILLER_0_250_593 ();
 DECAPx2_ASAP7_75t_R FILLER_0_250_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_607 ();
 DECAPx1_ASAP7_75t_R FILLER_0_250_616 ();
 DECAPx10_ASAP7_75t_R FILLER_0_250_630 ();
 DECAPx6_ASAP7_75t_R FILLER_0_250_652 ();
 DECAPx2_ASAP7_75t_R FILLER_0_250_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_680 ();
 DECAPx1_ASAP7_75t_R FILLER_0_250_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_691 ();
 FILLER_ASAP7_75t_R FILLER_0_250_700 ();
 DECAPx2_ASAP7_75t_R FILLER_0_250_710 ();
 FILLER_ASAP7_75t_R FILLER_0_250_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_718 ();
 DECAPx2_ASAP7_75t_R FILLER_0_250_729 ();
 DECAPx2_ASAP7_75t_R FILLER_0_250_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_752 ();
 FILLER_ASAP7_75t_R FILLER_0_250_759 ();
 FILLER_ASAP7_75t_R FILLER_0_250_766 ();
 FILLER_ASAP7_75t_R FILLER_0_250_775 ();
 DECAPx4_ASAP7_75t_R FILLER_0_250_787 ();
 FILLER_ASAP7_75t_R FILLER_0_250_797 ();
 FILLER_ASAP7_75t_R FILLER_0_250_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_250_813 ();
 FILLER_ASAP7_75t_R FILLER_0_250_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_829 ();
 DECAPx6_ASAP7_75t_R FILLER_0_250_840 ();
 DECAPx1_ASAP7_75t_R FILLER_0_250_854 ();
 FILLER_ASAP7_75t_R FILLER_0_250_864 ();
 DECAPx2_ASAP7_75t_R FILLER_0_250_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_882 ();
 FILLER_ASAP7_75t_R FILLER_0_250_897 ();
 FILLER_ASAP7_75t_R FILLER_0_250_909 ();
 FILLER_ASAP7_75t_R FILLER_0_250_917 ();
 FILLER_ASAP7_75t_R FILLER_0_250_924 ();
 FILLER_ASAP7_75t_R FILLER_0_250_931 ();
 FILLER_ASAP7_75t_R FILLER_0_250_936 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_938 ();
 DECAPx6_ASAP7_75t_R FILLER_0_250_945 ();
 FILLER_ASAP7_75t_R FILLER_0_250_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_961 ();
 FILLER_ASAP7_75t_R FILLER_0_250_967 ();
 DECAPx4_ASAP7_75t_R FILLER_0_250_975 ();
 FILLER_ASAP7_75t_R FILLER_0_250_985 ();
 DECAPx1_ASAP7_75t_R FILLER_0_250_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_997 ();
 FILLER_ASAP7_75t_R FILLER_0_250_1004 ();
 FILLER_ASAP7_75t_R FILLER_0_250_1012 ();
 DECAPx2_ASAP7_75t_R FILLER_0_250_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_1024 ();
 FILLER_ASAP7_75t_R FILLER_0_250_1031 ();
 FILLER_ASAP7_75t_R FILLER_0_250_1043 ();
 FILLER_ASAP7_75t_R FILLER_0_250_1050 ();
 DECAPx4_ASAP7_75t_R FILLER_0_250_1057 ();
 FILLER_ASAP7_75t_R FILLER_0_250_1073 ();
 FILLER_ASAP7_75t_R FILLER_0_250_1081 ();
 DECAPx1_ASAP7_75t_R FILLER_0_250_1089 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_1093 ();
 DECAPx6_ASAP7_75t_R FILLER_0_250_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_1114 ();
 DECAPx2_ASAP7_75t_R FILLER_0_250_1125 ();
 FILLER_ASAP7_75t_R FILLER_0_250_1131 ();
 DECAPx2_ASAP7_75t_R FILLER_0_250_1137 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_1143 ();
 DECAPx1_ASAP7_75t_R FILLER_0_250_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_1158 ();
 DECAPx1_ASAP7_75t_R FILLER_0_250_1165 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_1169 ();
 FILLER_ASAP7_75t_R FILLER_0_250_1180 ();
 FILLER_ASAP7_75t_R FILLER_0_250_1192 ();
 FILLER_ASAP7_75t_R FILLER_0_250_1200 ();
 FILLER_ASAP7_75t_R FILLER_0_250_1208 ();
 FILLER_ASAP7_75t_R FILLER_0_250_1216 ();
 FILLER_ASAP7_75t_R FILLER_0_250_1224 ();
 FILLER_ASAP7_75t_R FILLER_0_250_1232 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_1234 ();
 FILLER_ASAP7_75t_R FILLER_0_250_1243 ();
 DECAPx2_ASAP7_75t_R FILLER_0_250_1251 ();
 FILLER_ASAP7_75t_R FILLER_0_250_1265 ();
 DECAPx6_ASAP7_75t_R FILLER_0_250_1285 ();
 FILLER_ASAP7_75t_R FILLER_0_250_1299 ();
 DECAPx1_ASAP7_75t_R FILLER_0_250_1311 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_1315 ();
 DECAPx2_ASAP7_75t_R FILLER_0_250_1328 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_1334 ();
 FILLER_ASAP7_75t_R FILLER_0_250_1339 ();
 FILLER_ASAP7_75t_R FILLER_0_250_1349 ();
 FILLER_ASAP7_75t_R FILLER_0_250_1357 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_1359 ();
 FILLER_ASAP7_75t_R FILLER_0_250_1368 ();
 DECAPx2_ASAP7_75t_R FILLER_0_250_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_251_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_251_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_251_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_251_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_251_90 ();
 DECAPx4_ASAP7_75t_R FILLER_0_251_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_251_143 ();
 DECAPx10_ASAP7_75t_R FILLER_0_251_165 ();
 DECAPx10_ASAP7_75t_R FILLER_0_251_187 ();
 DECAPx4_ASAP7_75t_R FILLER_0_251_209 ();
 FILLER_ASAP7_75t_R FILLER_0_251_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_221 ();
 FILLER_ASAP7_75t_R FILLER_0_251_227 ();
 FILLER_ASAP7_75t_R FILLER_0_251_234 ();
 FILLER_ASAP7_75t_R FILLER_0_251_241 ();
 FILLER_ASAP7_75t_R FILLER_0_251_253 ();
 FILLER_ASAP7_75t_R FILLER_0_251_265 ();
 DECAPx2_ASAP7_75t_R FILLER_0_251_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_283 ();
 FILLER_ASAP7_75t_R FILLER_0_251_294 ();
 FILLER_ASAP7_75t_R FILLER_0_251_306 ();
 DECAPx2_ASAP7_75t_R FILLER_0_251_314 ();
 FILLER_ASAP7_75t_R FILLER_0_251_325 ();
 DECAPx1_ASAP7_75t_R FILLER_0_251_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_338 ();
 DECAPx2_ASAP7_75t_R FILLER_0_251_349 ();
 FILLER_ASAP7_75t_R FILLER_0_251_355 ();
 FILLER_ASAP7_75t_R FILLER_0_251_363 ();
 FILLER_ASAP7_75t_R FILLER_0_251_372 ();
 DECAPx4_ASAP7_75t_R FILLER_0_251_379 ();
 DECAPx1_ASAP7_75t_R FILLER_0_251_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_401 ();
 DECAPx2_ASAP7_75t_R FILLER_0_251_412 ();
 FILLER_ASAP7_75t_R FILLER_0_251_424 ();
 DECAPx6_ASAP7_75t_R FILLER_0_251_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_446 ();
 DECAPx2_ASAP7_75t_R FILLER_0_251_453 ();
 FILLER_ASAP7_75t_R FILLER_0_251_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_251_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_490 ();
 DECAPx6_ASAP7_75t_R FILLER_0_251_497 ();
 DECAPx4_ASAP7_75t_R FILLER_0_251_532 ();
 FILLER_ASAP7_75t_R FILLER_0_251_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_544 ();
 DECAPx2_ASAP7_75t_R FILLER_0_251_549 ();
 FILLER_ASAP7_75t_R FILLER_0_251_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_563 ();
 DECAPx6_ASAP7_75t_R FILLER_0_251_567 ();
 FILLER_ASAP7_75t_R FILLER_0_251_589 ();
 DECAPx2_ASAP7_75t_R FILLER_0_251_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_603 ();
 DECAPx2_ASAP7_75t_R FILLER_0_251_614 ();
 FILLER_ASAP7_75t_R FILLER_0_251_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_622 ();
 DECAPx6_ASAP7_75t_R FILLER_0_251_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_643 ();
 DECAPx2_ASAP7_75t_R FILLER_0_251_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_658 ();
 FILLER_ASAP7_75t_R FILLER_0_251_665 ();
 DECAPx2_ASAP7_75t_R FILLER_0_251_673 ();
 FILLER_ASAP7_75t_R FILLER_0_251_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_681 ();
 DECAPx1_ASAP7_75t_R FILLER_0_251_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_698 ();
 DECAPx6_ASAP7_75t_R FILLER_0_251_704 ();
 DECAPx1_ASAP7_75t_R FILLER_0_251_718 ();
 DECAPx1_ASAP7_75t_R FILLER_0_251_728 ();
 DECAPx1_ASAP7_75t_R FILLER_0_251_742 ();
 DECAPx6_ASAP7_75t_R FILLER_0_251_757 ();
 DECAPx2_ASAP7_75t_R FILLER_0_251_781 ();
 FILLER_ASAP7_75t_R FILLER_0_251_794 ();
 FILLER_ASAP7_75t_R FILLER_0_251_806 ();
 FILLER_ASAP7_75t_R FILLER_0_251_814 ();
 DECAPx4_ASAP7_75t_R FILLER_0_251_822 ();
 DECAPx4_ASAP7_75t_R FILLER_0_251_842 ();
 FILLER_ASAP7_75t_R FILLER_0_251_852 ();
 FILLER_ASAP7_75t_R FILLER_0_251_864 ();
 FILLER_ASAP7_75t_R FILLER_0_251_871 ();
 FILLER_ASAP7_75t_R FILLER_0_251_891 ();
 FILLER_ASAP7_75t_R FILLER_0_251_903 ();
 FILLER_ASAP7_75t_R FILLER_0_251_911 ();
 DECAPx2_ASAP7_75t_R FILLER_0_251_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_924 ();
 DECAPx1_ASAP7_75t_R FILLER_0_251_927 ();
 DECAPx2_ASAP7_75t_R FILLER_0_251_938 ();
 FILLER_ASAP7_75t_R FILLER_0_251_944 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_946 ();
 DECAPx2_ASAP7_75t_R FILLER_0_251_957 ();
 DECAPx10_ASAP7_75t_R FILLER_0_251_968 ();
 DECAPx2_ASAP7_75t_R FILLER_0_251_990 ();
 FILLER_ASAP7_75t_R FILLER_0_251_996 ();
 FILLER_ASAP7_75t_R FILLER_0_251_1008 ();
 FILLER_ASAP7_75t_R FILLER_0_251_1020 ();
 FILLER_ASAP7_75t_R FILLER_0_251_1030 ();
 DECAPx4_ASAP7_75t_R FILLER_0_251_1038 ();
 FILLER_ASAP7_75t_R FILLER_0_251_1054 ();
 DECAPx4_ASAP7_75t_R FILLER_0_251_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_1072 ();
 FILLER_ASAP7_75t_R FILLER_0_251_1083 ();
 DECAPx1_ASAP7_75t_R FILLER_0_251_1091 ();
 DECAPx6_ASAP7_75t_R FILLER_0_251_1105 ();
 FILLER_ASAP7_75t_R FILLER_0_251_1119 ();
 DECAPx6_ASAP7_75t_R FILLER_0_251_1131 ();
 DECAPx2_ASAP7_75t_R FILLER_0_251_1145 ();
 FILLER_ASAP7_75t_R FILLER_0_251_1161 ();
 FILLER_ASAP7_75t_R FILLER_0_251_1168 ();
 FILLER_ASAP7_75t_R FILLER_0_251_1178 ();
 FILLER_ASAP7_75t_R FILLER_0_251_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_251_1194 ();
 FILLER_ASAP7_75t_R FILLER_0_251_1202 ();
 FILLER_ASAP7_75t_R FILLER_0_251_1210 ();
 FILLER_ASAP7_75t_R FILLER_0_251_1218 ();
 DECAPx2_ASAP7_75t_R FILLER_0_251_1226 ();
 FILLER_ASAP7_75t_R FILLER_0_251_1239 ();
 DECAPx2_ASAP7_75t_R FILLER_0_251_1247 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_1253 ();
 DECAPx1_ASAP7_75t_R FILLER_0_251_1264 ();
 FILLER_ASAP7_75t_R FILLER_0_251_1278 ();
 DECAPx2_ASAP7_75t_R FILLER_0_251_1292 ();
 FILLER_ASAP7_75t_R FILLER_0_251_1298 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_1300 ();
 FILLER_ASAP7_75t_R FILLER_0_251_1311 ();
 DECAPx1_ASAP7_75t_R FILLER_0_251_1318 ();
 FILLER_ASAP7_75t_R FILLER_0_251_1334 ();
 DECAPx2_ASAP7_75t_R FILLER_0_251_1341 ();
 FILLER_ASAP7_75t_R FILLER_0_251_1357 ();
 DECAPx2_ASAP7_75t_R FILLER_0_251_1365 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_1371 ();
 DECAPx1_ASAP7_75t_R FILLER_0_251_1378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_252_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_252_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_252_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_252_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_252_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_252_112 ();
 DECAPx2_ASAP7_75t_R FILLER_0_252_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_252_140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_252_144 ();
 DECAPx10_ASAP7_75t_R FILLER_0_252_166 ();
 DECAPx10_ASAP7_75t_R FILLER_0_252_188 ();
 DECAPx6_ASAP7_75t_R FILLER_0_252_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_252_224 ();
 FILLER_ASAP7_75t_R FILLER_0_252_230 ();
 FILLER_ASAP7_75t_R FILLER_0_252_237 ();
 FILLER_ASAP7_75t_R FILLER_0_252_251 ();
 DECAPx1_ASAP7_75t_R FILLER_0_252_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_252_267 ();
 FILLER_ASAP7_75t_R FILLER_0_252_278 ();
 FILLER_ASAP7_75t_R FILLER_0_252_290 ();
 FILLER_ASAP7_75t_R FILLER_0_252_302 ();
 FILLER_ASAP7_75t_R FILLER_0_252_310 ();
 DECAPx2_ASAP7_75t_R FILLER_0_252_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_252_323 ();
 FILLER_ASAP7_75t_R FILLER_0_252_329 ();
 DECAPx2_ASAP7_75t_R FILLER_0_252_335 ();
 FILLER_ASAP7_75t_R FILLER_0_252_347 ();
 DECAPx1_ASAP7_75t_R FILLER_0_252_356 ();
 FILLER_ASAP7_75t_R FILLER_0_252_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_252_367 ();
 FILLER_ASAP7_75t_R FILLER_0_252_378 ();
 FILLER_ASAP7_75t_R FILLER_0_252_390 ();
 DECAPx2_ASAP7_75t_R FILLER_0_252_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_252_403 ();
 DECAPx6_ASAP7_75t_R FILLER_0_252_409 ();
 FILLER_ASAP7_75t_R FILLER_0_252_423 ();
 FILLER_ASAP7_75t_R FILLER_0_252_431 ();
 FILLER_ASAP7_75t_R FILLER_0_252_439 ();
 FILLER_ASAP7_75t_R FILLER_0_252_447 ();
 FILLER_ASAP7_75t_R FILLER_0_252_460 ();
 DECAPx1_ASAP7_75t_R FILLER_0_252_464 ();
 DECAPx2_ASAP7_75t_R FILLER_0_252_476 ();
 FILLER_ASAP7_75t_R FILLER_0_252_482 ();
 FILLER_ASAP7_75t_R FILLER_0_252_490 ();
 FILLER_ASAP7_75t_R FILLER_0_252_498 ();
 DECAPx1_ASAP7_75t_R FILLER_0_252_506 ();
 DECAPx2_ASAP7_75t_R FILLER_0_252_516 ();
 FILLER_ASAP7_75t_R FILLER_0_252_533 ();
 FILLER_ASAP7_75t_R FILLER_0_252_556 ();
 FILLER_ASAP7_75t_R FILLER_0_252_564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_252_574 ();
 DECAPx2_ASAP7_75t_R FILLER_0_252_596 ();
 FILLER_ASAP7_75t_R FILLER_0_252_612 ();
 FILLER_ASAP7_75t_R FILLER_0_252_622 ();
 FILLER_ASAP7_75t_R FILLER_0_252_634 ();
 FILLER_ASAP7_75t_R FILLER_0_252_644 ();
 FILLER_ASAP7_75t_R FILLER_0_252_652 ();
 DECAPx2_ASAP7_75t_R FILLER_0_252_660 ();
 FILLER_ASAP7_75t_R FILLER_0_252_666 ();
 DECAPx4_ASAP7_75t_R FILLER_0_252_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_252_681 ();
 DECAPx10_ASAP7_75t_R FILLER_0_252_688 ();
 DECAPx4_ASAP7_75t_R FILLER_0_252_710 ();
 FILLER_ASAP7_75t_R FILLER_0_252_720 ();
 FILLER_ASAP7_75t_R FILLER_0_252_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_252_732 ();
 DECAPx2_ASAP7_75t_R FILLER_0_252_755 ();
 DECAPx1_ASAP7_75t_R FILLER_0_252_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_252_785 ();
 DECAPx2_ASAP7_75t_R FILLER_0_252_806 ();
 FILLER_ASAP7_75t_R FILLER_0_252_820 ();
 FILLER_ASAP7_75t_R FILLER_0_252_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_252_830 ();
 DECAPx2_ASAP7_75t_R FILLER_0_252_852 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_252_858 ();
 FILLER_ASAP7_75t_R FILLER_0_252_873 ();
 FILLER_ASAP7_75t_R FILLER_0_252_886 ();
 FILLER_ASAP7_75t_R FILLER_0_252_898 ();
 DECAPx2_ASAP7_75t_R FILLER_0_252_906 ();
 FILLER_ASAP7_75t_R FILLER_0_252_912 ();
 DECAPx2_ASAP7_75t_R FILLER_0_252_924 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_252_930 ();
 FILLER_ASAP7_75t_R FILLER_0_252_945 ();
 DECAPx4_ASAP7_75t_R FILLER_0_252_953 ();
 DECAPx1_ASAP7_75t_R FILLER_0_252_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_252_973 ();
 FILLER_ASAP7_75t_R FILLER_0_252_984 ();
 FILLER_ASAP7_75t_R FILLER_0_252_996 ();
 FILLER_ASAP7_75t_R FILLER_0_252_1008 ();
 FILLER_ASAP7_75t_R FILLER_0_252_1020 ();
 FILLER_ASAP7_75t_R FILLER_0_252_1032 ();
 DECAPx1_ASAP7_75t_R FILLER_0_252_1039 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_252_1043 ();
 FILLER_ASAP7_75t_R FILLER_0_252_1050 ();
 FILLER_ASAP7_75t_R FILLER_0_252_1060 ();
 DECAPx2_ASAP7_75t_R FILLER_0_252_1068 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_252_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_0_252_1081 ();
 FILLER_ASAP7_75t_R FILLER_0_252_1087 ();
 FILLER_ASAP7_75t_R FILLER_0_252_1099 ();
 DECAPx6_ASAP7_75t_R FILLER_0_252_1104 ();
 DECAPx2_ASAP7_75t_R FILLER_0_252_1118 ();
 DECAPx6_ASAP7_75t_R FILLER_0_252_1134 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_252_1148 ();
 FILLER_ASAP7_75t_R FILLER_0_252_1152 ();
 FILLER_ASAP7_75t_R FILLER_0_252_1160 ();
 DECAPx1_ASAP7_75t_R FILLER_0_252_1172 ();
 DECAPx2_ASAP7_75t_R FILLER_0_252_1184 ();
 FILLER_ASAP7_75t_R FILLER_0_252_1190 ();
 FILLER_ASAP7_75t_R FILLER_0_252_1206 ();
 DECAPx1_ASAP7_75t_R FILLER_0_252_1214 ();
 FILLER_ASAP7_75t_R FILLER_0_252_1228 ();
 FILLER_ASAP7_75t_R FILLER_0_252_1237 ();
 DECAPx2_ASAP7_75t_R FILLER_0_252_1249 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_252_1255 ();
 FILLER_ASAP7_75t_R FILLER_0_252_1268 ();
 DECAPx4_ASAP7_75t_R FILLER_0_252_1275 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_252_1285 ();
 DECAPx2_ASAP7_75t_R FILLER_0_252_1292 ();
 FILLER_ASAP7_75t_R FILLER_0_252_1298 ();
 FILLER_ASAP7_75t_R FILLER_0_252_1303 ();
 FILLER_ASAP7_75t_R FILLER_0_252_1315 ();
 FILLER_ASAP7_75t_R FILLER_0_252_1322 ();
 FILLER_ASAP7_75t_R FILLER_0_252_1336 ();
 DECAPx1_ASAP7_75t_R FILLER_0_252_1343 ();
 DECAPx4_ASAP7_75t_R FILLER_0_252_1353 ();
 DECAPx2_ASAP7_75t_R FILLER_0_252_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_252_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_252_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_253_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_253_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_253_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_253_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_253_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_253_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_253_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_253_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_253_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_253_200 ();
 DECAPx1_ASAP7_75t_R FILLER_0_253_222 ();
 FILLER_ASAP7_75t_R FILLER_0_253_231 ();
 FILLER_ASAP7_75t_R FILLER_0_253_239 ();
 FILLER_ASAP7_75t_R FILLER_0_253_251 ();
 DECAPx2_ASAP7_75t_R FILLER_0_253_263 ();
 FILLER_ASAP7_75t_R FILLER_0_253_269 ();
 DECAPx1_ASAP7_75t_R FILLER_0_253_281 ();
 FILLER_ASAP7_75t_R FILLER_0_253_291 ();
 FILLER_ASAP7_75t_R FILLER_0_253_303 ();
 DECAPx2_ASAP7_75t_R FILLER_0_253_313 ();
 FILLER_ASAP7_75t_R FILLER_0_253_329 ();
 FILLER_ASAP7_75t_R FILLER_0_253_341 ();
 FILLER_ASAP7_75t_R FILLER_0_253_353 ();
 FILLER_ASAP7_75t_R FILLER_0_253_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_253_367 ();
 FILLER_ASAP7_75t_R FILLER_0_253_378 ();
 FILLER_ASAP7_75t_R FILLER_0_253_390 ();
 FILLER_ASAP7_75t_R FILLER_0_253_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_253_404 ();
 DECAPx6_ASAP7_75t_R FILLER_0_253_411 ();
 DECAPx1_ASAP7_75t_R FILLER_0_253_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_253_429 ();
 FILLER_ASAP7_75t_R FILLER_0_253_440 ();
 DECAPx1_ASAP7_75t_R FILLER_0_253_448 ();
 FILLER_ASAP7_75t_R FILLER_0_253_458 ();
 FILLER_ASAP7_75t_R FILLER_0_253_466 ();
 DECAPx4_ASAP7_75t_R FILLER_0_253_474 ();
 DECAPx2_ASAP7_75t_R FILLER_0_253_490 ();
 FILLER_ASAP7_75t_R FILLER_0_253_496 ();
 FILLER_ASAP7_75t_R FILLER_0_253_520 ();
 FILLER_ASAP7_75t_R FILLER_0_253_534 ();
 FILLER_ASAP7_75t_R FILLER_0_253_542 ();
 FILLER_ASAP7_75t_R FILLER_0_253_550 ();
 DECAPx1_ASAP7_75t_R FILLER_0_253_557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_253_573 ();
 DECAPx2_ASAP7_75t_R FILLER_0_253_591 ();
 FILLER_ASAP7_75t_R FILLER_0_253_597 ();
 FILLER_ASAP7_75t_R FILLER_0_253_602 ();
 FILLER_ASAP7_75t_R FILLER_0_253_612 ();
 FILLER_ASAP7_75t_R FILLER_0_253_624 ();
 DECAPx2_ASAP7_75t_R FILLER_0_253_636 ();
 FILLER_ASAP7_75t_R FILLER_0_253_642 ();
 FILLER_ASAP7_75t_R FILLER_0_253_650 ();
 FILLER_ASAP7_75t_R FILLER_0_253_664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_253_678 ();
 DECAPx2_ASAP7_75t_R FILLER_0_253_700 ();
 FILLER_ASAP7_75t_R FILLER_0_253_706 ();
 FILLER_ASAP7_75t_R FILLER_0_253_714 ();
 FILLER_ASAP7_75t_R FILLER_0_253_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_253_721 ();
 FILLER_ASAP7_75t_R FILLER_0_253_730 ();
 DECAPx2_ASAP7_75t_R FILLER_0_253_740 ();
 FILLER_ASAP7_75t_R FILLER_0_253_757 ();
 FILLER_ASAP7_75t_R FILLER_0_253_769 ();
 FILLER_ASAP7_75t_R FILLER_0_253_779 ();
 FILLER_ASAP7_75t_R FILLER_0_253_789 ();
 FILLER_ASAP7_75t_R FILLER_0_253_801 ();
 DECAPx6_ASAP7_75t_R FILLER_0_253_809 ();
 FILLER_ASAP7_75t_R FILLER_0_253_823 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_253_825 ();
 FILLER_ASAP7_75t_R FILLER_0_253_832 ();
 FILLER_ASAP7_75t_R FILLER_0_253_839 ();
 DECAPx6_ASAP7_75t_R FILLER_0_253_844 ();
 FILLER_ASAP7_75t_R FILLER_0_253_863 ();
 FILLER_ASAP7_75t_R FILLER_0_253_881 ();
 FILLER_ASAP7_75t_R FILLER_0_253_891 ();
 FILLER_ASAP7_75t_R FILLER_0_253_899 ();
 DECAPx2_ASAP7_75t_R FILLER_0_253_907 ();
 FILLER_ASAP7_75t_R FILLER_0_253_923 ();
 FILLER_ASAP7_75t_R FILLER_0_253_927 ();
 FILLER_ASAP7_75t_R FILLER_0_253_937 ();
 DECAPx2_ASAP7_75t_R FILLER_0_253_945 ();
 FILLER_ASAP7_75t_R FILLER_0_253_951 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_253_953 ();
 DECAPx2_ASAP7_75t_R FILLER_0_253_964 ();
 DECAPx1_ASAP7_75t_R FILLER_0_253_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_253_980 ();
 FILLER_ASAP7_75t_R FILLER_0_253_988 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_253_990 ();
 FILLER_ASAP7_75t_R FILLER_0_253_1005 ();
 FILLER_ASAP7_75t_R FILLER_0_253_1017 ();
 FILLER_ASAP7_75t_R FILLER_0_253_1029 ();
 FILLER_ASAP7_75t_R FILLER_0_253_1041 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_253_1043 ();
 FILLER_ASAP7_75t_R FILLER_0_253_1064 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_253_1066 ();
 FILLER_ASAP7_75t_R FILLER_0_253_1070 ();
 FILLER_ASAP7_75t_R FILLER_0_253_1092 ();
 DECAPx1_ASAP7_75t_R FILLER_0_253_1099 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_253_1103 ();
 DECAPx6_ASAP7_75t_R FILLER_0_253_1110 ();
 FILLER_ASAP7_75t_R FILLER_0_253_1124 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_253_1126 ();
 FILLER_ASAP7_75t_R FILLER_0_253_1137 ();
 FILLER_ASAP7_75t_R FILLER_0_253_1151 ();
 DECAPx1_ASAP7_75t_R FILLER_0_253_1167 ();
 FILLER_ASAP7_75t_R FILLER_0_253_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_253_1183 ();
 FILLER_ASAP7_75t_R FILLER_0_253_1194 ();
 FILLER_ASAP7_75t_R FILLER_0_253_1202 ();
 FILLER_ASAP7_75t_R FILLER_0_253_1209 ();
 FILLER_ASAP7_75t_R FILLER_0_253_1219 ();
 FILLER_ASAP7_75t_R FILLER_0_253_1226 ();
 DECAPx4_ASAP7_75t_R FILLER_0_253_1232 ();
 DECAPx2_ASAP7_75t_R FILLER_0_253_1248 ();
 FILLER_ASAP7_75t_R FILLER_0_253_1254 ();
 FILLER_ASAP7_75t_R FILLER_0_253_1268 ();
 FILLER_ASAP7_75t_R FILLER_0_253_1276 ();
 FILLER_ASAP7_75t_R FILLER_0_253_1285 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_253_1287 ();
 DECAPx1_ASAP7_75t_R FILLER_0_253_1299 ();
 FILLER_ASAP7_75t_R FILLER_0_253_1308 ();
 FILLER_ASAP7_75t_R FILLER_0_253_1322 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_253_1324 ();
 DECAPx1_ASAP7_75t_R FILLER_0_253_1333 ();
 FILLER_ASAP7_75t_R FILLER_0_253_1348 ();
 FILLER_ASAP7_75t_R FILLER_0_253_1353 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_253_1355 ();
 DECAPx2_ASAP7_75t_R FILLER_0_253_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_254_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_254_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_254_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_254_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_254_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_254_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_254_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_254_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_254_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_254_200 ();
 FILLER_ASAP7_75t_R FILLER_0_254_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_224 ();
 FILLER_ASAP7_75t_R FILLER_0_254_230 ();
 FILLER_ASAP7_75t_R FILLER_0_254_238 ();
 DECAPx2_ASAP7_75t_R FILLER_0_254_250 ();
 FILLER_ASAP7_75t_R FILLER_0_254_266 ();
 FILLER_ASAP7_75t_R FILLER_0_254_275 ();
 FILLER_ASAP7_75t_R FILLER_0_254_283 ();
 FILLER_ASAP7_75t_R FILLER_0_254_291 ();
 FILLER_ASAP7_75t_R FILLER_0_254_298 ();
 FILLER_ASAP7_75t_R FILLER_0_254_305 ();
 FILLER_ASAP7_75t_R FILLER_0_254_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_315 ();
 DECAPx2_ASAP7_75t_R FILLER_0_254_322 ();
 FILLER_ASAP7_75t_R FILLER_0_254_338 ();
 DECAPx1_ASAP7_75t_R FILLER_0_254_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_354 ();
 FILLER_ASAP7_75t_R FILLER_0_254_360 ();
 FILLER_ASAP7_75t_R FILLER_0_254_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_370 ();
 FILLER_ASAP7_75t_R FILLER_0_254_381 ();
 DECAPx2_ASAP7_75t_R FILLER_0_254_393 ();
 FILLER_ASAP7_75t_R FILLER_0_254_405 ();
 FILLER_ASAP7_75t_R FILLER_0_254_413 ();
 DECAPx2_ASAP7_75t_R FILLER_0_254_421 ();
 FILLER_ASAP7_75t_R FILLER_0_254_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_429 ();
 FILLER_ASAP7_75t_R FILLER_0_254_433 ();
 FILLER_ASAP7_75t_R FILLER_0_254_441 ();
 FILLER_ASAP7_75t_R FILLER_0_254_449 ();
 DECAPx2_ASAP7_75t_R FILLER_0_254_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_461 ();
 DECAPx2_ASAP7_75t_R FILLER_0_254_464 ();
 FILLER_ASAP7_75t_R FILLER_0_254_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_472 ();
 DECAPx2_ASAP7_75t_R FILLER_0_254_480 ();
 FILLER_ASAP7_75t_R FILLER_0_254_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_254_505 ();
 DECAPx2_ASAP7_75t_R FILLER_0_254_527 ();
 FILLER_ASAP7_75t_R FILLER_0_254_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_535 ();
 FILLER_ASAP7_75t_R FILLER_0_254_539 ();
 DECAPx6_ASAP7_75t_R FILLER_0_254_546 ();
 DECAPx1_ASAP7_75t_R FILLER_0_254_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_564 ();
 DECAPx6_ASAP7_75t_R FILLER_0_254_586 ();
 DECAPx1_ASAP7_75t_R FILLER_0_254_600 ();
 FILLER_ASAP7_75t_R FILLER_0_254_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_614 ();
 DECAPx1_ASAP7_75t_R FILLER_0_254_625 ();
 DECAPx6_ASAP7_75t_R FILLER_0_254_641 ();
 DECAPx1_ASAP7_75t_R FILLER_0_254_655 ();
 DECAPx10_ASAP7_75t_R FILLER_0_254_680 ();
 FILLER_ASAP7_75t_R FILLER_0_254_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_704 ();
 FILLER_ASAP7_75t_R FILLER_0_254_717 ();
 DECAPx2_ASAP7_75t_R FILLER_0_254_725 ();
 FILLER_ASAP7_75t_R FILLER_0_254_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_733 ();
 DECAPx4_ASAP7_75t_R FILLER_0_254_737 ();
 FILLER_ASAP7_75t_R FILLER_0_254_747 ();
 DECAPx6_ASAP7_75t_R FILLER_0_254_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_254_777 ();
 DECAPx1_ASAP7_75t_R FILLER_0_254_799 ();
 DECAPx6_ASAP7_75t_R FILLER_0_254_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_825 ();
 DECAPx6_ASAP7_75t_R FILLER_0_254_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_852 ();
 FILLER_ASAP7_75t_R FILLER_0_254_858 ();
 FILLER_ASAP7_75t_R FILLER_0_254_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_872 ();
 FILLER_ASAP7_75t_R FILLER_0_254_891 ();
 FILLER_ASAP7_75t_R FILLER_0_254_899 ();
 FILLER_ASAP7_75t_R FILLER_0_254_907 ();
 FILLER_ASAP7_75t_R FILLER_0_254_917 ();
 DECAPx2_ASAP7_75t_R FILLER_0_254_929 ();
 FILLER_ASAP7_75t_R FILLER_0_254_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_937 ();
 FILLER_ASAP7_75t_R FILLER_0_254_948 ();
 FILLER_ASAP7_75t_R FILLER_0_254_956 ();
 DECAPx1_ASAP7_75t_R FILLER_0_254_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_968 ();
 FILLER_ASAP7_75t_R FILLER_0_254_972 ();
 FILLER_ASAP7_75t_R FILLER_0_254_980 ();
 FILLER_ASAP7_75t_R FILLER_0_254_992 ();
 FILLER_ASAP7_75t_R FILLER_0_254_1004 ();
 FILLER_ASAP7_75t_R FILLER_0_254_1016 ();
 FILLER_ASAP7_75t_R FILLER_0_254_1024 ();
 FILLER_ASAP7_75t_R FILLER_0_254_1032 ();
 DECAPx6_ASAP7_75t_R FILLER_0_254_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_1054 ();
 FILLER_ASAP7_75t_R FILLER_0_254_1060 ();
 FILLER_ASAP7_75t_R FILLER_0_254_1072 ();
 FILLER_ASAP7_75t_R FILLER_0_254_1080 ();
 FILLER_ASAP7_75t_R FILLER_0_254_1088 ();
 FILLER_ASAP7_75t_R FILLER_0_254_1100 ();
 DECAPx6_ASAP7_75t_R FILLER_0_254_1105 ();
 DECAPx2_ASAP7_75t_R FILLER_0_254_1119 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_1125 ();
 DECAPx4_ASAP7_75t_R FILLER_0_254_1132 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_1142 ();
 FILLER_ASAP7_75t_R FILLER_0_254_1148 ();
 FILLER_ASAP7_75t_R FILLER_0_254_1156 ();
 DECAPx2_ASAP7_75t_R FILLER_0_254_1164 ();
 FILLER_ASAP7_75t_R FILLER_0_254_1178 ();
 FILLER_ASAP7_75t_R FILLER_0_254_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_254_1194 ();
 FILLER_ASAP7_75t_R FILLER_0_254_1202 ();
 FILLER_ASAP7_75t_R FILLER_0_254_1210 ();
 FILLER_ASAP7_75t_R FILLER_0_254_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_1217 ();
 DECAPx1_ASAP7_75t_R FILLER_0_254_1228 ();
 DECAPx6_ASAP7_75t_R FILLER_0_254_1238 ();
 FILLER_ASAP7_75t_R FILLER_0_254_1252 ();
 FILLER_ASAP7_75t_R FILLER_0_254_1260 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_1262 ();
 DECAPx6_ASAP7_75t_R FILLER_0_254_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_1283 ();
 FILLER_ASAP7_75t_R FILLER_0_254_1292 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_1294 ();
 DECAPx1_ASAP7_75t_R FILLER_0_254_1301 ();
 DECAPx6_ASAP7_75t_R FILLER_0_254_1315 ();
 FILLER_ASAP7_75t_R FILLER_0_254_1329 ();
 FILLER_ASAP7_75t_R FILLER_0_254_1339 ();
 DECAPx1_ASAP7_75t_R FILLER_0_254_1347 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_1351 ();
 FILLER_ASAP7_75t_R FILLER_0_254_1358 ();
 FILLER_ASAP7_75t_R FILLER_0_254_1367 ();
 DECAPx2_ASAP7_75t_R FILLER_0_254_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_255_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_255_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_255_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_255_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_255_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_255_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_255_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_255_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_255_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_255_200 ();
 DECAPx4_ASAP7_75t_R FILLER_0_255_222 ();
 FILLER_ASAP7_75t_R FILLER_0_255_237 ();
 FILLER_ASAP7_75t_R FILLER_0_255_245 ();
 FILLER_ASAP7_75t_R FILLER_0_255_257 ();
 DECAPx2_ASAP7_75t_R FILLER_0_255_275 ();
 DECAPx2_ASAP7_75t_R FILLER_0_255_287 ();
 DECAPx2_ASAP7_75t_R FILLER_0_255_301 ();
 FILLER_ASAP7_75t_R FILLER_0_255_307 ();
 DECAPx1_ASAP7_75t_R FILLER_0_255_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_255_319 ();
 DECAPx2_ASAP7_75t_R FILLER_0_255_326 ();
 FILLER_ASAP7_75t_R FILLER_0_255_340 ();
 FILLER_ASAP7_75t_R FILLER_0_255_350 ();
 FILLER_ASAP7_75t_R FILLER_0_255_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_255_362 ();
 FILLER_ASAP7_75t_R FILLER_0_255_369 ();
 FILLER_ASAP7_75t_R FILLER_0_255_381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_255_393 ();
 DECAPx4_ASAP7_75t_R FILLER_0_255_415 ();
 DECAPx1_ASAP7_75t_R FILLER_0_255_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_255_439 ();
 DECAPx10_ASAP7_75t_R FILLER_0_255_445 ();
 DECAPx1_ASAP7_75t_R FILLER_0_255_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_255_471 ();
 DECAPx6_ASAP7_75t_R FILLER_0_255_478 ();
 FILLER_ASAP7_75t_R FILLER_0_255_492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_255_498 ();
 DECAPx4_ASAP7_75t_R FILLER_0_255_520 ();
 DECAPx4_ASAP7_75t_R FILLER_0_255_552 ();
 FILLER_ASAP7_75t_R FILLER_0_255_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_255_564 ();
 FILLER_ASAP7_75t_R FILLER_0_255_571 ();
 DECAPx2_ASAP7_75t_R FILLER_0_255_576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_255_603 ();
 DECAPx10_ASAP7_75t_R FILLER_0_255_625 ();
 DECAPx4_ASAP7_75t_R FILLER_0_255_647 ();
 FILLER_ASAP7_75t_R FILLER_0_255_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_255_659 ();
 FILLER_ASAP7_75t_R FILLER_0_255_666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_255_671 ();
 DECAPx10_ASAP7_75t_R FILLER_0_255_693 ();
 DECAPx4_ASAP7_75t_R FILLER_0_255_715 ();
 FILLER_ASAP7_75t_R FILLER_0_255_731 ();
 DECAPx2_ASAP7_75t_R FILLER_0_255_741 ();
 FILLER_ASAP7_75t_R FILLER_0_255_753 ();
 FILLER_ASAP7_75t_R FILLER_0_255_761 ();
 DECAPx10_ASAP7_75t_R FILLER_0_255_774 ();
 DECAPx6_ASAP7_75t_R FILLER_0_255_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_255_810 ();
 DECAPx4_ASAP7_75t_R FILLER_0_255_817 ();
 DECAPx2_ASAP7_75t_R FILLER_0_255_839 ();
 FILLER_ASAP7_75t_R FILLER_0_255_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_255_847 ();
 FILLER_ASAP7_75t_R FILLER_0_255_852 ();
 FILLER_ASAP7_75t_R FILLER_0_255_859 ();
 FILLER_ASAP7_75t_R FILLER_0_255_866 ();
 FILLER_ASAP7_75t_R FILLER_0_255_878 ();
 FILLER_ASAP7_75t_R FILLER_0_255_890 ();
 FILLER_ASAP7_75t_R FILLER_0_255_902 ();
 FILLER_ASAP7_75t_R FILLER_0_255_914 ();
 FILLER_ASAP7_75t_R FILLER_0_255_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_255_924 ();
 FILLER_ASAP7_75t_R FILLER_0_255_927 ();
 FILLER_ASAP7_75t_R FILLER_0_255_935 ();
 FILLER_ASAP7_75t_R FILLER_0_255_947 ();
 DECAPx2_ASAP7_75t_R FILLER_0_255_955 ();
 DECAPx2_ASAP7_75t_R FILLER_0_255_966 ();
 FILLER_ASAP7_75t_R FILLER_0_255_977 ();
 FILLER_ASAP7_75t_R FILLER_0_255_985 ();
 DECAPx2_ASAP7_75t_R FILLER_0_255_997 ();
 FILLER_ASAP7_75t_R FILLER_0_255_1011 ();
 FILLER_ASAP7_75t_R FILLER_0_255_1023 ();
 DECAPx1_ASAP7_75t_R FILLER_0_255_1031 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_255_1035 ();
 DECAPx4_ASAP7_75t_R FILLER_0_255_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_255_1054 ();
 DECAPx2_ASAP7_75t_R FILLER_0_255_1061 ();
 FILLER_ASAP7_75t_R FILLER_0_255_1077 ();
 FILLER_ASAP7_75t_R FILLER_0_255_1085 ();
 FILLER_ASAP7_75t_R FILLER_0_255_1095 ();
 FILLER_ASAP7_75t_R FILLER_0_255_1102 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_255_1104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_255_1111 ();
 DECAPx6_ASAP7_75t_R FILLER_0_255_1133 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_255_1147 ();
 FILLER_ASAP7_75t_R FILLER_0_255_1158 ();
 FILLER_ASAP7_75t_R FILLER_0_255_1166 ();
 DECAPx2_ASAP7_75t_R FILLER_0_255_1178 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_255_1184 ();
 FILLER_ASAP7_75t_R FILLER_0_255_1193 ();
 FILLER_ASAP7_75t_R FILLER_0_255_1201 ();
 FILLER_ASAP7_75t_R FILLER_0_255_1209 ();
 DECAPx2_ASAP7_75t_R FILLER_0_255_1217 ();
 DECAPx1_ASAP7_75t_R FILLER_0_255_1230 ();
 DECAPx6_ASAP7_75t_R FILLER_0_255_1242 ();
 FILLER_ASAP7_75t_R FILLER_0_255_1266 ();
 DECAPx4_ASAP7_75t_R FILLER_0_255_1274 ();
 FILLER_ASAP7_75t_R FILLER_0_255_1284 ();
 DECAPx6_ASAP7_75t_R FILLER_0_255_1295 ();
 DECAPx2_ASAP7_75t_R FILLER_0_255_1309 ();
 DECAPx1_ASAP7_75t_R FILLER_0_255_1322 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_255_1326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_255_1334 ();
 DECAPx2_ASAP7_75t_R FILLER_0_255_1356 ();
 DECAPx6_ASAP7_75t_R FILLER_0_255_1368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_256_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_256_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_256_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_256_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_256_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_256_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_256_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_256_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_256_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_256_200 ();
 DECAPx6_ASAP7_75t_R FILLER_0_256_222 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_242 ();
 FILLER_ASAP7_75t_R FILLER_0_256_251 ();
 FILLER_ASAP7_75t_R FILLER_0_256_271 ();
 FILLER_ASAP7_75t_R FILLER_0_256_279 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_287 ();
 FILLER_ASAP7_75t_R FILLER_0_256_301 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_309 ();
 FILLER_ASAP7_75t_R FILLER_0_256_321 ();
 FILLER_ASAP7_75t_R FILLER_0_256_328 ();
 FILLER_ASAP7_75t_R FILLER_0_256_336 ();
 FILLER_ASAP7_75t_R FILLER_0_256_341 ();
 FILLER_ASAP7_75t_R FILLER_0_256_348 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_362 ();
 FILLER_ASAP7_75t_R FILLER_0_256_368 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_382 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_389 ();
 FILLER_ASAP7_75t_R FILLER_0_256_395 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_403 ();
 FILLER_ASAP7_75t_R FILLER_0_256_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_411 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_418 ();
 FILLER_ASAP7_75t_R FILLER_0_256_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_426 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_433 ();
 FILLER_ASAP7_75t_R FILLER_0_256_439 ();
 FILLER_ASAP7_75t_R FILLER_0_256_448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_456 ();
 FILLER_ASAP7_75t_R FILLER_0_256_464 ();
 FILLER_ASAP7_75t_R FILLER_0_256_472 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_256_496 ();
 DECAPx1_ASAP7_75t_R FILLER_0_256_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_522 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_526 ();
 DECAPx1_ASAP7_75t_R FILLER_0_256_535 ();
 FILLER_ASAP7_75t_R FILLER_0_256_551 ();
 DECAPx1_ASAP7_75t_R FILLER_0_256_556 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_567 ();
 FILLER_ASAP7_75t_R FILLER_0_256_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_575 ();
 FILLER_ASAP7_75t_R FILLER_0_256_587 ();
 DECAPx1_ASAP7_75t_R FILLER_0_256_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_596 ();
 DECAPx1_ASAP7_75t_R FILLER_0_256_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_607 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_626 ();
 DECAPx1_ASAP7_75t_R FILLER_0_256_639 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_661 ();
 DECAPx4_ASAP7_75t_R FILLER_0_256_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_684 ();
 FILLER_ASAP7_75t_R FILLER_0_256_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_698 ();
 DECAPx6_ASAP7_75t_R FILLER_0_256_707 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_721 ();
 DECAPx4_ASAP7_75t_R FILLER_0_256_733 ();
 FILLER_ASAP7_75t_R FILLER_0_256_751 ();
 FILLER_ASAP7_75t_R FILLER_0_256_761 ();
 DECAPx6_ASAP7_75t_R FILLER_0_256_769 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_783 ();
 DECAPx6_ASAP7_75t_R FILLER_0_256_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_256_819 ();
 DECAPx6_ASAP7_75t_R FILLER_0_256_841 ();
 FILLER_ASAP7_75t_R FILLER_0_256_855 ();
 FILLER_ASAP7_75t_R FILLER_0_256_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_869 ();
 FILLER_ASAP7_75t_R FILLER_0_256_880 ();
 DECAPx1_ASAP7_75t_R FILLER_0_256_892 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_920 ();
 FILLER_ASAP7_75t_R FILLER_0_256_928 ();
 FILLER_ASAP7_75t_R FILLER_0_256_936 ();
 DECAPx1_ASAP7_75t_R FILLER_0_256_948 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_952 ();
 FILLER_ASAP7_75t_R FILLER_0_256_956 ();
 FILLER_ASAP7_75t_R FILLER_0_256_964 ();
 FILLER_ASAP7_75t_R FILLER_0_256_976 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_978 ();
 FILLER_ASAP7_75t_R FILLER_0_256_984 ();
 FILLER_ASAP7_75t_R FILLER_0_256_994 ();
 FILLER_ASAP7_75t_R FILLER_0_256_1004 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_1006 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_1014 ();
 FILLER_ASAP7_75t_R FILLER_0_256_1030 ();
 FILLER_ASAP7_75t_R FILLER_0_256_1038 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_1046 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_1062 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_1068 ();
 FILLER_ASAP7_75t_R FILLER_0_256_1076 ();
 FILLER_ASAP7_75t_R FILLER_0_256_1084 ();
 FILLER_ASAP7_75t_R FILLER_0_256_1092 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_1114 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_1120 ();
 FILLER_ASAP7_75t_R FILLER_0_256_1141 ();
 DECAPx4_ASAP7_75t_R FILLER_0_256_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_1163 ();
 FILLER_ASAP7_75t_R FILLER_0_256_1174 ();
 FILLER_ASAP7_75t_R FILLER_0_256_1181 ();
 FILLER_ASAP7_75t_R FILLER_0_256_1188 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_1190 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_1199 ();
 FILLER_ASAP7_75t_R FILLER_0_256_1205 ();
 DECAPx1_ASAP7_75t_R FILLER_0_256_1214 ();
 FILLER_ASAP7_75t_R FILLER_0_256_1223 ();
 FILLER_ASAP7_75t_R FILLER_0_256_1231 ();
 FILLER_ASAP7_75t_R FILLER_0_256_1239 ();
 DECAPx1_ASAP7_75t_R FILLER_0_256_1248 ();
 FILLER_ASAP7_75t_R FILLER_0_256_1259 ();
 FILLER_ASAP7_75t_R FILLER_0_256_1271 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_1281 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_1287 ();
 DECAPx2_ASAP7_75t_R FILLER_0_256_1294 ();
 FILLER_ASAP7_75t_R FILLER_0_256_1308 ();
 FILLER_ASAP7_75t_R FILLER_0_256_1322 ();
 DECAPx6_ASAP7_75t_R FILLER_0_256_1329 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_1343 ();
 FILLER_ASAP7_75t_R FILLER_0_256_1354 ();
 FILLER_ASAP7_75t_R FILLER_0_256_1364 ();
 DECAPx1_ASAP7_75t_R FILLER_0_256_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_257_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_257_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_257_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_257_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_257_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_257_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_257_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_257_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_257_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_257_200 ();
 DECAPx6_ASAP7_75t_R FILLER_0_257_222 ();
 DECAPx2_ASAP7_75t_R FILLER_0_257_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_242 ();
 FILLER_ASAP7_75t_R FILLER_0_257_255 ();
 FILLER_ASAP7_75t_R FILLER_0_257_263 ();
 DECAPx1_ASAP7_75t_R FILLER_0_257_276 ();
 FILLER_ASAP7_75t_R FILLER_0_257_286 ();
 DECAPx2_ASAP7_75t_R FILLER_0_257_298 ();
 FILLER_ASAP7_75t_R FILLER_0_257_304 ();
 DECAPx4_ASAP7_75t_R FILLER_0_257_312 ();
 DECAPx1_ASAP7_75t_R FILLER_0_257_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_332 ();
 FILLER_ASAP7_75t_R FILLER_0_257_344 ();
 FILLER_ASAP7_75t_R FILLER_0_257_349 ();
 DECAPx2_ASAP7_75t_R FILLER_0_257_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_367 ();
 DECAPx2_ASAP7_75t_R FILLER_0_257_378 ();
 FILLER_ASAP7_75t_R FILLER_0_257_391 ();
 DECAPx2_ASAP7_75t_R FILLER_0_257_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_410 ();
 FILLER_ASAP7_75t_R FILLER_0_257_417 ();
 FILLER_ASAP7_75t_R FILLER_0_257_425 ();
 FILLER_ASAP7_75t_R FILLER_0_257_433 ();
 DECAPx4_ASAP7_75t_R FILLER_0_257_445 ();
 FILLER_ASAP7_75t_R FILLER_0_257_455 ();
 FILLER_ASAP7_75t_R FILLER_0_257_463 ();
 FILLER_ASAP7_75t_R FILLER_0_257_475 ();
 DECAPx6_ASAP7_75t_R FILLER_0_257_483 ();
 FILLER_ASAP7_75t_R FILLER_0_257_497 ();
 DECAPx1_ASAP7_75t_R FILLER_0_257_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_506 ();
 FILLER_ASAP7_75t_R FILLER_0_257_513 ();
 FILLER_ASAP7_75t_R FILLER_0_257_518 ();
 FILLER_ASAP7_75t_R FILLER_0_257_542 ();
 FILLER_ASAP7_75t_R FILLER_0_257_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_551 ();
 FILLER_ASAP7_75t_R FILLER_0_257_558 ();
 FILLER_ASAP7_75t_R FILLER_0_257_566 ();
 DECAPx2_ASAP7_75t_R FILLER_0_257_571 ();
 FILLER_ASAP7_75t_R FILLER_0_257_580 ();
 DECAPx6_ASAP7_75t_R FILLER_0_257_585 ();
 DECAPx1_ASAP7_75t_R FILLER_0_257_599 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_603 ();
 DECAPx1_ASAP7_75t_R FILLER_0_257_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_614 ();
 DECAPx2_ASAP7_75t_R FILLER_0_257_637 ();
 DECAPx2_ASAP7_75t_R FILLER_0_257_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_661 ();
 DECAPx2_ASAP7_75t_R FILLER_0_257_674 ();
 FILLER_ASAP7_75t_R FILLER_0_257_701 ();
 DECAPx1_ASAP7_75t_R FILLER_0_257_711 ();
 DECAPx6_ASAP7_75t_R FILLER_0_257_723 ();
 DECAPx2_ASAP7_75t_R FILLER_0_257_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_743 ();
 DECAPx6_ASAP7_75t_R FILLER_0_257_756 ();
 FILLER_ASAP7_75t_R FILLER_0_257_770 ();
 DECAPx2_ASAP7_75t_R FILLER_0_257_776 ();
 FILLER_ASAP7_75t_R FILLER_0_257_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_784 ();
 FILLER_ASAP7_75t_R FILLER_0_257_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_793 ();
 FILLER_ASAP7_75t_R FILLER_0_257_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_257_817 ();
 DECAPx1_ASAP7_75t_R FILLER_0_257_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_843 ();
 FILLER_ASAP7_75t_R FILLER_0_257_865 ();
 DECAPx1_ASAP7_75t_R FILLER_0_257_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_881 ();
 FILLER_ASAP7_75t_R FILLER_0_257_892 ();
 FILLER_ASAP7_75t_R FILLER_0_257_904 ();
 FILLER_ASAP7_75t_R FILLER_0_257_916 ();
 FILLER_ASAP7_75t_R FILLER_0_257_923 ();
 FILLER_ASAP7_75t_R FILLER_0_257_927 ();
 FILLER_ASAP7_75t_R FILLER_0_257_935 ();
 FILLER_ASAP7_75t_R FILLER_0_257_943 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_945 ();
 DECAPx1_ASAP7_75t_R FILLER_0_257_954 ();
 FILLER_ASAP7_75t_R FILLER_0_257_964 ();
 FILLER_ASAP7_75t_R FILLER_0_257_976 ();
 FILLER_ASAP7_75t_R FILLER_0_257_982 ();
 DECAPx1_ASAP7_75t_R FILLER_0_257_994 ();
 DECAPx2_ASAP7_75t_R FILLER_0_257_1010 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_1016 ();
 DECAPx1_ASAP7_75t_R FILLER_0_257_1027 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_1031 ();
 DECAPx1_ASAP7_75t_R FILLER_0_257_1040 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_1044 ();
 FILLER_ASAP7_75t_R FILLER_0_257_1050 ();
 DECAPx1_ASAP7_75t_R FILLER_0_257_1060 ();
 FILLER_ASAP7_75t_R FILLER_0_257_1074 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_1076 ();
 FILLER_ASAP7_75t_R FILLER_0_257_1080 ();
 FILLER_ASAP7_75t_R FILLER_0_257_1092 ();
 FILLER_ASAP7_75t_R FILLER_0_257_1104 ();
 FILLER_ASAP7_75t_R FILLER_0_257_1116 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_1118 ();
 FILLER_ASAP7_75t_R FILLER_0_257_1122 ();
 FILLER_ASAP7_75t_R FILLER_0_257_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_1132 ();
 DECAPx1_ASAP7_75t_R FILLER_0_257_1139 ();
 DECAPx1_ASAP7_75t_R FILLER_0_257_1149 ();
 DECAPx1_ASAP7_75t_R FILLER_0_257_1173 ();
 FILLER_ASAP7_75t_R FILLER_0_257_1184 ();
 FILLER_ASAP7_75t_R FILLER_0_257_1191 ();
 DECAPx2_ASAP7_75t_R FILLER_0_257_1198 ();
 FILLER_ASAP7_75t_R FILLER_0_257_1204 ();
 DECAPx1_ASAP7_75t_R FILLER_0_257_1213 ();
 FILLER_ASAP7_75t_R FILLER_0_257_1225 ();
 FILLER_ASAP7_75t_R FILLER_0_257_1234 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_1236 ();
 DECAPx4_ASAP7_75t_R FILLER_0_257_1243 ();
 FILLER_ASAP7_75t_R FILLER_0_257_1253 ();
 FILLER_ASAP7_75t_R FILLER_0_257_1260 ();
 FILLER_ASAP7_75t_R FILLER_0_257_1272 ();
 FILLER_ASAP7_75t_R FILLER_0_257_1279 ();
 DECAPx10_ASAP7_75t_R FILLER_0_257_1288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_257_1310 ();
 FILLER_ASAP7_75t_R FILLER_0_257_1332 ();
 FILLER_ASAP7_75t_R FILLER_0_257_1340 ();
 DECAPx1_ASAP7_75t_R FILLER_0_257_1348 ();
 FILLER_ASAP7_75t_R FILLER_0_257_1362 ();
 DECAPx2_ASAP7_75t_R FILLER_0_257_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_258_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_258_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_258_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_258_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_258_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_258_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_258_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_258_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_258_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_258_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_258_222 ();
 FILLER_ASAP7_75t_R FILLER_0_258_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_246 ();
 FILLER_ASAP7_75t_R FILLER_0_258_253 ();
 FILLER_ASAP7_75t_R FILLER_0_258_275 ();
 FILLER_ASAP7_75t_R FILLER_0_258_288 ();
 DECAPx4_ASAP7_75t_R FILLER_0_258_296 ();
 DECAPx2_ASAP7_75t_R FILLER_0_258_317 ();
 FILLER_ASAP7_75t_R FILLER_0_258_323 ();
 DECAPx6_ASAP7_75t_R FILLER_0_258_331 ();
 DECAPx2_ASAP7_75t_R FILLER_0_258_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_351 ();
 FILLER_ASAP7_75t_R FILLER_0_258_358 ();
 DECAPx2_ASAP7_75t_R FILLER_0_258_367 ();
 FILLER_ASAP7_75t_R FILLER_0_258_383 ();
 DECAPx2_ASAP7_75t_R FILLER_0_258_390 ();
 DECAPx1_ASAP7_75t_R FILLER_0_258_402 ();
 FILLER_ASAP7_75t_R FILLER_0_258_412 ();
 FILLER_ASAP7_75t_R FILLER_0_258_420 ();
 FILLER_ASAP7_75t_R FILLER_0_258_428 ();
 FILLER_ASAP7_75t_R FILLER_0_258_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_442 ();
 DECAPx1_ASAP7_75t_R FILLER_0_258_449 ();
 FILLER_ASAP7_75t_R FILLER_0_258_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_461 ();
 FILLER_ASAP7_75t_R FILLER_0_258_464 ();
 FILLER_ASAP7_75t_R FILLER_0_258_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_475 ();
 DECAPx2_ASAP7_75t_R FILLER_0_258_482 ();
 FILLER_ASAP7_75t_R FILLER_0_258_488 ();
 FILLER_ASAP7_75t_R FILLER_0_258_495 ();
 FILLER_ASAP7_75t_R FILLER_0_258_500 ();
 FILLER_ASAP7_75t_R FILLER_0_258_508 ();
 DECAPx1_ASAP7_75t_R FILLER_0_258_515 ();
 FILLER_ASAP7_75t_R FILLER_0_258_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_533 ();
 FILLER_ASAP7_75t_R FILLER_0_258_546 ();
 FILLER_ASAP7_75t_R FILLER_0_258_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_553 ();
 FILLER_ASAP7_75t_R FILLER_0_258_566 ();
 DECAPx2_ASAP7_75t_R FILLER_0_258_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_595 ();
 FILLER_ASAP7_75t_R FILLER_0_258_602 ();
 DECAPx2_ASAP7_75t_R FILLER_0_258_607 ();
 FILLER_ASAP7_75t_R FILLER_0_258_619 ();
 DECAPx2_ASAP7_75t_R FILLER_0_258_624 ();
 DECAPx2_ASAP7_75t_R FILLER_0_258_642 ();
 FILLER_ASAP7_75t_R FILLER_0_258_648 ();
 DECAPx2_ASAP7_75t_R FILLER_0_258_671 ();
 FILLER_ASAP7_75t_R FILLER_0_258_677 ();
 FILLER_ASAP7_75t_R FILLER_0_258_685 ();
 DECAPx6_ASAP7_75t_R FILLER_0_258_690 ();
 FILLER_ASAP7_75t_R FILLER_0_258_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_706 ();
 FILLER_ASAP7_75t_R FILLER_0_258_715 ();
 DECAPx10_ASAP7_75t_R FILLER_0_258_725 ();
 DECAPx6_ASAP7_75t_R FILLER_0_258_747 ();
 FILLER_ASAP7_75t_R FILLER_0_258_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_763 ();
 FILLER_ASAP7_75t_R FILLER_0_258_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_771 ();
 DECAPx2_ASAP7_75t_R FILLER_0_258_782 ();
 DECAPx2_ASAP7_75t_R FILLER_0_258_800 ();
 FILLER_ASAP7_75t_R FILLER_0_258_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_811 ();
 DECAPx2_ASAP7_75t_R FILLER_0_258_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_826 ();
 FILLER_ASAP7_75t_R FILLER_0_258_839 ();
 FILLER_ASAP7_75t_R FILLER_0_258_853 ();
 DECAPx4_ASAP7_75t_R FILLER_0_258_858 ();
 FILLER_ASAP7_75t_R FILLER_0_258_868 ();
 FILLER_ASAP7_75t_R FILLER_0_258_875 ();
 FILLER_ASAP7_75t_R FILLER_0_258_883 ();
 FILLER_ASAP7_75t_R FILLER_0_258_909 ();
 FILLER_ASAP7_75t_R FILLER_0_258_921 ();
 DECAPx2_ASAP7_75t_R FILLER_0_258_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_935 ();
 DECAPx10_ASAP7_75t_R FILLER_0_258_947 ();
 FILLER_ASAP7_75t_R FILLER_0_258_969 ();
 FILLER_ASAP7_75t_R FILLER_0_258_989 ();
 FILLER_ASAP7_75t_R FILLER_0_258_996 ();
 FILLER_ASAP7_75t_R FILLER_0_258_1018 ();
 DECAPx1_ASAP7_75t_R FILLER_0_258_1028 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_1032 ();
 FILLER_ASAP7_75t_R FILLER_0_258_1039 ();
 DECAPx2_ASAP7_75t_R FILLER_0_258_1046 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_1052 ();
 FILLER_ASAP7_75t_R FILLER_0_258_1063 ();
 FILLER_ASAP7_75t_R FILLER_0_258_1071 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_1073 ();
 FILLER_ASAP7_75t_R FILLER_0_258_1084 ();
 FILLER_ASAP7_75t_R FILLER_0_258_1098 ();
 FILLER_ASAP7_75t_R FILLER_0_258_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_0_258_1122 ();
 FILLER_ASAP7_75t_R FILLER_0_258_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_1146 ();
 FILLER_ASAP7_75t_R FILLER_0_258_1153 ();
 DECAPx2_ASAP7_75t_R FILLER_0_258_1158 ();
 FILLER_ASAP7_75t_R FILLER_0_258_1164 ();
 FILLER_ASAP7_75t_R FILLER_0_258_1172 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_1174 ();
 FILLER_ASAP7_75t_R FILLER_0_258_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_1183 ();
 DECAPx2_ASAP7_75t_R FILLER_0_258_1195 ();
 FILLER_ASAP7_75t_R FILLER_0_258_1207 ();
 FILLER_ASAP7_75t_R FILLER_0_258_1215 ();
 DECAPx6_ASAP7_75t_R FILLER_0_258_1223 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_1237 ();
 DECAPx6_ASAP7_75t_R FILLER_0_258_1244 ();
 FILLER_ASAP7_75t_R FILLER_0_258_1258 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_1260 ();
 DECAPx2_ASAP7_75t_R FILLER_0_258_1269 ();
 DECAPx2_ASAP7_75t_R FILLER_0_258_1281 ();
 FILLER_ASAP7_75t_R FILLER_0_258_1295 ();
 FILLER_ASAP7_75t_R FILLER_0_258_1303 ();
 FILLER_ASAP7_75t_R FILLER_0_258_1311 ();
 FILLER_ASAP7_75t_R FILLER_0_258_1320 ();
 FILLER_ASAP7_75t_R FILLER_0_258_1328 ();
 FILLER_ASAP7_75t_R FILLER_0_258_1337 ();
 DECAPx4_ASAP7_75t_R FILLER_0_258_1349 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_1359 ();
 DECAPx6_ASAP7_75t_R FILLER_0_258_1366 ();
 FILLER_ASAP7_75t_R FILLER_0_258_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_259_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_259_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_259_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_259_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_259_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_259_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_259_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_259_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_259_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_259_200 ();
 DECAPx6_ASAP7_75t_R FILLER_0_259_222 ();
 DECAPx2_ASAP7_75t_R FILLER_0_259_236 ();
 FILLER_ASAP7_75t_R FILLER_0_259_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_259_256 ();
 DECAPx2_ASAP7_75t_R FILLER_0_259_263 ();
 FILLER_ASAP7_75t_R FILLER_0_259_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_259_271 ();
 FILLER_ASAP7_75t_R FILLER_0_259_280 ();
 DECAPx6_ASAP7_75t_R FILLER_0_259_287 ();
 FILLER_ASAP7_75t_R FILLER_0_259_307 ();
 DECAPx1_ASAP7_75t_R FILLER_0_259_329 ();
 FILLER_ASAP7_75t_R FILLER_0_259_337 ();
 DECAPx4_ASAP7_75t_R FILLER_0_259_346 ();
 FILLER_ASAP7_75t_R FILLER_0_259_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_259_358 ();
 DECAPx2_ASAP7_75t_R FILLER_0_259_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_259_372 ();
 FILLER_ASAP7_75t_R FILLER_0_259_385 ();
 FILLER_ASAP7_75t_R FILLER_0_259_392 ();
 FILLER_ASAP7_75t_R FILLER_0_259_399 ();
 FILLER_ASAP7_75t_R FILLER_0_259_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_259_406 ();
 FILLER_ASAP7_75t_R FILLER_0_259_413 ();
 DECAPx2_ASAP7_75t_R FILLER_0_259_421 ();
 FILLER_ASAP7_75t_R FILLER_0_259_432 ();
 DECAPx1_ASAP7_75t_R FILLER_0_259_440 ();
 FILLER_ASAP7_75t_R FILLER_0_259_454 ();
 DECAPx6_ASAP7_75t_R FILLER_0_259_461 ();
 DECAPx1_ASAP7_75t_R FILLER_0_259_475 ();
 FILLER_ASAP7_75t_R FILLER_0_259_485 ();
 FILLER_ASAP7_75t_R FILLER_0_259_497 ();
 DECAPx1_ASAP7_75t_R FILLER_0_259_504 ();
 FILLER_ASAP7_75t_R FILLER_0_259_513 ();
 FILLER_ASAP7_75t_R FILLER_0_259_520 ();
 FILLER_ASAP7_75t_R FILLER_0_259_528 ();
 FILLER_ASAP7_75t_R FILLER_0_259_533 ();
 DECAPx1_ASAP7_75t_R FILLER_0_259_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_259_551 ();
 FILLER_ASAP7_75t_R FILLER_0_259_557 ();
 FILLER_ASAP7_75t_R FILLER_0_259_570 ();
 DECAPx2_ASAP7_75t_R FILLER_0_259_578 ();
 FILLER_ASAP7_75t_R FILLER_0_259_605 ();
 FILLER_ASAP7_75t_R FILLER_0_259_610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_259_615 ();
 DECAPx6_ASAP7_75t_R FILLER_0_259_637 ();
 FILLER_ASAP7_75t_R FILLER_0_259_657 ();
 DECAPx6_ASAP7_75t_R FILLER_0_259_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_259_676 ();
 DECAPx4_ASAP7_75t_R FILLER_0_259_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_259_693 ();
 DECAPx6_ASAP7_75t_R FILLER_0_259_700 ();
 FILLER_ASAP7_75t_R FILLER_0_259_714 ();
 FILLER_ASAP7_75t_R FILLER_0_259_724 ();
 DECAPx2_ASAP7_75t_R FILLER_0_259_734 ();
 FILLER_ASAP7_75t_R FILLER_0_259_740 ();
 DECAPx4_ASAP7_75t_R FILLER_0_259_746 ();
 FILLER_ASAP7_75t_R FILLER_0_259_756 ();
 FILLER_ASAP7_75t_R FILLER_0_259_770 ();
 DECAPx4_ASAP7_75t_R FILLER_0_259_778 ();
 FILLER_ASAP7_75t_R FILLER_0_259_788 ();
 FILLER_ASAP7_75t_R FILLER_0_259_796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_259_804 ();
 DECAPx10_ASAP7_75t_R FILLER_0_259_826 ();
 DECAPx2_ASAP7_75t_R FILLER_0_259_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_259_860 ();
 DECAPx2_ASAP7_75t_R FILLER_0_259_871 ();
 FILLER_ASAP7_75t_R FILLER_0_259_882 ();
 DECAPx1_ASAP7_75t_R FILLER_0_259_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_259_893 ();
 FILLER_ASAP7_75t_R FILLER_0_259_900 ();
 DECAPx1_ASAP7_75t_R FILLER_0_259_907 ();
 DECAPx2_ASAP7_75t_R FILLER_0_259_917 ();
 FILLER_ASAP7_75t_R FILLER_0_259_923 ();
 FILLER_ASAP7_75t_R FILLER_0_259_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_259_929 ();
 FILLER_ASAP7_75t_R FILLER_0_259_941 ();
 FILLER_ASAP7_75t_R FILLER_0_259_949 ();
 FILLER_ASAP7_75t_R FILLER_0_259_957 ();
 DECAPx1_ASAP7_75t_R FILLER_0_259_965 ();
 FILLER_ASAP7_75t_R FILLER_0_259_975 ();
 DECAPx4_ASAP7_75t_R FILLER_0_259_984 ();
 FILLER_ASAP7_75t_R FILLER_0_259_1001 ();
 FILLER_ASAP7_75t_R FILLER_0_259_1013 ();
 FILLER_ASAP7_75t_R FILLER_0_259_1020 ();
 FILLER_ASAP7_75t_R FILLER_0_259_1046 ();
 FILLER_ASAP7_75t_R FILLER_0_259_1068 ();
 FILLER_ASAP7_75t_R FILLER_0_259_1076 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_259_1078 ();
 FILLER_ASAP7_75t_R FILLER_0_259_1089 ();
 FILLER_ASAP7_75t_R FILLER_0_259_1099 ();
 FILLER_ASAP7_75t_R FILLER_0_259_1122 ();
 DECAPx4_ASAP7_75t_R FILLER_0_259_1134 ();
 FILLER_ASAP7_75t_R FILLER_0_259_1144 ();
 FILLER_ASAP7_75t_R FILLER_0_259_1152 ();
 DECAPx4_ASAP7_75t_R FILLER_0_259_1160 ();
 FILLER_ASAP7_75t_R FILLER_0_259_1170 ();
 DECAPx1_ASAP7_75t_R FILLER_0_259_1178 ();
 FILLER_ASAP7_75t_R FILLER_0_259_1192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_259_1200 ();
 FILLER_ASAP7_75t_R FILLER_0_259_1220 ();
 DECAPx6_ASAP7_75t_R FILLER_0_259_1228 ();
 FILLER_ASAP7_75t_R FILLER_0_259_1252 ();
 DECAPx1_ASAP7_75t_R FILLER_0_259_1260 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_259_1264 ();
 DECAPx1_ASAP7_75t_R FILLER_0_259_1271 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_259_1275 ();
 FILLER_ASAP7_75t_R FILLER_0_259_1281 ();
 FILLER_ASAP7_75t_R FILLER_0_259_1295 ();
 DECAPx2_ASAP7_75t_R FILLER_0_259_1305 ();
 FILLER_ASAP7_75t_R FILLER_0_259_1311 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_259_1313 ();
 FILLER_ASAP7_75t_R FILLER_0_259_1326 ();
 DECAPx1_ASAP7_75t_R FILLER_0_259_1334 ();
 DECAPx4_ASAP7_75t_R FILLER_0_259_1348 ();
 FILLER_ASAP7_75t_R FILLER_0_259_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_260_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_260_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_260_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_260_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_260_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_260_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_260_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_260_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_260_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_260_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_260_222 ();
 DECAPx2_ASAP7_75t_R FILLER_0_260_244 ();
 FILLER_ASAP7_75t_R FILLER_0_260_258 ();
 DECAPx1_ASAP7_75t_R FILLER_0_260_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_260_270 ();
 DECAPx6_ASAP7_75t_R FILLER_0_260_277 ();
 FILLER_ASAP7_75t_R FILLER_0_260_291 ();
 DECAPx4_ASAP7_75t_R FILLER_0_260_301 ();
 FILLER_ASAP7_75t_R FILLER_0_260_323 ();
 FILLER_ASAP7_75t_R FILLER_0_260_331 ();
 FILLER_ASAP7_75t_R FILLER_0_260_338 ();
 DECAPx1_ASAP7_75t_R FILLER_0_260_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_260_354 ();
 FILLER_ASAP7_75t_R FILLER_0_260_365 ();
 FILLER_ASAP7_75t_R FILLER_0_260_379 ();
 DECAPx6_ASAP7_75t_R FILLER_0_260_393 ();
 FILLER_ASAP7_75t_R FILLER_0_260_407 ();
 DECAPx6_ASAP7_75t_R FILLER_0_260_415 ();
 FILLER_ASAP7_75t_R FILLER_0_260_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_260_437 ();
 DECAPx4_ASAP7_75t_R FILLER_0_260_444 ();
 FILLER_ASAP7_75t_R FILLER_0_260_460 ();
 DECAPx2_ASAP7_75t_R FILLER_0_260_464 ();
 FILLER_ASAP7_75t_R FILLER_0_260_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_260_472 ();
 FILLER_ASAP7_75t_R FILLER_0_260_478 ();
 FILLER_ASAP7_75t_R FILLER_0_260_486 ();
 DECAPx1_ASAP7_75t_R FILLER_0_260_498 ();
 FILLER_ASAP7_75t_R FILLER_0_260_508 ();
 FILLER_ASAP7_75t_R FILLER_0_260_513 ();
 FILLER_ASAP7_75t_R FILLER_0_260_537 ();
 FILLER_ASAP7_75t_R FILLER_0_260_551 ();
 FILLER_ASAP7_75t_R FILLER_0_260_558 ();
 DECAPx1_ASAP7_75t_R FILLER_0_260_565 ();
 FILLER_ASAP7_75t_R FILLER_0_260_575 ();
 FILLER_ASAP7_75t_R FILLER_0_260_582 ();
 FILLER_ASAP7_75t_R FILLER_0_260_590 ();
 FILLER_ASAP7_75t_R FILLER_0_260_597 ();
 FILLER_ASAP7_75t_R FILLER_0_260_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_260_605 ();
 FILLER_ASAP7_75t_R FILLER_0_260_616 ();
 FILLER_ASAP7_75t_R FILLER_0_260_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_260_623 ();
 DECAPx6_ASAP7_75t_R FILLER_0_260_630 ();
 DECAPx4_ASAP7_75t_R FILLER_0_260_650 ();
 DECAPx4_ASAP7_75t_R FILLER_0_260_666 ();
 DECAPx6_ASAP7_75t_R FILLER_0_260_682 ();
 FILLER_ASAP7_75t_R FILLER_0_260_696 ();
 FILLER_ASAP7_75t_R FILLER_0_260_708 ();
 DECAPx4_ASAP7_75t_R FILLER_0_260_720 ();
 FILLER_ASAP7_75t_R FILLER_0_260_738 ();
 FILLER_ASAP7_75t_R FILLER_0_260_743 ();
 FILLER_ASAP7_75t_R FILLER_0_260_756 ();
 FILLER_ASAP7_75t_R FILLER_0_260_770 ();
 DECAPx2_ASAP7_75t_R FILLER_0_260_778 ();
 FILLER_ASAP7_75t_R FILLER_0_260_784 ();
 FILLER_ASAP7_75t_R FILLER_0_260_794 ();
 FILLER_ASAP7_75t_R FILLER_0_260_800 ();
 DECAPx1_ASAP7_75t_R FILLER_0_260_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_260_814 ();
 DECAPx2_ASAP7_75t_R FILLER_0_260_821 ();
 FILLER_ASAP7_75t_R FILLER_0_260_849 ();
 DECAPx2_ASAP7_75t_R FILLER_0_260_854 ();
 FILLER_ASAP7_75t_R FILLER_0_260_860 ();
 FILLER_ASAP7_75t_R FILLER_0_260_872 ();
 FILLER_ASAP7_75t_R FILLER_0_260_880 ();
 FILLER_ASAP7_75t_R FILLER_0_260_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_260_890 ();
 FILLER_ASAP7_75t_R FILLER_0_260_897 ();
 FILLER_ASAP7_75t_R FILLER_0_260_905 ();
 FILLER_ASAP7_75t_R FILLER_0_260_913 ();
 FILLER_ASAP7_75t_R FILLER_0_260_921 ();
 FILLER_ASAP7_75t_R FILLER_0_260_929 ();
 DECAPx2_ASAP7_75t_R FILLER_0_260_937 ();
 FILLER_ASAP7_75t_R FILLER_0_260_949 ();
 DECAPx2_ASAP7_75t_R FILLER_0_260_959 ();
 DECAPx4_ASAP7_75t_R FILLER_0_260_977 ();
 FILLER_ASAP7_75t_R FILLER_0_260_990 ();
 FILLER_ASAP7_75t_R FILLER_0_260_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_260_1014 ();
 FILLER_ASAP7_75t_R FILLER_0_260_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_260_1023 ();
 DECAPx2_ASAP7_75t_R FILLER_0_260_1031 ();
 FILLER_ASAP7_75t_R FILLER_0_260_1037 ();
 FILLER_ASAP7_75t_R FILLER_0_260_1049 ();
 FILLER_ASAP7_75t_R FILLER_0_260_1061 ();
 FILLER_ASAP7_75t_R FILLER_0_260_1068 ();
 FILLER_ASAP7_75t_R FILLER_0_260_1077 ();
 FILLER_ASAP7_75t_R FILLER_0_260_1089 ();
 FILLER_ASAP7_75t_R FILLER_0_260_1101 ();
 FILLER_ASAP7_75t_R FILLER_0_260_1113 ();
 DECAPx1_ASAP7_75t_R FILLER_0_260_1120 ();
 FILLER_ASAP7_75t_R FILLER_0_260_1134 ();
 DECAPx1_ASAP7_75t_R FILLER_0_260_1139 ();
 FILLER_ASAP7_75t_R FILLER_0_260_1150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_260_1158 ();
 DECAPx6_ASAP7_75t_R FILLER_0_260_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_260_1194 ();
 DECAPx1_ASAP7_75t_R FILLER_0_260_1201 ();
 DECAPx1_ASAP7_75t_R FILLER_0_260_1215 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_260_1219 ();
 DECAPx4_ASAP7_75t_R FILLER_0_260_1223 ();
 FILLER_ASAP7_75t_R FILLER_0_260_1233 ();
 FILLER_ASAP7_75t_R FILLER_0_260_1245 ();
 FILLER_ASAP7_75t_R FILLER_0_260_1253 ();
 DECAPx1_ASAP7_75t_R FILLER_0_260_1261 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_260_1265 ();
 FILLER_ASAP7_75t_R FILLER_0_260_1272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_260_1278 ();
 FILLER_ASAP7_75t_R FILLER_0_260_1306 ();
 DECAPx2_ASAP7_75t_R FILLER_0_260_1319 ();
 FILLER_ASAP7_75t_R FILLER_0_260_1325 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_260_1327 ();
 FILLER_ASAP7_75t_R FILLER_0_260_1338 ();
 FILLER_ASAP7_75t_R FILLER_0_260_1348 ();
 FILLER_ASAP7_75t_R FILLER_0_260_1356 ();
 DECAPx6_ASAP7_75t_R FILLER_0_260_1368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_261_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_261_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_261_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_261_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_261_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_261_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_261_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_261_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_261_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_261_200 ();
 DECAPx6_ASAP7_75t_R FILLER_0_261_222 ();
 FILLER_ASAP7_75t_R FILLER_0_261_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_238 ();
 DECAPx4_ASAP7_75t_R FILLER_0_261_250 ();
 DECAPx4_ASAP7_75t_R FILLER_0_261_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_276 ();
 DECAPx1_ASAP7_75t_R FILLER_0_261_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_287 ();
 FILLER_ASAP7_75t_R FILLER_0_261_294 ();
 FILLER_ASAP7_75t_R FILLER_0_261_302 ();
 FILLER_ASAP7_75t_R FILLER_0_261_314 ();
 FILLER_ASAP7_75t_R FILLER_0_261_322 ();
 DECAPx2_ASAP7_75t_R FILLER_0_261_330 ();
 FILLER_ASAP7_75t_R FILLER_0_261_336 ();
 DECAPx2_ASAP7_75t_R FILLER_0_261_345 ();
 DECAPx1_ASAP7_75t_R FILLER_0_261_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_375 ();
 DECAPx6_ASAP7_75t_R FILLER_0_261_388 ();
 FILLER_ASAP7_75t_R FILLER_0_261_402 ();
 DECAPx2_ASAP7_75t_R FILLER_0_261_411 ();
 FILLER_ASAP7_75t_R FILLER_0_261_417 ();
 DECAPx6_ASAP7_75t_R FILLER_0_261_425 ();
 DECAPx4_ASAP7_75t_R FILLER_0_261_445 ();
 FILLER_ASAP7_75t_R FILLER_0_261_462 ();
 FILLER_ASAP7_75t_R FILLER_0_261_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_472 ();
 DECAPx1_ASAP7_75t_R FILLER_0_261_479 ();
 FILLER_ASAP7_75t_R FILLER_0_261_489 ();
 FILLER_ASAP7_75t_R FILLER_0_261_494 ();
 FILLER_ASAP7_75t_R FILLER_0_261_501 ();
 FILLER_ASAP7_75t_R FILLER_0_261_509 ();
 FILLER_ASAP7_75t_R FILLER_0_261_514 ();
 FILLER_ASAP7_75t_R FILLER_0_261_537 ();
 FILLER_ASAP7_75t_R FILLER_0_261_551 ();
 FILLER_ASAP7_75t_R FILLER_0_261_558 ();
 FILLER_ASAP7_75t_R FILLER_0_261_565 ();
 DECAPx1_ASAP7_75t_R FILLER_0_261_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_583 ();
 FILLER_ASAP7_75t_R FILLER_0_261_589 ();
 FILLER_ASAP7_75t_R FILLER_0_261_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_598 ();
 FILLER_ASAP7_75t_R FILLER_0_261_619 ();
 FILLER_ASAP7_75t_R FILLER_0_261_642 ();
 FILLER_ASAP7_75t_R FILLER_0_261_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_656 ();
 FILLER_ASAP7_75t_R FILLER_0_261_678 ();
 DECAPx2_ASAP7_75t_R FILLER_0_261_701 ();
 FILLER_ASAP7_75t_R FILLER_0_261_711 ();
 FILLER_ASAP7_75t_R FILLER_0_261_723 ();
 FILLER_ASAP7_75t_R FILLER_0_261_733 ();
 FILLER_ASAP7_75t_R FILLER_0_261_743 ();
 DECAPx4_ASAP7_75t_R FILLER_0_261_757 ();
 FILLER_ASAP7_75t_R FILLER_0_261_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_769 ();
 DECAPx2_ASAP7_75t_R FILLER_0_261_778 ();
 FILLER_ASAP7_75t_R FILLER_0_261_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_786 ();
 FILLER_ASAP7_75t_R FILLER_0_261_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_797 ();
 DECAPx4_ASAP7_75t_R FILLER_0_261_806 ();
 FILLER_ASAP7_75t_R FILLER_0_261_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_818 ();
 FILLER_ASAP7_75t_R FILLER_0_261_827 ();
 FILLER_ASAP7_75t_R FILLER_0_261_832 ();
 FILLER_ASAP7_75t_R FILLER_0_261_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_839 ();
 FILLER_ASAP7_75t_R FILLER_0_261_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_845 ();
 DECAPx2_ASAP7_75t_R FILLER_0_261_857 ();
 FILLER_ASAP7_75t_R FILLER_0_261_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_865 ();
 FILLER_ASAP7_75t_R FILLER_0_261_884 ();
 DECAPx2_ASAP7_75t_R FILLER_0_261_894 ();
 FILLER_ASAP7_75t_R FILLER_0_261_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_902 ();
 FILLER_ASAP7_75t_R FILLER_0_261_914 ();
 FILLER_ASAP7_75t_R FILLER_0_261_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_924 ();
 FILLER_ASAP7_75t_R FILLER_0_261_927 ();
 FILLER_ASAP7_75t_R FILLER_0_261_935 ();
 DECAPx2_ASAP7_75t_R FILLER_0_261_943 ();
 FILLER_ASAP7_75t_R FILLER_0_261_969 ();
 FILLER_ASAP7_75t_R FILLER_0_261_981 ();
 FILLER_ASAP7_75t_R FILLER_0_261_989 ();
 FILLER_ASAP7_75t_R FILLER_0_261_997 ();
 FILLER_ASAP7_75t_R FILLER_0_261_1005 ();
 FILLER_ASAP7_75t_R FILLER_0_261_1013 ();
 FILLER_ASAP7_75t_R FILLER_0_261_1021 ();
 FILLER_ASAP7_75t_R FILLER_0_261_1029 ();
 FILLER_ASAP7_75t_R FILLER_0_261_1037 ();
 DECAPx2_ASAP7_75t_R FILLER_0_261_1044 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_1050 ();
 DECAPx2_ASAP7_75t_R FILLER_0_261_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_1063 ();
 FILLER_ASAP7_75t_R FILLER_0_261_1070 ();
 FILLER_ASAP7_75t_R FILLER_0_261_1078 ();
 FILLER_ASAP7_75t_R FILLER_0_261_1090 ();
 FILLER_ASAP7_75t_R FILLER_0_261_1102 ();
 FILLER_ASAP7_75t_R FILLER_0_261_1112 ();
 DECAPx1_ASAP7_75t_R FILLER_0_261_1117 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_1121 ();
 FILLER_ASAP7_75t_R FILLER_0_261_1128 ();
 DECAPx2_ASAP7_75t_R FILLER_0_261_1133 ();
 FILLER_ASAP7_75t_R FILLER_0_261_1139 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_1141 ();
 DECAPx6_ASAP7_75t_R FILLER_0_261_1148 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_1162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_261_1169 ();
 DECAPx1_ASAP7_75t_R FILLER_0_261_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_1195 ();
 DECAPx6_ASAP7_75t_R FILLER_0_261_1202 ();
 FILLER_ASAP7_75t_R FILLER_0_261_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_1218 ();
 DECAPx10_ASAP7_75t_R FILLER_0_261_1229 ();
 DECAPx6_ASAP7_75t_R FILLER_0_261_1251 ();
 FILLER_ASAP7_75t_R FILLER_0_261_1275 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_1277 ();
 FILLER_ASAP7_75t_R FILLER_0_261_1288 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_1290 ();
 DECAPx4_ASAP7_75t_R FILLER_0_261_1301 ();
 FILLER_ASAP7_75t_R FILLER_0_261_1311 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_1313 ();
 DECAPx1_ASAP7_75t_R FILLER_0_261_1320 ();
 FILLER_ASAP7_75t_R FILLER_0_261_1334 ();
 DECAPx2_ASAP7_75t_R FILLER_0_261_1346 ();
 FILLER_ASAP7_75t_R FILLER_0_261_1352 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_1354 ();
 FILLER_ASAP7_75t_R FILLER_0_261_1366 ();
 FILLER_ASAP7_75t_R FILLER_0_261_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_262_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_262_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_262_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_262_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_262_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_262_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_262_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_262_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_262_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_262_200 ();
 DECAPx6_ASAP7_75t_R FILLER_0_262_222 ();
 DECAPx1_ASAP7_75t_R FILLER_0_262_236 ();
 DECAPx2_ASAP7_75t_R FILLER_0_262_250 ();
 FILLER_ASAP7_75t_R FILLER_0_262_256 ();
 FILLER_ASAP7_75t_R FILLER_0_262_264 ();
 FILLER_ASAP7_75t_R FILLER_0_262_272 ();
 FILLER_ASAP7_75t_R FILLER_0_262_285 ();
 DECAPx10_ASAP7_75t_R FILLER_0_262_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_315 ();
 DECAPx1_ASAP7_75t_R FILLER_0_262_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_331 ();
 DECAPx1_ASAP7_75t_R FILLER_0_262_352 ();
 DECAPx1_ASAP7_75t_R FILLER_0_262_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_370 ();
 FILLER_ASAP7_75t_R FILLER_0_262_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_393 ();
 DECAPx1_ASAP7_75t_R FILLER_0_262_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_406 ();
 DECAPx2_ASAP7_75t_R FILLER_0_262_413 ();
 DECAPx2_ASAP7_75t_R FILLER_0_262_425 ();
 FILLER_ASAP7_75t_R FILLER_0_262_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_433 ();
 FILLER_ASAP7_75t_R FILLER_0_262_444 ();
 DECAPx1_ASAP7_75t_R FILLER_0_262_449 ();
 FILLER_ASAP7_75t_R FILLER_0_262_460 ();
 FILLER_ASAP7_75t_R FILLER_0_262_464 ();
 FILLER_ASAP7_75t_R FILLER_0_262_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_474 ();
 FILLER_ASAP7_75t_R FILLER_0_262_480 ();
 FILLER_ASAP7_75t_R FILLER_0_262_502 ();
 DECAPx1_ASAP7_75t_R FILLER_0_262_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_513 ();
 FILLER_ASAP7_75t_R FILLER_0_262_519 ();
 FILLER_ASAP7_75t_R FILLER_0_262_526 ();
 FILLER_ASAP7_75t_R FILLER_0_262_533 ();
 FILLER_ASAP7_75t_R FILLER_0_262_545 ();
 FILLER_ASAP7_75t_R FILLER_0_262_559 ();
 FILLER_ASAP7_75t_R FILLER_0_262_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_568 ();
 DECAPx1_ASAP7_75t_R FILLER_0_262_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_594 ();
 FILLER_ASAP7_75t_R FILLER_0_262_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_602 ();
 DECAPx1_ASAP7_75t_R FILLER_0_262_611 ();
 FILLER_ASAP7_75t_R FILLER_0_262_620 ();
 DECAPx2_ASAP7_75t_R FILLER_0_262_628 ();
 DECAPx1_ASAP7_75t_R FILLER_0_262_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_659 ();
 FILLER_ASAP7_75t_R FILLER_0_262_666 ();
 FILLER_ASAP7_75t_R FILLER_0_262_673 ();
 FILLER_ASAP7_75t_R FILLER_0_262_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_680 ();
 FILLER_ASAP7_75t_R FILLER_0_262_687 ();
 DECAPx4_ASAP7_75t_R FILLER_0_262_695 ();
 FILLER_ASAP7_75t_R FILLER_0_262_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_707 ();
 DECAPx2_ASAP7_75t_R FILLER_0_262_718 ();
 FILLER_ASAP7_75t_R FILLER_0_262_724 ();
 DECAPx1_ASAP7_75t_R FILLER_0_262_734 ();
 DECAPx10_ASAP7_75t_R FILLER_0_262_746 ();
 DECAPx4_ASAP7_75t_R FILLER_0_262_768 ();
 DECAPx10_ASAP7_75t_R FILLER_0_262_783 ();
 DECAPx2_ASAP7_75t_R FILLER_0_262_805 ();
 FILLER_ASAP7_75t_R FILLER_0_262_819 ();
 DECAPx2_ASAP7_75t_R FILLER_0_262_833 ();
 FILLER_ASAP7_75t_R FILLER_0_262_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_841 ();
 DECAPx2_ASAP7_75t_R FILLER_0_262_850 ();
 FILLER_ASAP7_75t_R FILLER_0_262_856 ();
 FILLER_ASAP7_75t_R FILLER_0_262_864 ();
 FILLER_ASAP7_75t_R FILLER_0_262_876 ();
 FILLER_ASAP7_75t_R FILLER_0_262_884 ();
 DECAPx1_ASAP7_75t_R FILLER_0_262_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_896 ();
 DECAPx1_ASAP7_75t_R FILLER_0_262_904 ();
 FILLER_ASAP7_75t_R FILLER_0_262_914 ();
 FILLER_ASAP7_75t_R FILLER_0_262_921 ();
 DECAPx6_ASAP7_75t_R FILLER_0_262_934 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_948 ();
 DECAPx2_ASAP7_75t_R FILLER_0_262_955 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_961 ();
 DECAPx2_ASAP7_75t_R FILLER_0_262_968 ();
 FILLER_ASAP7_75t_R FILLER_0_262_974 ();
 DECAPx6_ASAP7_75t_R FILLER_0_262_981 ();
 DECAPx2_ASAP7_75t_R FILLER_0_262_995 ();
 DECAPx1_ASAP7_75t_R FILLER_0_262_1011 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_1015 ();
 DECAPx1_ASAP7_75t_R FILLER_0_262_1020 ();
 FILLER_ASAP7_75t_R FILLER_0_262_1030 ();
 FILLER_ASAP7_75t_R FILLER_0_262_1038 ();
 DECAPx1_ASAP7_75t_R FILLER_0_262_1045 ();
 FILLER_ASAP7_75t_R FILLER_0_262_1055 ();
 FILLER_ASAP7_75t_R FILLER_0_262_1063 ();
 FILLER_ASAP7_75t_R FILLER_0_262_1085 ();
 FILLER_ASAP7_75t_R FILLER_0_262_1103 ();
 DECAPx6_ASAP7_75t_R FILLER_0_262_1108 ();
 DECAPx1_ASAP7_75t_R FILLER_0_262_1122 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_1126 ();
 DECAPx2_ASAP7_75t_R FILLER_0_262_1133 ();
 DECAPx2_ASAP7_75t_R FILLER_0_262_1142 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_1148 ();
 DECAPx1_ASAP7_75t_R FILLER_0_262_1159 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_1163 ();
 FILLER_ASAP7_75t_R FILLER_0_262_1170 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_1172 ();
 FILLER_ASAP7_75t_R FILLER_0_262_1179 ();
 DECAPx2_ASAP7_75t_R FILLER_0_262_1187 ();
 FILLER_ASAP7_75t_R FILLER_0_262_1199 ();
 DECAPx1_ASAP7_75t_R FILLER_0_262_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_1211 ();
 DECAPx2_ASAP7_75t_R FILLER_0_262_1232 ();
 DECAPx2_ASAP7_75t_R FILLER_0_262_1248 ();
 FILLER_ASAP7_75t_R FILLER_0_262_1260 ();
 DECAPx2_ASAP7_75t_R FILLER_0_262_1273 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_1279 ();
 DECAPx4_ASAP7_75t_R FILLER_0_262_1300 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_1310 ();
 FILLER_ASAP7_75t_R FILLER_0_262_1331 ();
 FILLER_ASAP7_75t_R FILLER_0_262_1343 ();
 FILLER_ASAP7_75t_R FILLER_0_262_1351 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_1353 ();
 DECAPx2_ASAP7_75t_R FILLER_0_262_1360 ();
 FILLER_ASAP7_75t_R FILLER_0_262_1366 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_1368 ();
 DECAPx1_ASAP7_75t_R FILLER_0_262_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_263_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_263_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_263_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_263_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_263_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_263_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_263_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_263_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_263_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_263_200 ();
 DECAPx6_ASAP7_75t_R FILLER_0_263_222 ();
 FILLER_ASAP7_75t_R FILLER_0_263_248 ();
 FILLER_ASAP7_75t_R FILLER_0_263_255 ();
 DECAPx1_ASAP7_75t_R FILLER_0_263_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_267 ();
 FILLER_ASAP7_75t_R FILLER_0_263_274 ();
 FILLER_ASAP7_75t_R FILLER_0_263_282 ();
 FILLER_ASAP7_75t_R FILLER_0_263_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_291 ();
 DECAPx6_ASAP7_75t_R FILLER_0_263_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_312 ();
 FILLER_ASAP7_75t_R FILLER_0_263_319 ();
 DECAPx2_ASAP7_75t_R FILLER_0_263_331 ();
 DECAPx6_ASAP7_75t_R FILLER_0_263_343 ();
 DECAPx1_ASAP7_75t_R FILLER_0_263_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_361 ();
 DECAPx6_ASAP7_75t_R FILLER_0_263_368 ();
 DECAPx1_ASAP7_75t_R FILLER_0_263_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_386 ();
 DECAPx10_ASAP7_75t_R FILLER_0_263_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_416 ();
 DECAPx6_ASAP7_75t_R FILLER_0_263_423 ();
 DECAPx1_ASAP7_75t_R FILLER_0_263_437 ();
 DECAPx2_ASAP7_75t_R FILLER_0_263_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_453 ();
 FILLER_ASAP7_75t_R FILLER_0_263_459 ();
 FILLER_ASAP7_75t_R FILLER_0_263_467 ();
 FILLER_ASAP7_75t_R FILLER_0_263_480 ();
 DECAPx2_ASAP7_75t_R FILLER_0_263_492 ();
 FILLER_ASAP7_75t_R FILLER_0_263_503 ();
 FILLER_ASAP7_75t_R FILLER_0_263_511 ();
 FILLER_ASAP7_75t_R FILLER_0_263_517 ();
 FILLER_ASAP7_75t_R FILLER_0_263_525 ();
 DECAPx2_ASAP7_75t_R FILLER_0_263_533 ();
 FILLER_ASAP7_75t_R FILLER_0_263_544 ();
 FILLER_ASAP7_75t_R FILLER_0_263_551 ();
 DECAPx2_ASAP7_75t_R FILLER_0_263_565 ();
 FILLER_ASAP7_75t_R FILLER_0_263_579 ();
 FILLER_ASAP7_75t_R FILLER_0_263_586 ();
 FILLER_ASAP7_75t_R FILLER_0_263_591 ();
 FILLER_ASAP7_75t_R FILLER_0_263_598 ();
 FILLER_ASAP7_75t_R FILLER_0_263_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_614 ();
 FILLER_ASAP7_75t_R FILLER_0_263_618 ();
 DECAPx2_ASAP7_75t_R FILLER_0_263_630 ();
 FILLER_ASAP7_75t_R FILLER_0_263_642 ();
 FILLER_ASAP7_75t_R FILLER_0_263_650 ();
 FILLER_ASAP7_75t_R FILLER_0_263_658 ();
 DECAPx6_ASAP7_75t_R FILLER_0_263_665 ();
 FILLER_ASAP7_75t_R FILLER_0_263_679 ();
 FILLER_ASAP7_75t_R FILLER_0_263_684 ();
 DECAPx2_ASAP7_75t_R FILLER_0_263_691 ();
 FILLER_ASAP7_75t_R FILLER_0_263_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_699 ();
 FILLER_ASAP7_75t_R FILLER_0_263_706 ();
 DECAPx6_ASAP7_75t_R FILLER_0_263_718 ();
 FILLER_ASAP7_75t_R FILLER_0_263_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_734 ();
 FILLER_ASAP7_75t_R FILLER_0_263_743 ();
 DECAPx10_ASAP7_75t_R FILLER_0_263_753 ();
 DECAPx2_ASAP7_75t_R FILLER_0_263_775 ();
 FILLER_ASAP7_75t_R FILLER_0_263_781 ();
 DECAPx6_ASAP7_75t_R FILLER_0_263_793 ();
 DECAPx1_ASAP7_75t_R FILLER_0_263_807 ();
 FILLER_ASAP7_75t_R FILLER_0_263_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_819 ();
 DECAPx4_ASAP7_75t_R FILLER_0_263_826 ();
 FILLER_ASAP7_75t_R FILLER_0_263_836 ();
 DECAPx6_ASAP7_75t_R FILLER_0_263_850 ();
 DECAPx2_ASAP7_75t_R FILLER_0_263_864 ();
 FILLER_ASAP7_75t_R FILLER_0_263_878 ();
 FILLER_ASAP7_75t_R FILLER_0_263_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_888 ();
 DECAPx1_ASAP7_75t_R FILLER_0_263_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_899 ();
 DECAPx1_ASAP7_75t_R FILLER_0_263_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_911 ();
 FILLER_ASAP7_75t_R FILLER_0_263_923 ();
 DECAPx4_ASAP7_75t_R FILLER_0_263_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_937 ();
 FILLER_ASAP7_75t_R FILLER_0_263_948 ();
 FILLER_ASAP7_75t_R FILLER_0_263_956 ();
 DECAPx2_ASAP7_75t_R FILLER_0_263_964 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_970 ();
 DECAPx2_ASAP7_75t_R FILLER_0_263_981 ();
 FILLER_ASAP7_75t_R FILLER_0_263_987 ();
 DECAPx2_ASAP7_75t_R FILLER_0_263_992 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_998 ();
 FILLER_ASAP7_75t_R FILLER_0_263_1005 ();
 FILLER_ASAP7_75t_R FILLER_0_263_1013 ();
 DECAPx2_ASAP7_75t_R FILLER_0_263_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_1027 ();
 DECAPx1_ASAP7_75t_R FILLER_0_263_1035 ();
 FILLER_ASAP7_75t_R FILLER_0_263_1049 ();
 FILLER_ASAP7_75t_R FILLER_0_263_1057 ();
 FILLER_ASAP7_75t_R FILLER_0_263_1066 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_1068 ();
 FILLER_ASAP7_75t_R FILLER_0_263_1074 ();
 DECAPx2_ASAP7_75t_R FILLER_0_263_1086 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_1092 ();
 FILLER_ASAP7_75t_R FILLER_0_263_1099 ();
 DECAPx6_ASAP7_75t_R FILLER_0_263_1112 ();
 DECAPx1_ASAP7_75t_R FILLER_0_263_1126 ();
 FILLER_ASAP7_75t_R FILLER_0_263_1136 ();
 DECAPx2_ASAP7_75t_R FILLER_0_263_1144 ();
 DECAPx2_ASAP7_75t_R FILLER_0_263_1156 ();
 FILLER_ASAP7_75t_R FILLER_0_263_1168 ();
 DECAPx4_ASAP7_75t_R FILLER_0_263_1176 ();
 FILLER_ASAP7_75t_R FILLER_0_263_1192 ();
 DECAPx1_ASAP7_75t_R FILLER_0_263_1199 ();
 FILLER_ASAP7_75t_R FILLER_0_263_1213 ();
 DECAPx6_ASAP7_75t_R FILLER_0_263_1222 ();
 DECAPx1_ASAP7_75t_R FILLER_0_263_1236 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_1240 ();
 FILLER_ASAP7_75t_R FILLER_0_263_1244 ();
 DECAPx4_ASAP7_75t_R FILLER_0_263_1252 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_1262 ();
 DECAPx2_ASAP7_75t_R FILLER_0_263_1269 ();
 FILLER_ASAP7_75t_R FILLER_0_263_1275 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_1277 ();
 DECAPx1_ASAP7_75t_R FILLER_0_263_1286 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_1290 ();
 FILLER_ASAP7_75t_R FILLER_0_263_1297 ();
 DECAPx1_ASAP7_75t_R FILLER_0_263_1305 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_1309 ();
 DECAPx4_ASAP7_75t_R FILLER_0_263_1326 ();
 FILLER_ASAP7_75t_R FILLER_0_263_1336 ();
 FILLER_ASAP7_75t_R FILLER_0_263_1344 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_1346 ();
 FILLER_ASAP7_75t_R FILLER_0_263_1353 ();
 FILLER_ASAP7_75t_R FILLER_0_263_1361 ();
 FILLER_ASAP7_75t_R FILLER_0_263_1369 ();
 DECAPx1_ASAP7_75t_R FILLER_0_263_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_264_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_264_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_264_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_264_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_264_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_264_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_264_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_264_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_264_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_264_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_264_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_244 ();
 FILLER_ASAP7_75t_R FILLER_0_264_251 ();
 FILLER_ASAP7_75t_R FILLER_0_264_259 ();
 DECAPx2_ASAP7_75t_R FILLER_0_264_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_273 ();
 DECAPx6_ASAP7_75t_R FILLER_0_264_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_293 ();
 DECAPx4_ASAP7_75t_R FILLER_0_264_300 ();
 FILLER_ASAP7_75t_R FILLER_0_264_310 ();
 FILLER_ASAP7_75t_R FILLER_0_264_318 ();
 DECAPx2_ASAP7_75t_R FILLER_0_264_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_331 ();
 FILLER_ASAP7_75t_R FILLER_0_264_338 ();
 FILLER_ASAP7_75t_R FILLER_0_264_350 ();
 DECAPx1_ASAP7_75t_R FILLER_0_264_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_364 ();
 FILLER_ASAP7_75t_R FILLER_0_264_373 ();
 DECAPx1_ASAP7_75t_R FILLER_0_264_381 ();
 DECAPx1_ASAP7_75t_R FILLER_0_264_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_395 ();
 FILLER_ASAP7_75t_R FILLER_0_264_401 ();
 DECAPx2_ASAP7_75t_R FILLER_0_264_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_415 ();
 FILLER_ASAP7_75t_R FILLER_0_264_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_424 ();
 FILLER_ASAP7_75t_R FILLER_0_264_431 ();
 FILLER_ASAP7_75t_R FILLER_0_264_438 ();
 FILLER_ASAP7_75t_R FILLER_0_264_446 ();
 FILLER_ASAP7_75t_R FILLER_0_264_453 ();
 FILLER_ASAP7_75t_R FILLER_0_264_460 ();
 FILLER_ASAP7_75t_R FILLER_0_264_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_466 ();
 FILLER_ASAP7_75t_R FILLER_0_264_473 ();
 FILLER_ASAP7_75t_R FILLER_0_264_478 ();
 FILLER_ASAP7_75t_R FILLER_0_264_486 ();
 DECAPx1_ASAP7_75t_R FILLER_0_264_494 ();
 FILLER_ASAP7_75t_R FILLER_0_264_503 ();
 FILLER_ASAP7_75t_R FILLER_0_264_510 ();
 FILLER_ASAP7_75t_R FILLER_0_264_517 ();
 FILLER_ASAP7_75t_R FILLER_0_264_527 ();
 FILLER_ASAP7_75t_R FILLER_0_264_532 ();
 FILLER_ASAP7_75t_R FILLER_0_264_539 ();
 FILLER_ASAP7_75t_R FILLER_0_264_552 ();
 DECAPx1_ASAP7_75t_R FILLER_0_264_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_563 ();
 FILLER_ASAP7_75t_R FILLER_0_264_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_587 ();
 FILLER_ASAP7_75t_R FILLER_0_264_591 ();
 FILLER_ASAP7_75t_R FILLER_0_264_599 ();
 FILLER_ASAP7_75t_R FILLER_0_264_606 ();
 FILLER_ASAP7_75t_R FILLER_0_264_611 ();
 FILLER_ASAP7_75t_R FILLER_0_264_635 ();
 FILLER_ASAP7_75t_R FILLER_0_264_659 ();
 FILLER_ASAP7_75t_R FILLER_0_264_664 ();
 FILLER_ASAP7_75t_R FILLER_0_264_669 ();
 FILLER_ASAP7_75t_R FILLER_0_264_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_676 ();
 FILLER_ASAP7_75t_R FILLER_0_264_683 ();
 DECAPx4_ASAP7_75t_R FILLER_0_264_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_264_722 ();
 FILLER_ASAP7_75t_R FILLER_0_264_744 ();
 FILLER_ASAP7_75t_R FILLER_0_264_767 ();
 DECAPx10_ASAP7_75t_R FILLER_0_264_775 ();
 DECAPx6_ASAP7_75t_R FILLER_0_264_797 ();
 DECAPx4_ASAP7_75t_R FILLER_0_264_817 ();
 FILLER_ASAP7_75t_R FILLER_0_264_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_829 ();
 DECAPx6_ASAP7_75t_R FILLER_0_264_852 ();
 DECAPx1_ASAP7_75t_R FILLER_0_264_866 ();
 DECAPx2_ASAP7_75t_R FILLER_0_264_873 ();
 FILLER_ASAP7_75t_R FILLER_0_264_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_881 ();
 FILLER_ASAP7_75t_R FILLER_0_264_888 ();
 DECAPx2_ASAP7_75t_R FILLER_0_264_897 ();
 FILLER_ASAP7_75t_R FILLER_0_264_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_905 ();
 FILLER_ASAP7_75t_R FILLER_0_264_912 ();
 DECAPx2_ASAP7_75t_R FILLER_0_264_920 ();
 FILLER_ASAP7_75t_R FILLER_0_264_926 ();
 DECAPx4_ASAP7_75t_R FILLER_0_264_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_945 ();
 DECAPx6_ASAP7_75t_R FILLER_0_264_956 ();
 FILLER_ASAP7_75t_R FILLER_0_264_970 ();
 DECAPx1_ASAP7_75t_R FILLER_0_264_979 ();
 FILLER_ASAP7_75t_R FILLER_0_264_991 ();
 DECAPx1_ASAP7_75t_R FILLER_0_264_999 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_1003 ();
 FILLER_ASAP7_75t_R FILLER_0_264_1010 ();
 DECAPx2_ASAP7_75t_R FILLER_0_264_1018 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_1024 ();
 DECAPx2_ASAP7_75t_R FILLER_0_264_1037 ();
 FILLER_ASAP7_75t_R FILLER_0_264_1043 ();
 FILLER_ASAP7_75t_R FILLER_0_264_1052 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_1054 ();
 FILLER_ASAP7_75t_R FILLER_0_264_1061 ();
 FILLER_ASAP7_75t_R FILLER_0_264_1073 ();
 FILLER_ASAP7_75t_R FILLER_0_264_1081 ();
 FILLER_ASAP7_75t_R FILLER_0_264_1089 ();
 FILLER_ASAP7_75t_R FILLER_0_264_1097 ();
 FILLER_ASAP7_75t_R FILLER_0_264_1104 ();
 DECAPx6_ASAP7_75t_R FILLER_0_264_1112 ();
 DECAPx2_ASAP7_75t_R FILLER_0_264_1126 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_1132 ();
 FILLER_ASAP7_75t_R FILLER_0_264_1139 ();
 FILLER_ASAP7_75t_R FILLER_0_264_1147 ();
 DECAPx2_ASAP7_75t_R FILLER_0_264_1155 ();
 FILLER_ASAP7_75t_R FILLER_0_264_1167 ();
 DECAPx4_ASAP7_75t_R FILLER_0_264_1175 ();
 DECAPx2_ASAP7_75t_R FILLER_0_264_1191 ();
 FILLER_ASAP7_75t_R FILLER_0_264_1197 ();
 DECAPx2_ASAP7_75t_R FILLER_0_264_1205 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_1211 ();
 DECAPx6_ASAP7_75t_R FILLER_0_264_1218 ();
 DECAPx1_ASAP7_75t_R FILLER_0_264_1232 ();
 DECAPx2_ASAP7_75t_R FILLER_0_264_1256 ();
 FILLER_ASAP7_75t_R FILLER_0_264_1262 ();
 DECAPx2_ASAP7_75t_R FILLER_0_264_1267 ();
 FILLER_ASAP7_75t_R FILLER_0_264_1273 ();
 FILLER_ASAP7_75t_R FILLER_0_264_1280 ();
 DECAPx2_ASAP7_75t_R FILLER_0_264_1292 ();
 FILLER_ASAP7_75t_R FILLER_0_264_1305 ();
 DECAPx6_ASAP7_75t_R FILLER_0_264_1313 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_1327 ();
 DECAPx4_ASAP7_75t_R FILLER_0_264_1335 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_1345 ();
 DECAPx10_ASAP7_75t_R FILLER_0_264_1351 ();
 DECAPx2_ASAP7_75t_R FILLER_0_264_1373 ();
 FILLER_ASAP7_75t_R FILLER_0_264_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_265_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_265_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_265_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_265_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_265_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_265_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_265_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_265_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_265_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_265_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_265_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_265_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_265_266 ();
 DECAPx1_ASAP7_75t_R FILLER_0_265_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_292 ();
 DECAPx6_ASAP7_75t_R FILLER_0_265_299 ();
 FILLER_ASAP7_75t_R FILLER_0_265_313 ();
 DECAPx1_ASAP7_75t_R FILLER_0_265_322 ();
 DECAPx6_ASAP7_75t_R FILLER_0_265_332 ();
 FILLER_ASAP7_75t_R FILLER_0_265_366 ();
 DECAPx1_ASAP7_75t_R FILLER_0_265_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_380 ();
 DECAPx1_ASAP7_75t_R FILLER_0_265_392 ();
 FILLER_ASAP7_75t_R FILLER_0_265_402 ();
 DECAPx2_ASAP7_75t_R FILLER_0_265_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_418 ();
 DECAPx2_ASAP7_75t_R FILLER_0_265_425 ();
 FILLER_ASAP7_75t_R FILLER_0_265_431 ();
 FILLER_ASAP7_75t_R FILLER_0_265_439 ();
 FILLER_ASAP7_75t_R FILLER_0_265_452 ();
 FILLER_ASAP7_75t_R FILLER_0_265_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_462 ();
 FILLER_ASAP7_75t_R FILLER_0_265_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_476 ();
 FILLER_ASAP7_75t_R FILLER_0_265_480 ();
 FILLER_ASAP7_75t_R FILLER_0_265_488 ();
 FILLER_ASAP7_75t_R FILLER_0_265_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_503 ();
 FILLER_ASAP7_75t_R FILLER_0_265_509 ();
 FILLER_ASAP7_75t_R FILLER_0_265_516 ();
 FILLER_ASAP7_75t_R FILLER_0_265_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_528 ();
 FILLER_ASAP7_75t_R FILLER_0_265_534 ();
 FILLER_ASAP7_75t_R FILLER_0_265_541 ();
 FILLER_ASAP7_75t_R FILLER_0_265_548 ();
 FILLER_ASAP7_75t_R FILLER_0_265_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_564 ();
 FILLER_ASAP7_75t_R FILLER_0_265_570 ();
 FILLER_ASAP7_75t_R FILLER_0_265_577 ();
 FILLER_ASAP7_75t_R FILLER_0_265_584 ();
 DECAPx1_ASAP7_75t_R FILLER_0_265_591 ();
 FILLER_ASAP7_75t_R FILLER_0_265_601 ();
 FILLER_ASAP7_75t_R FILLER_0_265_625 ();
 DECAPx1_ASAP7_75t_R FILLER_0_265_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_636 ();
 FILLER_ASAP7_75t_R FILLER_0_265_658 ();
 FILLER_ASAP7_75t_R FILLER_0_265_666 ();
 FILLER_ASAP7_75t_R FILLER_0_265_671 ();
 FILLER_ASAP7_75t_R FILLER_0_265_676 ();
 FILLER_ASAP7_75t_R FILLER_0_265_683 ();
 FILLER_ASAP7_75t_R FILLER_0_265_691 ();
 FILLER_ASAP7_75t_R FILLER_0_265_699 ();
 DECAPx2_ASAP7_75t_R FILLER_0_265_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_728 ();
 FILLER_ASAP7_75t_R FILLER_0_265_751 ();
 DECAPx6_ASAP7_75t_R FILLER_0_265_756 ();
 FILLER_ASAP7_75t_R FILLER_0_265_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_772 ();
 DECAPx1_ASAP7_75t_R FILLER_0_265_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_783 ();
 FILLER_ASAP7_75t_R FILLER_0_265_790 ();
 DECAPx1_ASAP7_75t_R FILLER_0_265_813 ();
 FILLER_ASAP7_75t_R FILLER_0_265_823 ();
 FILLER_ASAP7_75t_R FILLER_0_265_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_832 ();
 FILLER_ASAP7_75t_R FILLER_0_265_853 ();
 FILLER_ASAP7_75t_R FILLER_0_265_868 ();
 DECAPx4_ASAP7_75t_R FILLER_0_265_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_883 ();
 FILLER_ASAP7_75t_R FILLER_0_265_890 ();
 FILLER_ASAP7_75t_R FILLER_0_265_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_900 ();
 DECAPx2_ASAP7_75t_R FILLER_0_265_907 ();
 FILLER_ASAP7_75t_R FILLER_0_265_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_915 ();
 FILLER_ASAP7_75t_R FILLER_0_265_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_924 ();
 FILLER_ASAP7_75t_R FILLER_0_265_927 ();
 DECAPx2_ASAP7_75t_R FILLER_0_265_935 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_941 ();
 DECAPx1_ASAP7_75t_R FILLER_0_265_962 ();
 DECAPx1_ASAP7_75t_R FILLER_0_265_972 ();
 DECAPx1_ASAP7_75t_R FILLER_0_265_987 ();
 DECAPx1_ASAP7_75t_R FILLER_0_265_1002 ();
 DECAPx4_ASAP7_75t_R FILLER_0_265_1016 ();
 FILLER_ASAP7_75t_R FILLER_0_265_1026 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_1028 ();
 DECAPx4_ASAP7_75t_R FILLER_0_265_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_1045 ();
 DECAPx6_ASAP7_75t_R FILLER_0_265_1051 ();
 DECAPx2_ASAP7_75t_R FILLER_0_265_1071 ();
 FILLER_ASAP7_75t_R FILLER_0_265_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_1085 ();
 FILLER_ASAP7_75t_R FILLER_0_265_1092 ();
 DECAPx1_ASAP7_75t_R FILLER_0_265_1100 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_1104 ();
 DECAPx6_ASAP7_75t_R FILLER_0_265_1115 ();
 FILLER_ASAP7_75t_R FILLER_0_265_1132 ();
 DECAPx10_ASAP7_75t_R FILLER_0_265_1145 ();
 DECAPx4_ASAP7_75t_R FILLER_0_265_1167 ();
 FILLER_ASAP7_75t_R FILLER_0_265_1177 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_1179 ();
 FILLER_ASAP7_75t_R FILLER_0_265_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_265_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_0_265_1203 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_1225 ();
 FILLER_ASAP7_75t_R FILLER_0_265_1236 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_1238 ();
 FILLER_ASAP7_75t_R FILLER_0_265_1245 ();
 DECAPx2_ASAP7_75t_R FILLER_0_265_1253 ();
 FILLER_ASAP7_75t_R FILLER_0_265_1279 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_1281 ();
 FILLER_ASAP7_75t_R FILLER_0_265_1288 ();
 FILLER_ASAP7_75t_R FILLER_0_265_1295 ();
 DECAPx2_ASAP7_75t_R FILLER_0_265_1317 ();
 FILLER_ASAP7_75t_R FILLER_0_265_1326 ();
 DECAPx2_ASAP7_75t_R FILLER_0_265_1334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_265_1346 ();
 DECAPx6_ASAP7_75t_R FILLER_0_265_1368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_266_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_266_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_266_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_266_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_266_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_266_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_266_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_266_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_266_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_266_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_266_222 ();
 DECAPx4_ASAP7_75t_R FILLER_0_266_244 ();
 DECAPx1_ASAP7_75t_R FILLER_0_266_260 ();
 FILLER_ASAP7_75t_R FILLER_0_266_269 ();
 FILLER_ASAP7_75t_R FILLER_0_266_277 ();
 DECAPx2_ASAP7_75t_R FILLER_0_266_285 ();
 DECAPx1_ASAP7_75t_R FILLER_0_266_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_305 ();
 FILLER_ASAP7_75t_R FILLER_0_266_312 ();
 DECAPx2_ASAP7_75t_R FILLER_0_266_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_326 ();
 FILLER_ASAP7_75t_R FILLER_0_266_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_336 ();
 DECAPx1_ASAP7_75t_R FILLER_0_266_343 ();
 FILLER_ASAP7_75t_R FILLER_0_266_353 ();
 FILLER_ASAP7_75t_R FILLER_0_266_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_377 ();
 FILLER_ASAP7_75t_R FILLER_0_266_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_386 ();
 FILLER_ASAP7_75t_R FILLER_0_266_393 ();
 DECAPx2_ASAP7_75t_R FILLER_0_266_405 ();
 FILLER_ASAP7_75t_R FILLER_0_266_411 ();
 DECAPx1_ASAP7_75t_R FILLER_0_266_419 ();
 FILLER_ASAP7_75t_R FILLER_0_266_428 ();
 FILLER_ASAP7_75t_R FILLER_0_266_435 ();
 FILLER_ASAP7_75t_R FILLER_0_266_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_445 ();
 FILLER_ASAP7_75t_R FILLER_0_266_451 ();
 FILLER_ASAP7_75t_R FILLER_0_266_460 ();
 FILLER_ASAP7_75t_R FILLER_0_266_464 ();
 FILLER_ASAP7_75t_R FILLER_0_266_482 ();
 FILLER_ASAP7_75t_R FILLER_0_266_490 ();
 FILLER_ASAP7_75t_R FILLER_0_266_498 ();
 FILLER_ASAP7_75t_R FILLER_0_266_510 ();
 FILLER_ASAP7_75t_R FILLER_0_266_515 ();
 FILLER_ASAP7_75t_R FILLER_0_266_539 ();
 DECAPx1_ASAP7_75t_R FILLER_0_266_553 ();
 FILLER_ASAP7_75t_R FILLER_0_266_563 ();
 FILLER_ASAP7_75t_R FILLER_0_266_570 ();
 FILLER_ASAP7_75t_R FILLER_0_266_577 ();
 FILLER_ASAP7_75t_R FILLER_0_266_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_587 ();
 FILLER_ASAP7_75t_R FILLER_0_266_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_596 ();
 FILLER_ASAP7_75t_R FILLER_0_266_600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_266_624 ();
 FILLER_ASAP7_75t_R FILLER_0_266_652 ();
 FILLER_ASAP7_75t_R FILLER_0_266_660 ();
 FILLER_ASAP7_75t_R FILLER_0_266_667 ();
 FILLER_ASAP7_75t_R FILLER_0_266_672 ();
 FILLER_ASAP7_75t_R FILLER_0_266_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_679 ();
 DECAPx1_ASAP7_75t_R FILLER_0_266_686 ();
 DECAPx2_ASAP7_75t_R FILLER_0_266_695 ();
 FILLER_ASAP7_75t_R FILLER_0_266_707 ();
 DECAPx1_ASAP7_75t_R FILLER_0_266_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_718 ();
 DECAPx4_ASAP7_75t_R FILLER_0_266_741 ();
 DECAPx4_ASAP7_75t_R FILLER_0_266_754 ();
 FILLER_ASAP7_75t_R FILLER_0_266_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_766 ();
 FILLER_ASAP7_75t_R FILLER_0_266_788 ();
 DECAPx1_ASAP7_75t_R FILLER_0_266_795 ();
 FILLER_ASAP7_75t_R FILLER_0_266_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_807 ();
 FILLER_ASAP7_75t_R FILLER_0_266_811 ();
 FILLER_ASAP7_75t_R FILLER_0_266_834 ();
 FILLER_ASAP7_75t_R FILLER_0_266_839 ();
 FILLER_ASAP7_75t_R FILLER_0_266_844 ();
 FILLER_ASAP7_75t_R FILLER_0_266_849 ();
 FILLER_ASAP7_75t_R FILLER_0_266_854 ();
 DECAPx1_ASAP7_75t_R FILLER_0_266_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_863 ();
 FILLER_ASAP7_75t_R FILLER_0_266_872 ();
 FILLER_ASAP7_75t_R FILLER_0_266_880 ();
 DECAPx2_ASAP7_75t_R FILLER_0_266_888 ();
 FILLER_ASAP7_75t_R FILLER_0_266_894 ();
 FILLER_ASAP7_75t_R FILLER_0_266_902 ();
 DECAPx1_ASAP7_75t_R FILLER_0_266_910 ();
 DECAPx2_ASAP7_75t_R FILLER_0_266_925 ();
 FILLER_ASAP7_75t_R FILLER_0_266_931 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_933 ();
 FILLER_ASAP7_75t_R FILLER_0_266_940 ();
 FILLER_ASAP7_75t_R FILLER_0_266_948 ();
 DECAPx2_ASAP7_75t_R FILLER_0_266_956 ();
 FILLER_ASAP7_75t_R FILLER_0_266_962 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_964 ();
 DECAPx2_ASAP7_75t_R FILLER_0_266_970 ();
 DECAPx1_ASAP7_75t_R FILLER_0_266_981 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_985 ();
 FILLER_ASAP7_75t_R FILLER_0_266_992 ();
 DECAPx1_ASAP7_75t_R FILLER_0_266_1004 ();
 FILLER_ASAP7_75t_R FILLER_0_266_1014 ();
 DECAPx1_ASAP7_75t_R FILLER_0_266_1021 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_1025 ();
 FILLER_ASAP7_75t_R FILLER_0_266_1032 ();
 DECAPx10_ASAP7_75t_R FILLER_0_266_1040 ();
 DECAPx2_ASAP7_75t_R FILLER_0_266_1062 ();
 FILLER_ASAP7_75t_R FILLER_0_266_1068 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_1070 ();
 FILLER_ASAP7_75t_R FILLER_0_266_1077 ();
 DECAPx6_ASAP7_75t_R FILLER_0_266_1083 ();
 DECAPx1_ASAP7_75t_R FILLER_0_266_1097 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_1101 ();
 DECAPx10_ASAP7_75t_R FILLER_0_266_1108 ();
 DECAPx2_ASAP7_75t_R FILLER_0_266_1130 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_1136 ();
 DECAPx2_ASAP7_75t_R FILLER_0_266_1143 ();
 DECAPx4_ASAP7_75t_R FILLER_0_266_1152 ();
 FILLER_ASAP7_75t_R FILLER_0_266_1172 ();
 FILLER_ASAP7_75t_R FILLER_0_266_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_1182 ();
 DECAPx2_ASAP7_75t_R FILLER_0_266_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_1195 ();
 DECAPx6_ASAP7_75t_R FILLER_0_266_1202 ();
 DECAPx2_ASAP7_75t_R FILLER_0_266_1219 ();
 FILLER_ASAP7_75t_R FILLER_0_266_1225 ();
 DECAPx4_ASAP7_75t_R FILLER_0_266_1233 ();
 FILLER_ASAP7_75t_R FILLER_0_266_1243 ();
 FILLER_ASAP7_75t_R FILLER_0_266_1255 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_1257 ();
 FILLER_ASAP7_75t_R FILLER_0_266_1264 ();
 DECAPx2_ASAP7_75t_R FILLER_0_266_1272 ();
 DECAPx1_ASAP7_75t_R FILLER_0_266_1284 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_1288 ();
 DECAPx2_ASAP7_75t_R FILLER_0_266_1295 ();
 FILLER_ASAP7_75t_R FILLER_0_266_1301 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_1303 ();
 DECAPx1_ASAP7_75t_R FILLER_0_266_1314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_266_1324 ();
 DECAPx1_ASAP7_75t_R FILLER_0_266_1346 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_1350 ();
 DECAPx10_ASAP7_75t_R FILLER_0_266_1357 ();
 FILLER_ASAP7_75t_R FILLER_0_266_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_267_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_267_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_267_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_267_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_267_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_267_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_267_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_267_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_267_178 ();
 DECAPx1_ASAP7_75t_R FILLER_0_267_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_204 ();
 FILLER_ASAP7_75t_R FILLER_0_267_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_228 ();
 DECAPx2_ASAP7_75t_R FILLER_0_267_250 ();
 FILLER_ASAP7_75t_R FILLER_0_267_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_258 ();
 DECAPx2_ASAP7_75t_R FILLER_0_267_265 ();
 FILLER_ASAP7_75t_R FILLER_0_267_271 ();
 FILLER_ASAP7_75t_R FILLER_0_267_279 ();
 FILLER_ASAP7_75t_R FILLER_0_267_287 ();
 FILLER_ASAP7_75t_R FILLER_0_267_295 ();
 DECAPx2_ASAP7_75t_R FILLER_0_267_302 ();
 FILLER_ASAP7_75t_R FILLER_0_267_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_310 ();
 DECAPx4_ASAP7_75t_R FILLER_0_267_317 ();
 FILLER_ASAP7_75t_R FILLER_0_267_333 ();
 DECAPx6_ASAP7_75t_R FILLER_0_267_340 ();
 DECAPx1_ASAP7_75t_R FILLER_0_267_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_358 ();
 DECAPx6_ASAP7_75t_R FILLER_0_267_367 ();
 DECAPx2_ASAP7_75t_R FILLER_0_267_381 ();
 DECAPx1_ASAP7_75t_R FILLER_0_267_407 ();
 FILLER_ASAP7_75t_R FILLER_0_267_416 ();
 FILLER_ASAP7_75t_R FILLER_0_267_424 ();
 FILLER_ASAP7_75t_R FILLER_0_267_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_438 ();
 FILLER_ASAP7_75t_R FILLER_0_267_445 ();
 FILLER_ASAP7_75t_R FILLER_0_267_450 ();
 FILLER_ASAP7_75t_R FILLER_0_267_457 ();
 FILLER_ASAP7_75t_R FILLER_0_267_464 ();
 FILLER_ASAP7_75t_R FILLER_0_267_471 ();
 FILLER_ASAP7_75t_R FILLER_0_267_478 ();
 FILLER_ASAP7_75t_R FILLER_0_267_485 ();
 FILLER_ASAP7_75t_R FILLER_0_267_492 ();
 FILLER_ASAP7_75t_R FILLER_0_267_499 ();
 FILLER_ASAP7_75t_R FILLER_0_267_506 ();
 FILLER_ASAP7_75t_R FILLER_0_267_513 ();
 FILLER_ASAP7_75t_R FILLER_0_267_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_523 ();
 FILLER_ASAP7_75t_R FILLER_0_267_527 ();
 FILLER_ASAP7_75t_R FILLER_0_267_534 ();
 FILLER_ASAP7_75t_R FILLER_0_267_541 ();
 FILLER_ASAP7_75t_R FILLER_0_267_548 ();
 FILLER_ASAP7_75t_R FILLER_0_267_571 ();
 FILLER_ASAP7_75t_R FILLER_0_267_576 ();
 FILLER_ASAP7_75t_R FILLER_0_267_599 ();
 FILLER_ASAP7_75t_R FILLER_0_267_606 ();
 DECAPx1_ASAP7_75t_R FILLER_0_267_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_619 ();
 FILLER_ASAP7_75t_R FILLER_0_267_625 ();
 FILLER_ASAP7_75t_R FILLER_0_267_632 ();
 DECAPx1_ASAP7_75t_R FILLER_0_267_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_643 ();
 FILLER_ASAP7_75t_R FILLER_0_267_649 ();
 DECAPx1_ASAP7_75t_R FILLER_0_267_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_660 ();
 FILLER_ASAP7_75t_R FILLER_0_267_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_668 ();
 FILLER_ASAP7_75t_R FILLER_0_267_691 ();
 DECAPx2_ASAP7_75t_R FILLER_0_267_696 ();
 FILLER_ASAP7_75t_R FILLER_0_267_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_704 ();
 FILLER_ASAP7_75t_R FILLER_0_267_708 ();
 FILLER_ASAP7_75t_R FILLER_0_267_731 ();
 FILLER_ASAP7_75t_R FILLER_0_267_736 ();
 FILLER_ASAP7_75t_R FILLER_0_267_741 ();
 DECAPx6_ASAP7_75t_R FILLER_0_267_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_760 ();
 DECAPx2_ASAP7_75t_R FILLER_0_267_783 ();
 FILLER_ASAP7_75t_R FILLER_0_267_792 ();
 FILLER_ASAP7_75t_R FILLER_0_267_797 ();
 FILLER_ASAP7_75t_R FILLER_0_267_805 ();
 FILLER_ASAP7_75t_R FILLER_0_267_812 ();
 FILLER_ASAP7_75t_R FILLER_0_267_817 ();
 FILLER_ASAP7_75t_R FILLER_0_267_825 ();
 FILLER_ASAP7_75t_R FILLER_0_267_830 ();
 DECAPx2_ASAP7_75t_R FILLER_0_267_835 ();
 FILLER_ASAP7_75t_R FILLER_0_267_847 ();
 FILLER_ASAP7_75t_R FILLER_0_267_852 ();
 FILLER_ASAP7_75t_R FILLER_0_267_857 ();
 DECAPx1_ASAP7_75t_R FILLER_0_267_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_870 ();
 FILLER_ASAP7_75t_R FILLER_0_267_879 ();
 FILLER_ASAP7_75t_R FILLER_0_267_887 ();
 DECAPx4_ASAP7_75t_R FILLER_0_267_895 ();
 DECAPx6_ASAP7_75t_R FILLER_0_267_911 ();
 FILLER_ASAP7_75t_R FILLER_0_267_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_929 ();
 DECAPx10_ASAP7_75t_R FILLER_0_267_936 ();
 DECAPx4_ASAP7_75t_R FILLER_0_267_958 ();
 FILLER_ASAP7_75t_R FILLER_0_267_968 ();
 FILLER_ASAP7_75t_R FILLER_0_267_980 ();
 FILLER_ASAP7_75t_R FILLER_0_267_985 ();
 FILLER_ASAP7_75t_R FILLER_0_267_993 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_995 ();
 FILLER_ASAP7_75t_R FILLER_0_267_1002 ();
 DECAPx2_ASAP7_75t_R FILLER_0_267_1011 ();
 DECAPx10_ASAP7_75t_R FILLER_0_267_1029 ();
 FILLER_ASAP7_75t_R FILLER_0_267_1051 ();
 FILLER_ASAP7_75t_R FILLER_0_267_1065 ();
 DECAPx2_ASAP7_75t_R FILLER_0_267_1077 ();
 FILLER_ASAP7_75t_R FILLER_0_267_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_1085 ();
 FILLER_ASAP7_75t_R FILLER_0_267_1098 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_1100 ();
 DECAPx10_ASAP7_75t_R FILLER_0_267_1107 ();
 DECAPx4_ASAP7_75t_R FILLER_0_267_1129 ();
 FILLER_ASAP7_75t_R FILLER_0_267_1139 ();
 FILLER_ASAP7_75t_R FILLER_0_267_1144 ();
 DECAPx2_ASAP7_75t_R FILLER_0_267_1152 ();
 FILLER_ASAP7_75t_R FILLER_0_267_1158 ();
 DECAPx2_ASAP7_75t_R FILLER_0_267_1163 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_1169 ();
 FILLER_ASAP7_75t_R FILLER_0_267_1176 ();
 DECAPx1_ASAP7_75t_R FILLER_0_267_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_1185 ();
 DECAPx4_ASAP7_75t_R FILLER_0_267_1192 ();
 FILLER_ASAP7_75t_R FILLER_0_267_1208 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_1210 ();
 DECAPx1_ASAP7_75t_R FILLER_0_267_1217 ();
 DECAPx6_ASAP7_75t_R FILLER_0_267_1232 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_1246 ();
 DECAPx4_ASAP7_75t_R FILLER_0_267_1250 ();
 FILLER_ASAP7_75t_R FILLER_0_267_1260 ();
 FILLER_ASAP7_75t_R FILLER_0_267_1268 ();
 DECAPx1_ASAP7_75t_R FILLER_0_267_1276 ();
 FILLER_ASAP7_75t_R FILLER_0_267_1286 ();
 DECAPx1_ASAP7_75t_R FILLER_0_267_1294 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_1298 ();
 FILLER_ASAP7_75t_R FILLER_0_267_1305 ();
 FILLER_ASAP7_75t_R FILLER_0_267_1313 ();
 DECAPx2_ASAP7_75t_R FILLER_0_267_1321 ();
 FILLER_ASAP7_75t_R FILLER_0_267_1327 ();
 DECAPx2_ASAP7_75t_R FILLER_0_267_1335 ();
 FILLER_ASAP7_75t_R FILLER_0_267_1341 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_1343 ();
 FILLER_ASAP7_75t_R FILLER_0_267_1350 ();
 DECAPx10_ASAP7_75t_R FILLER_0_267_1360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_268_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_268_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_268_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_268_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_268_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_268_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_268_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_268_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_268_178 ();
 DECAPx2_ASAP7_75t_R FILLER_0_268_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_206 ();
 FILLER_ASAP7_75t_R FILLER_0_268_210 ();
 FILLER_ASAP7_75t_R FILLER_0_268_224 ();
 DECAPx1_ASAP7_75t_R FILLER_0_268_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_236 ();
 FILLER_ASAP7_75t_R FILLER_0_268_246 ();
 DECAPx1_ASAP7_75t_R FILLER_0_268_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_255 ();
 DECAPx10_ASAP7_75t_R FILLER_0_268_262 ();
 DECAPx10_ASAP7_75t_R FILLER_0_268_284 ();
 DECAPx4_ASAP7_75t_R FILLER_0_268_306 ();
 FILLER_ASAP7_75t_R FILLER_0_268_316 ();
 DECAPx4_ASAP7_75t_R FILLER_0_268_324 ();
 FILLER_ASAP7_75t_R FILLER_0_268_340 ();
 DECAPx4_ASAP7_75t_R FILLER_0_268_347 ();
 FILLER_ASAP7_75t_R FILLER_0_268_357 ();
 DECAPx1_ASAP7_75t_R FILLER_0_268_365 ();
 FILLER_ASAP7_75t_R FILLER_0_268_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_377 ();
 FILLER_ASAP7_75t_R FILLER_0_268_384 ();
 FILLER_ASAP7_75t_R FILLER_0_268_393 ();
 FILLER_ASAP7_75t_R FILLER_0_268_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_403 ();
 FILLER_ASAP7_75t_R FILLER_0_268_412 ();
 FILLER_ASAP7_75t_R FILLER_0_268_417 ();
 FILLER_ASAP7_75t_R FILLER_0_268_424 ();
 FILLER_ASAP7_75t_R FILLER_0_268_431 ();
 FILLER_ASAP7_75t_R FILLER_0_268_453 ();
 FILLER_ASAP7_75t_R FILLER_0_268_460 ();
 DECAPx1_ASAP7_75t_R FILLER_0_268_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_468 ();
 FILLER_ASAP7_75t_R FILLER_0_268_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_477 ();
 FILLER_ASAP7_75t_R FILLER_0_268_481 ();
 FILLER_ASAP7_75t_R FILLER_0_268_488 ();
 FILLER_ASAP7_75t_R FILLER_0_268_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_502 ();
 FILLER_ASAP7_75t_R FILLER_0_268_506 ();
 FILLER_ASAP7_75t_R FILLER_0_268_513 ();
 FILLER_ASAP7_75t_R FILLER_0_268_520 ();
 FILLER_ASAP7_75t_R FILLER_0_268_527 ();
 FILLER_ASAP7_75t_R FILLER_0_268_534 ();
 FILLER_ASAP7_75t_R FILLER_0_268_541 ();
 FILLER_ASAP7_75t_R FILLER_0_268_548 ();
 FILLER_ASAP7_75t_R FILLER_0_268_556 ();
 FILLER_ASAP7_75t_R FILLER_0_268_563 ();
 FILLER_ASAP7_75t_R FILLER_0_268_570 ();
 FILLER_ASAP7_75t_R FILLER_0_268_577 ();
 FILLER_ASAP7_75t_R FILLER_0_268_584 ();
 DECAPx1_ASAP7_75t_R FILLER_0_268_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_596 ();
 FILLER_ASAP7_75t_R FILLER_0_268_602 ();
 FILLER_ASAP7_75t_R FILLER_0_268_609 ();
 FILLER_ASAP7_75t_R FILLER_0_268_621 ();
 FILLER_ASAP7_75t_R FILLER_0_268_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_630 ();
 FILLER_ASAP7_75t_R FILLER_0_268_637 ();
 DECAPx1_ASAP7_75t_R FILLER_0_268_649 ();
 FILLER_ASAP7_75t_R FILLER_0_268_658 ();
 FILLER_ASAP7_75t_R FILLER_0_268_682 ();
 FILLER_ASAP7_75t_R FILLER_0_268_687 ();
 FILLER_ASAP7_75t_R FILLER_0_268_692 ();
 FILLER_ASAP7_75t_R FILLER_0_268_697 ();
 FILLER_ASAP7_75t_R FILLER_0_268_702 ();
 DECAPx1_ASAP7_75t_R FILLER_0_268_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_711 ();
 DECAPx2_ASAP7_75t_R FILLER_0_268_715 ();
 FILLER_ASAP7_75t_R FILLER_0_268_724 ();
 DECAPx2_ASAP7_75t_R FILLER_0_268_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_753 ();
 FILLER_ASAP7_75t_R FILLER_0_268_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_762 ();
 FILLER_ASAP7_75t_R FILLER_0_268_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_768 ();
 DECAPx2_ASAP7_75t_R FILLER_0_268_772 ();
 FILLER_ASAP7_75t_R FILLER_0_268_778 ();
 DECAPx1_ASAP7_75t_R FILLER_0_268_783 ();
 DECAPx2_ASAP7_75t_R FILLER_0_268_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_796 ();
 FILLER_ASAP7_75t_R FILLER_0_268_800 ();
 DECAPx2_ASAP7_75t_R FILLER_0_268_807 ();
 DECAPx2_ASAP7_75t_R FILLER_0_268_833 ();
 FILLER_ASAP7_75t_R FILLER_0_268_844 ();
 DECAPx1_ASAP7_75t_R FILLER_0_268_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_855 ();
 FILLER_ASAP7_75t_R FILLER_0_268_886 ();
 FILLER_ASAP7_75t_R FILLER_0_268_894 ();
 FILLER_ASAP7_75t_R FILLER_0_268_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_901 ();
 FILLER_ASAP7_75t_R FILLER_0_268_908 ();
 DECAPx1_ASAP7_75t_R FILLER_0_268_916 ();
 FILLER_ASAP7_75t_R FILLER_0_268_926 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_928 ();
 DECAPx2_ASAP7_75t_R FILLER_0_268_935 ();
 FILLER_ASAP7_75t_R FILLER_0_268_941 ();
 FILLER_ASAP7_75t_R FILLER_0_268_949 ();
 DECAPx1_ASAP7_75t_R FILLER_0_268_961 ();
 DECAPx6_ASAP7_75t_R FILLER_0_268_971 ();
 DECAPx1_ASAP7_75t_R FILLER_0_268_985 ();
 FILLER_ASAP7_75t_R FILLER_0_268_995 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1002 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1014 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_1021 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1028 ();
 DECAPx1_ASAP7_75t_R FILLER_0_268_1035 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_1039 ();
 DECAPx4_ASAP7_75t_R FILLER_0_268_1046 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1056 ();
 DECAPx4_ASAP7_75t_R FILLER_0_268_1070 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1080 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1087 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1097 ();
 DECAPx10_ASAP7_75t_R FILLER_0_268_1107 ();
 DECAPx2_ASAP7_75t_R FILLER_0_268_1129 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_1135 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1144 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_1146 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1153 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_1155 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1163 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_1173 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1180 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1188 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1196 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1204 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1212 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1222 ();
 DECAPx1_ASAP7_75t_R FILLER_0_268_1230 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_1234 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_0_268_1249 ();
 DECAPx1_ASAP7_75t_R FILLER_0_268_1271 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_1275 ();
 DECAPx2_ASAP7_75t_R FILLER_0_268_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_1288 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1295 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_1297 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1304 ();
 DECAPx4_ASAP7_75t_R FILLER_0_268_1312 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1322 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_1324 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1331 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1339 ();
 FILLER_ASAP7_75t_R FILLER_0_268_1347 ();
 DECAPx10_ASAP7_75t_R FILLER_0_268_1355 ();
 DECAPx1_ASAP7_75t_R FILLER_0_268_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_269_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_269_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_269_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_269_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_269_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_269_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_269_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_269_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_269_178 ();
 DECAPx4_ASAP7_75t_R FILLER_0_269_200 ();
 FILLER_ASAP7_75t_R FILLER_0_269_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_212 ();
 FILLER_ASAP7_75t_R FILLER_0_269_221 ();
 DECAPx1_ASAP7_75t_R FILLER_0_269_229 ();
 DECAPx2_ASAP7_75t_R FILLER_0_269_240 ();
 FILLER_ASAP7_75t_R FILLER_0_269_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_248 ();
 FILLER_ASAP7_75t_R FILLER_0_269_255 ();
 FILLER_ASAP7_75t_R FILLER_0_269_263 ();
 DECAPx4_ASAP7_75t_R FILLER_0_269_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_281 ();
 DECAPx1_ASAP7_75t_R FILLER_0_269_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_292 ();
 DECAPx2_ASAP7_75t_R FILLER_0_269_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_310 ();
 DECAPx1_ASAP7_75t_R FILLER_0_269_317 ();
 DECAPx2_ASAP7_75t_R FILLER_0_269_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_337 ();
 FILLER_ASAP7_75t_R FILLER_0_269_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_346 ();
 FILLER_ASAP7_75t_R FILLER_0_269_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_359 ();
 DECAPx2_ASAP7_75t_R FILLER_0_269_366 ();
 FILLER_ASAP7_75t_R FILLER_0_269_372 ();
 FILLER_ASAP7_75t_R FILLER_0_269_379 ();
 FILLER_ASAP7_75t_R FILLER_0_269_386 ();
 DECAPx1_ASAP7_75t_R FILLER_0_269_394 ();
 FILLER_ASAP7_75t_R FILLER_0_269_404 ();
 DECAPx2_ASAP7_75t_R FILLER_0_269_412 ();
 FILLER_ASAP7_75t_R FILLER_0_269_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_430 ();
 FILLER_ASAP7_75t_R FILLER_0_269_434 ();
 FILLER_ASAP7_75t_R FILLER_0_269_442 ();
 FILLER_ASAP7_75t_R FILLER_0_269_450 ();
 FILLER_ASAP7_75t_R FILLER_0_269_455 ();
 DECAPx1_ASAP7_75t_R FILLER_0_269_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_467 ();
 DECAPx1_ASAP7_75t_R FILLER_0_269_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_478 ();
 FILLER_ASAP7_75t_R FILLER_0_269_485 ();
 FILLER_ASAP7_75t_R FILLER_0_269_493 ();
 FILLER_ASAP7_75t_R FILLER_0_269_498 ();
 FILLER_ASAP7_75t_R FILLER_0_269_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_523 ();
 FILLER_ASAP7_75t_R FILLER_0_269_545 ();
 FILLER_ASAP7_75t_R FILLER_0_269_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_555 ();
 DECAPx1_ASAP7_75t_R FILLER_0_269_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_566 ();
 FILLER_ASAP7_75t_R FILLER_0_269_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_575 ();
 FILLER_ASAP7_75t_R FILLER_0_269_579 ();
 FILLER_ASAP7_75t_R FILLER_0_269_586 ();
 DECAPx1_ASAP7_75t_R FILLER_0_269_594 ();
 FILLER_ASAP7_75t_R FILLER_0_269_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_621 ();
 FILLER_ASAP7_75t_R FILLER_0_269_625 ();
 FILLER_ASAP7_75t_R FILLER_0_269_632 ();
 FILLER_ASAP7_75t_R FILLER_0_269_639 ();
 FILLER_ASAP7_75t_R FILLER_0_269_646 ();
 FILLER_ASAP7_75t_R FILLER_0_269_651 ();
 FILLER_ASAP7_75t_R FILLER_0_269_658 ();
 FILLER_ASAP7_75t_R FILLER_0_269_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_667 ();
 FILLER_ASAP7_75t_R FILLER_0_269_671 ();
 FILLER_ASAP7_75t_R FILLER_0_269_679 ();
 FILLER_ASAP7_75t_R FILLER_0_269_686 ();
 DECAPx1_ASAP7_75t_R FILLER_0_269_710 ();
 FILLER_ASAP7_75t_R FILLER_0_269_720 ();
 DECAPx2_ASAP7_75t_R FILLER_0_269_727 ();
 DECAPx2_ASAP7_75t_R FILLER_0_269_739 ();
 DECAPx6_ASAP7_75t_R FILLER_0_269_748 ();
 FILLER_ASAP7_75t_R FILLER_0_269_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_764 ();
 FILLER_ASAP7_75t_R FILLER_0_269_787 ();
 FILLER_ASAP7_75t_R FILLER_0_269_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_797 ();
 FILLER_ASAP7_75t_R FILLER_0_269_820 ();
 FILLER_ASAP7_75t_R FILLER_0_269_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_829 ();
 FILLER_ASAP7_75t_R FILLER_0_269_852 ();
 FILLER_ASAP7_75t_R FILLER_0_269_857 ();
 DECAPx2_ASAP7_75t_R FILLER_0_269_865 ();
 FILLER_ASAP7_75t_R FILLER_0_269_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_879 ();
 FILLER_ASAP7_75t_R FILLER_0_269_888 ();
 FILLER_ASAP7_75t_R FILLER_0_269_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_895 ();
 DECAPx2_ASAP7_75t_R FILLER_0_269_906 ();
 FILLER_ASAP7_75t_R FILLER_0_269_923 ();
 DECAPx2_ASAP7_75t_R FILLER_0_269_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_933 ();
 DECAPx10_ASAP7_75t_R FILLER_0_269_944 ();
 DECAPx4_ASAP7_75t_R FILLER_0_269_966 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_976 ();
 DECAPx4_ASAP7_75t_R FILLER_0_269_983 ();
 FILLER_ASAP7_75t_R FILLER_0_269_999 ();
 DECAPx4_ASAP7_75t_R FILLER_0_269_1011 ();
 DECAPx2_ASAP7_75t_R FILLER_0_269_1027 ();
 FILLER_ASAP7_75t_R FILLER_0_269_1033 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_1035 ();
 FILLER_ASAP7_75t_R FILLER_0_269_1042 ();
 FILLER_ASAP7_75t_R FILLER_0_269_1054 ();
 DECAPx2_ASAP7_75t_R FILLER_0_269_1067 ();
 DECAPx4_ASAP7_75t_R FILLER_0_269_1079 ();
 FILLER_ASAP7_75t_R FILLER_0_269_1095 ();
 DECAPx10_ASAP7_75t_R FILLER_0_269_1103 ();
 DECAPx4_ASAP7_75t_R FILLER_0_269_1125 ();
 FILLER_ASAP7_75t_R FILLER_0_269_1135 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_1137 ();
 FILLER_ASAP7_75t_R FILLER_0_269_1144 ();
 DECAPx10_ASAP7_75t_R FILLER_0_269_1152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_269_1174 ();
 DECAPx6_ASAP7_75t_R FILLER_0_269_1196 ();
 FILLER_ASAP7_75t_R FILLER_0_269_1210 ();
 DECAPx6_ASAP7_75t_R FILLER_0_269_1218 ();
 DECAPx2_ASAP7_75t_R FILLER_0_269_1232 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_1238 ();
 DECAPx1_ASAP7_75t_R FILLER_0_269_1245 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_1249 ();
 DECAPx10_ASAP7_75t_R FILLER_0_269_1256 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_1278 ();
 FILLER_ASAP7_75t_R FILLER_0_269_1284 ();
 FILLER_ASAP7_75t_R FILLER_0_269_1289 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_1291 ();
 FILLER_ASAP7_75t_R FILLER_0_269_1298 ();
 DECAPx6_ASAP7_75t_R FILLER_0_269_1305 ();
 DECAPx2_ASAP7_75t_R FILLER_0_269_1319 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_1325 ();
 FILLER_ASAP7_75t_R FILLER_0_269_1332 ();
 DECAPx2_ASAP7_75t_R FILLER_0_269_1340 ();
 FILLER_ASAP7_75t_R FILLER_0_269_1346 ();
 FILLER_ASAP7_75t_R FILLER_0_269_1355 ();
 DECAPx6_ASAP7_75t_R FILLER_0_269_1363 ();
 DECAPx1_ASAP7_75t_R FILLER_0_269_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_270_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_270_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_270_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_270_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_270_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_270_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_270_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_270_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_270_178 ();
 DECAPx4_ASAP7_75t_R FILLER_0_270_200 ();
 FILLER_ASAP7_75t_R FILLER_0_270_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_212 ();
 DECAPx2_ASAP7_75t_R FILLER_0_270_221 ();
 FILLER_ASAP7_75t_R FILLER_0_270_227 ();
 FILLER_ASAP7_75t_R FILLER_0_270_232 ();
 DECAPx6_ASAP7_75t_R FILLER_0_270_240 ();
 DECAPx1_ASAP7_75t_R FILLER_0_270_254 ();
 DECAPx2_ASAP7_75t_R FILLER_0_270_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_270 ();
 FILLER_ASAP7_75t_R FILLER_0_270_277 ();
 FILLER_ASAP7_75t_R FILLER_0_270_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_292 ();
 FILLER_ASAP7_75t_R FILLER_0_270_299 ();
 DECAPx2_ASAP7_75t_R FILLER_0_270_307 ();
 FILLER_ASAP7_75t_R FILLER_0_270_313 ();
 FILLER_ASAP7_75t_R FILLER_0_270_321 ();
 DECAPx2_ASAP7_75t_R FILLER_0_270_329 ();
 FILLER_ASAP7_75t_R FILLER_0_270_342 ();
 FILLER_ASAP7_75t_R FILLER_0_270_364 ();
 DECAPx1_ASAP7_75t_R FILLER_0_270_370 ();
 FILLER_ASAP7_75t_R FILLER_0_270_379 ();
 FILLER_ASAP7_75t_R FILLER_0_270_386 ();
 FILLER_ASAP7_75t_R FILLER_0_270_393 ();
 FILLER_ASAP7_75t_R FILLER_0_270_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_403 ();
 FILLER_ASAP7_75t_R FILLER_0_270_407 ();
 FILLER_ASAP7_75t_R FILLER_0_270_414 ();
 FILLER_ASAP7_75t_R FILLER_0_270_422 ();
 FILLER_ASAP7_75t_R FILLER_0_270_427 ();
 FILLER_ASAP7_75t_R FILLER_0_270_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_437 ();
 FILLER_ASAP7_75t_R FILLER_0_270_443 ();
 FILLER_ASAP7_75t_R FILLER_0_270_450 ();
 DECAPx1_ASAP7_75t_R FILLER_0_270_458 ();
 FILLER_ASAP7_75t_R FILLER_0_270_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_466 ();
 FILLER_ASAP7_75t_R FILLER_0_270_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_475 ();
 FILLER_ASAP7_75t_R FILLER_0_270_481 ();
 DECAPx1_ASAP7_75t_R FILLER_0_270_489 ();
 FILLER_ASAP7_75t_R FILLER_0_270_498 ();
 DECAPx1_ASAP7_75t_R FILLER_0_270_510 ();
 FILLER_ASAP7_75t_R FILLER_0_270_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_522 ();
 DECAPx1_ASAP7_75t_R FILLER_0_270_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_548 ();
 FILLER_ASAP7_75t_R FILLER_0_270_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_557 ();
 FILLER_ASAP7_75t_R FILLER_0_270_561 ();
 FILLER_ASAP7_75t_R FILLER_0_270_568 ();
 FILLER_ASAP7_75t_R FILLER_0_270_575 ();
 DECAPx1_ASAP7_75t_R FILLER_0_270_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_602 ();
 FILLER_ASAP7_75t_R FILLER_0_270_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_611 ();
 DECAPx1_ASAP7_75t_R FILLER_0_270_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_622 ();
 DECAPx1_ASAP7_75t_R FILLER_0_270_644 ();
 DECAPx2_ASAP7_75t_R FILLER_0_270_669 ();
 DECAPx1_ASAP7_75t_R FILLER_0_270_680 ();
 DECAPx1_ASAP7_75t_R FILLER_0_270_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_693 ();
 FILLER_ASAP7_75t_R FILLER_0_270_704 ();
 DECAPx1_ASAP7_75t_R FILLER_0_270_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_713 ();
 DECAPx2_ASAP7_75t_R FILLER_0_270_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_726 ();
 FILLER_ASAP7_75t_R FILLER_0_270_733 ();
 FILLER_ASAP7_75t_R FILLER_0_270_741 ();
 FILLER_ASAP7_75t_R FILLER_0_270_764 ();
 FILLER_ASAP7_75t_R FILLER_0_270_776 ();
 FILLER_ASAP7_75t_R FILLER_0_270_783 ();
 DECAPx2_ASAP7_75t_R FILLER_0_270_807 ();
 FILLER_ASAP7_75t_R FILLER_0_270_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_820 ();
 FILLER_ASAP7_75t_R FILLER_0_270_826 ();
 FILLER_ASAP7_75t_R FILLER_0_270_834 ();
 FILLER_ASAP7_75t_R FILLER_0_270_842 ();
 FILLER_ASAP7_75t_R FILLER_0_270_849 ();
 DECAPx1_ASAP7_75t_R FILLER_0_270_856 ();
 FILLER_ASAP7_75t_R FILLER_0_270_866 ();
 DECAPx1_ASAP7_75t_R FILLER_0_270_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_878 ();
 FILLER_ASAP7_75t_R FILLER_0_270_885 ();
 FILLER_ASAP7_75t_R FILLER_0_270_893 ();
 DECAPx1_ASAP7_75t_R FILLER_0_270_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_905 ();
 FILLER_ASAP7_75t_R FILLER_0_270_912 ();
 FILLER_ASAP7_75t_R FILLER_0_270_920 ();
 FILLER_ASAP7_75t_R FILLER_0_270_927 ();
 FILLER_ASAP7_75t_R FILLER_0_270_935 ();
 DECAPx4_ASAP7_75t_R FILLER_0_270_940 ();
 FILLER_ASAP7_75t_R FILLER_0_270_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_952 ();
 DECAPx2_ASAP7_75t_R FILLER_0_270_959 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_965 ();
 DECAPx6_ASAP7_75t_R FILLER_0_270_971 ();
 DECAPx2_ASAP7_75t_R FILLER_0_270_985 ();
 FILLER_ASAP7_75t_R FILLER_0_270_997 ();
 FILLER_ASAP7_75t_R FILLER_0_270_1019 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_1021 ();
 DECAPx1_ASAP7_75t_R FILLER_0_270_1028 ();
 FILLER_ASAP7_75t_R FILLER_0_270_1038 ();
 DECAPx1_ASAP7_75t_R FILLER_0_270_1047 ();
 DECAPx1_ASAP7_75t_R FILLER_0_270_1057 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_1061 ();
 DECAPx1_ASAP7_75t_R FILLER_0_270_1068 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_1072 ();
 DECAPx2_ASAP7_75t_R FILLER_0_270_1079 ();
 FILLER_ASAP7_75t_R FILLER_0_270_1085 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_1087 ();
 DECAPx10_ASAP7_75t_R FILLER_0_270_1101 ();
 DECAPx10_ASAP7_75t_R FILLER_0_270_1123 ();
 DECAPx4_ASAP7_75t_R FILLER_0_270_1145 ();
 FILLER_ASAP7_75t_R FILLER_0_270_1155 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_1157 ();
 DECAPx6_ASAP7_75t_R FILLER_0_270_1164 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_1178 ();
 DECAPx4_ASAP7_75t_R FILLER_0_270_1185 ();
 FILLER_ASAP7_75t_R FILLER_0_270_1195 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_1197 ();
 FILLER_ASAP7_75t_R FILLER_0_270_1204 ();
 FILLER_ASAP7_75t_R FILLER_0_270_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_1214 ();
 DECAPx1_ASAP7_75t_R FILLER_0_270_1221 ();
 FILLER_ASAP7_75t_R FILLER_0_270_1231 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_1233 ();
 DECAPx2_ASAP7_75t_R FILLER_0_270_1240 ();
 FILLER_ASAP7_75t_R FILLER_0_270_1252 ();
 FILLER_ASAP7_75t_R FILLER_0_270_1264 ();
 FILLER_ASAP7_75t_R FILLER_0_270_1274 ();
 FILLER_ASAP7_75t_R FILLER_0_270_1284 ();
 FILLER_ASAP7_75t_R FILLER_0_270_1292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_270_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_270_1322 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_1344 ();
 FILLER_ASAP7_75t_R FILLER_0_270_1351 ();
 DECAPx10_ASAP7_75t_R FILLER_0_270_1359 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_271_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_271_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_271_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_271_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_271_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_271_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_271_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_271_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_271_178 ();
 DECAPx4_ASAP7_75t_R FILLER_0_271_200 ();
 FILLER_ASAP7_75t_R FILLER_0_271_210 ();
 FILLER_ASAP7_75t_R FILLER_0_271_233 ();
 DECAPx6_ASAP7_75t_R FILLER_0_271_241 ();
 DECAPx1_ASAP7_75t_R FILLER_0_271_255 ();
 DECAPx10_ASAP7_75t_R FILLER_0_271_265 ();
 FILLER_ASAP7_75t_R FILLER_0_271_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_295 ();
 DECAPx10_ASAP7_75t_R FILLER_0_271_302 ();
 FILLER_ASAP7_75t_R FILLER_0_271_324 ();
 FILLER_ASAP7_75t_R FILLER_0_271_332 ();
 DECAPx2_ASAP7_75t_R FILLER_0_271_344 ();
 DECAPx1_ASAP7_75t_R FILLER_0_271_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_360 ();
 FILLER_ASAP7_75t_R FILLER_0_271_366 ();
 FILLER_ASAP7_75t_R FILLER_0_271_374 ();
 FILLER_ASAP7_75t_R FILLER_0_271_381 ();
 FILLER_ASAP7_75t_R FILLER_0_271_388 ();
 FILLER_ASAP7_75t_R FILLER_0_271_395 ();
 FILLER_ASAP7_75t_R FILLER_0_271_403 ();
 FILLER_ASAP7_75t_R FILLER_0_271_411 ();
 FILLER_ASAP7_75t_R FILLER_0_271_418 ();
 FILLER_ASAP7_75t_R FILLER_0_271_425 ();
 DECAPx1_ASAP7_75t_R FILLER_0_271_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_437 ();
 FILLER_ASAP7_75t_R FILLER_0_271_443 ();
 DECAPx2_ASAP7_75t_R FILLER_0_271_451 ();
 FILLER_ASAP7_75t_R FILLER_0_271_464 ();
 FILLER_ASAP7_75t_R FILLER_0_271_477 ();
 FILLER_ASAP7_75t_R FILLER_0_271_482 ();
 FILLER_ASAP7_75t_R FILLER_0_271_489 ();
 FILLER_ASAP7_75t_R FILLER_0_271_497 ();
 FILLER_ASAP7_75t_R FILLER_0_271_504 ();
 FILLER_ASAP7_75t_R FILLER_0_271_512 ();
 DECAPx1_ASAP7_75t_R FILLER_0_271_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_524 ();
 FILLER_ASAP7_75t_R FILLER_0_271_530 ();
 FILLER_ASAP7_75t_R FILLER_0_271_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_540 ();
 FILLER_ASAP7_75t_R FILLER_0_271_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_549 ();
 FILLER_ASAP7_75t_R FILLER_0_271_555 ();
 DECAPx1_ASAP7_75t_R FILLER_0_271_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_583 ();
 FILLER_ASAP7_75t_R FILLER_0_271_589 ();
 FILLER_ASAP7_75t_R FILLER_0_271_596 ();
 FILLER_ASAP7_75t_R FILLER_0_271_603 ();
 FILLER_ASAP7_75t_R FILLER_0_271_610 ();
 FILLER_ASAP7_75t_R FILLER_0_271_617 ();
 FILLER_ASAP7_75t_R FILLER_0_271_624 ();
 FILLER_ASAP7_75t_R FILLER_0_271_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_634 ();
 FILLER_ASAP7_75t_R FILLER_0_271_640 ();
 FILLER_ASAP7_75t_R FILLER_0_271_647 ();
 FILLER_ASAP7_75t_R FILLER_0_271_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_657 ();
 DECAPx2_ASAP7_75t_R FILLER_0_271_664 ();
 DECAPx2_ASAP7_75t_R FILLER_0_271_675 ();
 FILLER_ASAP7_75t_R FILLER_0_271_686 ();
 FILLER_ASAP7_75t_R FILLER_0_271_693 ();
 FILLER_ASAP7_75t_R FILLER_0_271_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_702 ();
 FILLER_ASAP7_75t_R FILLER_0_271_708 ();
 FILLER_ASAP7_75t_R FILLER_0_271_713 ();
 DECAPx1_ASAP7_75t_R FILLER_0_271_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_722 ();
 DECAPx2_ASAP7_75t_R FILLER_0_271_728 ();
 FILLER_ASAP7_75t_R FILLER_0_271_734 ();
 DECAPx2_ASAP7_75t_R FILLER_0_271_741 ();
 FILLER_ASAP7_75t_R FILLER_0_271_747 ();
 FILLER_ASAP7_75t_R FILLER_0_271_752 ();
 FILLER_ASAP7_75t_R FILLER_0_271_760 ();
 FILLER_ASAP7_75t_R FILLER_0_271_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_767 ();
 DECAPx2_ASAP7_75t_R FILLER_0_271_773 ();
 FILLER_ASAP7_75t_R FILLER_0_271_784 ();
 DECAPx1_ASAP7_75t_R FILLER_0_271_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_795 ();
 FILLER_ASAP7_75t_R FILLER_0_271_801 ();
 FILLER_ASAP7_75t_R FILLER_0_271_808 ();
 FILLER_ASAP7_75t_R FILLER_0_271_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_817 ();
 FILLER_ASAP7_75t_R FILLER_0_271_823 ();
 FILLER_ASAP7_75t_R FILLER_0_271_846 ();
 FILLER_ASAP7_75t_R FILLER_0_271_853 ();
 DECAPx2_ASAP7_75t_R FILLER_0_271_860 ();
 DECAPx2_ASAP7_75t_R FILLER_0_271_872 ();
 FILLER_ASAP7_75t_R FILLER_0_271_884 ();
 FILLER_ASAP7_75t_R FILLER_0_271_891 ();
 FILLER_ASAP7_75t_R FILLER_0_271_899 ();
 FILLER_ASAP7_75t_R FILLER_0_271_906 ();
 FILLER_ASAP7_75t_R FILLER_0_271_913 ();
 DECAPx1_ASAP7_75t_R FILLER_0_271_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_924 ();
 FILLER_ASAP7_75t_R FILLER_0_271_927 ();
 FILLER_ASAP7_75t_R FILLER_0_271_932 ();
 DECAPx4_ASAP7_75t_R FILLER_0_271_940 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_950 ();
 FILLER_ASAP7_75t_R FILLER_0_271_957 ();
 FILLER_ASAP7_75t_R FILLER_0_271_965 ();
 FILLER_ASAP7_75t_R FILLER_0_271_978 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_980 ();
 DECAPx6_ASAP7_75t_R FILLER_0_271_987 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_1001 ();
 DECAPx4_ASAP7_75t_R FILLER_0_271_1008 ();
 FILLER_ASAP7_75t_R FILLER_0_271_1018 ();
 FILLER_ASAP7_75t_R FILLER_0_271_1026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_271_1034 ();
 DECAPx4_ASAP7_75t_R FILLER_0_271_1056 ();
 FILLER_ASAP7_75t_R FILLER_0_271_1072 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_1074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_271_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_0_271_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_0_271_1125 ();
 FILLER_ASAP7_75t_R FILLER_0_271_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_1149 ();
 FILLER_ASAP7_75t_R FILLER_0_271_1156 ();
 FILLER_ASAP7_75t_R FILLER_0_271_1166 ();
 FILLER_ASAP7_75t_R FILLER_0_271_1174 ();
 DECAPx1_ASAP7_75t_R FILLER_0_271_1182 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_1186 ();
 FILLER_ASAP7_75t_R FILLER_0_271_1193 ();
 FILLER_ASAP7_75t_R FILLER_0_271_1205 ();
 DECAPx2_ASAP7_75t_R FILLER_0_271_1213 ();
 FILLER_ASAP7_75t_R FILLER_0_271_1219 ();
 DECAPx4_ASAP7_75t_R FILLER_0_271_1227 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_1237 ();
 FILLER_ASAP7_75t_R FILLER_0_271_1248 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_1250 ();
 FILLER_ASAP7_75t_R FILLER_0_271_1261 ();
 FILLER_ASAP7_75t_R FILLER_0_271_1269 ();
 DECAPx1_ASAP7_75t_R FILLER_0_271_1277 ();
 FILLER_ASAP7_75t_R FILLER_0_271_1287 ();
 DECAPx10_ASAP7_75t_R FILLER_0_271_1295 ();
 DECAPx10_ASAP7_75t_R FILLER_0_271_1317 ();
 DECAPx10_ASAP7_75t_R FILLER_0_271_1339 ();
 DECAPx6_ASAP7_75t_R FILLER_0_271_1361 ();
 DECAPx2_ASAP7_75t_R FILLER_0_271_1375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_272_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_272_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_272_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_272_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_272_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_272_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_272_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_272_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_272_178 ();
 DECAPx6_ASAP7_75t_R FILLER_0_272_200 ();
 FILLER_ASAP7_75t_R FILLER_0_272_217 ();
 DECAPx4_ASAP7_75t_R FILLER_0_272_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_234 ();
 FILLER_ASAP7_75t_R FILLER_0_272_243 ();
 DECAPx2_ASAP7_75t_R FILLER_0_272_248 ();
 FILLER_ASAP7_75t_R FILLER_0_272_260 ();
 FILLER_ASAP7_75t_R FILLER_0_272_268 ();
 DECAPx4_ASAP7_75t_R FILLER_0_272_276 ();
 FILLER_ASAP7_75t_R FILLER_0_272_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_288 ();
 DECAPx4_ASAP7_75t_R FILLER_0_272_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_305 ();
 FILLER_ASAP7_75t_R FILLER_0_272_312 ();
 DECAPx4_ASAP7_75t_R FILLER_0_272_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_330 ();
 FILLER_ASAP7_75t_R FILLER_0_272_337 ();
 FILLER_ASAP7_75t_R FILLER_0_272_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_347 ();
 DECAPx1_ASAP7_75t_R FILLER_0_272_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_358 ();
 FILLER_ASAP7_75t_R FILLER_0_272_364 ();
 DECAPx2_ASAP7_75t_R FILLER_0_272_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_378 ();
 FILLER_ASAP7_75t_R FILLER_0_272_385 ();
 FILLER_ASAP7_75t_R FILLER_0_272_393 ();
 DECAPx2_ASAP7_75t_R FILLER_0_272_401 ();
 FILLER_ASAP7_75t_R FILLER_0_272_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_415 ();
 FILLER_ASAP7_75t_R FILLER_0_272_421 ();
 FILLER_ASAP7_75t_R FILLER_0_272_429 ();
 FILLER_ASAP7_75t_R FILLER_0_272_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_439 ();
 FILLER_ASAP7_75t_R FILLER_0_272_445 ();
 FILLER_ASAP7_75t_R FILLER_0_272_453 ();
 FILLER_ASAP7_75t_R FILLER_0_272_460 ();
 FILLER_ASAP7_75t_R FILLER_0_272_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_466 ();
 FILLER_ASAP7_75t_R FILLER_0_272_473 ();
 DECAPx1_ASAP7_75t_R FILLER_0_272_485 ();
 FILLER_ASAP7_75t_R FILLER_0_272_494 ();
 FILLER_ASAP7_75t_R FILLER_0_272_501 ();
 FILLER_ASAP7_75t_R FILLER_0_272_508 ();
 FILLER_ASAP7_75t_R FILLER_0_272_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_518 ();
 FILLER_ASAP7_75t_R FILLER_0_272_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_527 ();
 FILLER_ASAP7_75t_R FILLER_0_272_534 ();
 FILLER_ASAP7_75t_R FILLER_0_272_541 ();
 FILLER_ASAP7_75t_R FILLER_0_272_548 ();
 FILLER_ASAP7_75t_R FILLER_0_272_555 ();
 FILLER_ASAP7_75t_R FILLER_0_272_562 ();
 FILLER_ASAP7_75t_R FILLER_0_272_569 ();
 FILLER_ASAP7_75t_R FILLER_0_272_577 ();
 FILLER_ASAP7_75t_R FILLER_0_272_584 ();
 FILLER_ASAP7_75t_R FILLER_0_272_592 ();
 FILLER_ASAP7_75t_R FILLER_0_272_597 ();
 FILLER_ASAP7_75t_R FILLER_0_272_604 ();
 FILLER_ASAP7_75t_R FILLER_0_272_611 ();
 FILLER_ASAP7_75t_R FILLER_0_272_618 ();
 FILLER_ASAP7_75t_R FILLER_0_272_625 ();
 FILLER_ASAP7_75t_R FILLER_0_272_632 ();
 FILLER_ASAP7_75t_R FILLER_0_272_639 ();
 FILLER_ASAP7_75t_R FILLER_0_272_646 ();
 FILLER_ASAP7_75t_R FILLER_0_272_653 ();
 FILLER_ASAP7_75t_R FILLER_0_272_660 ();
 FILLER_ASAP7_75t_R FILLER_0_272_667 ();
 DECAPx2_ASAP7_75t_R FILLER_0_272_690 ();
 FILLER_ASAP7_75t_R FILLER_0_272_702 ();
 FILLER_ASAP7_75t_R FILLER_0_272_709 ();
 FILLER_ASAP7_75t_R FILLER_0_272_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_718 ();
 DECAPx1_ASAP7_75t_R FILLER_0_272_725 ();
 DECAPx4_ASAP7_75t_R FILLER_0_272_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_749 ();
 FILLER_ASAP7_75t_R FILLER_0_272_755 ();
 FILLER_ASAP7_75t_R FILLER_0_272_763 ();
 FILLER_ASAP7_75t_R FILLER_0_272_770 ();
 FILLER_ASAP7_75t_R FILLER_0_272_778 ();
 FILLER_ASAP7_75t_R FILLER_0_272_785 ();
 DECAPx2_ASAP7_75t_R FILLER_0_272_792 ();
 FILLER_ASAP7_75t_R FILLER_0_272_803 ();
 FILLER_ASAP7_75t_R FILLER_0_272_810 ();
 FILLER_ASAP7_75t_R FILLER_0_272_817 ();
 FILLER_ASAP7_75t_R FILLER_0_272_824 ();
 FILLER_ASAP7_75t_R FILLER_0_272_832 ();
 FILLER_ASAP7_75t_R FILLER_0_272_837 ();
 FILLER_ASAP7_75t_R FILLER_0_272_861 ();
 DECAPx1_ASAP7_75t_R FILLER_0_272_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_872 ();
 FILLER_ASAP7_75t_R FILLER_0_272_889 ();
 DECAPx2_ASAP7_75t_R FILLER_0_272_896 ();
 FILLER_ASAP7_75t_R FILLER_0_272_908 ();
 FILLER_ASAP7_75t_R FILLER_0_272_916 ();
 FILLER_ASAP7_75t_R FILLER_0_272_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_925 ();
 FILLER_ASAP7_75t_R FILLER_0_272_937 ();
 FILLER_ASAP7_75t_R FILLER_0_272_945 ();
 FILLER_ASAP7_75t_R FILLER_0_272_953 ();
 DECAPx2_ASAP7_75t_R FILLER_0_272_961 ();
 FILLER_ASAP7_75t_R FILLER_0_272_967 ();
 DECAPx6_ASAP7_75t_R FILLER_0_272_975 ();
 DECAPx2_ASAP7_75t_R FILLER_0_272_989 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_995 ();
 DECAPx6_ASAP7_75t_R FILLER_0_272_1012 ();
 DECAPx2_ASAP7_75t_R FILLER_0_272_1026 ();
 DECAPx2_ASAP7_75t_R FILLER_0_272_1038 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_1044 ();
 DECAPx2_ASAP7_75t_R FILLER_0_272_1051 ();
 FILLER_ASAP7_75t_R FILLER_0_272_1063 ();
 FILLER_ASAP7_75t_R FILLER_0_272_1072 ();
 FILLER_ASAP7_75t_R FILLER_0_272_1080 ();
 FILLER_ASAP7_75t_R FILLER_0_272_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_0_272_1100 ();
 DECAPx10_ASAP7_75t_R FILLER_0_272_1122 ();
 DECAPx10_ASAP7_75t_R FILLER_0_272_1144 ();
 DECAPx6_ASAP7_75t_R FILLER_0_272_1166 ();
 FILLER_ASAP7_75t_R FILLER_0_272_1180 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_1182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_272_1189 ();
 DECAPx10_ASAP7_75t_R FILLER_0_272_1211 ();
 DECAPx2_ASAP7_75t_R FILLER_0_272_1233 ();
 FILLER_ASAP7_75t_R FILLER_0_272_1239 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_1241 ();
 DECAPx10_ASAP7_75t_R FILLER_0_272_1245 ();
 DECAPx10_ASAP7_75t_R FILLER_0_272_1267 ();
 DECAPx10_ASAP7_75t_R FILLER_0_272_1289 ();
 DECAPx10_ASAP7_75t_R FILLER_0_272_1311 ();
 DECAPx10_ASAP7_75t_R FILLER_0_272_1333 ();
 DECAPx10_ASAP7_75t_R FILLER_0_272_1355 ();
 DECAPx1_ASAP7_75t_R FILLER_0_272_1377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_1381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273_200 ();
 DECAPx2_ASAP7_75t_R FILLER_0_273_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_273_228 ();
 FILLER_ASAP7_75t_R FILLER_0_273_232 ();
 FILLER_ASAP7_75t_R FILLER_0_273_240 ();
 DECAPx6_ASAP7_75t_R FILLER_0_273_249 ();
 FILLER_ASAP7_75t_R FILLER_0_273_269 ();
 DECAPx1_ASAP7_75t_R FILLER_0_273_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_273_283 ();
 FILLER_ASAP7_75t_R FILLER_0_273_290 ();
 DECAPx1_ASAP7_75t_R FILLER_0_273_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_273_306 ();
 FILLER_ASAP7_75t_R FILLER_0_273_318 ();
 DECAPx1_ASAP7_75t_R FILLER_0_273_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_273_330 ();
 FILLER_ASAP7_75t_R FILLER_0_273_336 ();
 DECAPx1_ASAP7_75t_R FILLER_0_273_344 ();
 DECAPx1_ASAP7_75t_R FILLER_0_273_354 ();
 DECAPx2_ASAP7_75t_R FILLER_0_273_364 ();
 DECAPx1_ASAP7_75t_R FILLER_0_273_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_273_380 ();
 FILLER_ASAP7_75t_R FILLER_0_273_387 ();
 FILLER_ASAP7_75t_R FILLER_0_273_395 ();
 DECAPx1_ASAP7_75t_R FILLER_0_273_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_273_407 ();
 FILLER_ASAP7_75t_R FILLER_0_273_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_273_416 ();
 FILLER_ASAP7_75t_R FILLER_0_273_423 ();
 FILLER_ASAP7_75t_R FILLER_0_273_431 ();
 FILLER_ASAP7_75t_R FILLER_0_273_443 ();
 DECAPx1_ASAP7_75t_R FILLER_0_273_456 ();
 FILLER_ASAP7_75t_R FILLER_0_273_466 ();
 FILLER_ASAP7_75t_R FILLER_0_273_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_273_476 ();
 FILLER_ASAP7_75t_R FILLER_0_273_482 ();
 FILLER_ASAP7_75t_R FILLER_0_273_489 ();
 DECAPx1_ASAP7_75t_R FILLER_0_273_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_273_501 ();
 FILLER_ASAP7_75t_R FILLER_0_273_507 ();
 FILLER_ASAP7_75t_R FILLER_0_273_530 ();
 FILLER_ASAP7_75t_R FILLER_0_273_553 ();
 FILLER_ASAP7_75t_R FILLER_0_273_558 ();
 FILLER_ASAP7_75t_R FILLER_0_273_582 ();
 FILLER_ASAP7_75t_R FILLER_0_273_587 ();
 FILLER_ASAP7_75t_R FILLER_0_273_610 ();
 FILLER_ASAP7_75t_R FILLER_0_273_634 ();
 DECAPx1_ASAP7_75t_R FILLER_0_273_642 ();
 FILLER_ASAP7_75t_R FILLER_0_273_668 ();
 FILLER_ASAP7_75t_R FILLER_0_273_673 ();
 FILLER_ASAP7_75t_R FILLER_0_273_681 ();
 FILLER_ASAP7_75t_R FILLER_0_273_689 ();
 FILLER_ASAP7_75t_R FILLER_0_273_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_273_715 ();
 DECAPx1_ASAP7_75t_R FILLER_0_273_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_273_741 ();
 FILLER_ASAP7_75t_R FILLER_0_273_747 ();
 DECAPx2_ASAP7_75t_R FILLER_0_273_754 ();
 FILLER_ASAP7_75t_R FILLER_0_273_760 ();
 FILLER_ASAP7_75t_R FILLER_0_273_783 ();
 FILLER_ASAP7_75t_R FILLER_0_273_806 ();
 FILLER_ASAP7_75t_R FILLER_0_273_814 ();
 FILLER_ASAP7_75t_R FILLER_0_273_821 ();
 FILLER_ASAP7_75t_R FILLER_0_273_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_273_828 ();
 FILLER_ASAP7_75t_R FILLER_0_273_850 ();
 FILLER_ASAP7_75t_R FILLER_0_273_857 ();
 DECAPx2_ASAP7_75t_R FILLER_0_273_864 ();
 FILLER_ASAP7_75t_R FILLER_0_273_876 ();
 FILLER_ASAP7_75t_R FILLER_0_273_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_273_891 ();
 FILLER_ASAP7_75t_R FILLER_0_273_898 ();
 FILLER_ASAP7_75t_R FILLER_0_273_906 ();
 FILLER_ASAP7_75t_R FILLER_0_273_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_273_916 ();
 FILLER_ASAP7_75t_R FILLER_0_273_923 ();
 FILLER_ASAP7_75t_R FILLER_0_273_927 ();
 FILLER_ASAP7_75t_R FILLER_0_273_932 ();
 FILLER_ASAP7_75t_R FILLER_0_273_942 ();
 DECAPx1_ASAP7_75t_R FILLER_0_273_950 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_273_954 ();
 FILLER_ASAP7_75t_R FILLER_0_273_961 ();
 FILLER_ASAP7_75t_R FILLER_0_273_969 ();
 DECAPx1_ASAP7_75t_R FILLER_0_273_974 ();
 DECAPx2_ASAP7_75t_R FILLER_0_273_984 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_273_990 ();
 FILLER_ASAP7_75t_R FILLER_0_273_997 ();
 DECAPx1_ASAP7_75t_R FILLER_0_273_1019 ();
 FILLER_ASAP7_75t_R FILLER_0_273_1029 ();
 FILLER_ASAP7_75t_R FILLER_0_273_1042 ();
 DECAPx2_ASAP7_75t_R FILLER_0_273_1050 ();
 FILLER_ASAP7_75t_R FILLER_0_273_1056 ();
 FILLER_ASAP7_75t_R FILLER_0_273_1065 ();
 DECAPx1_ASAP7_75t_R FILLER_0_273_1083 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_273_1087 ();
 FILLER_ASAP7_75t_R FILLER_0_273_1094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_273_1366 ();
 FILLER_ASAP7_75t_R FILLER_0_273_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_200 ();
 DECAPx1_ASAP7_75t_R FILLER_0_274_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_274_226 ();
 FILLER_ASAP7_75t_R FILLER_0_274_248 ();
 DECAPx2_ASAP7_75t_R FILLER_0_274_272 ();
 FILLER_ASAP7_75t_R FILLER_0_274_278 ();
 DECAPx1_ASAP7_75t_R FILLER_0_274_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_274_287 ();
 DECAPx6_ASAP7_75t_R FILLER_0_274_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_274_308 ();
 FILLER_ASAP7_75t_R FILLER_0_274_315 ();
 DECAPx1_ASAP7_75t_R FILLER_0_274_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_274_327 ();
 FILLER_ASAP7_75t_R FILLER_0_274_331 ();
 DECAPx1_ASAP7_75t_R FILLER_0_274_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_274_343 ();
 FILLER_ASAP7_75t_R FILLER_0_274_349 ();
 DECAPx1_ASAP7_75t_R FILLER_0_274_357 ();
 FILLER_ASAP7_75t_R FILLER_0_274_366 ();
 FILLER_ASAP7_75t_R FILLER_0_274_378 ();
 DECAPx1_ASAP7_75t_R FILLER_0_274_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_274_390 ();
 DECAPx2_ASAP7_75t_R FILLER_0_274_397 ();
 FILLER_ASAP7_75t_R FILLER_0_274_408 ();
 FILLER_ASAP7_75t_R FILLER_0_274_416 ();
 FILLER_ASAP7_75t_R FILLER_0_274_424 ();
 FILLER_ASAP7_75t_R FILLER_0_274_429 ();
 FILLER_ASAP7_75t_R FILLER_0_274_436 ();
 FILLER_ASAP7_75t_R FILLER_0_274_443 ();
 DECAPx1_ASAP7_75t_R FILLER_0_274_451 ();
 FILLER_ASAP7_75t_R FILLER_0_274_460 ();
 FILLER_ASAP7_75t_R FILLER_0_274_464 ();
 FILLER_ASAP7_75t_R FILLER_0_274_472 ();
 FILLER_ASAP7_75t_R FILLER_0_274_495 ();
 DECAPx1_ASAP7_75t_R FILLER_0_274_503 ();
 FILLER_ASAP7_75t_R FILLER_0_274_512 ();
 FILLER_ASAP7_75t_R FILLER_0_274_520 ();
 FILLER_ASAP7_75t_R FILLER_0_274_532 ();
 FILLER_ASAP7_75t_R FILLER_0_274_539 ();
 FILLER_ASAP7_75t_R FILLER_0_274_547 ();
 FILLER_ASAP7_75t_R FILLER_0_274_555 ();
 FILLER_ASAP7_75t_R FILLER_0_274_567 ();
 DECAPx1_ASAP7_75t_R FILLER_0_274_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_274_583 ();
 FILLER_ASAP7_75t_R FILLER_0_274_589 ();
 FILLER_ASAP7_75t_R FILLER_0_274_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_274_599 ();
 FILLER_ASAP7_75t_R FILLER_0_274_605 ();
 FILLER_ASAP7_75t_R FILLER_0_274_613 ();
 DECAPx1_ASAP7_75t_R FILLER_0_274_621 ();
 FILLER_ASAP7_75t_R FILLER_0_274_630 ();
 FILLER_ASAP7_75t_R FILLER_0_274_638 ();
 DECAPx2_ASAP7_75t_R FILLER_0_274_646 ();
 FILLER_ASAP7_75t_R FILLER_0_274_657 ();
 FILLER_ASAP7_75t_R FILLER_0_274_664 ();
 FILLER_ASAP7_75t_R FILLER_0_274_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_274_674 ();
 FILLER_ASAP7_75t_R FILLER_0_274_680 ();
 FILLER_ASAP7_75t_R FILLER_0_274_687 ();
 FILLER_ASAP7_75t_R FILLER_0_274_694 ();
 FILLER_ASAP7_75t_R FILLER_0_274_701 ();
 FILLER_ASAP7_75t_R FILLER_0_274_708 ();
 FILLER_ASAP7_75t_R FILLER_0_274_715 ();
 FILLER_ASAP7_75t_R FILLER_0_274_723 ();
 FILLER_ASAP7_75t_R FILLER_0_274_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_274_732 ();
 FILLER_ASAP7_75t_R FILLER_0_274_738 ();
 FILLER_ASAP7_75t_R FILLER_0_274_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_274_747 ();
 FILLER_ASAP7_75t_R FILLER_0_274_758 ();
 FILLER_ASAP7_75t_R FILLER_0_274_765 ();
 FILLER_ASAP7_75t_R FILLER_0_274_770 ();
 FILLER_ASAP7_75t_R FILLER_0_274_778 ();
 FILLER_ASAP7_75t_R FILLER_0_274_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_274_787 ();
 FILLER_ASAP7_75t_R FILLER_0_274_794 ();
 FILLER_ASAP7_75t_R FILLER_0_274_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_274_801 ();
 FILLER_ASAP7_75t_R FILLER_0_274_823 ();
 FILLER_ASAP7_75t_R FILLER_0_274_830 ();
 FILLER_ASAP7_75t_R FILLER_0_274_837 ();
 FILLER_ASAP7_75t_R FILLER_0_274_844 ();
 FILLER_ASAP7_75t_R FILLER_0_274_868 ();
 FILLER_ASAP7_75t_R FILLER_0_274_875 ();
 FILLER_ASAP7_75t_R FILLER_0_274_882 ();
 DECAPx2_ASAP7_75t_R FILLER_0_274_889 ();
 FILLER_ASAP7_75t_R FILLER_0_274_906 ();
 FILLER_ASAP7_75t_R FILLER_0_274_913 ();
 DECAPx1_ASAP7_75t_R FILLER_0_274_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_274_924 ();
 DECAPx2_ASAP7_75t_R FILLER_0_274_931 ();
 FILLER_ASAP7_75t_R FILLER_0_274_943 ();
 FILLER_ASAP7_75t_R FILLER_0_274_950 ();
 DECAPx6_ASAP7_75t_R FILLER_0_274_955 ();
 DECAPx2_ASAP7_75t_R FILLER_0_274_969 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_274_975 ();
 FILLER_ASAP7_75t_R FILLER_0_274_997 ();
 FILLER_ASAP7_75t_R FILLER_0_274_1004 ();
 DECAPx2_ASAP7_75t_R FILLER_0_274_1012 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_274_1018 ();
 FILLER_ASAP7_75t_R FILLER_0_274_1025 ();
 FILLER_ASAP7_75t_R FILLER_0_274_1033 ();
 FILLER_ASAP7_75t_R FILLER_0_274_1038 ();
 DECAPx4_ASAP7_75t_R FILLER_0_274_1051 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_274_1061 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_1068 ();
 FILLER_ASAP7_75t_R FILLER_0_274_1090 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_1098 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_1120 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_1142 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_1164 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_1186 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_1208 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_1230 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_1252 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_1274 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_1296 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_1318 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_1340 ();
 DECAPx6_ASAP7_75t_R FILLER_0_274_1362 ();
 DECAPx2_ASAP7_75t_R FILLER_0_274_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_178 ();
 DECAPx6_ASAP7_75t_R FILLER_0_275_200 ();
 DECAPx2_ASAP7_75t_R FILLER_0_275_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_275_220 ();
 FILLER_ASAP7_75t_R FILLER_0_275_224 ();
 FILLER_ASAP7_75t_R FILLER_0_275_231 ();
 FILLER_ASAP7_75t_R FILLER_0_275_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_275_241 ();
 FILLER_ASAP7_75t_R FILLER_0_275_245 ();
 DECAPx1_ASAP7_75t_R FILLER_0_275_252 ();
 FILLER_ASAP7_75t_R FILLER_0_275_261 ();
 FILLER_ASAP7_75t_R FILLER_0_275_268 ();
 DECAPx2_ASAP7_75t_R FILLER_0_275_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_275_281 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_287 ();
 DECAPx6_ASAP7_75t_R FILLER_0_275_309 ();
 DECAPx1_ASAP7_75t_R FILLER_0_275_323 ();
 FILLER_ASAP7_75t_R FILLER_0_275_332 ();
 FILLER_ASAP7_75t_R FILLER_0_275_339 ();
 FILLER_ASAP7_75t_R FILLER_0_275_346 ();
 FILLER_ASAP7_75t_R FILLER_0_275_353 ();
 FILLER_ASAP7_75t_R FILLER_0_275_360 ();
 FILLER_ASAP7_75t_R FILLER_0_275_367 ();
 FILLER_ASAP7_75t_R FILLER_0_275_374 ();
 FILLER_ASAP7_75t_R FILLER_0_275_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_275_384 ();
 FILLER_ASAP7_75t_R FILLER_0_275_388 ();
 FILLER_ASAP7_75t_R FILLER_0_275_395 ();
 FILLER_ASAP7_75t_R FILLER_0_275_402 ();
 FILLER_ASAP7_75t_R FILLER_0_275_409 ();
 FILLER_ASAP7_75t_R FILLER_0_275_416 ();
 FILLER_ASAP7_75t_R FILLER_0_275_423 ();
 FILLER_ASAP7_75t_R FILLER_0_275_430 ();
 FILLER_ASAP7_75t_R FILLER_0_275_437 ();
 FILLER_ASAP7_75t_R FILLER_0_275_444 ();
 FILLER_ASAP7_75t_R FILLER_0_275_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_275_454 ();
 FILLER_ASAP7_75t_R FILLER_0_275_460 ();
 FILLER_ASAP7_75t_R FILLER_0_275_464 ();
 FILLER_ASAP7_75t_R FILLER_0_275_469 ();
 FILLER_ASAP7_75t_R FILLER_0_275_476 ();
 FILLER_ASAP7_75t_R FILLER_0_275_483 ();
 FILLER_ASAP7_75t_R FILLER_0_275_490 ();
 FILLER_ASAP7_75t_R FILLER_0_275_497 ();
 FILLER_ASAP7_75t_R FILLER_0_275_504 ();
 FILLER_ASAP7_75t_R FILLER_0_275_511 ();
 FILLER_ASAP7_75t_R FILLER_0_275_519 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_275_521 ();
 FILLER_ASAP7_75t_R FILLER_0_275_527 ();
 FILLER_ASAP7_75t_R FILLER_0_275_534 ();
 FILLER_ASAP7_75t_R FILLER_0_275_541 ();
 FILLER_ASAP7_75t_R FILLER_0_275_548 ();
 FILLER_ASAP7_75t_R FILLER_0_275_555 ();
 FILLER_ASAP7_75t_R FILLER_0_275_562 ();
 FILLER_ASAP7_75t_R FILLER_0_275_569 ();
 FILLER_ASAP7_75t_R FILLER_0_275_576 ();
 FILLER_ASAP7_75t_R FILLER_0_275_584 ();
 FILLER_ASAP7_75t_R FILLER_0_275_590 ();
 FILLER_ASAP7_75t_R FILLER_0_275_597 ();
 FILLER_ASAP7_75t_R FILLER_0_275_604 ();
 FILLER_ASAP7_75t_R FILLER_0_275_611 ();
 FILLER_ASAP7_75t_R FILLER_0_275_618 ();
 FILLER_ASAP7_75t_R FILLER_0_275_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_275_628 ();
 FILLER_ASAP7_75t_R FILLER_0_275_634 ();
 FILLER_ASAP7_75t_R FILLER_0_275_641 ();
 FILLER_ASAP7_75t_R FILLER_0_275_648 ();
 FILLER_ASAP7_75t_R FILLER_0_275_655 ();
 FILLER_ASAP7_75t_R FILLER_0_275_662 ();
 FILLER_ASAP7_75t_R FILLER_0_275_669 ();
 FILLER_ASAP7_75t_R FILLER_0_275_676 ();
 FILLER_ASAP7_75t_R FILLER_0_275_683 ();
 FILLER_ASAP7_75t_R FILLER_0_275_690 ();
 FILLER_ASAP7_75t_R FILLER_0_275_697 ();
 FILLER_ASAP7_75t_R FILLER_0_275_704 ();
 FILLER_ASAP7_75t_R FILLER_0_275_711 ();
 FILLER_ASAP7_75t_R FILLER_0_275_718 ();
 FILLER_ASAP7_75t_R FILLER_0_275_730 ();
 FILLER_ASAP7_75t_R FILLER_0_275_737 ();
 FILLER_ASAP7_75t_R FILLER_0_275_744 ();
 FILLER_ASAP7_75t_R FILLER_0_275_751 ();
 FILLER_ASAP7_75t_R FILLER_0_275_758 ();
 FILLER_ASAP7_75t_R FILLER_0_275_765 ();
 FILLER_ASAP7_75t_R FILLER_0_275_772 ();
 FILLER_ASAP7_75t_R FILLER_0_275_779 ();
 FILLER_ASAP7_75t_R FILLER_0_275_786 ();
 DECAPx1_ASAP7_75t_R FILLER_0_275_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_275_797 ();
 FILLER_ASAP7_75t_R FILLER_0_275_804 ();
 FILLER_ASAP7_75t_R FILLER_0_275_811 ();
 FILLER_ASAP7_75t_R FILLER_0_275_818 ();
 FILLER_ASAP7_75t_R FILLER_0_275_823 ();
 FILLER_ASAP7_75t_R FILLER_0_275_831 ();
 FILLER_ASAP7_75t_R FILLER_0_275_838 ();
 DECAPx2_ASAP7_75t_R FILLER_0_275_845 ();
 FILLER_ASAP7_75t_R FILLER_0_275_857 ();
 FILLER_ASAP7_75t_R FILLER_0_275_864 ();
 FILLER_ASAP7_75t_R FILLER_0_275_871 ();
 FILLER_ASAP7_75t_R FILLER_0_275_878 ();
 FILLER_ASAP7_75t_R FILLER_0_275_885 ();
 FILLER_ASAP7_75t_R FILLER_0_275_892 ();
 FILLER_ASAP7_75t_R FILLER_0_275_899 ();
 FILLER_ASAP7_75t_R FILLER_0_275_906 ();
 FILLER_ASAP7_75t_R FILLER_0_275_913 ();
 DECAPx1_ASAP7_75t_R FILLER_0_275_920 ();
 FILLER_ASAP7_75t_R FILLER_0_275_926 ();
 FILLER_ASAP7_75t_R FILLER_0_275_933 ();
 FILLER_ASAP7_75t_R FILLER_0_275_940 ();
 FILLER_ASAP7_75t_R FILLER_0_275_947 ();
 DECAPx4_ASAP7_75t_R FILLER_0_275_954 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_275_964 ();
 FILLER_ASAP7_75t_R FILLER_0_275_968 ();
 FILLER_ASAP7_75t_R FILLER_0_275_975 ();
 FILLER_ASAP7_75t_R FILLER_0_275_982 ();
 FILLER_ASAP7_75t_R FILLER_0_275_990 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_997 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_1019 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_1041 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_1063 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_1085 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_1107 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_1129 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_1151 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_1173 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_1195 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_1217 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_1239 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_1261 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_1283 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_1305 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_1327 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_1349 ();
 DECAPx4_ASAP7_75t_R FILLER_0_275_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_275_1381 ();
endmodule
