VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeregfile_64x64
  FOREIGN fakeregfile_64x64 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 8.360 BY 28.000 ;
  CLASS BLOCK ;
  PIN rdata_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.096 0.024 0.120 ;
    END
  END rdata_out[0]
  PIN rdata_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.192 0.024 0.216 ;
    END
  END rdata_out[1]
  PIN rdata_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.288 0.024 0.312 ;
    END
  END rdata_out[2]
  PIN rdata_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.384 0.024 0.408 ;
    END
  END rdata_out[3]
  PIN rdata_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.480 0.024 0.504 ;
    END
  END rdata_out[4]
  PIN rdata_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.576 0.024 0.600 ;
    END
  END rdata_out[5]
  PIN rdata_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.672 0.024 0.696 ;
    END
  END rdata_out[6]
  PIN rdata_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.768 0.024 0.792 ;
    END
  END rdata_out[7]
  PIN rdata_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.864 0.024 0.888 ;
    END
  END rdata_out[8]
  PIN rdata_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.960 0.024 0.984 ;
    END
  END rdata_out[9]
  PIN rdata_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.056 0.024 1.080 ;
    END
  END rdata_out[10]
  PIN rdata_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.152 0.024 1.176 ;
    END
  END rdata_out[11]
  PIN rdata_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.248 0.024 1.272 ;
    END
  END rdata_out[12]
  PIN rdata_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.344 0.024 1.368 ;
    END
  END rdata_out[13]
  PIN rdata_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.440 0.024 1.464 ;
    END
  END rdata_out[14]
  PIN rdata_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.536 0.024 1.560 ;
    END
  END rdata_out[15]
  PIN rdata_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.632 0.024 1.656 ;
    END
  END rdata_out[16]
  PIN rdata_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.728 0.024 1.752 ;
    END
  END rdata_out[17]
  PIN rdata_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.824 0.024 1.848 ;
    END
  END rdata_out[18]
  PIN rdata_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.920 0.024 1.944 ;
    END
  END rdata_out[19]
  PIN rdata_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.016 0.024 2.040 ;
    END
  END rdata_out[20]
  PIN rdata_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.112 0.024 2.136 ;
    END
  END rdata_out[21]
  PIN rdata_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.208 0.024 2.232 ;
    END
  END rdata_out[22]
  PIN rdata_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.304 0.024 2.328 ;
    END
  END rdata_out[23]
  PIN rdata_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.400 0.024 2.424 ;
    END
  END rdata_out[24]
  PIN rdata_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.496 0.024 2.520 ;
    END
  END rdata_out[25]
  PIN rdata_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.592 0.024 2.616 ;
    END
  END rdata_out[26]
  PIN rdata_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.688 0.024 2.712 ;
    END
  END rdata_out[27]
  PIN rdata_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.784 0.024 2.808 ;
    END
  END rdata_out[28]
  PIN rdata_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.880 0.024 2.904 ;
    END
  END rdata_out[29]
  PIN rdata_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.976 0.024 3.000 ;
    END
  END rdata_out[30]
  PIN rdata_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.072 0.024 3.096 ;
    END
  END rdata_out[31]
  PIN rdata_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.168 0.024 3.192 ;
    END
  END rdata_out[32]
  PIN rdata_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.264 0.024 3.288 ;
    END
  END rdata_out[33]
  PIN rdata_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.360 0.024 3.384 ;
    END
  END rdata_out[34]
  PIN rdata_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.456 0.024 3.480 ;
    END
  END rdata_out[35]
  PIN rdata_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.552 0.024 3.576 ;
    END
  END rdata_out[36]
  PIN rdata_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.648 0.024 3.672 ;
    END
  END rdata_out[37]
  PIN rdata_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.744 0.024 3.768 ;
    END
  END rdata_out[38]
  PIN rdata_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.840 0.024 3.864 ;
    END
  END rdata_out[39]
  PIN rdata_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.936 0.024 3.960 ;
    END
  END rdata_out[40]
  PIN rdata_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.032 0.024 4.056 ;
    END
  END rdata_out[41]
  PIN rdata_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.128 0.024 4.152 ;
    END
  END rdata_out[42]
  PIN rdata_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.224 0.024 4.248 ;
    END
  END rdata_out[43]
  PIN rdata_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.320 0.024 4.344 ;
    END
  END rdata_out[44]
  PIN rdata_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.416 0.024 4.440 ;
    END
  END rdata_out[45]
  PIN rdata_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.512 0.024 4.536 ;
    END
  END rdata_out[46]
  PIN rdata_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.608 0.024 4.632 ;
    END
  END rdata_out[47]
  PIN rdata_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.704 0.024 4.728 ;
    END
  END rdata_out[48]
  PIN rdata_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.800 0.024 4.824 ;
    END
  END rdata_out[49]
  PIN rdata_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.896 0.024 4.920 ;
    END
  END rdata_out[50]
  PIN rdata_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.992 0.024 5.016 ;
    END
  END rdata_out[51]
  PIN rdata_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.088 0.024 5.112 ;
    END
  END rdata_out[52]
  PIN rdata_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.184 0.024 5.208 ;
    END
  END rdata_out[53]
  PIN rdata_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.280 0.024 5.304 ;
    END
  END rdata_out[54]
  PIN rdata_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.376 0.024 5.400 ;
    END
  END rdata_out[55]
  PIN rdata_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.472 0.024 5.496 ;
    END
  END rdata_out[56]
  PIN rdata_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.568 0.024 5.592 ;
    END
  END rdata_out[57]
  PIN rdata_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.664 0.024 5.688 ;
    END
  END rdata_out[58]
  PIN rdata_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.760 0.024 5.784 ;
    END
  END rdata_out[59]
  PIN rdata_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.856 0.024 5.880 ;
    END
  END rdata_out[60]
  PIN rdata_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.952 0.024 5.976 ;
    END
  END rdata_out[61]
  PIN rdata_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.048 0.024 6.072 ;
    END
  END rdata_out[62]
  PIN rdata_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.144 0.024 6.168 ;
    END
  END rdata_out[63]
  PIN wdata_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.392 0.024 7.416 ;
    END
  END wdata_in[0]
  PIN wdata_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.488 0.024 7.512 ;
    END
  END wdata_in[1]
  PIN wdata_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.584 0.024 7.608 ;
    END
  END wdata_in[2]
  PIN wdata_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.680 0.024 7.704 ;
    END
  END wdata_in[3]
  PIN wdata_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.776 0.024 7.800 ;
    END
  END wdata_in[4]
  PIN wdata_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.872 0.024 7.896 ;
    END
  END wdata_in[5]
  PIN wdata_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.968 0.024 7.992 ;
    END
  END wdata_in[6]
  PIN wdata_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.064 0.024 8.088 ;
    END
  END wdata_in[7]
  PIN wdata_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.160 0.024 8.184 ;
    END
  END wdata_in[8]
  PIN wdata_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.256 0.024 8.280 ;
    END
  END wdata_in[9]
  PIN wdata_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.352 0.024 8.376 ;
    END
  END wdata_in[10]
  PIN wdata_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.448 0.024 8.472 ;
    END
  END wdata_in[11]
  PIN wdata_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.544 0.024 8.568 ;
    END
  END wdata_in[12]
  PIN wdata_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.640 0.024 8.664 ;
    END
  END wdata_in[13]
  PIN wdata_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.736 0.024 8.760 ;
    END
  END wdata_in[14]
  PIN wdata_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.832 0.024 8.856 ;
    END
  END wdata_in[15]
  PIN wdata_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.928 0.024 8.952 ;
    END
  END wdata_in[16]
  PIN wdata_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.024 0.024 9.048 ;
    END
  END wdata_in[17]
  PIN wdata_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.120 0.024 9.144 ;
    END
  END wdata_in[18]
  PIN wdata_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.216 0.024 9.240 ;
    END
  END wdata_in[19]
  PIN wdata_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.312 0.024 9.336 ;
    END
  END wdata_in[20]
  PIN wdata_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.408 0.024 9.432 ;
    END
  END wdata_in[21]
  PIN wdata_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.504 0.024 9.528 ;
    END
  END wdata_in[22]
  PIN wdata_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.600 0.024 9.624 ;
    END
  END wdata_in[23]
  PIN wdata_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.696 0.024 9.720 ;
    END
  END wdata_in[24]
  PIN wdata_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.792 0.024 9.816 ;
    END
  END wdata_in[25]
  PIN wdata_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.888 0.024 9.912 ;
    END
  END wdata_in[26]
  PIN wdata_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.984 0.024 10.008 ;
    END
  END wdata_in[27]
  PIN wdata_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.080 0.024 10.104 ;
    END
  END wdata_in[28]
  PIN wdata_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.176 0.024 10.200 ;
    END
  END wdata_in[29]
  PIN wdata_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.272 0.024 10.296 ;
    END
  END wdata_in[30]
  PIN wdata_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.368 0.024 10.392 ;
    END
  END wdata_in[31]
  PIN wdata_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.464 0.024 10.488 ;
    END
  END wdata_in[32]
  PIN wdata_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.560 0.024 10.584 ;
    END
  END wdata_in[33]
  PIN wdata_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.656 0.024 10.680 ;
    END
  END wdata_in[34]
  PIN wdata_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.752 0.024 10.776 ;
    END
  END wdata_in[35]
  PIN wdata_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.848 0.024 10.872 ;
    END
  END wdata_in[36]
  PIN wdata_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.944 0.024 10.968 ;
    END
  END wdata_in[37]
  PIN wdata_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.040 0.024 11.064 ;
    END
  END wdata_in[38]
  PIN wdata_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.136 0.024 11.160 ;
    END
  END wdata_in[39]
  PIN wdata_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.232 0.024 11.256 ;
    END
  END wdata_in[40]
  PIN wdata_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.328 0.024 11.352 ;
    END
  END wdata_in[41]
  PIN wdata_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.424 0.024 11.448 ;
    END
  END wdata_in[42]
  PIN wdata_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.520 0.024 11.544 ;
    END
  END wdata_in[43]
  PIN wdata_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.616 0.024 11.640 ;
    END
  END wdata_in[44]
  PIN wdata_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.712 0.024 11.736 ;
    END
  END wdata_in[45]
  PIN wdata_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.808 0.024 11.832 ;
    END
  END wdata_in[46]
  PIN wdata_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.904 0.024 11.928 ;
    END
  END wdata_in[47]
  PIN wdata_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.000 0.024 12.024 ;
    END
  END wdata_in[48]
  PIN wdata_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.096 0.024 12.120 ;
    END
  END wdata_in[49]
  PIN wdata_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.192 0.024 12.216 ;
    END
  END wdata_in[50]
  PIN wdata_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.288 0.024 12.312 ;
    END
  END wdata_in[51]
  PIN wdata_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.384 0.024 12.408 ;
    END
  END wdata_in[52]
  PIN wdata_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.480 0.024 12.504 ;
    END
  END wdata_in[53]
  PIN wdata_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.576 0.024 12.600 ;
    END
  END wdata_in[54]
  PIN wdata_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.672 0.024 12.696 ;
    END
  END wdata_in[55]
  PIN wdata_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.768 0.024 12.792 ;
    END
  END wdata_in[56]
  PIN wdata_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.864 0.024 12.888 ;
    END
  END wdata_in[57]
  PIN wdata_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.960 0.024 12.984 ;
    END
  END wdata_in[58]
  PIN wdata_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.056 0.024 13.080 ;
    END
  END wdata_in[59]
  PIN wdata_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.152 0.024 13.176 ;
    END
  END wdata_in[60]
  PIN wdata_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.248 0.024 13.272 ;
    END
  END wdata_in[61]
  PIN wdata_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.344 0.024 13.368 ;
    END
  END wdata_in[62]
  PIN wdata_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.440 0.024 13.464 ;
    END
  END wdata_in[63]
  PIN raddr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.688 0.024 14.712 ;
    END
  END raddr_in[0]
  PIN raddr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.784 0.024 14.808 ;
    END
  END raddr_in[1]
  PIN raddr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.880 0.024 14.904 ;
    END
  END raddr_in[2]
  PIN raddr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.976 0.024 15.000 ;
    END
  END raddr_in[3]
  PIN raddr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.072 0.024 15.096 ;
    END
  END raddr_in[4]
  PIN raddr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.168 0.024 15.192 ;
    END
  END raddr_in[5]
  PIN waddr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.416 0.024 16.440 ;
    END
  END waddr_in[0]
  PIN waddr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.512 0.024 16.536 ;
    END
  END waddr_in[1]
  PIN waddr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.608 0.024 16.632 ;
    END
  END waddr_in[2]
  PIN waddr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.704 0.024 16.728 ;
    END
  END waddr_in[3]
  PIN waddr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.800 0.024 16.824 ;
    END
  END waddr_in[4]
  PIN waddr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.896 0.024 16.920 ;
    END
  END waddr_in[5]
  PIN wmask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.144 0.024 18.168 ;
    END
  END wmask_in[0]
  PIN wmask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.240 0.024 18.264 ;
    END
  END wmask_in[1]
  PIN wmask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.336 0.024 18.360 ;
    END
  END wmask_in[2]
  PIN wmask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.432 0.024 18.456 ;
    END
  END wmask_in[3]
  PIN wmask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.528 0.024 18.552 ;
    END
  END wmask_in[4]
  PIN wmask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.624 0.024 18.648 ;
    END
  END wmask_in[5]
  PIN wmask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.720 0.024 18.744 ;
    END
  END wmask_in[6]
  PIN wmask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.816 0.024 18.840 ;
    END
  END wmask_in[7]
  PIN wmask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.912 0.024 18.936 ;
    END
  END wmask_in[8]
  PIN wmask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.008 0.024 19.032 ;
    END
  END wmask_in[9]
  PIN wmask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.104 0.024 19.128 ;
    END
  END wmask_in[10]
  PIN wmask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.200 0.024 19.224 ;
    END
  END wmask_in[11]
  PIN wmask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.296 0.024 19.320 ;
    END
  END wmask_in[12]
  PIN wmask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.392 0.024 19.416 ;
    END
  END wmask_in[13]
  PIN wmask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.488 0.024 19.512 ;
    END
  END wmask_in[14]
  PIN wmask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.584 0.024 19.608 ;
    END
  END wmask_in[15]
  PIN wmask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.680 0.024 19.704 ;
    END
  END wmask_in[16]
  PIN wmask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.776 0.024 19.800 ;
    END
  END wmask_in[17]
  PIN wmask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.872 0.024 19.896 ;
    END
  END wmask_in[18]
  PIN wmask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.968 0.024 19.992 ;
    END
  END wmask_in[19]
  PIN wmask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.064 0.024 20.088 ;
    END
  END wmask_in[20]
  PIN wmask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.160 0.024 20.184 ;
    END
  END wmask_in[21]
  PIN wmask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.256 0.024 20.280 ;
    END
  END wmask_in[22]
  PIN wmask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.352 0.024 20.376 ;
    END
  END wmask_in[23]
  PIN wmask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.448 0.024 20.472 ;
    END
  END wmask_in[24]
  PIN wmask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.544 0.024 20.568 ;
    END
  END wmask_in[25]
  PIN wmask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.640 0.024 20.664 ;
    END
  END wmask_in[26]
  PIN wmask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.736 0.024 20.760 ;
    END
  END wmask_in[27]
  PIN wmask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.832 0.024 20.856 ;
    END
  END wmask_in[28]
  PIN wmask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.928 0.024 20.952 ;
    END
  END wmask_in[29]
  PIN wmask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.024 0.024 21.048 ;
    END
  END wmask_in[30]
  PIN wmask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.120 0.024 21.144 ;
    END
  END wmask_in[31]
  PIN wmask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.216 0.024 21.240 ;
    END
  END wmask_in[32]
  PIN wmask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.312 0.024 21.336 ;
    END
  END wmask_in[33]
  PIN wmask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.408 0.024 21.432 ;
    END
  END wmask_in[34]
  PIN wmask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.504 0.024 21.528 ;
    END
  END wmask_in[35]
  PIN wmask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.600 0.024 21.624 ;
    END
  END wmask_in[36]
  PIN wmask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.696 0.024 21.720 ;
    END
  END wmask_in[37]
  PIN wmask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.792 0.024 21.816 ;
    END
  END wmask_in[38]
  PIN wmask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.888 0.024 21.912 ;
    END
  END wmask_in[39]
  PIN wmask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.984 0.024 22.008 ;
    END
  END wmask_in[40]
  PIN wmask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.080 0.024 22.104 ;
    END
  END wmask_in[41]
  PIN wmask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.176 0.024 22.200 ;
    END
  END wmask_in[42]
  PIN wmask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.272 0.024 22.296 ;
    END
  END wmask_in[43]
  PIN wmask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.368 0.024 22.392 ;
    END
  END wmask_in[44]
  PIN wmask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.464 0.024 22.488 ;
    END
  END wmask_in[45]
  PIN wmask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.560 0.024 22.584 ;
    END
  END wmask_in[46]
  PIN wmask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.656 0.024 22.680 ;
    END
  END wmask_in[47]
  PIN wmask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.752 0.024 22.776 ;
    END
  END wmask_in[48]
  PIN wmask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.848 0.024 22.872 ;
    END
  END wmask_in[49]
  PIN wmask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.944 0.024 22.968 ;
    END
  END wmask_in[50]
  PIN wmask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.040 0.024 23.064 ;
    END
  END wmask_in[51]
  PIN wmask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.136 0.024 23.160 ;
    END
  END wmask_in[52]
  PIN wmask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.232 0.024 23.256 ;
    END
  END wmask_in[53]
  PIN wmask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.328 0.024 23.352 ;
    END
  END wmask_in[54]
  PIN wmask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.424 0.024 23.448 ;
    END
  END wmask_in[55]
  PIN wmask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.520 0.024 23.544 ;
    END
  END wmask_in[56]
  PIN wmask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.616 0.024 23.640 ;
    END
  END wmask_in[57]
  PIN wmask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.712 0.024 23.736 ;
    END
  END wmask_in[58]
  PIN wmask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.808 0.024 23.832 ;
    END
  END wmask_in[59]
  PIN wmask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.904 0.024 23.928 ;
    END
  END wmask_in[60]
  PIN wmask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.000 0.024 24.024 ;
    END
  END wmask_in[61]
  PIN wmask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.096 0.024 24.120 ;
    END
  END wmask_in[62]
  PIN wmask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.192 0.024 24.216 ;
    END
  END wmask_in[63]
  PIN wen_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.440 0.024 25.464 ;
    END
  END wen_in
  PIN ren_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.536 0.024 25.560 ;
    END
  END ren_in
  PIN wclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.632 0.024 25.656 ;
    END
  END wclk
  PIN rclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.728 0.024 25.752 ;
    END
  END rclk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.096 0.048 8.264 0.144 ;
      RECT 0.096 1.584 8.264 1.680 ;
      RECT 0.096 3.120 8.264 3.216 ;
      RECT 0.096 4.656 8.264 4.752 ;
      RECT 0.096 6.192 8.264 6.288 ;
      RECT 0.096 7.728 8.264 7.824 ;
      RECT 0.096 9.264 8.264 9.360 ;
      RECT 0.096 10.800 8.264 10.896 ;
      RECT 0.096 12.336 8.264 12.432 ;
      RECT 0.096 13.872 8.264 13.968 ;
      RECT 0.096 15.408 8.264 15.504 ;
      RECT 0.096 16.944 8.264 17.040 ;
      RECT 0.096 18.480 8.264 18.576 ;
      RECT 0.096 20.016 8.264 20.112 ;
      RECT 0.096 21.552 8.264 21.648 ;
      RECT 0.096 23.088 8.264 23.184 ;
      RECT 0.096 24.624 8.264 24.720 ;
      RECT 0.096 26.160 8.264 26.256 ;
      RECT 0.096 27.696 8.264 27.792 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.096 0.816 8.264 0.912 ;
      RECT 0.096 2.352 8.264 2.448 ;
      RECT 0.096 3.888 8.264 3.984 ;
      RECT 0.096 5.424 8.264 5.520 ;
      RECT 0.096 6.960 8.264 7.056 ;
      RECT 0.096 8.496 8.264 8.592 ;
      RECT 0.096 10.032 8.264 10.128 ;
      RECT 0.096 11.568 8.264 11.664 ;
      RECT 0.096 13.104 8.264 13.200 ;
      RECT 0.096 14.640 8.264 14.736 ;
      RECT 0.096 16.176 8.264 16.272 ;
      RECT 0.096 17.712 8.264 17.808 ;
      RECT 0.096 19.248 8.264 19.344 ;
      RECT 0.096 20.784 8.264 20.880 ;
      RECT 0.096 22.320 8.264 22.416 ;
      RECT 0.096 23.856 8.264 23.952 ;
      RECT 0.096 25.392 8.264 25.488 ;
      RECT 0.096 26.928 8.264 27.024 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 8.360 28.000 ;
    LAYER M2 ;
    RECT 0 0 8.360 28.000 ;
    LAYER M3 ;
    RECT 0 0 8.360 28.000 ;
    LAYER M4 ;
    RECT 0.1 0 8.260 28.000 ;
  END
END fakeregfile_64x64

END LIBRARY
