../../nangate45/lef/fakeram45_64x7.lef