module MuxTest_width_1_inputs_1_outputs_16_pipeline_0( // @[:@3.2]
  input        clock, // @[:@4.4]
  input        reset, // @[:@5.4]
  input  [2:0] io_operation_0, // @[:@6.4]
  input  [2:0] io_operation_1, // @[:@6.4]
  input  [2:0] io_operation_2, // @[:@6.4]
  input  [2:0] io_operation_3, // @[:@6.4]
  input  [2:0] io_operation_4, // @[:@6.4]
  input  [2:0] io_operation_5, // @[:@6.4]
  input  [2:0] io_operation_6, // @[:@6.4]
  input  [2:0] io_operation_7, // @[:@6.4]
  input  [2:0] io_operation_8, // @[:@6.4]
  input  [2:0] io_operation_9, // @[:@6.4]
  input  [2:0] io_operation_10, // @[:@6.4]
  input  [2:0] io_operation_11, // @[:@6.4]
  input  [2:0] io_operation_12, // @[:@6.4]
  input  [2:0] io_operation_13, // @[:@6.4]
  input  [2:0] io_operation_14, // @[:@6.4]
  input  [2:0] io_operation_15, // @[:@6.4]
  input        io_inputs_0, // @[:@6.4]
  output       io_outputs_0, // @[:@6.4]
  output       io_outputs_1, // @[:@6.4]
  output       io_outputs_2, // @[:@6.4]
  output       io_outputs_3, // @[:@6.4]
  output       io_outputs_4, // @[:@6.4]
  output       io_outputs_5, // @[:@6.4]
  output       io_outputs_6, // @[:@6.4]
  output       io_outputs_7, // @[:@6.4]
  output       io_outputs_8, // @[:@6.4]
  output       io_outputs_9, // @[:@6.4]
  output       io_outputs_10, // @[:@6.4]
  output       io_outputs_11, // @[:@6.4]
  output       io_outputs_12, // @[:@6.4]
  output       io_outputs_13, // @[:@6.4]
  output       io_outputs_14, // @[:@6.4]
  output       io_outputs_15 // @[:@6.4]
);
  wire [1:0] _T_724; // @[MuxTest_width_1_inputs_1_outputs_16_pipeline_0s.scala 32:53:@8.4]
  wire  _T_725; // @[MuxTest_width_1_inputs_1_outputs_16_pipeline_0s.scala 32:53:@9.4]
  wire [1:0] _T_727; // @[MuxTest_width_1_inputs_1_outputs_16_pipeline_0s.scala 33:58:@10.4]
  wire  _T_729; // @[MuxTest_width_1_inputs_1_outputs_16_pipeline_0s.scala 34:56:@11.4]
  wire  _T_730; // @[Mux.scala 46:19:@12.4]
  wire  _T_731; // @[Mux.scala 46:16:@13.4]
  wire  _T_732; // @[Mux.scala 46:19:@14.4]
  wire [1:0] _T_733; // @[Mux.scala 46:16:@15.4]
  wire  _T_734; // @[Mux.scala 46:19:@16.4]
  wire [1:0] _T_735; // @[Mux.scala 46:16:@17.4]
  wire  _T_736; // @[Mux.scala 46:19:@18.4]
  wire [1:0] _T_737; // @[Mux.scala 46:16:@19.4]
  wire  _T_747; // @[Mux.scala 46:19:@24.4]
  wire  _T_748; // @[Mux.scala 46:16:@25.4]
  wire  _T_749; // @[Mux.scala 46:19:@26.4]
  wire [1:0] _T_750; // @[Mux.scala 46:16:@27.4]
  wire  _T_751; // @[Mux.scala 46:19:@28.4]
  wire [1:0] _T_752; // @[Mux.scala 46:16:@29.4]
  wire  _T_753; // @[Mux.scala 46:19:@30.4]
  wire [1:0] _T_754; // @[Mux.scala 46:16:@31.4]
  wire  _T_764; // @[Mux.scala 46:19:@36.4]
  wire  _T_765; // @[Mux.scala 46:16:@37.4]
  wire  _T_766; // @[Mux.scala 46:19:@38.4]
  wire [1:0] _T_767; // @[Mux.scala 46:16:@39.4]
  wire  _T_768; // @[Mux.scala 46:19:@40.4]
  wire [1:0] _T_769; // @[Mux.scala 46:16:@41.4]
  wire  _T_770; // @[Mux.scala 46:19:@42.4]
  wire [1:0] _T_771; // @[Mux.scala 46:16:@43.4]
  wire  _T_781; // @[Mux.scala 46:19:@48.4]
  wire  _T_782; // @[Mux.scala 46:16:@49.4]
  wire  _T_783; // @[Mux.scala 46:19:@50.4]
  wire [1:0] _T_784; // @[Mux.scala 46:16:@51.4]
  wire  _T_785; // @[Mux.scala 46:19:@52.4]
  wire [1:0] _T_786; // @[Mux.scala 46:16:@53.4]
  wire  _T_787; // @[Mux.scala 46:19:@54.4]
  wire [1:0] _T_788; // @[Mux.scala 46:16:@55.4]
  wire  _T_798; // @[Mux.scala 46:19:@60.4]
  wire  _T_799; // @[Mux.scala 46:16:@61.4]
  wire  _T_800; // @[Mux.scala 46:19:@62.4]
  wire [1:0] _T_801; // @[Mux.scala 46:16:@63.4]
  wire  _T_802; // @[Mux.scala 46:19:@64.4]
  wire [1:0] _T_803; // @[Mux.scala 46:16:@65.4]
  wire  _T_804; // @[Mux.scala 46:19:@66.4]
  wire [1:0] _T_805; // @[Mux.scala 46:16:@67.4]
  wire  _T_815; // @[Mux.scala 46:19:@72.4]
  wire  _T_816; // @[Mux.scala 46:16:@73.4]
  wire  _T_817; // @[Mux.scala 46:19:@74.4]
  wire [1:0] _T_818; // @[Mux.scala 46:16:@75.4]
  wire  _T_819; // @[Mux.scala 46:19:@76.4]
  wire [1:0] _T_820; // @[Mux.scala 46:16:@77.4]
  wire  _T_821; // @[Mux.scala 46:19:@78.4]
  wire [1:0] _T_822; // @[Mux.scala 46:16:@79.4]
  wire  _T_832; // @[Mux.scala 46:19:@84.4]
  wire  _T_833; // @[Mux.scala 46:16:@85.4]
  wire  _T_834; // @[Mux.scala 46:19:@86.4]
  wire [1:0] _T_835; // @[Mux.scala 46:16:@87.4]
  wire  _T_836; // @[Mux.scala 46:19:@88.4]
  wire [1:0] _T_837; // @[Mux.scala 46:16:@89.4]
  wire  _T_838; // @[Mux.scala 46:19:@90.4]
  wire [1:0] _T_839; // @[Mux.scala 46:16:@91.4]
  wire  _T_849; // @[Mux.scala 46:19:@96.4]
  wire  _T_850; // @[Mux.scala 46:16:@97.4]
  wire  _T_851; // @[Mux.scala 46:19:@98.4]
  wire [1:0] _T_852; // @[Mux.scala 46:16:@99.4]
  wire  _T_853; // @[Mux.scala 46:19:@100.4]
  wire [1:0] _T_854; // @[Mux.scala 46:16:@101.4]
  wire  _T_855; // @[Mux.scala 46:19:@102.4]
  wire [1:0] _T_856; // @[Mux.scala 46:16:@103.4]
  wire  _T_866; // @[Mux.scala 46:19:@108.4]
  wire  _T_867; // @[Mux.scala 46:16:@109.4]
  wire  _T_868; // @[Mux.scala 46:19:@110.4]
  wire [1:0] _T_869; // @[Mux.scala 46:16:@111.4]
  wire  _T_870; // @[Mux.scala 46:19:@112.4]
  wire [1:0] _T_871; // @[Mux.scala 46:16:@113.4]
  wire  _T_872; // @[Mux.scala 46:19:@114.4]
  wire [1:0] _T_873; // @[Mux.scala 46:16:@115.4]
  wire  _T_883; // @[Mux.scala 46:19:@120.4]
  wire  _T_884; // @[Mux.scala 46:16:@121.4]
  wire  _T_885; // @[Mux.scala 46:19:@122.4]
  wire [1:0] _T_886; // @[Mux.scala 46:16:@123.4]
  wire  _T_887; // @[Mux.scala 46:19:@124.4]
  wire [1:0] _T_888; // @[Mux.scala 46:16:@125.4]
  wire  _T_889; // @[Mux.scala 46:19:@126.4]
  wire [1:0] _T_890; // @[Mux.scala 46:16:@127.4]
  wire  _T_900; // @[Mux.scala 46:19:@132.4]
  wire  _T_901; // @[Mux.scala 46:16:@133.4]
  wire  _T_902; // @[Mux.scala 46:19:@134.4]
  wire [1:0] _T_903; // @[Mux.scala 46:16:@135.4]
  wire  _T_904; // @[Mux.scala 46:19:@136.4]
  wire [1:0] _T_905; // @[Mux.scala 46:16:@137.4]
  wire  _T_906; // @[Mux.scala 46:19:@138.4]
  wire [1:0] _T_907; // @[Mux.scala 46:16:@139.4]
  wire  _T_917; // @[Mux.scala 46:19:@144.4]
  wire  _T_918; // @[Mux.scala 46:16:@145.4]
  wire  _T_919; // @[Mux.scala 46:19:@146.4]
  wire [1:0] _T_920; // @[Mux.scala 46:16:@147.4]
  wire  _T_921; // @[Mux.scala 46:19:@148.4]
  wire [1:0] _T_922; // @[Mux.scala 46:16:@149.4]
  wire  _T_923; // @[Mux.scala 46:19:@150.4]
  wire [1:0] _T_924; // @[Mux.scala 46:16:@151.4]
  wire  _T_934; // @[Mux.scala 46:19:@156.4]
  wire  _T_935; // @[Mux.scala 46:16:@157.4]
  wire  _T_936; // @[Mux.scala 46:19:@158.4]
  wire [1:0] _T_937; // @[Mux.scala 46:16:@159.4]
  wire  _T_938; // @[Mux.scala 46:19:@160.4]
  wire [1:0] _T_939; // @[Mux.scala 46:16:@161.4]
  wire  _T_940; // @[Mux.scala 46:19:@162.4]
  wire [1:0] _T_941; // @[Mux.scala 46:16:@163.4]
  wire  _T_951; // @[Mux.scala 46:19:@168.4]
  wire  _T_952; // @[Mux.scala 46:16:@169.4]
  wire  _T_953; // @[Mux.scala 46:19:@170.4]
  wire [1:0] _T_954; // @[Mux.scala 46:16:@171.4]
  wire  _T_955; // @[Mux.scala 46:19:@172.4]
  wire [1:0] _T_956; // @[Mux.scala 46:16:@173.4]
  wire  _T_957; // @[Mux.scala 46:19:@174.4]
  wire [1:0] _T_958; // @[Mux.scala 46:16:@175.4]
  wire  _T_968; // @[Mux.scala 46:19:@180.4]
  wire  _T_969; // @[Mux.scala 46:16:@181.4]
  wire  _T_970; // @[Mux.scala 46:19:@182.4]
  wire [1:0] _T_971; // @[Mux.scala 46:16:@183.4]
  wire  _T_972; // @[Mux.scala 46:19:@184.4]
  wire [1:0] _T_973; // @[Mux.scala 46:16:@185.4]
  wire  _T_974; // @[Mux.scala 46:19:@186.4]
  wire [1:0] _T_975; // @[Mux.scala 46:16:@187.4]
  wire  _T_985; // @[Mux.scala 46:19:@192.4]
  wire  _T_986; // @[Mux.scala 46:16:@193.4]
  wire  _T_987; // @[Mux.scala 46:19:@194.4]
  wire [1:0] _T_988; // @[Mux.scala 46:16:@195.4]
  wire  _T_989; // @[Mux.scala 46:19:@196.4]
  wire [1:0] _T_990; // @[Mux.scala 46:16:@197.4]
  wire  _T_991; // @[Mux.scala 46:19:@198.4]
  wire [1:0] _T_992; // @[Mux.scala 46:16:@199.4]
  assign _T_724 = io_inputs_0 + io_inputs_0; // @[MuxTest_width_1_inputs_1_outputs_16_pipeline_0s.scala 32:53:@8.4]
  assign _T_725 = io_inputs_0 + io_inputs_0; // @[MuxTest_width_1_inputs_1_outputs_16_pipeline_0s.scala 32:53:@9.4]
  assign _T_727 = io_inputs_0 * io_inputs_0; // @[MuxTest_width_1_inputs_1_outputs_16_pipeline_0s.scala 33:58:@10.4]
  assign _T_729 = io_inputs_0 / io_inputs_0; // @[MuxTest_width_1_inputs_1_outputs_16_pipeline_0s.scala 34:56:@11.4]
  assign _T_730 = 3'h3 == io_operation_0; // @[Mux.scala 46:19:@12.4]
  assign _T_731 = _T_730 ? _T_729 : 1'h0; // @[Mux.scala 46:16:@13.4]
  assign _T_732 = 3'h2 == io_operation_0; // @[Mux.scala 46:19:@14.4]
  assign _T_733 = _T_732 ? _T_727 : {{1'd0}, _T_731}; // @[Mux.scala 46:16:@15.4]
  assign _T_734 = 3'h1 == io_operation_0; // @[Mux.scala 46:19:@16.4]
  assign _T_735 = _T_734 ? {{1'd0}, _T_725} : _T_733; // @[Mux.scala 46:16:@17.4]
  assign _T_736 = 3'h0 == io_operation_0; // @[Mux.scala 46:19:@18.4]
  assign _T_737 = _T_736 ? {{1'd0}, io_inputs_0} : _T_735; // @[Mux.scala 46:16:@19.4]
  assign _T_747 = 3'h3 == io_operation_1; // @[Mux.scala 46:19:@24.4]
  assign _T_748 = _T_747 ? _T_729 : 1'h0; // @[Mux.scala 46:16:@25.4]
  assign _T_749 = 3'h2 == io_operation_1; // @[Mux.scala 46:19:@26.4]
  assign _T_750 = _T_749 ? _T_727 : {{1'd0}, _T_748}; // @[Mux.scala 46:16:@27.4]
  assign _T_751 = 3'h1 == io_operation_1; // @[Mux.scala 46:19:@28.4]
  assign _T_752 = _T_751 ? {{1'd0}, _T_725} : _T_750; // @[Mux.scala 46:16:@29.4]
  assign _T_753 = 3'h0 == io_operation_1; // @[Mux.scala 46:19:@30.4]
  assign _T_754 = _T_753 ? {{1'd0}, io_inputs_0} : _T_752; // @[Mux.scala 46:16:@31.4]
  assign _T_764 = 3'h3 == io_operation_2; // @[Mux.scala 46:19:@36.4]
  assign _T_765 = _T_764 ? _T_729 : 1'h0; // @[Mux.scala 46:16:@37.4]
  assign _T_766 = 3'h2 == io_operation_2; // @[Mux.scala 46:19:@38.4]
  assign _T_767 = _T_766 ? _T_727 : {{1'd0}, _T_765}; // @[Mux.scala 46:16:@39.4]
  assign _T_768 = 3'h1 == io_operation_2; // @[Mux.scala 46:19:@40.4]
  assign _T_769 = _T_768 ? {{1'd0}, _T_725} : _T_767; // @[Mux.scala 46:16:@41.4]
  assign _T_770 = 3'h0 == io_operation_2; // @[Mux.scala 46:19:@42.4]
  assign _T_771 = _T_770 ? {{1'd0}, io_inputs_0} : _T_769; // @[Mux.scala 46:16:@43.4]
  assign _T_781 = 3'h3 == io_operation_3; // @[Mux.scala 46:19:@48.4]
  assign _T_782 = _T_781 ? _T_729 : 1'h0; // @[Mux.scala 46:16:@49.4]
  assign _T_783 = 3'h2 == io_operation_3; // @[Mux.scala 46:19:@50.4]
  assign _T_784 = _T_783 ? _T_727 : {{1'd0}, _T_782}; // @[Mux.scala 46:16:@51.4]
  assign _T_785 = 3'h1 == io_operation_3; // @[Mux.scala 46:19:@52.4]
  assign _T_786 = _T_785 ? {{1'd0}, _T_725} : _T_784; // @[Mux.scala 46:16:@53.4]
  assign _T_787 = 3'h0 == io_operation_3; // @[Mux.scala 46:19:@54.4]
  assign _T_788 = _T_787 ? {{1'd0}, io_inputs_0} : _T_786; // @[Mux.scala 46:16:@55.4]
  assign _T_798 = 3'h3 == io_operation_4; // @[Mux.scala 46:19:@60.4]
  assign _T_799 = _T_798 ? _T_729 : 1'h0; // @[Mux.scala 46:16:@61.4]
  assign _T_800 = 3'h2 == io_operation_4; // @[Mux.scala 46:19:@62.4]
  assign _T_801 = _T_800 ? _T_727 : {{1'd0}, _T_799}; // @[Mux.scala 46:16:@63.4]
  assign _T_802 = 3'h1 == io_operation_4; // @[Mux.scala 46:19:@64.4]
  assign _T_803 = _T_802 ? {{1'd0}, _T_725} : _T_801; // @[Mux.scala 46:16:@65.4]
  assign _T_804 = 3'h0 == io_operation_4; // @[Mux.scala 46:19:@66.4]
  assign _T_805 = _T_804 ? {{1'd0}, io_inputs_0} : _T_803; // @[Mux.scala 46:16:@67.4]
  assign _T_815 = 3'h3 == io_operation_5; // @[Mux.scala 46:19:@72.4]
  assign _T_816 = _T_815 ? _T_729 : 1'h0; // @[Mux.scala 46:16:@73.4]
  assign _T_817 = 3'h2 == io_operation_5; // @[Mux.scala 46:19:@74.4]
  assign _T_818 = _T_817 ? _T_727 : {{1'd0}, _T_816}; // @[Mux.scala 46:16:@75.4]
  assign _T_819 = 3'h1 == io_operation_5; // @[Mux.scala 46:19:@76.4]
  assign _T_820 = _T_819 ? {{1'd0}, _T_725} : _T_818; // @[Mux.scala 46:16:@77.4]
  assign _T_821 = 3'h0 == io_operation_5; // @[Mux.scala 46:19:@78.4]
  assign _T_822 = _T_821 ? {{1'd0}, io_inputs_0} : _T_820; // @[Mux.scala 46:16:@79.4]
  assign _T_832 = 3'h3 == io_operation_6; // @[Mux.scala 46:19:@84.4]
  assign _T_833 = _T_832 ? _T_729 : 1'h0; // @[Mux.scala 46:16:@85.4]
  assign _T_834 = 3'h2 == io_operation_6; // @[Mux.scala 46:19:@86.4]
  assign _T_835 = _T_834 ? _T_727 : {{1'd0}, _T_833}; // @[Mux.scala 46:16:@87.4]
  assign _T_836 = 3'h1 == io_operation_6; // @[Mux.scala 46:19:@88.4]
  assign _T_837 = _T_836 ? {{1'd0}, _T_725} : _T_835; // @[Mux.scala 46:16:@89.4]
  assign _T_838 = 3'h0 == io_operation_6; // @[Mux.scala 46:19:@90.4]
  assign _T_839 = _T_838 ? {{1'd0}, io_inputs_0} : _T_837; // @[Mux.scala 46:16:@91.4]
  assign _T_849 = 3'h3 == io_operation_7; // @[Mux.scala 46:19:@96.4]
  assign _T_850 = _T_849 ? _T_729 : 1'h0; // @[Mux.scala 46:16:@97.4]
  assign _T_851 = 3'h2 == io_operation_7; // @[Mux.scala 46:19:@98.4]
  assign _T_852 = _T_851 ? _T_727 : {{1'd0}, _T_850}; // @[Mux.scala 46:16:@99.4]
  assign _T_853 = 3'h1 == io_operation_7; // @[Mux.scala 46:19:@100.4]
  assign _T_854 = _T_853 ? {{1'd0}, _T_725} : _T_852; // @[Mux.scala 46:16:@101.4]
  assign _T_855 = 3'h0 == io_operation_7; // @[Mux.scala 46:19:@102.4]
  assign _T_856 = _T_855 ? {{1'd0}, io_inputs_0} : _T_854; // @[Mux.scala 46:16:@103.4]
  assign _T_866 = 3'h3 == io_operation_8; // @[Mux.scala 46:19:@108.4]
  assign _T_867 = _T_866 ? _T_729 : 1'h0; // @[Mux.scala 46:16:@109.4]
  assign _T_868 = 3'h2 == io_operation_8; // @[Mux.scala 46:19:@110.4]
  assign _T_869 = _T_868 ? _T_727 : {{1'd0}, _T_867}; // @[Mux.scala 46:16:@111.4]
  assign _T_870 = 3'h1 == io_operation_8; // @[Mux.scala 46:19:@112.4]
  assign _T_871 = _T_870 ? {{1'd0}, _T_725} : _T_869; // @[Mux.scala 46:16:@113.4]
  assign _T_872 = 3'h0 == io_operation_8; // @[Mux.scala 46:19:@114.4]
  assign _T_873 = _T_872 ? {{1'd0}, io_inputs_0} : _T_871; // @[Mux.scala 46:16:@115.4]
  assign _T_883 = 3'h3 == io_operation_9; // @[Mux.scala 46:19:@120.4]
  assign _T_884 = _T_883 ? _T_729 : 1'h0; // @[Mux.scala 46:16:@121.4]
  assign _T_885 = 3'h2 == io_operation_9; // @[Mux.scala 46:19:@122.4]
  assign _T_886 = _T_885 ? _T_727 : {{1'd0}, _T_884}; // @[Mux.scala 46:16:@123.4]
  assign _T_887 = 3'h1 == io_operation_9; // @[Mux.scala 46:19:@124.4]
  assign _T_888 = _T_887 ? {{1'd0}, _T_725} : _T_886; // @[Mux.scala 46:16:@125.4]
  assign _T_889 = 3'h0 == io_operation_9; // @[Mux.scala 46:19:@126.4]
  assign _T_890 = _T_889 ? {{1'd0}, io_inputs_0} : _T_888; // @[Mux.scala 46:16:@127.4]
  assign _T_900 = 3'h3 == io_operation_10; // @[Mux.scala 46:19:@132.4]
  assign _T_901 = _T_900 ? _T_729 : 1'h0; // @[Mux.scala 46:16:@133.4]
  assign _T_902 = 3'h2 == io_operation_10; // @[Mux.scala 46:19:@134.4]
  assign _T_903 = _T_902 ? _T_727 : {{1'd0}, _T_901}; // @[Mux.scala 46:16:@135.4]
  assign _T_904 = 3'h1 == io_operation_10; // @[Mux.scala 46:19:@136.4]
  assign _T_905 = _T_904 ? {{1'd0}, _T_725} : _T_903; // @[Mux.scala 46:16:@137.4]
  assign _T_906 = 3'h0 == io_operation_10; // @[Mux.scala 46:19:@138.4]
  assign _T_907 = _T_906 ? {{1'd0}, io_inputs_0} : _T_905; // @[Mux.scala 46:16:@139.4]
  assign _T_917 = 3'h3 == io_operation_11; // @[Mux.scala 46:19:@144.4]
  assign _T_918 = _T_917 ? _T_729 : 1'h0; // @[Mux.scala 46:16:@145.4]
  assign _T_919 = 3'h2 == io_operation_11; // @[Mux.scala 46:19:@146.4]
  assign _T_920 = _T_919 ? _T_727 : {{1'd0}, _T_918}; // @[Mux.scala 46:16:@147.4]
  assign _T_921 = 3'h1 == io_operation_11; // @[Mux.scala 46:19:@148.4]
  assign _T_922 = _T_921 ? {{1'd0}, _T_725} : _T_920; // @[Mux.scala 46:16:@149.4]
  assign _T_923 = 3'h0 == io_operation_11; // @[Mux.scala 46:19:@150.4]
  assign _T_924 = _T_923 ? {{1'd0}, io_inputs_0} : _T_922; // @[Mux.scala 46:16:@151.4]
  assign _T_934 = 3'h3 == io_operation_12; // @[Mux.scala 46:19:@156.4]
  assign _T_935 = _T_934 ? _T_729 : 1'h0; // @[Mux.scala 46:16:@157.4]
  assign _T_936 = 3'h2 == io_operation_12; // @[Mux.scala 46:19:@158.4]
  assign _T_937 = _T_936 ? _T_727 : {{1'd0}, _T_935}; // @[Mux.scala 46:16:@159.4]
  assign _T_938 = 3'h1 == io_operation_12; // @[Mux.scala 46:19:@160.4]
  assign _T_939 = _T_938 ? {{1'd0}, _T_725} : _T_937; // @[Mux.scala 46:16:@161.4]
  assign _T_940 = 3'h0 == io_operation_12; // @[Mux.scala 46:19:@162.4]
  assign _T_941 = _T_940 ? {{1'd0}, io_inputs_0} : _T_939; // @[Mux.scala 46:16:@163.4]
  assign _T_951 = 3'h3 == io_operation_13; // @[Mux.scala 46:19:@168.4]
  assign _T_952 = _T_951 ? _T_729 : 1'h0; // @[Mux.scala 46:16:@169.4]
  assign _T_953 = 3'h2 == io_operation_13; // @[Mux.scala 46:19:@170.4]
  assign _T_954 = _T_953 ? _T_727 : {{1'd0}, _T_952}; // @[Mux.scala 46:16:@171.4]
  assign _T_955 = 3'h1 == io_operation_13; // @[Mux.scala 46:19:@172.4]
  assign _T_956 = _T_955 ? {{1'd0}, _T_725} : _T_954; // @[Mux.scala 46:16:@173.4]
  assign _T_957 = 3'h0 == io_operation_13; // @[Mux.scala 46:19:@174.4]
  assign _T_958 = _T_957 ? {{1'd0}, io_inputs_0} : _T_956; // @[Mux.scala 46:16:@175.4]
  assign _T_968 = 3'h3 == io_operation_14; // @[Mux.scala 46:19:@180.4]
  assign _T_969 = _T_968 ? _T_729 : 1'h0; // @[Mux.scala 46:16:@181.4]
  assign _T_970 = 3'h2 == io_operation_14; // @[Mux.scala 46:19:@182.4]
  assign _T_971 = _T_970 ? _T_727 : {{1'd0}, _T_969}; // @[Mux.scala 46:16:@183.4]
  assign _T_972 = 3'h1 == io_operation_14; // @[Mux.scala 46:19:@184.4]
  assign _T_973 = _T_972 ? {{1'd0}, _T_725} : _T_971; // @[Mux.scala 46:16:@185.4]
  assign _T_974 = 3'h0 == io_operation_14; // @[Mux.scala 46:19:@186.4]
  assign _T_975 = _T_974 ? {{1'd0}, io_inputs_0} : _T_973; // @[Mux.scala 46:16:@187.4]
  assign _T_985 = 3'h3 == io_operation_15; // @[Mux.scala 46:19:@192.4]
  assign _T_986 = _T_985 ? _T_729 : 1'h0; // @[Mux.scala 46:16:@193.4]
  assign _T_987 = 3'h2 == io_operation_15; // @[Mux.scala 46:19:@194.4]
  assign _T_988 = _T_987 ? _T_727 : {{1'd0}, _T_986}; // @[Mux.scala 46:16:@195.4]
  assign _T_989 = 3'h1 == io_operation_15; // @[Mux.scala 46:19:@196.4]
  assign _T_990 = _T_989 ? {{1'd0}, _T_725} : _T_988; // @[Mux.scala 46:16:@197.4]
  assign _T_991 = 3'h0 == io_operation_15; // @[Mux.scala 46:19:@198.4]
  assign _T_992 = _T_991 ? {{1'd0}, io_inputs_0} : _T_990; // @[Mux.scala 46:16:@199.4]
  assign io_outputs_0 = _T_737[0]; // @[MuxTest_width_1_inputs_1_outputs_16_pipeline_0s.scala 23:14:@200.4]
  assign io_outputs_1 = _T_754[0]; // @[MuxTest_width_1_inputs_1_outputs_16_pipeline_0s.scala 23:14:@201.4]
  assign io_outputs_2 = _T_771[0]; // @[MuxTest_width_1_inputs_1_outputs_16_pipeline_0s.scala 23:14:@202.4]
  assign io_outputs_3 = _T_788[0]; // @[MuxTest_width_1_inputs_1_outputs_16_pipeline_0s.scala 23:14:@203.4]
  assign io_outputs_4 = _T_805[0]; // @[MuxTest_width_1_inputs_1_outputs_16_pipeline_0s.scala 23:14:@204.4]
  assign io_outputs_5 = _T_822[0]; // @[MuxTest_width_1_inputs_1_outputs_16_pipeline_0s.scala 23:14:@205.4]
  assign io_outputs_6 = _T_839[0]; // @[MuxTest_width_1_inputs_1_outputs_16_pipeline_0s.scala 23:14:@206.4]
  assign io_outputs_7 = _T_856[0]; // @[MuxTest_width_1_inputs_1_outputs_16_pipeline_0s.scala 23:14:@207.4]
  assign io_outputs_8 = _T_873[0]; // @[MuxTest_width_1_inputs_1_outputs_16_pipeline_0s.scala 23:14:@208.4]
  assign io_outputs_9 = _T_890[0]; // @[MuxTest_width_1_inputs_1_outputs_16_pipeline_0s.scala 23:14:@209.4]
  assign io_outputs_10 = _T_907[0]; // @[MuxTest_width_1_inputs_1_outputs_16_pipeline_0s.scala 23:14:@210.4]
  assign io_outputs_11 = _T_924[0]; // @[MuxTest_width_1_inputs_1_outputs_16_pipeline_0s.scala 23:14:@211.4]
  assign io_outputs_12 = _T_941[0]; // @[MuxTest_width_1_inputs_1_outputs_16_pipeline_0s.scala 23:14:@212.4]
  assign io_outputs_13 = _T_958[0]; // @[MuxTest_width_1_inputs_1_outputs_16_pipeline_0s.scala 23:14:@213.4]
  assign io_outputs_14 = _T_975[0]; // @[MuxTest_width_1_inputs_1_outputs_16_pipeline_0s.scala 23:14:@214.4]
  assign io_outputs_15 = _T_992[0]; // @[MuxTest_width_1_inputs_1_outputs_16_pipeline_0s.scala 23:14:@215.4]
endmodule
