module MockArray(
  input           clock,
  input           reset,
  input  [1023:0] io_insHorizontal_0_0,
  input  [1023:0] io_insHorizontal_0_1,
  input  [1023:0] io_insHorizontal_0_2,
  input  [1023:0] io_insHorizontal_0_3,
  input  [1023:0] io_insHorizontal_1_0,
  input  [1023:0] io_insHorizontal_1_1,
  input  [1023:0] io_insHorizontal_1_2,
  input  [1023:0] io_insHorizontal_1_3,
  output [1023:0] io_outsHorizontal_0_0,
  output [1023:0] io_outsHorizontal_0_1,
  output [1023:0] io_outsHorizontal_0_2,
  output [1023:0] io_outsHorizontal_0_3,
  output [1023:0] io_outsHorizontal_1_0,
  output [1023:0] io_outsHorizontal_1_1,
  output [1023:0] io_outsHorizontal_1_2,
  output [1023:0] io_outsHorizontal_1_3,
  input  [1023:0] io_insVertical_0_0,
  input  [1023:0] io_insVertical_0_1,
  input  [1023:0] io_insVertical_0_2,
  input  [1023:0] io_insVertical_0_3,
  input  [1023:0] io_insVertical_1_0,
  input  [1023:0] io_insVertical_1_1,
  input  [1023:0] io_insVertical_1_2,
  input  [1023:0] io_insVertical_1_3,
  output [1023:0] io_outsVertical_0_0,
  output [1023:0] io_outsVertical_0_1,
  output [1023:0] io_outsVertical_0_2,
  output [1023:0] io_outsVertical_0_3,
  output [1023:0] io_outsVertical_1_0,
  output [1023:0] io_outsVertical_1_1,
  output [1023:0] io_outsVertical_1_2,
  output [1023:0] io_outsVertical_1_3,
  output          io_lsbs_0,
  output          io_lsbs_1,
  output          io_lsbs_2,
  output          io_lsbs_3,
  output          io_lsbs_4,
  output          io_lsbs_5,
  output          io_lsbs_6,
  output          io_lsbs_7,
  output          io_lsbs_8,
  output          io_lsbs_9,
  output          io_lsbs_10,
  output          io_lsbs_11,
  output          io_lsbs_12,
  output          io_lsbs_13,
  output          io_lsbs_14,
  output          io_lsbs_15
);
  wire  ces_0_0_clock; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_1_clock; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_2_clock; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_3_clock; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_0_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_0_clock; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_1_clock; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_2_clock; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_3_clock; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_1_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_0_clock; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_1_clock; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_2_clock; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_3_clock; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_2_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_0_clock; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_1_clock; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_2_clock; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_3_clock; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [1023:0] ces_3_3_io_outs_3; // @[MockArray.scala 36:52]
  Element ces_0_0 ( // @[MockArray.scala 36:52]
    .clock(ces_0_0_clock),
    .io_ins_0(ces_0_0_io_ins_0),
    .io_ins_1(ces_0_0_io_ins_1),
    .io_ins_2(ces_0_0_io_ins_2),
    .io_ins_3(ces_0_0_io_ins_3),
    .io_outs_0(ces_0_0_io_outs_0),
    .io_outs_1(ces_0_0_io_outs_1),
    .io_outs_2(ces_0_0_io_outs_2),
    .io_outs_3(ces_0_0_io_outs_3)
  );
  Element ces_0_1 ( // @[MockArray.scala 36:52]
    .clock(ces_0_1_clock),
    .io_ins_0(ces_0_1_io_ins_0),
    .io_ins_1(ces_0_1_io_ins_1),
    .io_ins_2(ces_0_1_io_ins_2),
    .io_ins_3(ces_0_1_io_ins_3),
    .io_outs_0(ces_0_1_io_outs_0),
    .io_outs_1(ces_0_1_io_outs_1),
    .io_outs_2(ces_0_1_io_outs_2),
    .io_outs_3(ces_0_1_io_outs_3)
  );
  Element ces_0_2 ( // @[MockArray.scala 36:52]
    .clock(ces_0_2_clock),
    .io_ins_0(ces_0_2_io_ins_0),
    .io_ins_1(ces_0_2_io_ins_1),
    .io_ins_2(ces_0_2_io_ins_2),
    .io_ins_3(ces_0_2_io_ins_3),
    .io_outs_0(ces_0_2_io_outs_0),
    .io_outs_1(ces_0_2_io_outs_1),
    .io_outs_2(ces_0_2_io_outs_2),
    .io_outs_3(ces_0_2_io_outs_3)
  );
  Element ces_0_3 ( // @[MockArray.scala 36:52]
    .clock(ces_0_3_clock),
    .io_ins_0(ces_0_3_io_ins_0),
    .io_ins_1(ces_0_3_io_ins_1),
    .io_ins_2(ces_0_3_io_ins_2),
    .io_ins_3(ces_0_3_io_ins_3),
    .io_outs_0(ces_0_3_io_outs_0),
    .io_outs_1(ces_0_3_io_outs_1),
    .io_outs_2(ces_0_3_io_outs_2),
    .io_outs_3(ces_0_3_io_outs_3)
  );
  Element ces_1_0 ( // @[MockArray.scala 36:52]
    .clock(ces_1_0_clock),
    .io_ins_0(ces_1_0_io_ins_0),
    .io_ins_1(ces_1_0_io_ins_1),
    .io_ins_2(ces_1_0_io_ins_2),
    .io_ins_3(ces_1_0_io_ins_3),
    .io_outs_0(ces_1_0_io_outs_0),
    .io_outs_1(ces_1_0_io_outs_1),
    .io_outs_2(ces_1_0_io_outs_2),
    .io_outs_3(ces_1_0_io_outs_3)
  );
  Element ces_1_1 ( // @[MockArray.scala 36:52]
    .clock(ces_1_1_clock),
    .io_ins_0(ces_1_1_io_ins_0),
    .io_ins_1(ces_1_1_io_ins_1),
    .io_ins_2(ces_1_1_io_ins_2),
    .io_ins_3(ces_1_1_io_ins_3),
    .io_outs_0(ces_1_1_io_outs_0),
    .io_outs_1(ces_1_1_io_outs_1),
    .io_outs_2(ces_1_1_io_outs_2),
    .io_outs_3(ces_1_1_io_outs_3)
  );
  Element ces_1_2 ( // @[MockArray.scala 36:52]
    .clock(ces_1_2_clock),
    .io_ins_0(ces_1_2_io_ins_0),
    .io_ins_1(ces_1_2_io_ins_1),
    .io_ins_2(ces_1_2_io_ins_2),
    .io_ins_3(ces_1_2_io_ins_3),
    .io_outs_0(ces_1_2_io_outs_0),
    .io_outs_1(ces_1_2_io_outs_1),
    .io_outs_2(ces_1_2_io_outs_2),
    .io_outs_3(ces_1_2_io_outs_3)
  );
  Element ces_1_3 ( // @[MockArray.scala 36:52]
    .clock(ces_1_3_clock),
    .io_ins_0(ces_1_3_io_ins_0),
    .io_ins_1(ces_1_3_io_ins_1),
    .io_ins_2(ces_1_3_io_ins_2),
    .io_ins_3(ces_1_3_io_ins_3),
    .io_outs_0(ces_1_3_io_outs_0),
    .io_outs_1(ces_1_3_io_outs_1),
    .io_outs_2(ces_1_3_io_outs_2),
    .io_outs_3(ces_1_3_io_outs_3)
  );
  Element ces_2_0 ( // @[MockArray.scala 36:52]
    .clock(ces_2_0_clock),
    .io_ins_0(ces_2_0_io_ins_0),
    .io_ins_1(ces_2_0_io_ins_1),
    .io_ins_2(ces_2_0_io_ins_2),
    .io_ins_3(ces_2_0_io_ins_3),
    .io_outs_0(ces_2_0_io_outs_0),
    .io_outs_1(ces_2_0_io_outs_1),
    .io_outs_2(ces_2_0_io_outs_2),
    .io_outs_3(ces_2_0_io_outs_3)
  );
  Element ces_2_1 ( // @[MockArray.scala 36:52]
    .clock(ces_2_1_clock),
    .io_ins_0(ces_2_1_io_ins_0),
    .io_ins_1(ces_2_1_io_ins_1),
    .io_ins_2(ces_2_1_io_ins_2),
    .io_ins_3(ces_2_1_io_ins_3),
    .io_outs_0(ces_2_1_io_outs_0),
    .io_outs_1(ces_2_1_io_outs_1),
    .io_outs_2(ces_2_1_io_outs_2),
    .io_outs_3(ces_2_1_io_outs_3)
  );
  Element ces_2_2 ( // @[MockArray.scala 36:52]
    .clock(ces_2_2_clock),
    .io_ins_0(ces_2_2_io_ins_0),
    .io_ins_1(ces_2_2_io_ins_1),
    .io_ins_2(ces_2_2_io_ins_2),
    .io_ins_3(ces_2_2_io_ins_3),
    .io_outs_0(ces_2_2_io_outs_0),
    .io_outs_1(ces_2_2_io_outs_1),
    .io_outs_2(ces_2_2_io_outs_2),
    .io_outs_3(ces_2_2_io_outs_3)
  );
  Element ces_2_3 ( // @[MockArray.scala 36:52]
    .clock(ces_2_3_clock),
    .io_ins_0(ces_2_3_io_ins_0),
    .io_ins_1(ces_2_3_io_ins_1),
    .io_ins_2(ces_2_3_io_ins_2),
    .io_ins_3(ces_2_3_io_ins_3),
    .io_outs_0(ces_2_3_io_outs_0),
    .io_outs_1(ces_2_3_io_outs_1),
    .io_outs_2(ces_2_3_io_outs_2),
    .io_outs_3(ces_2_3_io_outs_3)
  );
  Element ces_3_0 ( // @[MockArray.scala 36:52]
    .clock(ces_3_0_clock),
    .io_ins_0(ces_3_0_io_ins_0),
    .io_ins_1(ces_3_0_io_ins_1),
    .io_ins_2(ces_3_0_io_ins_2),
    .io_ins_3(ces_3_0_io_ins_3),
    .io_outs_0(ces_3_0_io_outs_0),
    .io_outs_1(ces_3_0_io_outs_1),
    .io_outs_2(ces_3_0_io_outs_2),
    .io_outs_3(ces_3_0_io_outs_3)
  );
  Element ces_3_1 ( // @[MockArray.scala 36:52]
    .clock(ces_3_1_clock),
    .io_ins_0(ces_3_1_io_ins_0),
    .io_ins_1(ces_3_1_io_ins_1),
    .io_ins_2(ces_3_1_io_ins_2),
    .io_ins_3(ces_3_1_io_ins_3),
    .io_outs_0(ces_3_1_io_outs_0),
    .io_outs_1(ces_3_1_io_outs_1),
    .io_outs_2(ces_3_1_io_outs_2),
    .io_outs_3(ces_3_1_io_outs_3)
  );
  Element ces_3_2 ( // @[MockArray.scala 36:52]
    .clock(ces_3_2_clock),
    .io_ins_0(ces_3_2_io_ins_0),
    .io_ins_1(ces_3_2_io_ins_1),
    .io_ins_2(ces_3_2_io_ins_2),
    .io_ins_3(ces_3_2_io_ins_3),
    .io_outs_0(ces_3_2_io_outs_0),
    .io_outs_1(ces_3_2_io_outs_1),
    .io_outs_2(ces_3_2_io_outs_2),
    .io_outs_3(ces_3_2_io_outs_3)
  );
  Element ces_3_3 ( // @[MockArray.scala 36:52]
    .clock(ces_3_3_clock),
    .io_ins_0(ces_3_3_io_ins_0),
    .io_ins_1(ces_3_3_io_ins_1),
    .io_ins_2(ces_3_3_io_ins_2),
    .io_ins_3(ces_3_3_io_ins_3),
    .io_outs_0(ces_3_3_io_outs_0),
    .io_outs_1(ces_3_3_io_outs_1),
    .io_outs_2(ces_3_3_io_outs_2),
    .io_outs_3(ces_3_3_io_outs_3)
  );
  assign io_outsHorizontal_0_0 = ces_0_0_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_1 = ces_0_1_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_2 = ces_0_2_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_3 = ces_0_3_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_1_0 = ces_3_0_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_1 = ces_3_1_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_2 = ces_3_2_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_3 = ces_3_3_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_0 = ces_0_3_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_1 = ces_1_3_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_2 = ces_2_3_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_3 = ces_3_3_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_1_0 = ces_0_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_1 = ces_1_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_2 = ces_2_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_3 = ces_3_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_lsbs_0 = ces_0_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1 = ces_0_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_2 = ces_0_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_3 = ces_0_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_4 = ces_1_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_5 = ces_1_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_6 = ces_1_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_7 = ces_1_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_8 = ces_2_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_9 = ces_2_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_10 = ces_2_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_11 = ces_2_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_12 = ces_3_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_13 = ces_3_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_14 = ces_3_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_15 = ces_3_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign ces_0_0_clock = clock;
  assign ces_0_0_io_ins_0 = io_insHorizontal_0_0; // @[MockArray.scala 44:87]
  assign ces_0_0_io_ins_1 = ces_0_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_0_io_ins_2 = ces_1_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_0_io_ins_3 = io_insVertical_1_0; // @[MockArray.scala 47:87]
  assign ces_0_1_clock = clock;
  assign ces_0_1_io_ins_0 = io_insHorizontal_0_1; // @[MockArray.scala 44:87]
  assign ces_0_1_io_ins_1 = ces_0_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_1_io_ins_2 = ces_1_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_1_io_ins_3 = ces_0_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_2_clock = clock;
  assign ces_0_2_io_ins_0 = io_insHorizontal_0_2; // @[MockArray.scala 44:87]
  assign ces_0_2_io_ins_1 = ces_0_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_2_io_ins_2 = ces_1_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_2_io_ins_3 = ces_0_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_3_clock = clock;
  assign ces_0_3_io_ins_0 = io_insHorizontal_0_3; // @[MockArray.scala 44:87]
  assign ces_0_3_io_ins_1 = io_insVertical_0_0; // @[MockArray.scala 45:87]
  assign ces_0_3_io_ins_2 = ces_1_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_3_io_ins_3 = ces_0_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_0_clock = clock;
  assign ces_1_0_io_ins_0 = ces_0_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_0_io_ins_1 = ces_1_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_0_io_ins_2 = ces_2_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_0_io_ins_3 = io_insVertical_1_1; // @[MockArray.scala 47:87]
  assign ces_1_1_clock = clock;
  assign ces_1_1_io_ins_0 = ces_0_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_1_io_ins_1 = ces_1_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_1_io_ins_2 = ces_2_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_1_io_ins_3 = ces_1_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_2_clock = clock;
  assign ces_1_2_io_ins_0 = ces_0_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_2_io_ins_1 = ces_1_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_2_io_ins_2 = ces_2_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_2_io_ins_3 = ces_1_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_3_clock = clock;
  assign ces_1_3_io_ins_0 = ces_0_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_3_io_ins_1 = io_insVertical_0_1; // @[MockArray.scala 45:87]
  assign ces_1_3_io_ins_2 = ces_2_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_3_io_ins_3 = ces_1_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_0_clock = clock;
  assign ces_2_0_io_ins_0 = ces_1_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_0_io_ins_1 = ces_2_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_0_io_ins_2 = ces_3_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_0_io_ins_3 = io_insVertical_1_2; // @[MockArray.scala 47:87]
  assign ces_2_1_clock = clock;
  assign ces_2_1_io_ins_0 = ces_1_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_1_io_ins_1 = ces_2_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_1_io_ins_2 = ces_3_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_1_io_ins_3 = ces_2_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_2_clock = clock;
  assign ces_2_2_io_ins_0 = ces_1_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_2_io_ins_1 = ces_2_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_2_io_ins_2 = ces_3_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_2_io_ins_3 = ces_2_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_3_clock = clock;
  assign ces_2_3_io_ins_0 = ces_1_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_3_io_ins_1 = io_insVertical_0_2; // @[MockArray.scala 45:87]
  assign ces_2_3_io_ins_2 = ces_3_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_3_io_ins_3 = ces_2_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_0_clock = clock;
  assign ces_3_0_io_ins_0 = ces_2_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_0_io_ins_1 = ces_3_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_0_io_ins_2 = io_insHorizontal_1_0; // @[MockArray.scala 46:87]
  assign ces_3_0_io_ins_3 = io_insVertical_1_3; // @[MockArray.scala 47:87]
  assign ces_3_1_clock = clock;
  assign ces_3_1_io_ins_0 = ces_2_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_1_io_ins_1 = ces_3_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_1_io_ins_2 = io_insHorizontal_1_1; // @[MockArray.scala 46:87]
  assign ces_3_1_io_ins_3 = ces_3_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_2_clock = clock;
  assign ces_3_2_io_ins_0 = ces_2_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_2_io_ins_1 = ces_3_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_2_io_ins_2 = io_insHorizontal_1_2; // @[MockArray.scala 46:87]
  assign ces_3_2_io_ins_3 = ces_3_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_3_clock = clock;
  assign ces_3_3_io_ins_0 = ces_2_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_3_io_ins_1 = io_insVertical_0_3; // @[MockArray.scala 45:87]
  assign ces_3_3_io_ins_2 = io_insHorizontal_1_3; // @[MockArray.scala 46:87]
  assign ces_3_3_io_ins_3 = ces_3_2_io_outs_1; // @[MockArray.scala 63:19]
endmodule
