VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS
MACRO or1200_spram5
  FOREIGN or1200_spram5 0 0 ;
  CLASS BLOCK ;
  SIZE 108.84 BY 162.26 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal7 ;
        RECT  2.94 122.7 59.34 124.1 ;
        RECT  2.94 82.7 59.34 84.1 ;
        RECT  2.94 42.7 59.34 44.1 ;
        RECT  2.94 2.7 59.34 4.1 ;
      LAYER metal4 ;
        RECT  59.04 1.33 59.24 161.07 ;
        RECT  3.04 1.33 3.24 161.07 ;
      LAYER metal1 ;
        RECT  1.14 160.95 107.73 161.05 ;
        RECT  1.14 158.15 107.73 158.25 ;
        RECT  1.14 155.35 107.73 155.45 ;
        RECT  1.14 152.55 107.73 152.65 ;
        RECT  1.14 149.75 107.73 149.85 ;
        RECT  1.14 146.95 107.73 147.05 ;
        RECT  1.14 144.15 107.73 144.25 ;
        RECT  1.14 141.35 107.73 141.45 ;
        RECT  1.14 138.55 107.73 138.65 ;
        RECT  1.14 135.75 107.73 135.85 ;
        RECT  1.14 132.95 107.73 133.05 ;
        RECT  1.14 130.15 107.73 130.25 ;
        RECT  1.14 127.35 107.73 127.45 ;
        RECT  1.14 124.55 107.73 124.65 ;
        RECT  1.14 121.75 107.73 121.85 ;
        RECT  1.14 118.95 107.73 119.05 ;
        RECT  1.14 116.15 107.73 116.25 ;
        RECT  1.14 113.35 107.73 113.45 ;
        RECT  1.14 110.55 107.73 110.65 ;
        RECT  1.14 107.75 107.73 107.85 ;
        RECT  1.14 104.95 107.73 105.05 ;
        RECT  1.14 102.15 107.73 102.25 ;
        RECT  1.14 99.35 107.73 99.45 ;
        RECT  1.14 96.55 107.73 96.65 ;
        RECT  1.14 93.75 107.73 93.85 ;
        RECT  1.14 90.95 107.73 91.05 ;
        RECT  1.14 88.15 107.73 88.25 ;
        RECT  1.14 85.35 107.73 85.45 ;
        RECT  1.14 82.55 107.73 82.65 ;
        RECT  1.14 79.75 107.73 79.85 ;
        RECT  1.14 76.95 107.73 77.05 ;
        RECT  1.14 74.15 107.73 74.25 ;
        RECT  1.14 71.35 107.73 71.45 ;
        RECT  1.14 68.55 107.73 68.65 ;
        RECT  1.14 65.75 107.73 65.85 ;
        RECT  1.14 62.95 107.73 63.05 ;
        RECT  1.14 60.15 107.73 60.25 ;
        RECT  1.14 57.35 107.73 57.45 ;
        RECT  1.14 54.55 107.73 54.65 ;
        RECT  1.14 51.75 107.73 51.85 ;
        RECT  1.14 48.95 107.73 49.05 ;
        RECT  1.14 46.15 107.73 46.25 ;
        RECT  1.14 43.35 107.73 43.45 ;
        RECT  1.14 40.55 107.73 40.65 ;
        RECT  1.14 37.75 107.73 37.85 ;
        RECT  1.14 34.95 107.73 35.05 ;
        RECT  1.14 32.15 107.73 32.25 ;
        RECT  1.14 29.35 107.73 29.45 ;
        RECT  1.14 26.55 107.73 26.65 ;
        RECT  1.14 23.75 107.73 23.85 ;
        RECT  1.14 20.95 107.73 21.05 ;
        RECT  1.14 18.15 107.73 18.25 ;
        RECT  1.14 15.35 107.73 15.45 ;
        RECT  1.14 12.55 107.73 12.65 ;
        RECT  1.14 9.75 107.73 9.85 ;
        RECT  1.14 6.95 107.73 7.05 ;
        RECT  1.14 4.15 107.73 4.25 ;
        RECT  1.14 1.35 107.73 1.45 ;
      VIA 59.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 161 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 161 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 161 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 158.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 158.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 158.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 155.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 155.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 155.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 152.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 152.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 152.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 149.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 149.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 149.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 147 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 147 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 147 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 144.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 144.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 144.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 141.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 141.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 141.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 138.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 138.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 138.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 1.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 161 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 161 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 161 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 158.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 158.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 158.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 155.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 155.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 155.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 152.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 152.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 152.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 149.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 149.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 149.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 147 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 147 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 147 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 144.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 144.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 144.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 141.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 141.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 141.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 138.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 138.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 138.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 1.4 via1_2_400_200_1_1_300_300 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal7 ;
        RECT  30.94 142.7 87.34 144.1 ;
        RECT  30.94 102.7 87.34 104.1 ;
        RECT  30.94 62.7 87.34 64.1 ;
        RECT  30.94 22.7 87.34 24.1 ;
      LAYER metal4 ;
        RECT  87.04 2.73 87.24 159.67 ;
        RECT  31.04 2.73 31.24 159.67 ;
      LAYER metal1 ;
        RECT  1.14 159.55 107.73 159.65 ;
        RECT  1.14 156.75 107.73 156.85 ;
        RECT  1.14 153.95 107.73 154.05 ;
        RECT  1.14 151.15 107.73 151.25 ;
        RECT  1.14 148.35 107.73 148.45 ;
        RECT  1.14 145.55 107.73 145.65 ;
        RECT  1.14 142.75 107.73 142.85 ;
        RECT  1.14 139.95 107.73 140.05 ;
        RECT  1.14 137.15 107.73 137.25 ;
        RECT  1.14 134.35 107.73 134.45 ;
        RECT  1.14 131.55 107.73 131.65 ;
        RECT  1.14 128.75 107.73 128.85 ;
        RECT  1.14 125.95 107.73 126.05 ;
        RECT  1.14 123.15 107.73 123.25 ;
        RECT  1.14 120.35 107.73 120.45 ;
        RECT  1.14 117.55 107.73 117.65 ;
        RECT  1.14 114.75 107.73 114.85 ;
        RECT  1.14 111.95 107.73 112.05 ;
        RECT  1.14 109.15 107.73 109.25 ;
        RECT  1.14 106.35 107.73 106.45 ;
        RECT  1.14 103.55 107.73 103.65 ;
        RECT  1.14 100.75 107.73 100.85 ;
        RECT  1.14 97.95 107.73 98.05 ;
        RECT  1.14 95.15 107.73 95.25 ;
        RECT  1.14 92.35 107.73 92.45 ;
        RECT  1.14 89.55 107.73 89.65 ;
        RECT  1.14 86.75 107.73 86.85 ;
        RECT  1.14 83.95 107.73 84.05 ;
        RECT  1.14 81.15 107.73 81.25 ;
        RECT  1.14 78.35 107.73 78.45 ;
        RECT  1.14 75.55 107.73 75.65 ;
        RECT  1.14 72.75 107.73 72.85 ;
        RECT  1.14 69.95 107.73 70.05 ;
        RECT  1.14 67.15 107.73 67.25 ;
        RECT  1.14 64.35 107.73 64.45 ;
        RECT  1.14 61.55 107.73 61.65 ;
        RECT  1.14 58.75 107.73 58.85 ;
        RECT  1.14 55.95 107.73 56.05 ;
        RECT  1.14 53.15 107.73 53.25 ;
        RECT  1.14 50.35 107.73 50.45 ;
        RECT  1.14 47.55 107.73 47.65 ;
        RECT  1.14 44.75 107.73 44.85 ;
        RECT  1.14 41.95 107.73 42.05 ;
        RECT  1.14 39.15 107.73 39.25 ;
        RECT  1.14 36.35 107.73 36.45 ;
        RECT  1.14 33.55 107.73 33.65 ;
        RECT  1.14 30.75 107.73 30.85 ;
        RECT  1.14 27.95 107.73 28.05 ;
        RECT  1.14 25.15 107.73 25.25 ;
        RECT  1.14 22.35 107.73 22.45 ;
        RECT  1.14 19.55 107.73 19.65 ;
        RECT  1.14 16.75 107.73 16.85 ;
        RECT  1.14 13.95 107.73 14.05 ;
        RECT  1.14 11.15 107.73 11.25 ;
        RECT  1.14 8.35 107.73 8.45 ;
        RECT  1.14 5.55 107.73 5.65 ;
        RECT  1.14 2.75 107.73 2.85 ;
      VIA 87.14 143.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 143.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 143.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 103.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 103.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 103.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 63.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 63.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 63.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 23.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 23.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 23.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 143.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 143.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 143.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 103.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 103.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 103.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 63.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 63.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 63.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 23.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 23.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 23.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 159.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 159.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 159.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 156.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 156.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 156.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 154 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 154 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 154 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 151.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 151.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 151.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 148.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 148.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 148.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 145.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 145.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 145.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 142.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 142.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 142.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 140 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 140 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 140 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 137.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 137.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 137.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 134.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 134.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 134.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 131.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 131.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 131.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 128.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 128.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 128.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 126 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 126 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 126 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 123.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 123.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 123.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 120.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 120.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 120.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 117.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 117.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 117.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 114.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 114.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 114.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 112 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 112 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 112 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 109.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 109.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 109.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 106.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 106.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 106.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 103.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 103.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 103.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 100.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 100.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 100.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 98 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 98 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 98 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 95.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 95.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 95.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 92.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 92.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 92.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 89.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 89.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 89.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 86.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 86.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 86.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 84 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 84 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 84 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 81.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 81.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 81.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 78.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 78.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 78.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 75.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 75.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 75.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 72.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 72.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 72.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 70 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 70 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 70 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 67.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 67.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 67.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 64.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 64.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 64.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 61.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 61.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 61.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 58.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 58.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 58.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 56 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 56 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 56 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 53.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 53.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 53.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 50.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 50.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 50.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 47.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 47.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 47.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 44.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 44.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 44.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 42 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 42 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 42 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 39.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 39.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 39.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 36.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 36.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 36.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 33.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 33.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 33.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 30.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 30.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 30.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 28 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 28 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 28 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 25.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 25.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 25.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 22.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 22.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 22.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 19.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 19.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 19.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 16.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 16.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 16.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 14 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 14 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 14 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 11.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 11.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 11.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 8.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 8.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 8.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 5.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 5.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 5.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 2.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 2.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 2.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 159.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 159.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 159.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 156.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 156.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 156.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 154 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 154 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 154 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 151.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 151.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 151.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 148.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 148.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 148.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 145.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 145.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 145.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 142.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 142.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 142.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 140 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 140 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 140 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 137.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 137.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 137.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 134.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 134.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 134.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 131.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 131.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 131.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 128.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 128.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 128.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 126 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 126 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 126 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 123.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 123.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 123.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 120.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 120.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 120.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 117.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 117.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 117.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 114.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 114.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 114.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 112 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 112 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 112 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 109.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 109.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 109.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 106.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 106.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 106.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 103.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 103.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 103.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 100.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 100.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 100.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 98 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 98 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 98 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 95.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 95.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 95.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 92.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 92.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 92.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 89.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 89.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 89.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 86.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 86.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 86.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 84 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 84 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 84 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 81.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 81.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 81.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 78.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 78.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 78.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 75.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 75.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 75.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 72.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 72.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 72.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 70 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 70 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 70 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 67.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 67.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 67.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 64.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 64.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 64.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 61.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 61.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 61.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 58.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 58.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 58.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 56 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 56 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 56 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 53.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 53.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 53.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 50.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 50.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 50.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 47.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 47.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 47.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 44.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 44.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 44.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 42 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 42 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 42 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 39.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 39.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 39.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 36.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 36.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 36.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 33.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 33.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 33.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 30.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 30.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 30.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 28 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 28 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 28 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 25.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 25.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 25.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 22.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 22.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 22.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 19.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 19.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 19.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 16.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 16.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 16.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 14 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 14 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 14 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 11.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 11.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 11.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 8.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 8.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 8.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 5.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 5.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 5.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 2.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 2.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 2.8 via1_2_400_200_1_1_300_300 ;
    END
  END VDD
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  76.185 0 76.325 0.14 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  108.7 52.64 108.84 52.78 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  108.7 34.16 108.84 34.3 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  9.545 0 9.685 0.14 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  56.585 162.12 56.725 162.26 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  108.7 100.24 108.84 100.38 ;
    END
  END addr[5]
  PIN ce
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  108.7 62.16 108.84 62.3 ;
    END
  END ce
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  108.7 15.12 108.84 15.26 ;
    END
  END clk
  PIN di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  108.7 128.24 108.84 128.38 ;
    END
  END di[0]
  PIN di[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  108.7 109.76 108.84 109.9 ;
    END
  END di[10]
  PIN di[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  108.7 137.76 108.84 137.9 ;
    END
  END di[11]
  PIN di[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  104.185 0 104.325 0.14 ;
    END
  END di[12]
  PIN di[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  28.585 0 28.725 0.14 ;
    END
  END di[13]
  PIN di[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  108.7 71.68 108.84 71.82 ;
    END
  END di[14]
  PIN di[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  47.065 162.12 47.205 162.26 ;
    END
  END di[15]
  PIN di[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  84.585 162.12 84.725 162.26 ;
    END
  END di[16]
  PIN di[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  94.665 0 94.805 0.14 ;
    END
  END di[17]
  PIN di[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 132.72 0.14 132.86 ;
    END
  END di[18]
  PIN di[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  108.7 156.8 108.84 156.94 ;
    END
  END di[19]
  PIN di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 94.64 0.14 94.78 ;
    END
  END di[1]
  PIN di[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 38.08 0.14 38.22 ;
    END
  END di[20]
  PIN di[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 76.16 0.14 76.3 ;
    END
  END di[21]
  PIN di[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  108.7 5.6 108.84 5.74 ;
    END
  END di[22]
  PIN di[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 151.76 0.14 151.9 ;
    END
  END di[23]
  PIN di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 104.16 0.14 104.3 ;
    END
  END di[2]
  PIN di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  108.7 43.68 108.84 43.82 ;
    END
  END di[3]
  PIN di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 113.68 0.14 113.82 ;
    END
  END di[4]
  PIN di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  75.065 162.12 75.205 162.26 ;
    END
  END di[5]
  PIN di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  8.985 162.12 9.125 162.26 ;
    END
  END di[6]
  PIN di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  37.545 162.12 37.685 162.26 ;
    END
  END di[7]
  PIN di[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  57.145 0 57.285 0.14 ;
    END
  END di[8]
  PIN di[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 66.64 0.14 66.78 ;
    END
  END di[9]
  PIN doq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 28.56 0.14 28.7 ;
    END
  END doq[0]
  PIN doq[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 142.24 0.14 142.38 ;
    END
  END doq[10]
  PIN doq[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  66.105 162.12 66.245 162.26 ;
    END
  END doq[11]
  PIN doq[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 19.04 0.14 19.18 ;
    END
  END doq[12]
  PIN doq[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  0.585 0 0.725 0.14 ;
    END
  END doq[13]
  PIN doq[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 57.12 0.14 57.26 ;
    END
  END doq[14]
  PIN doq[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  108.7 147.28 108.84 147.42 ;
    END
  END doq[15]
  PIN doq[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  47.625 0 47.765 0.14 ;
    END
  END doq[16]
  PIN doq[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  108.7 119.28 108.84 119.42 ;
    END
  END doq[17]
  PIN doq[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  108.7 24.64 108.84 24.78 ;
    END
  END doq[18]
  PIN doq[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  28.025 162.12 28.165 162.26 ;
    END
  END doq[19]
  PIN doq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  108.7 81.2 108.84 81.34 ;
    END
  END doq[1]
  PIN doq[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  19.065 0 19.205 0.14 ;
    END
  END doq[20]
  PIN doq[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  38.105 0 38.245 0.14 ;
    END
  END doq[21]
  PIN doq[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 85.12 0.14 85.26 ;
    END
  END doq[22]
  PIN doq[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 9.52 0.14 9.66 ;
    END
  END doq[23]
  PIN doq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  66.665 0 66.805 0.14 ;
    END
  END doq[2]
  PIN doq[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  103.625 162.12 103.765 162.26 ;
    END
  END doq[3]
  PIN doq[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  94.105 162.12 94.245 162.26 ;
    END
  END doq[4]
  PIN doq[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 160.72 0.14 160.86 ;
    END
  END doq[5]
  PIN doq[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  18.505 162.12 18.645 162.26 ;
    END
  END doq[6]
  PIN doq[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  85.145 0 85.285 0.14 ;
    END
  END doq[7]
  PIN doq[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 47.6 0.14 47.74 ;
    END
  END doq[8]
  PIN doq[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 123.2 0.14 123.34 ;
    END
  END doq[9]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  108.7 90.72 108.84 90.86 ;
    END
  END we
  OBS
    LAYER metal1 ;
     RECT  0 0 108.84 162.26 ;
    LAYER metal2 ;
     RECT  0 0 108.84 162.26 ;
    LAYER metal3 ;
     RECT  0 0 108.84 162.26 ;
    LAYER metal4 ;
     RECT  0 0 108.84 162.26 ;
    LAYER metal5 ;
     RECT  0 0 108.84 162.26 ;
    LAYER metal6 ;
     RECT  0 0 108.84 162.26 ;
    LAYER metal7 ;
     RECT  0 0 108.84 162.26 ;
  END
END or1200_spram5
END LIBRARY
