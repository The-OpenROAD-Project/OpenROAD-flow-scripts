VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_1024x32
  FOREIGN fakeram45_1024x32 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 152.190 BY 107.800 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.400 0.070 1.470 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.240 0.070 2.310 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.080 0.070 3.150 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.920 0.070 3.990 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.760 0.070 4.830 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.600 0.070 5.670 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.440 0.070 6.510 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.280 0.070 7.350 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.120 0.070 8.190 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.960 0.070 9.030 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.800 0.070 9.870 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.640 0.070 10.710 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.480 0.070 11.550 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.320 0.070 12.390 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.160 0.070 13.230 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.000 0.070 14.070 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.840 0.070 14.910 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.680 0.070 15.750 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.520 0.070 16.590 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.360 0.070 17.430 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.200 0.070 18.270 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.040 0.070 19.110 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.880 0.070 19.950 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.720 0.070 20.790 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.560 0.070 21.630 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.400 0.070 22.470 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.240 0.070 23.310 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.080 0.070 24.150 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.920 0.070 24.990 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.760 0.070 25.830 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.600 0.070 26.670 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.440 0.070 27.510 ;
    END
  END w_mask_in[31]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.660 0.070 30.730 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.500 0.070 31.570 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.340 0.070 32.410 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.180 0.070 33.250 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.020 0.070 34.090 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.860 0.070 34.930 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.700 0.070 35.770 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.540 0.070 36.610 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.380 0.070 37.450 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.220 0.070 38.290 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.060 0.070 39.130 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.900 0.070 39.970 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.740 0.070 40.810 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.580 0.070 41.650 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.420 0.070 42.490 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.260 0.070 43.330 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.100 0.070 44.170 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.940 0.070 45.010 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.780 0.070 45.850 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.620 0.070 46.690 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.460 0.070 47.530 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.300 0.070 48.370 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.140 0.070 49.210 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.980 0.070 50.050 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.820 0.070 50.890 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.660 0.070 51.730 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.500 0.070 52.570 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.340 0.070 53.410 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.180 0.070 54.250 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.020 0.070 55.090 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.860 0.070 55.930 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.700 0.070 56.770 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.920 0.070 59.990 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.760 0.070 60.830 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.600 0.070 61.670 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.440 0.070 62.510 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.280 0.070 63.350 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.120 0.070 64.190 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.960 0.070 65.030 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.800 0.070 65.870 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.640 0.070 66.710 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.480 0.070 67.550 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.320 0.070 68.390 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.160 0.070 69.230 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.000 0.070 70.070 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.840 0.070 70.910 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.680 0.070 71.750 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.520 0.070 72.590 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.360 0.070 73.430 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.200 0.070 74.270 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.040 0.070 75.110 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.880 0.070 75.950 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.720 0.070 76.790 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.560 0.070 77.630 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.400 0.070 78.470 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.240 0.070 79.310 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.080 0.070 80.150 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.920 0.070 80.990 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.760 0.070 81.830 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.600 0.070 82.670 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.440 0.070 83.510 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.280 0.070 84.350 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.120 0.070 85.190 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.960 0.070 86.030 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.180 0.070 89.250 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.020 0.070 90.090 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.860 0.070 90.930 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.700 0.070 91.770 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.540 0.070 92.610 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.380 0.070 93.450 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.220 0.070 94.290 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.060 0.070 95.130 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.900 0.070 95.970 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.740 0.070 96.810 ;
    END
  END addr_in[9]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.960 0.070 100.030 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.800 0.070 100.870 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.640 0.070 101.710 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 106.400 ;
      RECT 3.500 1.400 3.780 106.400 ;
      RECT 5.740 1.400 6.020 106.400 ;
      RECT 7.980 1.400 8.260 106.400 ;
      RECT 10.220 1.400 10.500 106.400 ;
      RECT 12.460 1.400 12.740 106.400 ;
      RECT 14.700 1.400 14.980 106.400 ;
      RECT 16.940 1.400 17.220 106.400 ;
      RECT 19.180 1.400 19.460 106.400 ;
      RECT 21.420 1.400 21.700 106.400 ;
      RECT 23.660 1.400 23.940 106.400 ;
      RECT 25.900 1.400 26.180 106.400 ;
      RECT 28.140 1.400 28.420 106.400 ;
      RECT 30.380 1.400 30.660 106.400 ;
      RECT 32.620 1.400 32.900 106.400 ;
      RECT 34.860 1.400 35.140 106.400 ;
      RECT 37.100 1.400 37.380 106.400 ;
      RECT 39.340 1.400 39.620 106.400 ;
      RECT 41.580 1.400 41.860 106.400 ;
      RECT 43.820 1.400 44.100 106.400 ;
      RECT 46.060 1.400 46.340 106.400 ;
      RECT 48.300 1.400 48.580 106.400 ;
      RECT 50.540 1.400 50.820 106.400 ;
      RECT 52.780 1.400 53.060 106.400 ;
      RECT 55.020 1.400 55.300 106.400 ;
      RECT 57.260 1.400 57.540 106.400 ;
      RECT 59.500 1.400 59.780 106.400 ;
      RECT 61.740 1.400 62.020 106.400 ;
      RECT 63.980 1.400 64.260 106.400 ;
      RECT 66.220 1.400 66.500 106.400 ;
      RECT 68.460 1.400 68.740 106.400 ;
      RECT 70.700 1.400 70.980 106.400 ;
      RECT 72.940 1.400 73.220 106.400 ;
      RECT 75.180 1.400 75.460 106.400 ;
      RECT 77.420 1.400 77.700 106.400 ;
      RECT 79.660 1.400 79.940 106.400 ;
      RECT 81.900 1.400 82.180 106.400 ;
      RECT 84.140 1.400 84.420 106.400 ;
      RECT 86.380 1.400 86.660 106.400 ;
      RECT 88.620 1.400 88.900 106.400 ;
      RECT 90.860 1.400 91.140 106.400 ;
      RECT 93.100 1.400 93.380 106.400 ;
      RECT 95.340 1.400 95.620 106.400 ;
      RECT 97.580 1.400 97.860 106.400 ;
      RECT 99.820 1.400 100.100 106.400 ;
      RECT 102.060 1.400 102.340 106.400 ;
      RECT 104.300 1.400 104.580 106.400 ;
      RECT 106.540 1.400 106.820 106.400 ;
      RECT 108.780 1.400 109.060 106.400 ;
      RECT 111.020 1.400 111.300 106.400 ;
      RECT 113.260 1.400 113.540 106.400 ;
      RECT 115.500 1.400 115.780 106.400 ;
      RECT 117.740 1.400 118.020 106.400 ;
      RECT 119.980 1.400 120.260 106.400 ;
      RECT 122.220 1.400 122.500 106.400 ;
      RECT 124.460 1.400 124.740 106.400 ;
      RECT 126.700 1.400 126.980 106.400 ;
      RECT 128.940 1.400 129.220 106.400 ;
      RECT 131.180 1.400 131.460 106.400 ;
      RECT 133.420 1.400 133.700 106.400 ;
      RECT 135.660 1.400 135.940 106.400 ;
      RECT 137.900 1.400 138.180 106.400 ;
      RECT 140.140 1.400 140.420 106.400 ;
      RECT 142.380 1.400 142.660 106.400 ;
      RECT 144.620 1.400 144.900 106.400 ;
      RECT 146.860 1.400 147.140 106.400 ;
      RECT 149.100 1.400 149.380 106.400 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 106.400 ;
      RECT 4.620 1.400 4.900 106.400 ;
      RECT 6.860 1.400 7.140 106.400 ;
      RECT 9.100 1.400 9.380 106.400 ;
      RECT 11.340 1.400 11.620 106.400 ;
      RECT 13.580 1.400 13.860 106.400 ;
      RECT 15.820 1.400 16.100 106.400 ;
      RECT 18.060 1.400 18.340 106.400 ;
      RECT 20.300 1.400 20.580 106.400 ;
      RECT 22.540 1.400 22.820 106.400 ;
      RECT 24.780 1.400 25.060 106.400 ;
      RECT 27.020 1.400 27.300 106.400 ;
      RECT 29.260 1.400 29.540 106.400 ;
      RECT 31.500 1.400 31.780 106.400 ;
      RECT 33.740 1.400 34.020 106.400 ;
      RECT 35.980 1.400 36.260 106.400 ;
      RECT 38.220 1.400 38.500 106.400 ;
      RECT 40.460 1.400 40.740 106.400 ;
      RECT 42.700 1.400 42.980 106.400 ;
      RECT 44.940 1.400 45.220 106.400 ;
      RECT 47.180 1.400 47.460 106.400 ;
      RECT 49.420 1.400 49.700 106.400 ;
      RECT 51.660 1.400 51.940 106.400 ;
      RECT 53.900 1.400 54.180 106.400 ;
      RECT 56.140 1.400 56.420 106.400 ;
      RECT 58.380 1.400 58.660 106.400 ;
      RECT 60.620 1.400 60.900 106.400 ;
      RECT 62.860 1.400 63.140 106.400 ;
      RECT 65.100 1.400 65.380 106.400 ;
      RECT 67.340 1.400 67.620 106.400 ;
      RECT 69.580 1.400 69.860 106.400 ;
      RECT 71.820 1.400 72.100 106.400 ;
      RECT 74.060 1.400 74.340 106.400 ;
      RECT 76.300 1.400 76.580 106.400 ;
      RECT 78.540 1.400 78.820 106.400 ;
      RECT 80.780 1.400 81.060 106.400 ;
      RECT 83.020 1.400 83.300 106.400 ;
      RECT 85.260 1.400 85.540 106.400 ;
      RECT 87.500 1.400 87.780 106.400 ;
      RECT 89.740 1.400 90.020 106.400 ;
      RECT 91.980 1.400 92.260 106.400 ;
      RECT 94.220 1.400 94.500 106.400 ;
      RECT 96.460 1.400 96.740 106.400 ;
      RECT 98.700 1.400 98.980 106.400 ;
      RECT 100.940 1.400 101.220 106.400 ;
      RECT 103.180 1.400 103.460 106.400 ;
      RECT 105.420 1.400 105.700 106.400 ;
      RECT 107.660 1.400 107.940 106.400 ;
      RECT 109.900 1.400 110.180 106.400 ;
      RECT 112.140 1.400 112.420 106.400 ;
      RECT 114.380 1.400 114.660 106.400 ;
      RECT 116.620 1.400 116.900 106.400 ;
      RECT 118.860 1.400 119.140 106.400 ;
      RECT 121.100 1.400 121.380 106.400 ;
      RECT 123.340 1.400 123.620 106.400 ;
      RECT 125.580 1.400 125.860 106.400 ;
      RECT 127.820 1.400 128.100 106.400 ;
      RECT 130.060 1.400 130.340 106.400 ;
      RECT 132.300 1.400 132.580 106.400 ;
      RECT 134.540 1.400 134.820 106.400 ;
      RECT 136.780 1.400 137.060 106.400 ;
      RECT 139.020 1.400 139.300 106.400 ;
      RECT 141.260 1.400 141.540 106.400 ;
      RECT 143.500 1.400 143.780 106.400 ;
      RECT 145.740 1.400 146.020 106.400 ;
      RECT 147.980 1.400 148.260 106.400 ;
      RECT 150.220 1.400 150.500 106.400 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 152.190 107.800 ;
    LAYER metal2 ;
    RECT 0 0 152.190 107.800 ;
    LAYER metal3 ;
    RECT 0.070 0 152.190 107.800 ;
    RECT 0 0.000 0.070 1.400 ;
    RECT 0 1.470 0.070 2.240 ;
    RECT 0 2.310 0.070 3.080 ;
    RECT 0 3.150 0.070 3.920 ;
    RECT 0 3.990 0.070 4.760 ;
    RECT 0 4.830 0.070 5.600 ;
    RECT 0 5.670 0.070 6.440 ;
    RECT 0 6.510 0.070 7.280 ;
    RECT 0 7.350 0.070 8.120 ;
    RECT 0 8.190 0.070 8.960 ;
    RECT 0 9.030 0.070 9.800 ;
    RECT 0 9.870 0.070 10.640 ;
    RECT 0 10.710 0.070 11.480 ;
    RECT 0 11.550 0.070 12.320 ;
    RECT 0 12.390 0.070 13.160 ;
    RECT 0 13.230 0.070 14.000 ;
    RECT 0 14.070 0.070 14.840 ;
    RECT 0 14.910 0.070 15.680 ;
    RECT 0 15.750 0.070 16.520 ;
    RECT 0 16.590 0.070 17.360 ;
    RECT 0 17.430 0.070 18.200 ;
    RECT 0 18.270 0.070 19.040 ;
    RECT 0 19.110 0.070 19.880 ;
    RECT 0 19.950 0.070 20.720 ;
    RECT 0 20.790 0.070 21.560 ;
    RECT 0 21.630 0.070 22.400 ;
    RECT 0 22.470 0.070 23.240 ;
    RECT 0 23.310 0.070 24.080 ;
    RECT 0 24.150 0.070 24.920 ;
    RECT 0 24.990 0.070 25.760 ;
    RECT 0 25.830 0.070 26.600 ;
    RECT 0 26.670 0.070 27.440 ;
    RECT 0 27.510 0.070 30.660 ;
    RECT 0 30.730 0.070 31.500 ;
    RECT 0 31.570 0.070 32.340 ;
    RECT 0 32.410 0.070 33.180 ;
    RECT 0 33.250 0.070 34.020 ;
    RECT 0 34.090 0.070 34.860 ;
    RECT 0 34.930 0.070 35.700 ;
    RECT 0 35.770 0.070 36.540 ;
    RECT 0 36.610 0.070 37.380 ;
    RECT 0 37.450 0.070 38.220 ;
    RECT 0 38.290 0.070 39.060 ;
    RECT 0 39.130 0.070 39.900 ;
    RECT 0 39.970 0.070 40.740 ;
    RECT 0 40.810 0.070 41.580 ;
    RECT 0 41.650 0.070 42.420 ;
    RECT 0 42.490 0.070 43.260 ;
    RECT 0 43.330 0.070 44.100 ;
    RECT 0 44.170 0.070 44.940 ;
    RECT 0 45.010 0.070 45.780 ;
    RECT 0 45.850 0.070 46.620 ;
    RECT 0 46.690 0.070 47.460 ;
    RECT 0 47.530 0.070 48.300 ;
    RECT 0 48.370 0.070 49.140 ;
    RECT 0 49.210 0.070 49.980 ;
    RECT 0 50.050 0.070 50.820 ;
    RECT 0 50.890 0.070 51.660 ;
    RECT 0 51.730 0.070 52.500 ;
    RECT 0 52.570 0.070 53.340 ;
    RECT 0 53.410 0.070 54.180 ;
    RECT 0 54.250 0.070 55.020 ;
    RECT 0 55.090 0.070 55.860 ;
    RECT 0 55.930 0.070 56.700 ;
    RECT 0 56.770 0.070 59.920 ;
    RECT 0 59.990 0.070 60.760 ;
    RECT 0 60.830 0.070 61.600 ;
    RECT 0 61.670 0.070 62.440 ;
    RECT 0 62.510 0.070 63.280 ;
    RECT 0 63.350 0.070 64.120 ;
    RECT 0 64.190 0.070 64.960 ;
    RECT 0 65.030 0.070 65.800 ;
    RECT 0 65.870 0.070 66.640 ;
    RECT 0 66.710 0.070 67.480 ;
    RECT 0 67.550 0.070 68.320 ;
    RECT 0 68.390 0.070 69.160 ;
    RECT 0 69.230 0.070 70.000 ;
    RECT 0 70.070 0.070 70.840 ;
    RECT 0 70.910 0.070 71.680 ;
    RECT 0 71.750 0.070 72.520 ;
    RECT 0 72.590 0.070 73.360 ;
    RECT 0 73.430 0.070 74.200 ;
    RECT 0 74.270 0.070 75.040 ;
    RECT 0 75.110 0.070 75.880 ;
    RECT 0 75.950 0.070 76.720 ;
    RECT 0 76.790 0.070 77.560 ;
    RECT 0 77.630 0.070 78.400 ;
    RECT 0 78.470 0.070 79.240 ;
    RECT 0 79.310 0.070 80.080 ;
    RECT 0 80.150 0.070 80.920 ;
    RECT 0 80.990 0.070 81.760 ;
    RECT 0 81.830 0.070 82.600 ;
    RECT 0 82.670 0.070 83.440 ;
    RECT 0 83.510 0.070 84.280 ;
    RECT 0 84.350 0.070 85.120 ;
    RECT 0 85.190 0.070 85.960 ;
    RECT 0 86.030 0.070 89.180 ;
    RECT 0 89.250 0.070 90.020 ;
    RECT 0 90.090 0.070 90.860 ;
    RECT 0 90.930 0.070 91.700 ;
    RECT 0 91.770 0.070 92.540 ;
    RECT 0 92.610 0.070 93.380 ;
    RECT 0 93.450 0.070 94.220 ;
    RECT 0 94.290 0.070 95.060 ;
    RECT 0 95.130 0.070 95.900 ;
    RECT 0 95.970 0.070 96.740 ;
    RECT 0 96.810 0.070 99.960 ;
    RECT 0 100.030 0.070 100.800 ;
    RECT 0 100.870 0.070 101.640 ;
    RECT 0 101.710 0.070 107.800 ;
    LAYER metal4 ;
    RECT 0 0 152.190 1.400 ;
    RECT 0 106.400 152.190 107.800 ;
    RECT 0.000 1.400 1.260 106.400 ;
    RECT 1.540 1.400 2.380 106.400 ;
    RECT 2.660 1.400 3.500 106.400 ;
    RECT 3.780 1.400 4.620 106.400 ;
    RECT 4.900 1.400 5.740 106.400 ;
    RECT 6.020 1.400 6.860 106.400 ;
    RECT 7.140 1.400 7.980 106.400 ;
    RECT 8.260 1.400 9.100 106.400 ;
    RECT 9.380 1.400 10.220 106.400 ;
    RECT 10.500 1.400 11.340 106.400 ;
    RECT 11.620 1.400 12.460 106.400 ;
    RECT 12.740 1.400 13.580 106.400 ;
    RECT 13.860 1.400 14.700 106.400 ;
    RECT 14.980 1.400 15.820 106.400 ;
    RECT 16.100 1.400 16.940 106.400 ;
    RECT 17.220 1.400 18.060 106.400 ;
    RECT 18.340 1.400 19.180 106.400 ;
    RECT 19.460 1.400 20.300 106.400 ;
    RECT 20.580 1.400 21.420 106.400 ;
    RECT 21.700 1.400 22.540 106.400 ;
    RECT 22.820 1.400 23.660 106.400 ;
    RECT 23.940 1.400 24.780 106.400 ;
    RECT 25.060 1.400 25.900 106.400 ;
    RECT 26.180 1.400 27.020 106.400 ;
    RECT 27.300 1.400 28.140 106.400 ;
    RECT 28.420 1.400 29.260 106.400 ;
    RECT 29.540 1.400 30.380 106.400 ;
    RECT 30.660 1.400 31.500 106.400 ;
    RECT 31.780 1.400 32.620 106.400 ;
    RECT 32.900 1.400 33.740 106.400 ;
    RECT 34.020 1.400 34.860 106.400 ;
    RECT 35.140 1.400 35.980 106.400 ;
    RECT 36.260 1.400 37.100 106.400 ;
    RECT 37.380 1.400 38.220 106.400 ;
    RECT 38.500 1.400 39.340 106.400 ;
    RECT 39.620 1.400 40.460 106.400 ;
    RECT 40.740 1.400 41.580 106.400 ;
    RECT 41.860 1.400 42.700 106.400 ;
    RECT 42.980 1.400 43.820 106.400 ;
    RECT 44.100 1.400 44.940 106.400 ;
    RECT 45.220 1.400 46.060 106.400 ;
    RECT 46.340 1.400 47.180 106.400 ;
    RECT 47.460 1.400 48.300 106.400 ;
    RECT 48.580 1.400 49.420 106.400 ;
    RECT 49.700 1.400 50.540 106.400 ;
    RECT 50.820 1.400 51.660 106.400 ;
    RECT 51.940 1.400 52.780 106.400 ;
    RECT 53.060 1.400 53.900 106.400 ;
    RECT 54.180 1.400 55.020 106.400 ;
    RECT 55.300 1.400 56.140 106.400 ;
    RECT 56.420 1.400 57.260 106.400 ;
    RECT 57.540 1.400 58.380 106.400 ;
    RECT 58.660 1.400 59.500 106.400 ;
    RECT 59.780 1.400 60.620 106.400 ;
    RECT 60.900 1.400 61.740 106.400 ;
    RECT 62.020 1.400 62.860 106.400 ;
    RECT 63.140 1.400 63.980 106.400 ;
    RECT 64.260 1.400 65.100 106.400 ;
    RECT 65.380 1.400 66.220 106.400 ;
    RECT 66.500 1.400 67.340 106.400 ;
    RECT 67.620 1.400 68.460 106.400 ;
    RECT 68.740 1.400 69.580 106.400 ;
    RECT 69.860 1.400 70.700 106.400 ;
    RECT 70.980 1.400 71.820 106.400 ;
    RECT 72.100 1.400 72.940 106.400 ;
    RECT 73.220 1.400 74.060 106.400 ;
    RECT 74.340 1.400 75.180 106.400 ;
    RECT 75.460 1.400 76.300 106.400 ;
    RECT 76.580 1.400 77.420 106.400 ;
    RECT 77.700 1.400 78.540 106.400 ;
    RECT 78.820 1.400 79.660 106.400 ;
    RECT 79.940 1.400 80.780 106.400 ;
    RECT 81.060 1.400 81.900 106.400 ;
    RECT 82.180 1.400 83.020 106.400 ;
    RECT 83.300 1.400 84.140 106.400 ;
    RECT 84.420 1.400 85.260 106.400 ;
    RECT 85.540 1.400 86.380 106.400 ;
    RECT 86.660 1.400 87.500 106.400 ;
    RECT 87.780 1.400 88.620 106.400 ;
    RECT 88.900 1.400 89.740 106.400 ;
    RECT 90.020 1.400 90.860 106.400 ;
    RECT 91.140 1.400 91.980 106.400 ;
    RECT 92.260 1.400 93.100 106.400 ;
    RECT 93.380 1.400 94.220 106.400 ;
    RECT 94.500 1.400 95.340 106.400 ;
    RECT 95.620 1.400 96.460 106.400 ;
    RECT 96.740 1.400 97.580 106.400 ;
    RECT 97.860 1.400 98.700 106.400 ;
    RECT 98.980 1.400 99.820 106.400 ;
    RECT 100.100 1.400 100.940 106.400 ;
    RECT 101.220 1.400 102.060 106.400 ;
    RECT 102.340 1.400 103.180 106.400 ;
    RECT 103.460 1.400 104.300 106.400 ;
    RECT 104.580 1.400 105.420 106.400 ;
    RECT 105.700 1.400 106.540 106.400 ;
    RECT 106.820 1.400 107.660 106.400 ;
    RECT 107.940 1.400 108.780 106.400 ;
    RECT 109.060 1.400 109.900 106.400 ;
    RECT 110.180 1.400 111.020 106.400 ;
    RECT 111.300 1.400 112.140 106.400 ;
    RECT 112.420 1.400 113.260 106.400 ;
    RECT 113.540 1.400 114.380 106.400 ;
    RECT 114.660 1.400 115.500 106.400 ;
    RECT 115.780 1.400 116.620 106.400 ;
    RECT 116.900 1.400 117.740 106.400 ;
    RECT 118.020 1.400 118.860 106.400 ;
    RECT 119.140 1.400 119.980 106.400 ;
    RECT 120.260 1.400 121.100 106.400 ;
    RECT 121.380 1.400 122.220 106.400 ;
    RECT 122.500 1.400 123.340 106.400 ;
    RECT 123.620 1.400 124.460 106.400 ;
    RECT 124.740 1.400 125.580 106.400 ;
    RECT 125.860 1.400 126.700 106.400 ;
    RECT 126.980 1.400 127.820 106.400 ;
    RECT 128.100 1.400 128.940 106.400 ;
    RECT 129.220 1.400 130.060 106.400 ;
    RECT 130.340 1.400 131.180 106.400 ;
    RECT 131.460 1.400 132.300 106.400 ;
    RECT 132.580 1.400 133.420 106.400 ;
    RECT 133.700 1.400 134.540 106.400 ;
    RECT 134.820 1.400 135.660 106.400 ;
    RECT 135.940 1.400 136.780 106.400 ;
    RECT 137.060 1.400 137.900 106.400 ;
    RECT 138.180 1.400 139.020 106.400 ;
    RECT 139.300 1.400 140.140 106.400 ;
    RECT 140.420 1.400 141.260 106.400 ;
    RECT 141.540 1.400 142.380 106.400 ;
    RECT 142.660 1.400 143.500 106.400 ;
    RECT 143.780 1.400 144.620 106.400 ;
    RECT 144.900 1.400 145.740 106.400 ;
    RECT 146.020 1.400 146.860 106.400 ;
    RECT 147.140 1.400 147.980 106.400 ;
    RECT 148.260 1.400 149.100 106.400 ;
    RECT 149.380 1.400 150.220 106.400 ;
    RECT 150.500 1.400 152.190 106.400 ;
    LAYER OVERLAP ;
    RECT 0 0 152.190 107.800 ;
  END
END fakeram45_1024x32

END LIBRARY
