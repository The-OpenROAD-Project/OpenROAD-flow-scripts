module MockArray(
  input         clock,
  input         reset,
  input  [63:0] io_insHorizontal_0_0,
  input  [63:0] io_insHorizontal_0_1,
  input  [63:0] io_insHorizontal_0_2,
  input  [63:0] io_insHorizontal_0_3,
  input  [63:0] io_insHorizontal_0_4,
  input  [63:0] io_insHorizontal_0_5,
  input  [63:0] io_insHorizontal_0_6,
  input  [63:0] io_insHorizontal_0_7,
  input  [63:0] io_insHorizontal_1_0,
  input  [63:0] io_insHorizontal_1_1,
  input  [63:0] io_insHorizontal_1_2,
  input  [63:0] io_insHorizontal_1_3,
  input  [63:0] io_insHorizontal_1_4,
  input  [63:0] io_insHorizontal_1_5,
  input  [63:0] io_insHorizontal_1_6,
  input  [63:0] io_insHorizontal_1_7,
  output [63:0] io_outsHorizontal_0_0,
  output [63:0] io_outsHorizontal_0_1,
  output [63:0] io_outsHorizontal_0_2,
  output [63:0] io_outsHorizontal_0_3,
  output [63:0] io_outsHorizontal_0_4,
  output [63:0] io_outsHorizontal_0_5,
  output [63:0] io_outsHorizontal_0_6,
  output [63:0] io_outsHorizontal_0_7,
  output [63:0] io_outsHorizontal_1_0,
  output [63:0] io_outsHorizontal_1_1,
  output [63:0] io_outsHorizontal_1_2,
  output [63:0] io_outsHorizontal_1_3,
  output [63:0] io_outsHorizontal_1_4,
  output [63:0] io_outsHorizontal_1_5,
  output [63:0] io_outsHorizontal_1_6,
  output [63:0] io_outsHorizontal_1_7,
  input  [63:0] io_insVertical_0_0,
  input  [63:0] io_insVertical_0_1,
  input  [63:0] io_insVertical_0_2,
  input  [63:0] io_insVertical_0_3,
  input  [63:0] io_insVertical_0_4,
  input  [63:0] io_insVertical_0_5,
  input  [63:0] io_insVertical_0_6,
  input  [63:0] io_insVertical_0_7,
  input  [63:0] io_insVertical_1_0,
  input  [63:0] io_insVertical_1_1,
  input  [63:0] io_insVertical_1_2,
  input  [63:0] io_insVertical_1_3,
  input  [63:0] io_insVertical_1_4,
  input  [63:0] io_insVertical_1_5,
  input  [63:0] io_insVertical_1_6,
  input  [63:0] io_insVertical_1_7,
  output [63:0] io_outsVertical_0_0,
  output [63:0] io_outsVertical_0_1,
  output [63:0] io_outsVertical_0_2,
  output [63:0] io_outsVertical_0_3,
  output [63:0] io_outsVertical_0_4,
  output [63:0] io_outsVertical_0_5,
  output [63:0] io_outsVertical_0_6,
  output [63:0] io_outsVertical_0_7,
  output [63:0] io_outsVertical_1_0,
  output [63:0] io_outsVertical_1_1,
  output [63:0] io_outsVertical_1_2,
  output [63:0] io_outsVertical_1_3,
  output [63:0] io_outsVertical_1_4,
  output [63:0] io_outsVertical_1_5,
  output [63:0] io_outsVertical_1_6,
  output [63:0] io_outsVertical_1_7,
  output        io_lsbs_0,
  output        io_lsbs_1,
  output        io_lsbs_2,
  output        io_lsbs_3,
  output        io_lsbs_4,
  output        io_lsbs_5,
  output        io_lsbs_6,
  output        io_lsbs_7,
  output        io_lsbs_8,
  output        io_lsbs_9,
  output        io_lsbs_10,
  output        io_lsbs_11,
  output        io_lsbs_12,
  output        io_lsbs_13,
  output        io_lsbs_14,
  output        io_lsbs_15,
  output        io_lsbs_16,
  output        io_lsbs_17,
  output        io_lsbs_18,
  output        io_lsbs_19,
  output        io_lsbs_20,
  output        io_lsbs_21,
  output        io_lsbs_22,
  output        io_lsbs_23,
  output        io_lsbs_24,
  output        io_lsbs_25,
  output        io_lsbs_26,
  output        io_lsbs_27,
  output        io_lsbs_28,
  output        io_lsbs_29,
  output        io_lsbs_30,
  output        io_lsbs_31,
  output        io_lsbs_32,
  output        io_lsbs_33,
  output        io_lsbs_34,
  output        io_lsbs_35,
  output        io_lsbs_36,
  output        io_lsbs_37,
  output        io_lsbs_38,
  output        io_lsbs_39,
  output        io_lsbs_40,
  output        io_lsbs_41,
  output        io_lsbs_42,
  output        io_lsbs_43,
  output        io_lsbs_44,
  output        io_lsbs_45,
  output        io_lsbs_46,
  output        io_lsbs_47,
  output        io_lsbs_48,
  output        io_lsbs_49,
  output        io_lsbs_50,
  output        io_lsbs_51,
  output        io_lsbs_52,
  output        io_lsbs_53,
  output        io_lsbs_54,
  output        io_lsbs_55,
  output        io_lsbs_56,
  output        io_lsbs_57,
  output        io_lsbs_58,
  output        io_lsbs_59,
  output        io_lsbs_60,
  output        io_lsbs_61,
  output        io_lsbs_62,
  output        io_lsbs_63
);
  wire  ces_0_0_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_0_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_0_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_0_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_0_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_0_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_0_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_0_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_0_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_0_1_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_1_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_1_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_1_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_1_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_1_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_1_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_1_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_1_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_0_2_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_2_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_2_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_2_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_2_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_2_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_2_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_2_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_2_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_0_3_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_3_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_3_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_3_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_3_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_3_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_3_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_3_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_3_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_0_4_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_4_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_4_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_4_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_4_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_4_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_4_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_4_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_4_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_0_5_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_5_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_5_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_5_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_5_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_5_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_5_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_5_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_5_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_0_6_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_6_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_6_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_6_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_6_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_6_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_6_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_6_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_6_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_0_7_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_7_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_7_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_7_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_7_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_7_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_7_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_7_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_0_7_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_1_0_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_0_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_0_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_0_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_0_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_0_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_0_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_0_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_0_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_1_1_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_1_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_1_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_1_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_1_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_1_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_1_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_1_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_1_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_1_2_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_2_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_2_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_2_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_2_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_2_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_2_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_2_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_2_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_1_3_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_3_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_3_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_3_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_3_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_3_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_3_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_3_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_3_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_1_4_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_4_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_4_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_4_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_4_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_4_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_4_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_4_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_4_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_1_5_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_5_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_5_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_5_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_5_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_5_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_5_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_5_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_5_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_1_6_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_6_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_6_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_6_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_6_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_6_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_6_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_6_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_6_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_1_7_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_7_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_7_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_7_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_7_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_7_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_7_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_7_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_1_7_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_2_0_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_0_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_0_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_0_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_0_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_0_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_0_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_0_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_0_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_2_1_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_1_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_1_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_1_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_1_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_1_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_1_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_1_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_1_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_2_2_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_2_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_2_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_2_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_2_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_2_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_2_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_2_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_2_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_2_3_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_3_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_3_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_3_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_3_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_3_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_3_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_3_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_3_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_2_4_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_4_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_4_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_4_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_4_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_4_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_4_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_4_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_4_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_2_5_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_5_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_5_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_5_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_5_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_5_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_5_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_5_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_5_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_2_6_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_6_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_6_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_6_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_6_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_6_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_6_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_6_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_6_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_2_7_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_7_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_7_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_7_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_7_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_7_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_7_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_7_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_2_7_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_3_0_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_0_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_0_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_0_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_0_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_0_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_0_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_0_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_0_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_3_1_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_1_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_1_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_1_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_1_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_1_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_1_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_1_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_1_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_3_2_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_2_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_2_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_2_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_2_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_2_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_2_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_2_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_2_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_3_3_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_3_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_3_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_3_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_3_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_3_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_3_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_3_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_3_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_3_4_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_4_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_4_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_4_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_4_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_4_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_4_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_4_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_4_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_3_5_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_5_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_5_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_5_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_5_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_5_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_5_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_5_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_5_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_3_6_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_6_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_6_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_6_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_6_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_6_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_6_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_6_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_6_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_3_7_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_7_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_7_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_7_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_7_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_7_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_7_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_7_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_3_7_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_4_0_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_0_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_0_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_0_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_0_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_0_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_0_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_0_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_0_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_4_1_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_1_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_1_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_1_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_1_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_1_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_1_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_1_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_1_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_4_2_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_2_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_2_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_2_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_2_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_2_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_2_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_2_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_2_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_4_3_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_3_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_3_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_3_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_3_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_3_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_3_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_3_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_3_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_4_4_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_4_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_4_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_4_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_4_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_4_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_4_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_4_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_4_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_4_5_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_5_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_5_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_5_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_5_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_5_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_5_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_5_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_5_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_4_6_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_6_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_6_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_6_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_6_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_6_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_6_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_6_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_6_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_4_7_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_7_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_7_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_7_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_7_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_7_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_7_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_7_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_4_7_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_5_0_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_0_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_0_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_0_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_0_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_0_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_0_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_0_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_0_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_5_1_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_1_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_1_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_1_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_1_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_1_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_1_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_1_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_1_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_5_2_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_2_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_2_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_2_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_2_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_2_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_2_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_2_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_2_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_5_3_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_3_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_3_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_3_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_3_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_3_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_3_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_3_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_3_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_5_4_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_4_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_4_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_4_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_4_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_4_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_4_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_4_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_4_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_5_5_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_5_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_5_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_5_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_5_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_5_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_5_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_5_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_5_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_5_6_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_6_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_6_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_6_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_6_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_6_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_6_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_6_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_6_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_5_7_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_7_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_7_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_7_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_7_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_7_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_7_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_7_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_5_7_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_6_0_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_0_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_0_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_0_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_0_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_0_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_0_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_0_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_0_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_6_1_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_1_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_1_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_1_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_1_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_1_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_1_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_1_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_1_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_6_2_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_2_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_2_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_2_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_2_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_2_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_2_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_2_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_2_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_6_3_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_3_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_3_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_3_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_3_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_3_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_3_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_3_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_3_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_6_4_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_4_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_4_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_4_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_4_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_4_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_4_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_4_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_4_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_6_5_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_5_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_5_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_5_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_5_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_5_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_5_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_5_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_5_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_6_6_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_6_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_6_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_6_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_6_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_6_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_6_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_6_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_6_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_6_7_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_7_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_7_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_7_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_7_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_7_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_7_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_7_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_6_7_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_7_0_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_0_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_0_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_0_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_0_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_0_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_0_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_0_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_0_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_7_1_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_1_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_1_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_1_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_1_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_1_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_1_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_1_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_1_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_7_2_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_2_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_2_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_2_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_2_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_2_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_2_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_2_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_2_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_7_3_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_3_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_3_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_3_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_3_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_3_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_3_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_3_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_3_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_7_4_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_4_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_4_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_4_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_4_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_4_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_4_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_4_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_4_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_7_5_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_5_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_5_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_5_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_5_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_5_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_5_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_5_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_5_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_7_6_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_6_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_6_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_6_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_6_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_6_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_6_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_6_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_6_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_7_7_clock; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_7_io_ins_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_7_io_ins_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_7_io_ins_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_7_io_ins_3; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_7_io_outs_0; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_7_io_outs_1; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_7_io_outs_2; // @[MockArray.scala 37:53]
  wire [63:0] ces_7_7_io_outs_3; // @[MockArray.scala 37:53]
  Element ces_0_0 ( // @[MockArray.scala 37:53]
    .clock(ces_0_0_clock),
    .io_ins_0(ces_0_0_io_ins_0),
    .io_ins_1(ces_0_0_io_ins_1),
    .io_ins_2(ces_0_0_io_ins_2),
    .io_ins_3(ces_0_0_io_ins_3),
    .io_outs_0(ces_0_0_io_outs_0),
    .io_outs_1(ces_0_0_io_outs_1),
    .io_outs_2(ces_0_0_io_outs_2),
    .io_outs_3(ces_0_0_io_outs_3)
  );
  Element ces_0_1 ( // @[MockArray.scala 37:53]
    .clock(ces_0_1_clock),
    .io_ins_0(ces_0_1_io_ins_0),
    .io_ins_1(ces_0_1_io_ins_1),
    .io_ins_2(ces_0_1_io_ins_2),
    .io_ins_3(ces_0_1_io_ins_3),
    .io_outs_0(ces_0_1_io_outs_0),
    .io_outs_1(ces_0_1_io_outs_1),
    .io_outs_2(ces_0_1_io_outs_2),
    .io_outs_3(ces_0_1_io_outs_3)
  );
  Element ces_0_2 ( // @[MockArray.scala 37:53]
    .clock(ces_0_2_clock),
    .io_ins_0(ces_0_2_io_ins_0),
    .io_ins_1(ces_0_2_io_ins_1),
    .io_ins_2(ces_0_2_io_ins_2),
    .io_ins_3(ces_0_2_io_ins_3),
    .io_outs_0(ces_0_2_io_outs_0),
    .io_outs_1(ces_0_2_io_outs_1),
    .io_outs_2(ces_0_2_io_outs_2),
    .io_outs_3(ces_0_2_io_outs_3)
  );
  Element ces_0_3 ( // @[MockArray.scala 37:53]
    .clock(ces_0_3_clock),
    .io_ins_0(ces_0_3_io_ins_0),
    .io_ins_1(ces_0_3_io_ins_1),
    .io_ins_2(ces_0_3_io_ins_2),
    .io_ins_3(ces_0_3_io_ins_3),
    .io_outs_0(ces_0_3_io_outs_0),
    .io_outs_1(ces_0_3_io_outs_1),
    .io_outs_2(ces_0_3_io_outs_2),
    .io_outs_3(ces_0_3_io_outs_3)
  );
  Element ces_0_4 ( // @[MockArray.scala 37:53]
    .clock(ces_0_4_clock),
    .io_ins_0(ces_0_4_io_ins_0),
    .io_ins_1(ces_0_4_io_ins_1),
    .io_ins_2(ces_0_4_io_ins_2),
    .io_ins_3(ces_0_4_io_ins_3),
    .io_outs_0(ces_0_4_io_outs_0),
    .io_outs_1(ces_0_4_io_outs_1),
    .io_outs_2(ces_0_4_io_outs_2),
    .io_outs_3(ces_0_4_io_outs_3)
  );
  Element ces_0_5 ( // @[MockArray.scala 37:53]
    .clock(ces_0_5_clock),
    .io_ins_0(ces_0_5_io_ins_0),
    .io_ins_1(ces_0_5_io_ins_1),
    .io_ins_2(ces_0_5_io_ins_2),
    .io_ins_3(ces_0_5_io_ins_3),
    .io_outs_0(ces_0_5_io_outs_0),
    .io_outs_1(ces_0_5_io_outs_1),
    .io_outs_2(ces_0_5_io_outs_2),
    .io_outs_3(ces_0_5_io_outs_3)
  );
  Element ces_0_6 ( // @[MockArray.scala 37:53]
    .clock(ces_0_6_clock),
    .io_ins_0(ces_0_6_io_ins_0),
    .io_ins_1(ces_0_6_io_ins_1),
    .io_ins_2(ces_0_6_io_ins_2),
    .io_ins_3(ces_0_6_io_ins_3),
    .io_outs_0(ces_0_6_io_outs_0),
    .io_outs_1(ces_0_6_io_outs_1),
    .io_outs_2(ces_0_6_io_outs_2),
    .io_outs_3(ces_0_6_io_outs_3)
  );
  Element ces_0_7 ( // @[MockArray.scala 37:53]
    .clock(ces_0_7_clock),
    .io_ins_0(ces_0_7_io_ins_0),
    .io_ins_1(ces_0_7_io_ins_1),
    .io_ins_2(ces_0_7_io_ins_2),
    .io_ins_3(ces_0_7_io_ins_3),
    .io_outs_0(ces_0_7_io_outs_0),
    .io_outs_1(ces_0_7_io_outs_1),
    .io_outs_2(ces_0_7_io_outs_2),
    .io_outs_3(ces_0_7_io_outs_3)
  );
  Element ces_1_0 ( // @[MockArray.scala 37:53]
    .clock(ces_1_0_clock),
    .io_ins_0(ces_1_0_io_ins_0),
    .io_ins_1(ces_1_0_io_ins_1),
    .io_ins_2(ces_1_0_io_ins_2),
    .io_ins_3(ces_1_0_io_ins_3),
    .io_outs_0(ces_1_0_io_outs_0),
    .io_outs_1(ces_1_0_io_outs_1),
    .io_outs_2(ces_1_0_io_outs_2),
    .io_outs_3(ces_1_0_io_outs_3)
  );
  Element ces_1_1 ( // @[MockArray.scala 37:53]
    .clock(ces_1_1_clock),
    .io_ins_0(ces_1_1_io_ins_0),
    .io_ins_1(ces_1_1_io_ins_1),
    .io_ins_2(ces_1_1_io_ins_2),
    .io_ins_3(ces_1_1_io_ins_3),
    .io_outs_0(ces_1_1_io_outs_0),
    .io_outs_1(ces_1_1_io_outs_1),
    .io_outs_2(ces_1_1_io_outs_2),
    .io_outs_3(ces_1_1_io_outs_3)
  );
  Element ces_1_2 ( // @[MockArray.scala 37:53]
    .clock(ces_1_2_clock),
    .io_ins_0(ces_1_2_io_ins_0),
    .io_ins_1(ces_1_2_io_ins_1),
    .io_ins_2(ces_1_2_io_ins_2),
    .io_ins_3(ces_1_2_io_ins_3),
    .io_outs_0(ces_1_2_io_outs_0),
    .io_outs_1(ces_1_2_io_outs_1),
    .io_outs_2(ces_1_2_io_outs_2),
    .io_outs_3(ces_1_2_io_outs_3)
  );
  Element ces_1_3 ( // @[MockArray.scala 37:53]
    .clock(ces_1_3_clock),
    .io_ins_0(ces_1_3_io_ins_0),
    .io_ins_1(ces_1_3_io_ins_1),
    .io_ins_2(ces_1_3_io_ins_2),
    .io_ins_3(ces_1_3_io_ins_3),
    .io_outs_0(ces_1_3_io_outs_0),
    .io_outs_1(ces_1_3_io_outs_1),
    .io_outs_2(ces_1_3_io_outs_2),
    .io_outs_3(ces_1_3_io_outs_3)
  );
  Element ces_1_4 ( // @[MockArray.scala 37:53]
    .clock(ces_1_4_clock),
    .io_ins_0(ces_1_4_io_ins_0),
    .io_ins_1(ces_1_4_io_ins_1),
    .io_ins_2(ces_1_4_io_ins_2),
    .io_ins_3(ces_1_4_io_ins_3),
    .io_outs_0(ces_1_4_io_outs_0),
    .io_outs_1(ces_1_4_io_outs_1),
    .io_outs_2(ces_1_4_io_outs_2),
    .io_outs_3(ces_1_4_io_outs_3)
  );
  Element ces_1_5 ( // @[MockArray.scala 37:53]
    .clock(ces_1_5_clock),
    .io_ins_0(ces_1_5_io_ins_0),
    .io_ins_1(ces_1_5_io_ins_1),
    .io_ins_2(ces_1_5_io_ins_2),
    .io_ins_3(ces_1_5_io_ins_3),
    .io_outs_0(ces_1_5_io_outs_0),
    .io_outs_1(ces_1_5_io_outs_1),
    .io_outs_2(ces_1_5_io_outs_2),
    .io_outs_3(ces_1_5_io_outs_3)
  );
  Element ces_1_6 ( // @[MockArray.scala 37:53]
    .clock(ces_1_6_clock),
    .io_ins_0(ces_1_6_io_ins_0),
    .io_ins_1(ces_1_6_io_ins_1),
    .io_ins_2(ces_1_6_io_ins_2),
    .io_ins_3(ces_1_6_io_ins_3),
    .io_outs_0(ces_1_6_io_outs_0),
    .io_outs_1(ces_1_6_io_outs_1),
    .io_outs_2(ces_1_6_io_outs_2),
    .io_outs_3(ces_1_6_io_outs_3)
  );
  Element ces_1_7 ( // @[MockArray.scala 37:53]
    .clock(ces_1_7_clock),
    .io_ins_0(ces_1_7_io_ins_0),
    .io_ins_1(ces_1_7_io_ins_1),
    .io_ins_2(ces_1_7_io_ins_2),
    .io_ins_3(ces_1_7_io_ins_3),
    .io_outs_0(ces_1_7_io_outs_0),
    .io_outs_1(ces_1_7_io_outs_1),
    .io_outs_2(ces_1_7_io_outs_2),
    .io_outs_3(ces_1_7_io_outs_3)
  );
  Element ces_2_0 ( // @[MockArray.scala 37:53]
    .clock(ces_2_0_clock),
    .io_ins_0(ces_2_0_io_ins_0),
    .io_ins_1(ces_2_0_io_ins_1),
    .io_ins_2(ces_2_0_io_ins_2),
    .io_ins_3(ces_2_0_io_ins_3),
    .io_outs_0(ces_2_0_io_outs_0),
    .io_outs_1(ces_2_0_io_outs_1),
    .io_outs_2(ces_2_0_io_outs_2),
    .io_outs_3(ces_2_0_io_outs_3)
  );
  Element ces_2_1 ( // @[MockArray.scala 37:53]
    .clock(ces_2_1_clock),
    .io_ins_0(ces_2_1_io_ins_0),
    .io_ins_1(ces_2_1_io_ins_1),
    .io_ins_2(ces_2_1_io_ins_2),
    .io_ins_3(ces_2_1_io_ins_3),
    .io_outs_0(ces_2_1_io_outs_0),
    .io_outs_1(ces_2_1_io_outs_1),
    .io_outs_2(ces_2_1_io_outs_2),
    .io_outs_3(ces_2_1_io_outs_3)
  );
  Element ces_2_2 ( // @[MockArray.scala 37:53]
    .clock(ces_2_2_clock),
    .io_ins_0(ces_2_2_io_ins_0),
    .io_ins_1(ces_2_2_io_ins_1),
    .io_ins_2(ces_2_2_io_ins_2),
    .io_ins_3(ces_2_2_io_ins_3),
    .io_outs_0(ces_2_2_io_outs_0),
    .io_outs_1(ces_2_2_io_outs_1),
    .io_outs_2(ces_2_2_io_outs_2),
    .io_outs_3(ces_2_2_io_outs_3)
  );
  Element ces_2_3 ( // @[MockArray.scala 37:53]
    .clock(ces_2_3_clock),
    .io_ins_0(ces_2_3_io_ins_0),
    .io_ins_1(ces_2_3_io_ins_1),
    .io_ins_2(ces_2_3_io_ins_2),
    .io_ins_3(ces_2_3_io_ins_3),
    .io_outs_0(ces_2_3_io_outs_0),
    .io_outs_1(ces_2_3_io_outs_1),
    .io_outs_2(ces_2_3_io_outs_2),
    .io_outs_3(ces_2_3_io_outs_3)
  );
  Element ces_2_4 ( // @[MockArray.scala 37:53]
    .clock(ces_2_4_clock),
    .io_ins_0(ces_2_4_io_ins_0),
    .io_ins_1(ces_2_4_io_ins_1),
    .io_ins_2(ces_2_4_io_ins_2),
    .io_ins_3(ces_2_4_io_ins_3),
    .io_outs_0(ces_2_4_io_outs_0),
    .io_outs_1(ces_2_4_io_outs_1),
    .io_outs_2(ces_2_4_io_outs_2),
    .io_outs_3(ces_2_4_io_outs_3)
  );
  Element ces_2_5 ( // @[MockArray.scala 37:53]
    .clock(ces_2_5_clock),
    .io_ins_0(ces_2_5_io_ins_0),
    .io_ins_1(ces_2_5_io_ins_1),
    .io_ins_2(ces_2_5_io_ins_2),
    .io_ins_3(ces_2_5_io_ins_3),
    .io_outs_0(ces_2_5_io_outs_0),
    .io_outs_1(ces_2_5_io_outs_1),
    .io_outs_2(ces_2_5_io_outs_2),
    .io_outs_3(ces_2_5_io_outs_3)
  );
  Element ces_2_6 ( // @[MockArray.scala 37:53]
    .clock(ces_2_6_clock),
    .io_ins_0(ces_2_6_io_ins_0),
    .io_ins_1(ces_2_6_io_ins_1),
    .io_ins_2(ces_2_6_io_ins_2),
    .io_ins_3(ces_2_6_io_ins_3),
    .io_outs_0(ces_2_6_io_outs_0),
    .io_outs_1(ces_2_6_io_outs_1),
    .io_outs_2(ces_2_6_io_outs_2),
    .io_outs_3(ces_2_6_io_outs_3)
  );
  Element ces_2_7 ( // @[MockArray.scala 37:53]
    .clock(ces_2_7_clock),
    .io_ins_0(ces_2_7_io_ins_0),
    .io_ins_1(ces_2_7_io_ins_1),
    .io_ins_2(ces_2_7_io_ins_2),
    .io_ins_3(ces_2_7_io_ins_3),
    .io_outs_0(ces_2_7_io_outs_0),
    .io_outs_1(ces_2_7_io_outs_1),
    .io_outs_2(ces_2_7_io_outs_2),
    .io_outs_3(ces_2_7_io_outs_3)
  );
  Element ces_3_0 ( // @[MockArray.scala 37:53]
    .clock(ces_3_0_clock),
    .io_ins_0(ces_3_0_io_ins_0),
    .io_ins_1(ces_3_0_io_ins_1),
    .io_ins_2(ces_3_0_io_ins_2),
    .io_ins_3(ces_3_0_io_ins_3),
    .io_outs_0(ces_3_0_io_outs_0),
    .io_outs_1(ces_3_0_io_outs_1),
    .io_outs_2(ces_3_0_io_outs_2),
    .io_outs_3(ces_3_0_io_outs_3)
  );
  Element ces_3_1 ( // @[MockArray.scala 37:53]
    .clock(ces_3_1_clock),
    .io_ins_0(ces_3_1_io_ins_0),
    .io_ins_1(ces_3_1_io_ins_1),
    .io_ins_2(ces_3_1_io_ins_2),
    .io_ins_3(ces_3_1_io_ins_3),
    .io_outs_0(ces_3_1_io_outs_0),
    .io_outs_1(ces_3_1_io_outs_1),
    .io_outs_2(ces_3_1_io_outs_2),
    .io_outs_3(ces_3_1_io_outs_3)
  );
  Element ces_3_2 ( // @[MockArray.scala 37:53]
    .clock(ces_3_2_clock),
    .io_ins_0(ces_3_2_io_ins_0),
    .io_ins_1(ces_3_2_io_ins_1),
    .io_ins_2(ces_3_2_io_ins_2),
    .io_ins_3(ces_3_2_io_ins_3),
    .io_outs_0(ces_3_2_io_outs_0),
    .io_outs_1(ces_3_2_io_outs_1),
    .io_outs_2(ces_3_2_io_outs_2),
    .io_outs_3(ces_3_2_io_outs_3)
  );
  Element ces_3_3 ( // @[MockArray.scala 37:53]
    .clock(ces_3_3_clock),
    .io_ins_0(ces_3_3_io_ins_0),
    .io_ins_1(ces_3_3_io_ins_1),
    .io_ins_2(ces_3_3_io_ins_2),
    .io_ins_3(ces_3_3_io_ins_3),
    .io_outs_0(ces_3_3_io_outs_0),
    .io_outs_1(ces_3_3_io_outs_1),
    .io_outs_2(ces_3_3_io_outs_2),
    .io_outs_3(ces_3_3_io_outs_3)
  );
  Element ces_3_4 ( // @[MockArray.scala 37:53]
    .clock(ces_3_4_clock),
    .io_ins_0(ces_3_4_io_ins_0),
    .io_ins_1(ces_3_4_io_ins_1),
    .io_ins_2(ces_3_4_io_ins_2),
    .io_ins_3(ces_3_4_io_ins_3),
    .io_outs_0(ces_3_4_io_outs_0),
    .io_outs_1(ces_3_4_io_outs_1),
    .io_outs_2(ces_3_4_io_outs_2),
    .io_outs_3(ces_3_4_io_outs_3)
  );
  Element ces_3_5 ( // @[MockArray.scala 37:53]
    .clock(ces_3_5_clock),
    .io_ins_0(ces_3_5_io_ins_0),
    .io_ins_1(ces_3_5_io_ins_1),
    .io_ins_2(ces_3_5_io_ins_2),
    .io_ins_3(ces_3_5_io_ins_3),
    .io_outs_0(ces_3_5_io_outs_0),
    .io_outs_1(ces_3_5_io_outs_1),
    .io_outs_2(ces_3_5_io_outs_2),
    .io_outs_3(ces_3_5_io_outs_3)
  );
  Element ces_3_6 ( // @[MockArray.scala 37:53]
    .clock(ces_3_6_clock),
    .io_ins_0(ces_3_6_io_ins_0),
    .io_ins_1(ces_3_6_io_ins_1),
    .io_ins_2(ces_3_6_io_ins_2),
    .io_ins_3(ces_3_6_io_ins_3),
    .io_outs_0(ces_3_6_io_outs_0),
    .io_outs_1(ces_3_6_io_outs_1),
    .io_outs_2(ces_3_6_io_outs_2),
    .io_outs_3(ces_3_6_io_outs_3)
  );
  Element ces_3_7 ( // @[MockArray.scala 37:53]
    .clock(ces_3_7_clock),
    .io_ins_0(ces_3_7_io_ins_0),
    .io_ins_1(ces_3_7_io_ins_1),
    .io_ins_2(ces_3_7_io_ins_2),
    .io_ins_3(ces_3_7_io_ins_3),
    .io_outs_0(ces_3_7_io_outs_0),
    .io_outs_1(ces_3_7_io_outs_1),
    .io_outs_2(ces_3_7_io_outs_2),
    .io_outs_3(ces_3_7_io_outs_3)
  );
  Element ces_4_0 ( // @[MockArray.scala 37:53]
    .clock(ces_4_0_clock),
    .io_ins_0(ces_4_0_io_ins_0),
    .io_ins_1(ces_4_0_io_ins_1),
    .io_ins_2(ces_4_0_io_ins_2),
    .io_ins_3(ces_4_0_io_ins_3),
    .io_outs_0(ces_4_0_io_outs_0),
    .io_outs_1(ces_4_0_io_outs_1),
    .io_outs_2(ces_4_0_io_outs_2),
    .io_outs_3(ces_4_0_io_outs_3)
  );
  Element ces_4_1 ( // @[MockArray.scala 37:53]
    .clock(ces_4_1_clock),
    .io_ins_0(ces_4_1_io_ins_0),
    .io_ins_1(ces_4_1_io_ins_1),
    .io_ins_2(ces_4_1_io_ins_2),
    .io_ins_3(ces_4_1_io_ins_3),
    .io_outs_0(ces_4_1_io_outs_0),
    .io_outs_1(ces_4_1_io_outs_1),
    .io_outs_2(ces_4_1_io_outs_2),
    .io_outs_3(ces_4_1_io_outs_3)
  );
  Element ces_4_2 ( // @[MockArray.scala 37:53]
    .clock(ces_4_2_clock),
    .io_ins_0(ces_4_2_io_ins_0),
    .io_ins_1(ces_4_2_io_ins_1),
    .io_ins_2(ces_4_2_io_ins_2),
    .io_ins_3(ces_4_2_io_ins_3),
    .io_outs_0(ces_4_2_io_outs_0),
    .io_outs_1(ces_4_2_io_outs_1),
    .io_outs_2(ces_4_2_io_outs_2),
    .io_outs_3(ces_4_2_io_outs_3)
  );
  Element ces_4_3 ( // @[MockArray.scala 37:53]
    .clock(ces_4_3_clock),
    .io_ins_0(ces_4_3_io_ins_0),
    .io_ins_1(ces_4_3_io_ins_1),
    .io_ins_2(ces_4_3_io_ins_2),
    .io_ins_3(ces_4_3_io_ins_3),
    .io_outs_0(ces_4_3_io_outs_0),
    .io_outs_1(ces_4_3_io_outs_1),
    .io_outs_2(ces_4_3_io_outs_2),
    .io_outs_3(ces_4_3_io_outs_3)
  );
  Element ces_4_4 ( // @[MockArray.scala 37:53]
    .clock(ces_4_4_clock),
    .io_ins_0(ces_4_4_io_ins_0),
    .io_ins_1(ces_4_4_io_ins_1),
    .io_ins_2(ces_4_4_io_ins_2),
    .io_ins_3(ces_4_4_io_ins_3),
    .io_outs_0(ces_4_4_io_outs_0),
    .io_outs_1(ces_4_4_io_outs_1),
    .io_outs_2(ces_4_4_io_outs_2),
    .io_outs_3(ces_4_4_io_outs_3)
  );
  Element ces_4_5 ( // @[MockArray.scala 37:53]
    .clock(ces_4_5_clock),
    .io_ins_0(ces_4_5_io_ins_0),
    .io_ins_1(ces_4_5_io_ins_1),
    .io_ins_2(ces_4_5_io_ins_2),
    .io_ins_3(ces_4_5_io_ins_3),
    .io_outs_0(ces_4_5_io_outs_0),
    .io_outs_1(ces_4_5_io_outs_1),
    .io_outs_2(ces_4_5_io_outs_2),
    .io_outs_3(ces_4_5_io_outs_3)
  );
  Element ces_4_6 ( // @[MockArray.scala 37:53]
    .clock(ces_4_6_clock),
    .io_ins_0(ces_4_6_io_ins_0),
    .io_ins_1(ces_4_6_io_ins_1),
    .io_ins_2(ces_4_6_io_ins_2),
    .io_ins_3(ces_4_6_io_ins_3),
    .io_outs_0(ces_4_6_io_outs_0),
    .io_outs_1(ces_4_6_io_outs_1),
    .io_outs_2(ces_4_6_io_outs_2),
    .io_outs_3(ces_4_6_io_outs_3)
  );
  Element ces_4_7 ( // @[MockArray.scala 37:53]
    .clock(ces_4_7_clock),
    .io_ins_0(ces_4_7_io_ins_0),
    .io_ins_1(ces_4_7_io_ins_1),
    .io_ins_2(ces_4_7_io_ins_2),
    .io_ins_3(ces_4_7_io_ins_3),
    .io_outs_0(ces_4_7_io_outs_0),
    .io_outs_1(ces_4_7_io_outs_1),
    .io_outs_2(ces_4_7_io_outs_2),
    .io_outs_3(ces_4_7_io_outs_3)
  );
  Element ces_5_0 ( // @[MockArray.scala 37:53]
    .clock(ces_5_0_clock),
    .io_ins_0(ces_5_0_io_ins_0),
    .io_ins_1(ces_5_0_io_ins_1),
    .io_ins_2(ces_5_0_io_ins_2),
    .io_ins_3(ces_5_0_io_ins_3),
    .io_outs_0(ces_5_0_io_outs_0),
    .io_outs_1(ces_5_0_io_outs_1),
    .io_outs_2(ces_5_0_io_outs_2),
    .io_outs_3(ces_5_0_io_outs_3)
  );
  Element ces_5_1 ( // @[MockArray.scala 37:53]
    .clock(ces_5_1_clock),
    .io_ins_0(ces_5_1_io_ins_0),
    .io_ins_1(ces_5_1_io_ins_1),
    .io_ins_2(ces_5_1_io_ins_2),
    .io_ins_3(ces_5_1_io_ins_3),
    .io_outs_0(ces_5_1_io_outs_0),
    .io_outs_1(ces_5_1_io_outs_1),
    .io_outs_2(ces_5_1_io_outs_2),
    .io_outs_3(ces_5_1_io_outs_3)
  );
  Element ces_5_2 ( // @[MockArray.scala 37:53]
    .clock(ces_5_2_clock),
    .io_ins_0(ces_5_2_io_ins_0),
    .io_ins_1(ces_5_2_io_ins_1),
    .io_ins_2(ces_5_2_io_ins_2),
    .io_ins_3(ces_5_2_io_ins_3),
    .io_outs_0(ces_5_2_io_outs_0),
    .io_outs_1(ces_5_2_io_outs_1),
    .io_outs_2(ces_5_2_io_outs_2),
    .io_outs_3(ces_5_2_io_outs_3)
  );
  Element ces_5_3 ( // @[MockArray.scala 37:53]
    .clock(ces_5_3_clock),
    .io_ins_0(ces_5_3_io_ins_0),
    .io_ins_1(ces_5_3_io_ins_1),
    .io_ins_2(ces_5_3_io_ins_2),
    .io_ins_3(ces_5_3_io_ins_3),
    .io_outs_0(ces_5_3_io_outs_0),
    .io_outs_1(ces_5_3_io_outs_1),
    .io_outs_2(ces_5_3_io_outs_2),
    .io_outs_3(ces_5_3_io_outs_3)
  );
  Element ces_5_4 ( // @[MockArray.scala 37:53]
    .clock(ces_5_4_clock),
    .io_ins_0(ces_5_4_io_ins_0),
    .io_ins_1(ces_5_4_io_ins_1),
    .io_ins_2(ces_5_4_io_ins_2),
    .io_ins_3(ces_5_4_io_ins_3),
    .io_outs_0(ces_5_4_io_outs_0),
    .io_outs_1(ces_5_4_io_outs_1),
    .io_outs_2(ces_5_4_io_outs_2),
    .io_outs_3(ces_5_4_io_outs_3)
  );
  Element ces_5_5 ( // @[MockArray.scala 37:53]
    .clock(ces_5_5_clock),
    .io_ins_0(ces_5_5_io_ins_0),
    .io_ins_1(ces_5_5_io_ins_1),
    .io_ins_2(ces_5_5_io_ins_2),
    .io_ins_3(ces_5_5_io_ins_3),
    .io_outs_0(ces_5_5_io_outs_0),
    .io_outs_1(ces_5_5_io_outs_1),
    .io_outs_2(ces_5_5_io_outs_2),
    .io_outs_3(ces_5_5_io_outs_3)
  );
  Element ces_5_6 ( // @[MockArray.scala 37:53]
    .clock(ces_5_6_clock),
    .io_ins_0(ces_5_6_io_ins_0),
    .io_ins_1(ces_5_6_io_ins_1),
    .io_ins_2(ces_5_6_io_ins_2),
    .io_ins_3(ces_5_6_io_ins_3),
    .io_outs_0(ces_5_6_io_outs_0),
    .io_outs_1(ces_5_6_io_outs_1),
    .io_outs_2(ces_5_6_io_outs_2),
    .io_outs_3(ces_5_6_io_outs_3)
  );
  Element ces_5_7 ( // @[MockArray.scala 37:53]
    .clock(ces_5_7_clock),
    .io_ins_0(ces_5_7_io_ins_0),
    .io_ins_1(ces_5_7_io_ins_1),
    .io_ins_2(ces_5_7_io_ins_2),
    .io_ins_3(ces_5_7_io_ins_3),
    .io_outs_0(ces_5_7_io_outs_0),
    .io_outs_1(ces_5_7_io_outs_1),
    .io_outs_2(ces_5_7_io_outs_2),
    .io_outs_3(ces_5_7_io_outs_3)
  );
  Element ces_6_0 ( // @[MockArray.scala 37:53]
    .clock(ces_6_0_clock),
    .io_ins_0(ces_6_0_io_ins_0),
    .io_ins_1(ces_6_0_io_ins_1),
    .io_ins_2(ces_6_0_io_ins_2),
    .io_ins_3(ces_6_0_io_ins_3),
    .io_outs_0(ces_6_0_io_outs_0),
    .io_outs_1(ces_6_0_io_outs_1),
    .io_outs_2(ces_6_0_io_outs_2),
    .io_outs_3(ces_6_0_io_outs_3)
  );
  Element ces_6_1 ( // @[MockArray.scala 37:53]
    .clock(ces_6_1_clock),
    .io_ins_0(ces_6_1_io_ins_0),
    .io_ins_1(ces_6_1_io_ins_1),
    .io_ins_2(ces_6_1_io_ins_2),
    .io_ins_3(ces_6_1_io_ins_3),
    .io_outs_0(ces_6_1_io_outs_0),
    .io_outs_1(ces_6_1_io_outs_1),
    .io_outs_2(ces_6_1_io_outs_2),
    .io_outs_3(ces_6_1_io_outs_3)
  );
  Element ces_6_2 ( // @[MockArray.scala 37:53]
    .clock(ces_6_2_clock),
    .io_ins_0(ces_6_2_io_ins_0),
    .io_ins_1(ces_6_2_io_ins_1),
    .io_ins_2(ces_6_2_io_ins_2),
    .io_ins_3(ces_6_2_io_ins_3),
    .io_outs_0(ces_6_2_io_outs_0),
    .io_outs_1(ces_6_2_io_outs_1),
    .io_outs_2(ces_6_2_io_outs_2),
    .io_outs_3(ces_6_2_io_outs_3)
  );
  Element ces_6_3 ( // @[MockArray.scala 37:53]
    .clock(ces_6_3_clock),
    .io_ins_0(ces_6_3_io_ins_0),
    .io_ins_1(ces_6_3_io_ins_1),
    .io_ins_2(ces_6_3_io_ins_2),
    .io_ins_3(ces_6_3_io_ins_3),
    .io_outs_0(ces_6_3_io_outs_0),
    .io_outs_1(ces_6_3_io_outs_1),
    .io_outs_2(ces_6_3_io_outs_2),
    .io_outs_3(ces_6_3_io_outs_3)
  );
  Element ces_6_4 ( // @[MockArray.scala 37:53]
    .clock(ces_6_4_clock),
    .io_ins_0(ces_6_4_io_ins_0),
    .io_ins_1(ces_6_4_io_ins_1),
    .io_ins_2(ces_6_4_io_ins_2),
    .io_ins_3(ces_6_4_io_ins_3),
    .io_outs_0(ces_6_4_io_outs_0),
    .io_outs_1(ces_6_4_io_outs_1),
    .io_outs_2(ces_6_4_io_outs_2),
    .io_outs_3(ces_6_4_io_outs_3)
  );
  Element ces_6_5 ( // @[MockArray.scala 37:53]
    .clock(ces_6_5_clock),
    .io_ins_0(ces_6_5_io_ins_0),
    .io_ins_1(ces_6_5_io_ins_1),
    .io_ins_2(ces_6_5_io_ins_2),
    .io_ins_3(ces_6_5_io_ins_3),
    .io_outs_0(ces_6_5_io_outs_0),
    .io_outs_1(ces_6_5_io_outs_1),
    .io_outs_2(ces_6_5_io_outs_2),
    .io_outs_3(ces_6_5_io_outs_3)
  );
  Element ces_6_6 ( // @[MockArray.scala 37:53]
    .clock(ces_6_6_clock),
    .io_ins_0(ces_6_6_io_ins_0),
    .io_ins_1(ces_6_6_io_ins_1),
    .io_ins_2(ces_6_6_io_ins_2),
    .io_ins_3(ces_6_6_io_ins_3),
    .io_outs_0(ces_6_6_io_outs_0),
    .io_outs_1(ces_6_6_io_outs_1),
    .io_outs_2(ces_6_6_io_outs_2),
    .io_outs_3(ces_6_6_io_outs_3)
  );
  Element ces_6_7 ( // @[MockArray.scala 37:53]
    .clock(ces_6_7_clock),
    .io_ins_0(ces_6_7_io_ins_0),
    .io_ins_1(ces_6_7_io_ins_1),
    .io_ins_2(ces_6_7_io_ins_2),
    .io_ins_3(ces_6_7_io_ins_3),
    .io_outs_0(ces_6_7_io_outs_0),
    .io_outs_1(ces_6_7_io_outs_1),
    .io_outs_2(ces_6_7_io_outs_2),
    .io_outs_3(ces_6_7_io_outs_3)
  );
  Element ces_7_0 ( // @[MockArray.scala 37:53]
    .clock(ces_7_0_clock),
    .io_ins_0(ces_7_0_io_ins_0),
    .io_ins_1(ces_7_0_io_ins_1),
    .io_ins_2(ces_7_0_io_ins_2),
    .io_ins_3(ces_7_0_io_ins_3),
    .io_outs_0(ces_7_0_io_outs_0),
    .io_outs_1(ces_7_0_io_outs_1),
    .io_outs_2(ces_7_0_io_outs_2),
    .io_outs_3(ces_7_0_io_outs_3)
  );
  Element ces_7_1 ( // @[MockArray.scala 37:53]
    .clock(ces_7_1_clock),
    .io_ins_0(ces_7_1_io_ins_0),
    .io_ins_1(ces_7_1_io_ins_1),
    .io_ins_2(ces_7_1_io_ins_2),
    .io_ins_3(ces_7_1_io_ins_3),
    .io_outs_0(ces_7_1_io_outs_0),
    .io_outs_1(ces_7_1_io_outs_1),
    .io_outs_2(ces_7_1_io_outs_2),
    .io_outs_3(ces_7_1_io_outs_3)
  );
  Element ces_7_2 ( // @[MockArray.scala 37:53]
    .clock(ces_7_2_clock),
    .io_ins_0(ces_7_2_io_ins_0),
    .io_ins_1(ces_7_2_io_ins_1),
    .io_ins_2(ces_7_2_io_ins_2),
    .io_ins_3(ces_7_2_io_ins_3),
    .io_outs_0(ces_7_2_io_outs_0),
    .io_outs_1(ces_7_2_io_outs_1),
    .io_outs_2(ces_7_2_io_outs_2),
    .io_outs_3(ces_7_2_io_outs_3)
  );
  Element ces_7_3 ( // @[MockArray.scala 37:53]
    .clock(ces_7_3_clock),
    .io_ins_0(ces_7_3_io_ins_0),
    .io_ins_1(ces_7_3_io_ins_1),
    .io_ins_2(ces_7_3_io_ins_2),
    .io_ins_3(ces_7_3_io_ins_3),
    .io_outs_0(ces_7_3_io_outs_0),
    .io_outs_1(ces_7_3_io_outs_1),
    .io_outs_2(ces_7_3_io_outs_2),
    .io_outs_3(ces_7_3_io_outs_3)
  );
  Element ces_7_4 ( // @[MockArray.scala 37:53]
    .clock(ces_7_4_clock),
    .io_ins_0(ces_7_4_io_ins_0),
    .io_ins_1(ces_7_4_io_ins_1),
    .io_ins_2(ces_7_4_io_ins_2),
    .io_ins_3(ces_7_4_io_ins_3),
    .io_outs_0(ces_7_4_io_outs_0),
    .io_outs_1(ces_7_4_io_outs_1),
    .io_outs_2(ces_7_4_io_outs_2),
    .io_outs_3(ces_7_4_io_outs_3)
  );
  Element ces_7_5 ( // @[MockArray.scala 37:53]
    .clock(ces_7_5_clock),
    .io_ins_0(ces_7_5_io_ins_0),
    .io_ins_1(ces_7_5_io_ins_1),
    .io_ins_2(ces_7_5_io_ins_2),
    .io_ins_3(ces_7_5_io_ins_3),
    .io_outs_0(ces_7_5_io_outs_0),
    .io_outs_1(ces_7_5_io_outs_1),
    .io_outs_2(ces_7_5_io_outs_2),
    .io_outs_3(ces_7_5_io_outs_3)
  );
  Element ces_7_6 ( // @[MockArray.scala 37:53]
    .clock(ces_7_6_clock),
    .io_ins_0(ces_7_6_io_ins_0),
    .io_ins_1(ces_7_6_io_ins_1),
    .io_ins_2(ces_7_6_io_ins_2),
    .io_ins_3(ces_7_6_io_ins_3),
    .io_outs_0(ces_7_6_io_outs_0),
    .io_outs_1(ces_7_6_io_outs_1),
    .io_outs_2(ces_7_6_io_outs_2),
    .io_outs_3(ces_7_6_io_outs_3)
  );
  Element ces_7_7 ( // @[MockArray.scala 37:53]
    .clock(ces_7_7_clock),
    .io_ins_0(ces_7_7_io_ins_0),
    .io_ins_1(ces_7_7_io_ins_1),
    .io_ins_2(ces_7_7_io_ins_2),
    .io_ins_3(ces_7_7_io_ins_3),
    .io_outs_0(ces_7_7_io_outs_0),
    .io_outs_1(ces_7_7_io_outs_1),
    .io_outs_2(ces_7_7_io_outs_2),
    .io_outs_3(ces_7_7_io_outs_3)
  );
  assign io_outsHorizontal_0_0 = ces_0_0_io_outs_0; // @[MockArray.scala 50:89]
  assign io_outsHorizontal_0_1 = ces_0_1_io_outs_0; // @[MockArray.scala 50:89]
  assign io_outsHorizontal_0_2 = ces_0_2_io_outs_0; // @[MockArray.scala 50:89]
  assign io_outsHorizontal_0_3 = ces_0_3_io_outs_0; // @[MockArray.scala 50:89]
  assign io_outsHorizontal_0_4 = ces_0_4_io_outs_0; // @[MockArray.scala 50:89]
  assign io_outsHorizontal_0_5 = ces_0_5_io_outs_0; // @[MockArray.scala 50:89]
  assign io_outsHorizontal_0_6 = ces_0_6_io_outs_0; // @[MockArray.scala 50:89]
  assign io_outsHorizontal_0_7 = ces_0_7_io_outs_0; // @[MockArray.scala 50:89]
  assign io_outsHorizontal_1_0 = ces_7_0_io_outs_2; // @[MockArray.scala 52:89]
  assign io_outsHorizontal_1_1 = ces_7_1_io_outs_2; // @[MockArray.scala 52:89]
  assign io_outsHorizontal_1_2 = ces_7_2_io_outs_2; // @[MockArray.scala 52:89]
  assign io_outsHorizontal_1_3 = ces_7_3_io_outs_2; // @[MockArray.scala 52:89]
  assign io_outsHorizontal_1_4 = ces_7_4_io_outs_2; // @[MockArray.scala 52:89]
  assign io_outsHorizontal_1_5 = ces_7_5_io_outs_2; // @[MockArray.scala 52:89]
  assign io_outsHorizontal_1_6 = ces_7_6_io_outs_2; // @[MockArray.scala 52:89]
  assign io_outsHorizontal_1_7 = ces_7_7_io_outs_2; // @[MockArray.scala 52:89]
  assign io_outsVertical_0_0 = ces_0_7_io_outs_1; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_1 = ces_1_7_io_outs_1; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_2 = ces_2_7_io_outs_1; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_3 = ces_3_7_io_outs_1; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_4 = ces_4_7_io_outs_1; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_5 = ces_5_7_io_outs_1; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_6 = ces_6_7_io_outs_1; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_7 = ces_7_7_io_outs_1; // @[MockArray.scala 51:89]
  assign io_outsVertical_1_0 = ces_0_0_io_outs_3; // @[MockArray.scala 53:89]
  assign io_outsVertical_1_1 = ces_1_0_io_outs_3; // @[MockArray.scala 53:89]
  assign io_outsVertical_1_2 = ces_2_0_io_outs_3; // @[MockArray.scala 53:89]
  assign io_outsVertical_1_3 = ces_3_0_io_outs_3; // @[MockArray.scala 53:89]
  assign io_outsVertical_1_4 = ces_4_0_io_outs_3; // @[MockArray.scala 53:89]
  assign io_outsVertical_1_5 = ces_5_0_io_outs_3; // @[MockArray.scala 53:89]
  assign io_outsVertical_1_6 = ces_6_0_io_outs_3; // @[MockArray.scala 53:89]
  assign io_outsVertical_1_7 = ces_7_0_io_outs_3; // @[MockArray.scala 53:89]
  assign io_lsbs_0 = ces_0_0_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_1 = ces_0_1_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_2 = ces_0_2_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_3 = ces_0_3_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_4 = ces_0_4_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_5 = ces_0_5_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_6 = ces_0_6_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_7 = ces_0_7_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_8 = ces_1_0_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_9 = ces_1_1_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_10 = ces_1_2_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_11 = ces_1_3_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_12 = ces_1_4_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_13 = ces_1_5_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_14 = ces_1_6_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_15 = ces_1_7_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_16 = ces_2_0_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_17 = ces_2_1_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_18 = ces_2_2_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_19 = ces_2_3_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_20 = ces_2_4_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_21 = ces_2_5_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_22 = ces_2_6_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_23 = ces_2_7_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_24 = ces_3_0_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_25 = ces_3_1_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_26 = ces_3_2_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_27 = ces_3_3_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_28 = ces_3_4_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_29 = ces_3_5_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_30 = ces_3_6_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_31 = ces_3_7_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_32 = ces_4_0_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_33 = ces_4_1_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_34 = ces_4_2_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_35 = ces_4_3_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_36 = ces_4_4_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_37 = ces_4_5_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_38 = ces_4_6_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_39 = ces_4_7_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_40 = ces_5_0_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_41 = ces_5_1_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_42 = ces_5_2_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_43 = ces_5_3_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_44 = ces_5_4_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_45 = ces_5_5_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_46 = ces_5_6_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_47 = ces_5_7_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_48 = ces_6_0_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_49 = ces_6_1_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_50 = ces_6_2_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_51 = ces_6_3_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_52 = ces_6_4_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_53 = ces_6_5_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_54 = ces_6_6_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_55 = ces_6_7_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_56 = ces_7_0_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_57 = ces_7_1_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_58 = ces_7_2_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_59 = ces_7_3_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_60 = ces_7_4_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_61 = ces_7_5_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_62 = ces_7_6_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign io_lsbs_63 = ces_7_7_io_outs_0[0]; // @[MockArray.scala 39:44]
  assign ces_0_0_clock = clock;
  assign ces_0_0_io_ins_0 = io_insHorizontal_0_0; // @[MockArray.scala 45:87]
  assign ces_0_0_io_ins_1 = ces_0_1_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_0_0_io_ins_2 = ces_1_0_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_0_0_io_ins_3 = io_insVertical_1_0; // @[MockArray.scala 48:87]
  assign ces_0_1_clock = clock;
  assign ces_0_1_io_ins_0 = io_insHorizontal_0_1; // @[MockArray.scala 45:87]
  assign ces_0_1_io_ins_1 = ces_0_2_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_0_1_io_ins_2 = ces_1_1_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_0_1_io_ins_3 = ces_0_0_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_0_2_clock = clock;
  assign ces_0_2_io_ins_0 = io_insHorizontal_0_2; // @[MockArray.scala 45:87]
  assign ces_0_2_io_ins_1 = ces_0_3_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_0_2_io_ins_2 = ces_1_2_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_0_2_io_ins_3 = ces_0_1_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_0_3_clock = clock;
  assign ces_0_3_io_ins_0 = io_insHorizontal_0_3; // @[MockArray.scala 45:87]
  assign ces_0_3_io_ins_1 = ces_0_4_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_0_3_io_ins_2 = ces_1_3_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_0_3_io_ins_3 = ces_0_2_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_0_4_clock = clock;
  assign ces_0_4_io_ins_0 = io_insHorizontal_0_4; // @[MockArray.scala 45:87]
  assign ces_0_4_io_ins_1 = ces_0_5_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_0_4_io_ins_2 = ces_1_4_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_0_4_io_ins_3 = ces_0_3_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_0_5_clock = clock;
  assign ces_0_5_io_ins_0 = io_insHorizontal_0_5; // @[MockArray.scala 45:87]
  assign ces_0_5_io_ins_1 = ces_0_6_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_0_5_io_ins_2 = ces_1_5_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_0_5_io_ins_3 = ces_0_4_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_0_6_clock = clock;
  assign ces_0_6_io_ins_0 = io_insHorizontal_0_6; // @[MockArray.scala 45:87]
  assign ces_0_6_io_ins_1 = ces_0_7_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_0_6_io_ins_2 = ces_1_6_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_0_6_io_ins_3 = ces_0_5_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_0_7_clock = clock;
  assign ces_0_7_io_ins_0 = io_insHorizontal_0_7; // @[MockArray.scala 45:87]
  assign ces_0_7_io_ins_1 = io_insVertical_0_0; // @[MockArray.scala 46:87]
  assign ces_0_7_io_ins_2 = ces_1_7_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_0_7_io_ins_3 = ces_0_6_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_1_0_clock = clock;
  assign ces_1_0_io_ins_0 = ces_0_0_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_1_0_io_ins_1 = ces_1_1_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_1_0_io_ins_2 = ces_2_0_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_1_0_io_ins_3 = io_insVertical_1_1; // @[MockArray.scala 48:87]
  assign ces_1_1_clock = clock;
  assign ces_1_1_io_ins_0 = ces_0_1_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_1_1_io_ins_1 = ces_1_2_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_1_1_io_ins_2 = ces_2_1_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_1_1_io_ins_3 = ces_1_0_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_1_2_clock = clock;
  assign ces_1_2_io_ins_0 = ces_0_2_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_1_2_io_ins_1 = ces_1_3_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_1_2_io_ins_2 = ces_2_2_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_1_2_io_ins_3 = ces_1_1_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_1_3_clock = clock;
  assign ces_1_3_io_ins_0 = ces_0_3_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_1_3_io_ins_1 = ces_1_4_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_1_3_io_ins_2 = ces_2_3_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_1_3_io_ins_3 = ces_1_2_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_1_4_clock = clock;
  assign ces_1_4_io_ins_0 = ces_0_4_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_1_4_io_ins_1 = ces_1_5_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_1_4_io_ins_2 = ces_2_4_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_1_4_io_ins_3 = ces_1_3_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_1_5_clock = clock;
  assign ces_1_5_io_ins_0 = ces_0_5_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_1_5_io_ins_1 = ces_1_6_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_1_5_io_ins_2 = ces_2_5_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_1_5_io_ins_3 = ces_1_4_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_1_6_clock = clock;
  assign ces_1_6_io_ins_0 = ces_0_6_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_1_6_io_ins_1 = ces_1_7_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_1_6_io_ins_2 = ces_2_6_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_1_6_io_ins_3 = ces_1_5_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_1_7_clock = clock;
  assign ces_1_7_io_ins_0 = ces_0_7_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_1_7_io_ins_1 = io_insVertical_0_1; // @[MockArray.scala 46:87]
  assign ces_1_7_io_ins_2 = ces_2_7_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_1_7_io_ins_3 = ces_1_6_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_2_0_clock = clock;
  assign ces_2_0_io_ins_0 = ces_1_0_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_2_0_io_ins_1 = ces_2_1_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_2_0_io_ins_2 = ces_3_0_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_2_0_io_ins_3 = io_insVertical_1_2; // @[MockArray.scala 48:87]
  assign ces_2_1_clock = clock;
  assign ces_2_1_io_ins_0 = ces_1_1_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_2_1_io_ins_1 = ces_2_2_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_2_1_io_ins_2 = ces_3_1_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_2_1_io_ins_3 = ces_2_0_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_2_2_clock = clock;
  assign ces_2_2_io_ins_0 = ces_1_2_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_2_2_io_ins_1 = ces_2_3_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_2_2_io_ins_2 = ces_3_2_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_2_2_io_ins_3 = ces_2_1_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_2_3_clock = clock;
  assign ces_2_3_io_ins_0 = ces_1_3_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_2_3_io_ins_1 = ces_2_4_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_2_3_io_ins_2 = ces_3_3_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_2_3_io_ins_3 = ces_2_2_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_2_4_clock = clock;
  assign ces_2_4_io_ins_0 = ces_1_4_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_2_4_io_ins_1 = ces_2_5_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_2_4_io_ins_2 = ces_3_4_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_2_4_io_ins_3 = ces_2_3_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_2_5_clock = clock;
  assign ces_2_5_io_ins_0 = ces_1_5_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_2_5_io_ins_1 = ces_2_6_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_2_5_io_ins_2 = ces_3_5_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_2_5_io_ins_3 = ces_2_4_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_2_6_clock = clock;
  assign ces_2_6_io_ins_0 = ces_1_6_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_2_6_io_ins_1 = ces_2_7_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_2_6_io_ins_2 = ces_3_6_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_2_6_io_ins_3 = ces_2_5_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_2_7_clock = clock;
  assign ces_2_7_io_ins_0 = ces_1_7_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_2_7_io_ins_1 = io_insVertical_0_2; // @[MockArray.scala 46:87]
  assign ces_2_7_io_ins_2 = ces_3_7_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_2_7_io_ins_3 = ces_2_6_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_3_0_clock = clock;
  assign ces_3_0_io_ins_0 = ces_2_0_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_3_0_io_ins_1 = ces_3_1_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_3_0_io_ins_2 = ces_4_0_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_3_0_io_ins_3 = io_insVertical_1_3; // @[MockArray.scala 48:87]
  assign ces_3_1_clock = clock;
  assign ces_3_1_io_ins_0 = ces_2_1_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_3_1_io_ins_1 = ces_3_2_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_3_1_io_ins_2 = ces_4_1_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_3_1_io_ins_3 = ces_3_0_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_3_2_clock = clock;
  assign ces_3_2_io_ins_0 = ces_2_2_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_3_2_io_ins_1 = ces_3_3_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_3_2_io_ins_2 = ces_4_2_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_3_2_io_ins_3 = ces_3_1_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_3_3_clock = clock;
  assign ces_3_3_io_ins_0 = ces_2_3_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_3_3_io_ins_1 = ces_3_4_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_3_3_io_ins_2 = ces_4_3_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_3_3_io_ins_3 = ces_3_2_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_3_4_clock = clock;
  assign ces_3_4_io_ins_0 = ces_2_4_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_3_4_io_ins_1 = ces_3_5_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_3_4_io_ins_2 = ces_4_4_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_3_4_io_ins_3 = ces_3_3_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_3_5_clock = clock;
  assign ces_3_5_io_ins_0 = ces_2_5_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_3_5_io_ins_1 = ces_3_6_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_3_5_io_ins_2 = ces_4_5_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_3_5_io_ins_3 = ces_3_4_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_3_6_clock = clock;
  assign ces_3_6_io_ins_0 = ces_2_6_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_3_6_io_ins_1 = ces_3_7_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_3_6_io_ins_2 = ces_4_6_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_3_6_io_ins_3 = ces_3_5_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_3_7_clock = clock;
  assign ces_3_7_io_ins_0 = ces_2_7_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_3_7_io_ins_1 = io_insVertical_0_3; // @[MockArray.scala 46:87]
  assign ces_3_7_io_ins_2 = ces_4_7_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_3_7_io_ins_3 = ces_3_6_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_4_0_clock = clock;
  assign ces_4_0_io_ins_0 = ces_3_0_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_4_0_io_ins_1 = ces_4_1_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_4_0_io_ins_2 = ces_5_0_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_4_0_io_ins_3 = io_insVertical_1_4; // @[MockArray.scala 48:87]
  assign ces_4_1_clock = clock;
  assign ces_4_1_io_ins_0 = ces_3_1_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_4_1_io_ins_1 = ces_4_2_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_4_1_io_ins_2 = ces_5_1_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_4_1_io_ins_3 = ces_4_0_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_4_2_clock = clock;
  assign ces_4_2_io_ins_0 = ces_3_2_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_4_2_io_ins_1 = ces_4_3_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_4_2_io_ins_2 = ces_5_2_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_4_2_io_ins_3 = ces_4_1_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_4_3_clock = clock;
  assign ces_4_3_io_ins_0 = ces_3_3_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_4_3_io_ins_1 = ces_4_4_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_4_3_io_ins_2 = ces_5_3_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_4_3_io_ins_3 = ces_4_2_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_4_4_clock = clock;
  assign ces_4_4_io_ins_0 = ces_3_4_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_4_4_io_ins_1 = ces_4_5_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_4_4_io_ins_2 = ces_5_4_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_4_4_io_ins_3 = ces_4_3_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_4_5_clock = clock;
  assign ces_4_5_io_ins_0 = ces_3_5_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_4_5_io_ins_1 = ces_4_6_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_4_5_io_ins_2 = ces_5_5_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_4_5_io_ins_3 = ces_4_4_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_4_6_clock = clock;
  assign ces_4_6_io_ins_0 = ces_3_6_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_4_6_io_ins_1 = ces_4_7_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_4_6_io_ins_2 = ces_5_6_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_4_6_io_ins_3 = ces_4_5_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_4_7_clock = clock;
  assign ces_4_7_io_ins_0 = ces_3_7_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_4_7_io_ins_1 = io_insVertical_0_4; // @[MockArray.scala 46:87]
  assign ces_4_7_io_ins_2 = ces_5_7_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_4_7_io_ins_3 = ces_4_6_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_5_0_clock = clock;
  assign ces_5_0_io_ins_0 = ces_4_0_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_5_0_io_ins_1 = ces_5_1_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_5_0_io_ins_2 = ces_6_0_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_5_0_io_ins_3 = io_insVertical_1_5; // @[MockArray.scala 48:87]
  assign ces_5_1_clock = clock;
  assign ces_5_1_io_ins_0 = ces_4_1_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_5_1_io_ins_1 = ces_5_2_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_5_1_io_ins_2 = ces_6_1_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_5_1_io_ins_3 = ces_5_0_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_5_2_clock = clock;
  assign ces_5_2_io_ins_0 = ces_4_2_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_5_2_io_ins_1 = ces_5_3_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_5_2_io_ins_2 = ces_6_2_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_5_2_io_ins_3 = ces_5_1_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_5_3_clock = clock;
  assign ces_5_3_io_ins_0 = ces_4_3_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_5_3_io_ins_1 = ces_5_4_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_5_3_io_ins_2 = ces_6_3_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_5_3_io_ins_3 = ces_5_2_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_5_4_clock = clock;
  assign ces_5_4_io_ins_0 = ces_4_4_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_5_4_io_ins_1 = ces_5_5_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_5_4_io_ins_2 = ces_6_4_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_5_4_io_ins_3 = ces_5_3_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_5_5_clock = clock;
  assign ces_5_5_io_ins_0 = ces_4_5_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_5_5_io_ins_1 = ces_5_6_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_5_5_io_ins_2 = ces_6_5_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_5_5_io_ins_3 = ces_5_4_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_5_6_clock = clock;
  assign ces_5_6_io_ins_0 = ces_4_6_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_5_6_io_ins_1 = ces_5_7_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_5_6_io_ins_2 = ces_6_6_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_5_6_io_ins_3 = ces_5_5_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_5_7_clock = clock;
  assign ces_5_7_io_ins_0 = ces_4_7_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_5_7_io_ins_1 = io_insVertical_0_5; // @[MockArray.scala 46:87]
  assign ces_5_7_io_ins_2 = ces_6_7_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_5_7_io_ins_3 = ces_5_6_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_6_0_clock = clock;
  assign ces_6_0_io_ins_0 = ces_5_0_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_6_0_io_ins_1 = ces_6_1_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_6_0_io_ins_2 = ces_7_0_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_6_0_io_ins_3 = io_insVertical_1_6; // @[MockArray.scala 48:87]
  assign ces_6_1_clock = clock;
  assign ces_6_1_io_ins_0 = ces_5_1_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_6_1_io_ins_1 = ces_6_2_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_6_1_io_ins_2 = ces_7_1_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_6_1_io_ins_3 = ces_6_0_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_6_2_clock = clock;
  assign ces_6_2_io_ins_0 = ces_5_2_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_6_2_io_ins_1 = ces_6_3_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_6_2_io_ins_2 = ces_7_2_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_6_2_io_ins_3 = ces_6_1_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_6_3_clock = clock;
  assign ces_6_3_io_ins_0 = ces_5_3_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_6_3_io_ins_1 = ces_6_4_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_6_3_io_ins_2 = ces_7_3_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_6_3_io_ins_3 = ces_6_2_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_6_4_clock = clock;
  assign ces_6_4_io_ins_0 = ces_5_4_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_6_4_io_ins_1 = ces_6_5_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_6_4_io_ins_2 = ces_7_4_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_6_4_io_ins_3 = ces_6_3_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_6_5_clock = clock;
  assign ces_6_5_io_ins_0 = ces_5_5_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_6_5_io_ins_1 = ces_6_6_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_6_5_io_ins_2 = ces_7_5_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_6_5_io_ins_3 = ces_6_4_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_6_6_clock = clock;
  assign ces_6_6_io_ins_0 = ces_5_6_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_6_6_io_ins_1 = ces_6_7_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_6_6_io_ins_2 = ces_7_6_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_6_6_io_ins_3 = ces_6_5_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_6_7_clock = clock;
  assign ces_6_7_io_ins_0 = ces_5_7_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_6_7_io_ins_1 = io_insVertical_0_6; // @[MockArray.scala 46:87]
  assign ces_6_7_io_ins_2 = ces_7_7_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_6_7_io_ins_3 = ces_6_6_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_7_0_clock = clock;
  assign ces_7_0_io_ins_0 = ces_6_0_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_7_0_io_ins_1 = ces_7_1_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_7_0_io_ins_2 = io_insHorizontal_1_0; // @[MockArray.scala 47:87]
  assign ces_7_0_io_ins_3 = io_insVertical_1_7; // @[MockArray.scala 48:87]
  assign ces_7_1_clock = clock;
  assign ces_7_1_io_ins_0 = ces_6_1_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_7_1_io_ins_1 = ces_7_2_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_7_1_io_ins_2 = io_insHorizontal_1_1; // @[MockArray.scala 47:87]
  assign ces_7_1_io_ins_3 = ces_7_0_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_7_2_clock = clock;
  assign ces_7_2_io_ins_0 = ces_6_2_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_7_2_io_ins_1 = ces_7_3_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_7_2_io_ins_2 = io_insHorizontal_1_2; // @[MockArray.scala 47:87]
  assign ces_7_2_io_ins_3 = ces_7_1_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_7_3_clock = clock;
  assign ces_7_3_io_ins_0 = ces_6_3_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_7_3_io_ins_1 = ces_7_4_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_7_3_io_ins_2 = io_insHorizontal_1_3; // @[MockArray.scala 47:87]
  assign ces_7_3_io_ins_3 = ces_7_2_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_7_4_clock = clock;
  assign ces_7_4_io_ins_0 = ces_6_4_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_7_4_io_ins_1 = ces_7_5_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_7_4_io_ins_2 = io_insHorizontal_1_4; // @[MockArray.scala 47:87]
  assign ces_7_4_io_ins_3 = ces_7_3_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_7_5_clock = clock;
  assign ces_7_5_io_ins_0 = ces_6_5_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_7_5_io_ins_1 = ces_7_6_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_7_5_io_ins_2 = io_insHorizontal_1_5; // @[MockArray.scala 47:87]
  assign ces_7_5_io_ins_3 = ces_7_4_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_7_6_clock = clock;
  assign ces_7_6_io_ins_0 = ces_6_6_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_7_6_io_ins_1 = ces_7_7_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_7_6_io_ins_2 = io_insHorizontal_1_6; // @[MockArray.scala 47:87]
  assign ces_7_6_io_ins_3 = ces_7_5_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_7_7_clock = clock;
  assign ces_7_7_io_ins_0 = ces_6_7_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_7_7_io_ins_1 = io_insVertical_0_7; // @[MockArray.scala 46:87]
  assign ces_7_7_io_ins_2 = io_insHorizontal_1_7; // @[MockArray.scala 47:87]
  assign ces_7_7_io_ins_3 = ces_7_6_io_outs_1; // @[MockArray.scala 64:19]
endmodule
