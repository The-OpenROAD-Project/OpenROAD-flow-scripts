VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO DFFHQNV4Xx1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNV4Xx1_ASAP7_75t_L 0 0 ;
  SIZE 1.08 BY 1.08 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.126 0.29 0.144 ;
        RECT 0.234 0.225 0.271 0.243 ;
        RECT 0.234 0.027 0.271 0.045 ;
        RECT 0.234 0.027 0.252 0.243 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.396 0.29 0.414 ;
        RECT 0.234 0.495 0.271 0.513 ;
        RECT 0.234 0.297 0.271 0.315 ;
        RECT 0.234 0.297 0.252 0.513 ;
    END
  END D1
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.666 0.29 0.684 ;
        RECT 0.234 0.765 0.271 0.783 ;
        RECT 0.234 0.567 0.271 0.585 ;
        RECT 0.234 0.567 0.252 0.783 ;
    END
  END D2
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.936 0.29 0.954 ;
        RECT 0.234 1.035 0.271 1.053 ;
        RECT 0.234 0.837 0.271 0.855 ;
        RECT 0.234 0.837 0.252 1.053 ;
    END
  END D3
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.225 1.062 0.243 ;
        RECT 1.044 0.027 1.062 0.243 ;
        RECT 1.012 0.027 1.062 0.045 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.495 1.062 0.513 ;
        RECT 1.044 0.297 1.062 0.513 ;
        RECT 1.012 0.297 1.062 0.315 ;
    END
  END QN1
  PIN QN2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.765 1.062 0.783 ;
        RECT 1.044 0.567 1.062 0.783 ;
        RECT 1.012 0.567 1.062 0.585 ;
    END
  END QN2
  PIN QN3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 1.035 1.062 1.053 ;
        RECT 1.044 0.837 1.062 1.053 ;
        RECT 1.012 0.837 1.062 0.855 ;
    END
  END QN3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.08 0.279 ;
        RECT 0 0.801 1.08 0.819 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.08 0.009 ;
        RECT 0 0.531 1.08 0.549 ;
        RECT 0 1.071 1.08 1.089 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 0.04 0.07 0.122 0.088 ;
        RECT 0.04 0.452 0.122 0.47 ;
        RECT 0.04 0.61 0.122 0.628 ;
        RECT 0.04 0.992 0.122 1.01 ;
      LAYER M3 ;
        RECT 0.045 0.05 0.063 1.03 ;
      LAYER M1 ;
        RECT 0.099 0.164 0.117 0.236 ;
        RECT 0.072 0.07 0.117 0.106 ;
        RECT 0.099 0.034 0.117 0.106 ;
        RECT 0.072 0.164 0.117 0.2 ;
        RECT 0.072 0.07 0.09 0.2 ;
        RECT 0.099 0.434 0.117 0.506 ;
        RECT 0.072 0.34 0.117 0.376 ;
        RECT 0.099 0.304 0.117 0.376 ;
        RECT 0.072 0.434 0.117 0.47 ;
        RECT 0.072 0.34 0.09 0.47 ;
        RECT 0.099 0.704 0.117 0.776 ;
        RECT 0.072 0.61 0.117 0.646 ;
        RECT 0.099 0.574 0.117 0.646 ;
        RECT 0.072 0.704 0.117 0.74 ;
        RECT 0.072 0.61 0.09 0.74 ;
        RECT 0.099 0.974 0.117 1.046 ;
        RECT 0.072 0.88 0.117 0.916 ;
        RECT 0.099 0.844 0.117 0.916 ;
        RECT 0.072 0.974 0.117 1.01 ;
        RECT 0.072 0.88 0.09 1.01 ;
      LAYER V2 ;
        RECT 0.045 0.992 0.063 1.01 ;
        RECT 0.045 0.61 0.063 0.628 ;
        RECT 0.045 0.452 0.063 0.47 ;
        RECT 0.045 0.07 0.063 0.088 ;
      LAYER V1 ;
        RECT 0.099 0.992 0.117 1.01 ;
        RECT 0.099 0.61 0.117 0.628 ;
        RECT 0.099 0.452 0.117 0.47 ;
        RECT 0.099 0.07 0.117 0.088 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 0.85 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.774 0.027 0.792 0.119 ;
      RECT 0.774 0.027 0.954 0.045 ;
      RECT 0.774 0.495 0.954 0.513 ;
      RECT 0.936 0.297 0.954 0.513 ;
      RECT 0.774 0.421 0.792 0.513 ;
      RECT 0.85 0.297 0.954 0.315 ;
      RECT 0.85 0.765 0.954 0.783 ;
      RECT 0.936 0.567 0.954 0.783 ;
      RECT 0.774 0.567 0.792 0.659 ;
      RECT 0.774 0.567 0.954 0.585 ;
      RECT 0.774 1.035 0.954 1.053 ;
      RECT 0.936 0.837 0.954 1.053 ;
      RECT 0.774 0.961 0.792 1.053 ;
      RECT 0.85 0.837 0.954 0.855 ;
      RECT 0.688 0.224 0.738 0.242 ;
      RECT 0.72 0.027 0.738 0.242 ;
      RECT 0.72 0.153 0.9 0.171 ;
      RECT 0.882 0.117 0.9 0.171 ;
      RECT 0.828 0.117 0.846 0.171 ;
      RECT 0.634 0.027 0.738 0.045 ;
      RECT 0.634 0.495 0.738 0.513 ;
      RECT 0.72 0.298 0.738 0.513 ;
      RECT 0.882 0.369 0.9 0.423 ;
      RECT 0.828 0.369 0.846 0.423 ;
      RECT 0.72 0.369 0.9 0.387 ;
      RECT 0.688 0.298 0.738 0.316 ;
      RECT 0.688 0.764 0.738 0.782 ;
      RECT 0.72 0.567 0.738 0.782 ;
      RECT 0.72 0.693 0.9 0.711 ;
      RECT 0.882 0.657 0.9 0.711 ;
      RECT 0.828 0.657 0.846 0.711 ;
      RECT 0.634 0.567 0.738 0.585 ;
      RECT 0.634 1.035 0.738 1.053 ;
      RECT 0.72 0.838 0.738 1.053 ;
      RECT 0.882 0.909 0.9 0.963 ;
      RECT 0.828 0.909 0.846 0.963 ;
      RECT 0.72 0.909 0.9 0.927 ;
      RECT 0.688 0.838 0.738 0.856 ;
      RECT 0.576 0.225 0.63 0.243 ;
      RECT 0.612 0.081 0.63 0.243 ;
      RECT 0.496 0.081 0.63 0.099 ;
      RECT 0.585 0.045 0.603 0.099 ;
      RECT 0.585 0.441 0.603 0.495 ;
      RECT 0.496 0.441 0.63 0.459 ;
      RECT 0.612 0.297 0.63 0.459 ;
      RECT 0.576 0.297 0.63 0.315 ;
      RECT 0.576 0.765 0.63 0.783 ;
      RECT 0.612 0.621 0.63 0.783 ;
      RECT 0.496 0.621 0.63 0.639 ;
      RECT 0.585 0.585 0.603 0.639 ;
      RECT 0.585 0.981 0.603 1.035 ;
      RECT 0.496 0.981 0.63 0.999 ;
      RECT 0.612 0.837 0.63 0.999 ;
      RECT 0.576 0.837 0.63 0.855 ;
      RECT 0.364 0.225 0.468 0.243 ;
      RECT 0.45 0.027 0.468 0.243 ;
      RECT 0.45 0.122 0.576 0.14 ;
      RECT 0.418 0.027 0.468 0.045 ;
      RECT 0.418 0.495 0.468 0.513 ;
      RECT 0.45 0.297 0.468 0.513 ;
      RECT 0.45 0.4 0.576 0.418 ;
      RECT 0.364 0.297 0.468 0.315 ;
      RECT 0.364 0.765 0.468 0.783 ;
      RECT 0.45 0.567 0.468 0.783 ;
      RECT 0.45 0.662 0.576 0.68 ;
      RECT 0.418 0.567 0.468 0.585 ;
      RECT 0.418 1.035 0.468 1.053 ;
      RECT 0.45 0.837 0.468 1.053 ;
      RECT 0.45 0.94 0.576 0.958 ;
      RECT 0.364 0.837 0.468 0.855 ;
      RECT 0.315 0.126 0.333 0.203 ;
      RECT 0.315 0.126 0.367 0.144 ;
      RECT 0.315 0.396 0.367 0.414 ;
      RECT 0.315 0.337 0.333 0.414 ;
      RECT 0.315 0.666 0.333 0.743 ;
      RECT 0.315 0.666 0.367 0.684 ;
      RECT 0.315 0.936 0.367 0.954 ;
      RECT 0.315 0.877 0.333 0.954 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.148 0.495 0.198 0.513 ;
      RECT 0.18 0.297 0.198 0.513 ;
      RECT 0.148 0.297 0.198 0.315 ;
      RECT 0.148 0.765 0.198 0.783 ;
      RECT 0.18 0.567 0.198 0.783 ;
      RECT 0.148 0.567 0.198 0.585 ;
      RECT 0.148 1.035 0.198 1.053 ;
      RECT 0.18 0.837 0.198 1.053 ;
      RECT 0.148 0.837 0.198 0.855 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.144 0.047 0.162 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 0.009 0.495 0.068 0.513 ;
      RECT 0.009 0.297 0.027 0.513 ;
      RECT 0.009 0.378 0.047 0.396 ;
      RECT 0.009 0.297 0.068 0.315 ;
      RECT 0.009 0.765 0.068 0.783 ;
      RECT 0.009 0.567 0.027 0.783 ;
      RECT 0.009 0.684 0.047 0.702 ;
      RECT 0.009 0.567 0.068 0.585 ;
      RECT 0.009 1.035 0.068 1.053 ;
      RECT 0.009 0.837 0.027 1.053 ;
      RECT 0.009 0.918 0.047 0.936 ;
      RECT 0.009 0.837 0.068 0.855 ;
      RECT 0.99 0.09 1.008 0.167 ;
      RECT 0.99 0.373 1.008 0.45 ;
      RECT 0.99 0.63 1.008 0.707 ;
      RECT 0.99 0.913 1.008 0.99 ;
      RECT 0.666 0.101 0.684 0.167 ;
      RECT 0.666 0.373 0.684 0.439 ;
      RECT 0.666 0.641 0.684 0.707 ;
      RECT 0.666 0.913 0.684 0.979 ;
      RECT 0.504 0.165 0.522 0.203 ;
      RECT 0.504 0.337 0.522 0.375 ;
      RECT 0.504 0.705 0.522 0.743 ;
      RECT 0.504 0.877 0.522 0.915 ;
      RECT 0.396 0.106 0.414 0.167 ;
      RECT 0.396 0.373 0.414 0.434 ;
      RECT 0.396 0.646 0.414 0.707 ;
      RECT 0.396 0.913 0.414 0.974 ;
      RECT 0.142 0.106 0.16 0.167 ;
      RECT 0.142 0.373 0.16 0.434 ;
      RECT 0.142 0.646 0.16 0.707 ;
      RECT 0.142 0.913 0.16 0.974 ;
    LAYER M2 ;
      RECT 0.877 0.144 1.013 0.162 ;
      RECT 0.877 0.378 1.013 0.396 ;
      RECT 0.877 0.684 1.013 0.702 ;
      RECT 0.877 0.918 1.013 0.936 ;
      RECT 0.019 0.144 0.689 0.162 ;
      RECT 0.019 0.378 0.689 0.396 ;
      RECT 0.019 0.684 0.689 0.702 ;
      RECT 0.019 0.918 0.689 0.936 ;
      RECT 0.175 0.18 0.527 0.198 ;
      RECT 0.175 0.342 0.527 0.36 ;
      RECT 0.175 0.72 0.527 0.738 ;
      RECT 0.175 0.882 0.527 0.9 ;
    LAYER V1 ;
      RECT 0.99 0.144 1.008 0.162 ;
      RECT 0.99 0.378 1.008 0.396 ;
      RECT 0.99 0.684 1.008 0.702 ;
      RECT 0.99 0.918 1.008 0.936 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.882 0.378 0.9 0.396 ;
      RECT 0.882 0.684 0.9 0.702 ;
      RECT 0.882 0.918 0.9 0.936 ;
      RECT 0.666 0.144 0.684 0.162 ;
      RECT 0.666 0.378 0.684 0.396 ;
      RECT 0.666 0.684 0.684 0.702 ;
      RECT 0.666 0.918 0.684 0.936 ;
      RECT 0.504 0.18 0.522 0.198 ;
      RECT 0.504 0.342 0.522 0.36 ;
      RECT 0.504 0.72 0.522 0.738 ;
      RECT 0.504 0.882 0.522 0.9 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.396 0.378 0.414 0.396 ;
      RECT 0.396 0.684 0.414 0.702 ;
      RECT 0.396 0.918 0.414 0.936 ;
      RECT 0.315 0.18 0.333 0.198 ;
      RECT 0.315 0.342 0.333 0.36 ;
      RECT 0.315 0.72 0.333 0.738 ;
      RECT 0.315 0.882 0.333 0.9 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.18 0.342 0.198 0.36 ;
      RECT 0.18 0.72 0.198 0.738 ;
      RECT 0.18 0.882 0.198 0.9 ;
      RECT 0.142 0.144 0.16 0.162 ;
      RECT 0.142 0.378 0.16 0.396 ;
      RECT 0.142 0.684 0.16 0.702 ;
      RECT 0.142 0.918 0.16 0.936 ;
      RECT 0.024 0.144 0.042 0.162 ;
      RECT 0.024 0.378 0.042 0.396 ;
      RECT 0.024 0.684 0.042 0.702 ;
      RECT 0.024 0.918 0.042 0.936 ;
  END
END DFFHQNV4Xx1_ASAP7_75t_L

MACRO DFFHQNV4Xx1_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNV4Xx1_ASAP7_75t_R 0 0 ;
  SIZE 1.08 BY 1.08 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.126 0.29 0.144 ;
        RECT 0.234 0.225 0.271 0.243 ;
        RECT 0.234 0.027 0.271 0.045 ;
        RECT 0.234 0.027 0.252 0.243 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.396 0.29 0.414 ;
        RECT 0.234 0.495 0.271 0.513 ;
        RECT 0.234 0.297 0.271 0.315 ;
        RECT 0.234 0.297 0.252 0.513 ;
    END
  END D1
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.666 0.29 0.684 ;
        RECT 0.234 0.765 0.271 0.783 ;
        RECT 0.234 0.567 0.271 0.585 ;
        RECT 0.234 0.567 0.252 0.783 ;
    END
  END D2
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.936 0.29 0.954 ;
        RECT 0.234 1.035 0.271 1.053 ;
        RECT 0.234 0.837 0.271 0.855 ;
        RECT 0.234 0.837 0.252 1.053 ;
    END
  END D3
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.225 1.062 0.243 ;
        RECT 1.044 0.027 1.062 0.243 ;
        RECT 1.012 0.027 1.062 0.045 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.495 1.062 0.513 ;
        RECT 1.044 0.297 1.062 0.513 ;
        RECT 1.012 0.297 1.062 0.315 ;
    END
  END QN1
  PIN QN2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.765 1.062 0.783 ;
        RECT 1.044 0.567 1.062 0.783 ;
        RECT 1.012 0.567 1.062 0.585 ;
    END
  END QN2
  PIN QN3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 1.035 1.062 1.053 ;
        RECT 1.044 0.837 1.062 1.053 ;
        RECT 1.012 0.837 1.062 0.855 ;
    END
  END QN3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.08 0.279 ;
        RECT 0 0.801 1.08 0.819 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.08 0.009 ;
        RECT 0 0.531 1.08 0.549 ;
        RECT 0 1.071 1.08 1.089 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 0.04 0.07 0.122 0.088 ;
        RECT 0.04 0.452 0.122 0.47 ;
        RECT 0.04 0.61 0.122 0.628 ;
        RECT 0.04 0.992 0.122 1.01 ;
      LAYER M3 ;
        RECT 0.045 0.05 0.063 1.03 ;
      LAYER M1 ;
        RECT 0.099 0.164 0.117 0.236 ;
        RECT 0.072 0.07 0.117 0.106 ;
        RECT 0.099 0.034 0.117 0.106 ;
        RECT 0.072 0.164 0.117 0.2 ;
        RECT 0.072 0.07 0.09 0.2 ;
        RECT 0.099 0.434 0.117 0.506 ;
        RECT 0.072 0.34 0.117 0.376 ;
        RECT 0.099 0.304 0.117 0.376 ;
        RECT 0.072 0.434 0.117 0.47 ;
        RECT 0.072 0.34 0.09 0.47 ;
        RECT 0.099 0.704 0.117 0.776 ;
        RECT 0.072 0.61 0.117 0.646 ;
        RECT 0.099 0.574 0.117 0.646 ;
        RECT 0.072 0.704 0.117 0.74 ;
        RECT 0.072 0.61 0.09 0.74 ;
        RECT 0.099 0.974 0.117 1.046 ;
        RECT 0.072 0.88 0.117 0.916 ;
        RECT 0.099 0.844 0.117 0.916 ;
        RECT 0.072 0.974 0.117 1.01 ;
        RECT 0.072 0.88 0.09 1.01 ;
      LAYER V2 ;
        RECT 0.045 0.992 0.063 1.01 ;
        RECT 0.045 0.61 0.063 0.628 ;
        RECT 0.045 0.452 0.063 0.47 ;
        RECT 0.045 0.07 0.063 0.088 ;
      LAYER V1 ;
        RECT 0.099 0.992 0.117 1.01 ;
        RECT 0.099 0.61 0.117 0.628 ;
        RECT 0.099 0.452 0.117 0.47 ;
        RECT 0.099 0.07 0.117 0.088 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 0.85 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.774 0.027 0.792 0.119 ;
      RECT 0.774 0.027 0.954 0.045 ;
      RECT 0.774 0.495 0.954 0.513 ;
      RECT 0.936 0.297 0.954 0.513 ;
      RECT 0.774 0.421 0.792 0.513 ;
      RECT 0.85 0.297 0.954 0.315 ;
      RECT 0.85 0.765 0.954 0.783 ;
      RECT 0.936 0.567 0.954 0.783 ;
      RECT 0.774 0.567 0.792 0.659 ;
      RECT 0.774 0.567 0.954 0.585 ;
      RECT 0.774 1.035 0.954 1.053 ;
      RECT 0.936 0.837 0.954 1.053 ;
      RECT 0.774 0.961 0.792 1.053 ;
      RECT 0.85 0.837 0.954 0.855 ;
      RECT 0.688 0.224 0.738 0.242 ;
      RECT 0.72 0.027 0.738 0.242 ;
      RECT 0.72 0.153 0.9 0.171 ;
      RECT 0.882 0.117 0.9 0.171 ;
      RECT 0.828 0.117 0.846 0.171 ;
      RECT 0.634 0.027 0.738 0.045 ;
      RECT 0.634 0.495 0.738 0.513 ;
      RECT 0.72 0.298 0.738 0.513 ;
      RECT 0.882 0.369 0.9 0.423 ;
      RECT 0.828 0.369 0.846 0.423 ;
      RECT 0.72 0.369 0.9 0.387 ;
      RECT 0.688 0.298 0.738 0.316 ;
      RECT 0.688 0.764 0.738 0.782 ;
      RECT 0.72 0.567 0.738 0.782 ;
      RECT 0.72 0.693 0.9 0.711 ;
      RECT 0.882 0.657 0.9 0.711 ;
      RECT 0.828 0.657 0.846 0.711 ;
      RECT 0.634 0.567 0.738 0.585 ;
      RECT 0.634 1.035 0.738 1.053 ;
      RECT 0.72 0.838 0.738 1.053 ;
      RECT 0.882 0.909 0.9 0.963 ;
      RECT 0.828 0.909 0.846 0.963 ;
      RECT 0.72 0.909 0.9 0.927 ;
      RECT 0.688 0.838 0.738 0.856 ;
      RECT 0.576 0.225 0.63 0.243 ;
      RECT 0.612 0.081 0.63 0.243 ;
      RECT 0.496 0.081 0.63 0.099 ;
      RECT 0.585 0.045 0.603 0.099 ;
      RECT 0.585 0.441 0.603 0.495 ;
      RECT 0.496 0.441 0.63 0.459 ;
      RECT 0.612 0.297 0.63 0.459 ;
      RECT 0.576 0.297 0.63 0.315 ;
      RECT 0.576 0.765 0.63 0.783 ;
      RECT 0.612 0.621 0.63 0.783 ;
      RECT 0.496 0.621 0.63 0.639 ;
      RECT 0.585 0.585 0.603 0.639 ;
      RECT 0.585 0.981 0.603 1.035 ;
      RECT 0.496 0.981 0.63 0.999 ;
      RECT 0.612 0.837 0.63 0.999 ;
      RECT 0.576 0.837 0.63 0.855 ;
      RECT 0.364 0.225 0.468 0.243 ;
      RECT 0.45 0.027 0.468 0.243 ;
      RECT 0.45 0.122 0.576 0.14 ;
      RECT 0.418 0.027 0.468 0.045 ;
      RECT 0.418 0.495 0.468 0.513 ;
      RECT 0.45 0.297 0.468 0.513 ;
      RECT 0.45 0.4 0.576 0.418 ;
      RECT 0.364 0.297 0.468 0.315 ;
      RECT 0.364 0.765 0.468 0.783 ;
      RECT 0.45 0.567 0.468 0.783 ;
      RECT 0.45 0.662 0.576 0.68 ;
      RECT 0.418 0.567 0.468 0.585 ;
      RECT 0.418 1.035 0.468 1.053 ;
      RECT 0.45 0.837 0.468 1.053 ;
      RECT 0.45 0.94 0.576 0.958 ;
      RECT 0.364 0.837 0.468 0.855 ;
      RECT 0.315 0.126 0.333 0.203 ;
      RECT 0.315 0.126 0.367 0.144 ;
      RECT 0.315 0.396 0.367 0.414 ;
      RECT 0.315 0.337 0.333 0.414 ;
      RECT 0.315 0.666 0.333 0.743 ;
      RECT 0.315 0.666 0.367 0.684 ;
      RECT 0.315 0.936 0.367 0.954 ;
      RECT 0.315 0.877 0.333 0.954 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.148 0.495 0.198 0.513 ;
      RECT 0.18 0.297 0.198 0.513 ;
      RECT 0.148 0.297 0.198 0.315 ;
      RECT 0.148 0.765 0.198 0.783 ;
      RECT 0.18 0.567 0.198 0.783 ;
      RECT 0.148 0.567 0.198 0.585 ;
      RECT 0.148 1.035 0.198 1.053 ;
      RECT 0.18 0.837 0.198 1.053 ;
      RECT 0.148 0.837 0.198 0.855 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.144 0.047 0.162 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 0.009 0.495 0.068 0.513 ;
      RECT 0.009 0.297 0.027 0.513 ;
      RECT 0.009 0.378 0.047 0.396 ;
      RECT 0.009 0.297 0.068 0.315 ;
      RECT 0.009 0.765 0.068 0.783 ;
      RECT 0.009 0.567 0.027 0.783 ;
      RECT 0.009 0.684 0.047 0.702 ;
      RECT 0.009 0.567 0.068 0.585 ;
      RECT 0.009 1.035 0.068 1.053 ;
      RECT 0.009 0.837 0.027 1.053 ;
      RECT 0.009 0.918 0.047 0.936 ;
      RECT 0.009 0.837 0.068 0.855 ;
      RECT 0.99 0.09 1.008 0.167 ;
      RECT 0.99 0.373 1.008 0.45 ;
      RECT 0.99 0.63 1.008 0.707 ;
      RECT 0.99 0.913 1.008 0.99 ;
      RECT 0.666 0.101 0.684 0.167 ;
      RECT 0.666 0.373 0.684 0.439 ;
      RECT 0.666 0.641 0.684 0.707 ;
      RECT 0.666 0.913 0.684 0.979 ;
      RECT 0.504 0.165 0.522 0.203 ;
      RECT 0.504 0.337 0.522 0.375 ;
      RECT 0.504 0.705 0.522 0.743 ;
      RECT 0.504 0.877 0.522 0.915 ;
      RECT 0.396 0.106 0.414 0.167 ;
      RECT 0.396 0.373 0.414 0.434 ;
      RECT 0.396 0.646 0.414 0.707 ;
      RECT 0.396 0.913 0.414 0.974 ;
      RECT 0.142 0.106 0.16 0.167 ;
      RECT 0.142 0.373 0.16 0.434 ;
      RECT 0.142 0.646 0.16 0.707 ;
      RECT 0.142 0.913 0.16 0.974 ;
    LAYER M2 ;
      RECT 0.877 0.144 1.013 0.162 ;
      RECT 0.877 0.378 1.013 0.396 ;
      RECT 0.877 0.684 1.013 0.702 ;
      RECT 0.877 0.918 1.013 0.936 ;
      RECT 0.019 0.144 0.689 0.162 ;
      RECT 0.019 0.378 0.689 0.396 ;
      RECT 0.019 0.684 0.689 0.702 ;
      RECT 0.019 0.918 0.689 0.936 ;
      RECT 0.175 0.18 0.527 0.198 ;
      RECT 0.175 0.342 0.527 0.36 ;
      RECT 0.175 0.72 0.527 0.738 ;
      RECT 0.175 0.882 0.527 0.9 ;
    LAYER V1 ;
      RECT 0.99 0.144 1.008 0.162 ;
      RECT 0.99 0.378 1.008 0.396 ;
      RECT 0.99 0.684 1.008 0.702 ;
      RECT 0.99 0.918 1.008 0.936 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.882 0.378 0.9 0.396 ;
      RECT 0.882 0.684 0.9 0.702 ;
      RECT 0.882 0.918 0.9 0.936 ;
      RECT 0.666 0.144 0.684 0.162 ;
      RECT 0.666 0.378 0.684 0.396 ;
      RECT 0.666 0.684 0.684 0.702 ;
      RECT 0.666 0.918 0.684 0.936 ;
      RECT 0.504 0.18 0.522 0.198 ;
      RECT 0.504 0.342 0.522 0.36 ;
      RECT 0.504 0.72 0.522 0.738 ;
      RECT 0.504 0.882 0.522 0.9 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.396 0.378 0.414 0.396 ;
      RECT 0.396 0.684 0.414 0.702 ;
      RECT 0.396 0.918 0.414 0.936 ;
      RECT 0.315 0.18 0.333 0.198 ;
      RECT 0.315 0.342 0.333 0.36 ;
      RECT 0.315 0.72 0.333 0.738 ;
      RECT 0.315 0.882 0.333 0.9 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.18 0.342 0.198 0.36 ;
      RECT 0.18 0.72 0.198 0.738 ;
      RECT 0.18 0.882 0.198 0.9 ;
      RECT 0.142 0.144 0.16 0.162 ;
      RECT 0.142 0.378 0.16 0.396 ;
      RECT 0.142 0.684 0.16 0.702 ;
      RECT 0.142 0.918 0.16 0.936 ;
      RECT 0.024 0.144 0.042 0.162 ;
      RECT 0.024 0.378 0.042 0.396 ;
      RECT 0.024 0.684 0.042 0.702 ;
      RECT 0.024 0.918 0.042 0.936 ;
  END
END DFFHQNV4Xx1_ASAP7_75t_R

MACRO DFFHQNV4Xx1_ASAP7_75t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNV4Xx1_ASAP7_75t_SL 0 0 ;
  SIZE 1.08 BY 1.08 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.126 0.29 0.144 ;
        RECT 0.234 0.225 0.271 0.243 ;
        RECT 0.234 0.027 0.271 0.045 ;
        RECT 0.234 0.027 0.252 0.243 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.396 0.29 0.414 ;
        RECT 0.234 0.495 0.271 0.513 ;
        RECT 0.234 0.297 0.271 0.315 ;
        RECT 0.234 0.297 0.252 0.513 ;
    END
  END D1
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.666 0.29 0.684 ;
        RECT 0.234 0.765 0.271 0.783 ;
        RECT 0.234 0.567 0.271 0.585 ;
        RECT 0.234 0.567 0.252 0.783 ;
    END
  END D2
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.936 0.29 0.954 ;
        RECT 0.234 1.035 0.271 1.053 ;
        RECT 0.234 0.837 0.271 0.855 ;
        RECT 0.234 0.837 0.252 1.053 ;
    END
  END D3
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.225 1.062 0.243 ;
        RECT 1.044 0.027 1.062 0.243 ;
        RECT 1.012 0.027 1.062 0.045 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.495 1.062 0.513 ;
        RECT 1.044 0.297 1.062 0.513 ;
        RECT 1.012 0.297 1.062 0.315 ;
    END
  END QN1
  PIN QN2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.765 1.062 0.783 ;
        RECT 1.044 0.567 1.062 0.783 ;
        RECT 1.012 0.567 1.062 0.585 ;
    END
  END QN2
  PIN QN3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 1.035 1.062 1.053 ;
        RECT 1.044 0.837 1.062 1.053 ;
        RECT 1.012 0.837 1.062 0.855 ;
    END
  END QN3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.08 0.279 ;
        RECT 0 0.801 1.08 0.819 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.08 0.009 ;
        RECT 0 0.531 1.08 0.549 ;
        RECT 0 1.071 1.08 1.089 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 0.04 0.07 0.122 0.088 ;
        RECT 0.04 0.452 0.122 0.47 ;
        RECT 0.04 0.61 0.122 0.628 ;
        RECT 0.04 0.992 0.122 1.01 ;
      LAYER M3 ;
        RECT 0.045 0.05 0.063 1.03 ;
      LAYER M1 ;
        RECT 0.099 0.164 0.117 0.236 ;
        RECT 0.072 0.07 0.117 0.106 ;
        RECT 0.099 0.034 0.117 0.106 ;
        RECT 0.072 0.164 0.117 0.2 ;
        RECT 0.072 0.07 0.09 0.2 ;
        RECT 0.099 0.434 0.117 0.506 ;
        RECT 0.072 0.34 0.117 0.376 ;
        RECT 0.099 0.304 0.117 0.376 ;
        RECT 0.072 0.434 0.117 0.47 ;
        RECT 0.072 0.34 0.09 0.47 ;
        RECT 0.099 0.704 0.117 0.776 ;
        RECT 0.072 0.61 0.117 0.646 ;
        RECT 0.099 0.574 0.117 0.646 ;
        RECT 0.072 0.704 0.117 0.74 ;
        RECT 0.072 0.61 0.09 0.74 ;
        RECT 0.099 0.974 0.117 1.046 ;
        RECT 0.072 0.88 0.117 0.916 ;
        RECT 0.099 0.844 0.117 0.916 ;
        RECT 0.072 0.974 0.117 1.01 ;
        RECT 0.072 0.88 0.09 1.01 ;
      LAYER V2 ;
        RECT 0.045 0.992 0.063 1.01 ;
        RECT 0.045 0.61 0.063 0.628 ;
        RECT 0.045 0.452 0.063 0.47 ;
        RECT 0.045 0.07 0.063 0.088 ;
      LAYER V1 ;
        RECT 0.099 0.992 0.117 1.01 ;
        RECT 0.099 0.61 0.117 0.628 ;
        RECT 0.099 0.452 0.117 0.47 ;
        RECT 0.099 0.07 0.117 0.088 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 0.85 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.774 0.027 0.792 0.119 ;
      RECT 0.774 0.027 0.954 0.045 ;
      RECT 0.774 0.495 0.954 0.513 ;
      RECT 0.936 0.297 0.954 0.513 ;
      RECT 0.774 0.421 0.792 0.513 ;
      RECT 0.85 0.297 0.954 0.315 ;
      RECT 0.85 0.765 0.954 0.783 ;
      RECT 0.936 0.567 0.954 0.783 ;
      RECT 0.774 0.567 0.792 0.659 ;
      RECT 0.774 0.567 0.954 0.585 ;
      RECT 0.774 1.035 0.954 1.053 ;
      RECT 0.936 0.837 0.954 1.053 ;
      RECT 0.774 0.961 0.792 1.053 ;
      RECT 0.85 0.837 0.954 0.855 ;
      RECT 0.688 0.224 0.738 0.242 ;
      RECT 0.72 0.027 0.738 0.242 ;
      RECT 0.72 0.153 0.9 0.171 ;
      RECT 0.882 0.117 0.9 0.171 ;
      RECT 0.828 0.117 0.846 0.171 ;
      RECT 0.634 0.027 0.738 0.045 ;
      RECT 0.634 0.495 0.738 0.513 ;
      RECT 0.72 0.298 0.738 0.513 ;
      RECT 0.882 0.369 0.9 0.423 ;
      RECT 0.828 0.369 0.846 0.423 ;
      RECT 0.72 0.369 0.9 0.387 ;
      RECT 0.688 0.298 0.738 0.316 ;
      RECT 0.688 0.764 0.738 0.782 ;
      RECT 0.72 0.567 0.738 0.782 ;
      RECT 0.72 0.693 0.9 0.711 ;
      RECT 0.882 0.657 0.9 0.711 ;
      RECT 0.828 0.657 0.846 0.711 ;
      RECT 0.634 0.567 0.738 0.585 ;
      RECT 0.634 1.035 0.738 1.053 ;
      RECT 0.72 0.838 0.738 1.053 ;
      RECT 0.882 0.909 0.9 0.963 ;
      RECT 0.828 0.909 0.846 0.963 ;
      RECT 0.72 0.909 0.9 0.927 ;
      RECT 0.688 0.838 0.738 0.856 ;
      RECT 0.576 0.225 0.63 0.243 ;
      RECT 0.612 0.081 0.63 0.243 ;
      RECT 0.496 0.081 0.63 0.099 ;
      RECT 0.585 0.045 0.603 0.099 ;
      RECT 0.585 0.441 0.603 0.495 ;
      RECT 0.496 0.441 0.63 0.459 ;
      RECT 0.612 0.297 0.63 0.459 ;
      RECT 0.576 0.297 0.63 0.315 ;
      RECT 0.576 0.765 0.63 0.783 ;
      RECT 0.612 0.621 0.63 0.783 ;
      RECT 0.496 0.621 0.63 0.639 ;
      RECT 0.585 0.585 0.603 0.639 ;
      RECT 0.585 0.981 0.603 1.035 ;
      RECT 0.496 0.981 0.63 0.999 ;
      RECT 0.612 0.837 0.63 0.999 ;
      RECT 0.576 0.837 0.63 0.855 ;
      RECT 0.364 0.225 0.468 0.243 ;
      RECT 0.45 0.027 0.468 0.243 ;
      RECT 0.45 0.122 0.576 0.14 ;
      RECT 0.418 0.027 0.468 0.045 ;
      RECT 0.418 0.495 0.468 0.513 ;
      RECT 0.45 0.297 0.468 0.513 ;
      RECT 0.45 0.4 0.576 0.418 ;
      RECT 0.364 0.297 0.468 0.315 ;
      RECT 0.364 0.765 0.468 0.783 ;
      RECT 0.45 0.567 0.468 0.783 ;
      RECT 0.45 0.662 0.576 0.68 ;
      RECT 0.418 0.567 0.468 0.585 ;
      RECT 0.418 1.035 0.468 1.053 ;
      RECT 0.45 0.837 0.468 1.053 ;
      RECT 0.45 0.94 0.576 0.958 ;
      RECT 0.364 0.837 0.468 0.855 ;
      RECT 0.315 0.126 0.333 0.203 ;
      RECT 0.315 0.126 0.367 0.144 ;
      RECT 0.315 0.396 0.367 0.414 ;
      RECT 0.315 0.337 0.333 0.414 ;
      RECT 0.315 0.666 0.333 0.743 ;
      RECT 0.315 0.666 0.367 0.684 ;
      RECT 0.315 0.936 0.367 0.954 ;
      RECT 0.315 0.877 0.333 0.954 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.148 0.495 0.198 0.513 ;
      RECT 0.18 0.297 0.198 0.513 ;
      RECT 0.148 0.297 0.198 0.315 ;
      RECT 0.148 0.765 0.198 0.783 ;
      RECT 0.18 0.567 0.198 0.783 ;
      RECT 0.148 0.567 0.198 0.585 ;
      RECT 0.148 1.035 0.198 1.053 ;
      RECT 0.18 0.837 0.198 1.053 ;
      RECT 0.148 0.837 0.198 0.855 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.144 0.047 0.162 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 0.009 0.495 0.068 0.513 ;
      RECT 0.009 0.297 0.027 0.513 ;
      RECT 0.009 0.378 0.047 0.396 ;
      RECT 0.009 0.297 0.068 0.315 ;
      RECT 0.009 0.765 0.068 0.783 ;
      RECT 0.009 0.567 0.027 0.783 ;
      RECT 0.009 0.684 0.047 0.702 ;
      RECT 0.009 0.567 0.068 0.585 ;
      RECT 0.009 1.035 0.068 1.053 ;
      RECT 0.009 0.837 0.027 1.053 ;
      RECT 0.009 0.918 0.047 0.936 ;
      RECT 0.009 0.837 0.068 0.855 ;
      RECT 0.99 0.09 1.008 0.167 ;
      RECT 0.99 0.373 1.008 0.45 ;
      RECT 0.99 0.63 1.008 0.707 ;
      RECT 0.99 0.913 1.008 0.99 ;
      RECT 0.666 0.101 0.684 0.167 ;
      RECT 0.666 0.373 0.684 0.439 ;
      RECT 0.666 0.641 0.684 0.707 ;
      RECT 0.666 0.913 0.684 0.979 ;
      RECT 0.504 0.165 0.522 0.203 ;
      RECT 0.504 0.337 0.522 0.375 ;
      RECT 0.504 0.705 0.522 0.743 ;
      RECT 0.504 0.877 0.522 0.915 ;
      RECT 0.396 0.106 0.414 0.167 ;
      RECT 0.396 0.373 0.414 0.434 ;
      RECT 0.396 0.646 0.414 0.707 ;
      RECT 0.396 0.913 0.414 0.974 ;
      RECT 0.142 0.106 0.16 0.167 ;
      RECT 0.142 0.373 0.16 0.434 ;
      RECT 0.142 0.646 0.16 0.707 ;
      RECT 0.142 0.913 0.16 0.974 ;
    LAYER M2 ;
      RECT 0.877 0.144 1.013 0.162 ;
      RECT 0.877 0.378 1.013 0.396 ;
      RECT 0.877 0.684 1.013 0.702 ;
      RECT 0.877 0.918 1.013 0.936 ;
      RECT 0.019 0.144 0.689 0.162 ;
      RECT 0.019 0.378 0.689 0.396 ;
      RECT 0.019 0.684 0.689 0.702 ;
      RECT 0.019 0.918 0.689 0.936 ;
      RECT 0.175 0.18 0.527 0.198 ;
      RECT 0.175 0.342 0.527 0.36 ;
      RECT 0.175 0.72 0.527 0.738 ;
      RECT 0.175 0.882 0.527 0.9 ;
    LAYER V1 ;
      RECT 0.99 0.144 1.008 0.162 ;
      RECT 0.99 0.378 1.008 0.396 ;
      RECT 0.99 0.684 1.008 0.702 ;
      RECT 0.99 0.918 1.008 0.936 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.882 0.378 0.9 0.396 ;
      RECT 0.882 0.684 0.9 0.702 ;
      RECT 0.882 0.918 0.9 0.936 ;
      RECT 0.666 0.144 0.684 0.162 ;
      RECT 0.666 0.378 0.684 0.396 ;
      RECT 0.666 0.684 0.684 0.702 ;
      RECT 0.666 0.918 0.684 0.936 ;
      RECT 0.504 0.18 0.522 0.198 ;
      RECT 0.504 0.342 0.522 0.36 ;
      RECT 0.504 0.72 0.522 0.738 ;
      RECT 0.504 0.882 0.522 0.9 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.396 0.378 0.414 0.396 ;
      RECT 0.396 0.684 0.414 0.702 ;
      RECT 0.396 0.918 0.414 0.936 ;
      RECT 0.315 0.18 0.333 0.198 ;
      RECT 0.315 0.342 0.333 0.36 ;
      RECT 0.315 0.72 0.333 0.738 ;
      RECT 0.315 0.882 0.333 0.9 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.18 0.342 0.198 0.36 ;
      RECT 0.18 0.72 0.198 0.738 ;
      RECT 0.18 0.882 0.198 0.9 ;
      RECT 0.142 0.144 0.16 0.162 ;
      RECT 0.142 0.378 0.16 0.396 ;
      RECT 0.142 0.684 0.16 0.702 ;
      RECT 0.142 0.918 0.16 0.936 ;
      RECT 0.024 0.144 0.042 0.162 ;
      RECT 0.024 0.378 0.042 0.396 ;
      RECT 0.024 0.684 0.042 0.702 ;
      RECT 0.024 0.918 0.042 0.936 ;
  END
END DFFHQNV4Xx1_ASAP7_75t_SL

MACRO DFFHQNV4Xx2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNV4Xx2_ASAP7_75t_L 0 0 ;
  SIZE 1.134 BY 1.08 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.126 0.29 0.144 ;
        RECT 0.234 0.225 0.271 0.243 ;
        RECT 0.234 0.027 0.271 0.045 ;
        RECT 0.234 0.027 0.252 0.243 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.396 0.29 0.414 ;
        RECT 0.234 0.495 0.271 0.513 ;
        RECT 0.234 0.297 0.271 0.315 ;
        RECT 0.234 0.297 0.252 0.513 ;
    END
  END D1
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.666 0.29 0.684 ;
        RECT 0.234 0.765 0.271 0.783 ;
        RECT 0.234 0.567 0.271 0.585 ;
        RECT 0.234 0.567 0.252 0.783 ;
    END
  END D2
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.936 0.29 0.954 ;
        RECT 0.234 1.035 0.271 1.053 ;
        RECT 0.234 0.837 0.271 0.855 ;
        RECT 0.234 0.837 0.252 1.053 ;
    END
  END D3
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.216 1.117 0.234 ;
        RECT 1.099 0.036 1.117 0.234 ;
        RECT 1.012 0.036 1.117 0.054 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.486 1.117 0.504 ;
        RECT 1.099 0.306 1.117 0.504 ;
        RECT 1.012 0.306 1.117 0.324 ;
    END
  END QN1
  PIN QN2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.756 1.117 0.774 ;
        RECT 1.099 0.576 1.117 0.774 ;
        RECT 1.012 0.576 1.117 0.594 ;
    END
  END QN2
  PIN QN3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 1.026 1.117 1.044 ;
        RECT 1.099 0.846 1.117 1.044 ;
        RECT 1.012 0.846 1.117 0.864 ;
    END
  END QN3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.134 0.279 ;
        RECT 0 0.801 1.134 0.819 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.134 0.009 ;
        RECT 0 0.531 1.134 0.549 ;
        RECT 0 1.071 1.134 1.089 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 0.04 0.07 0.122 0.088 ;
        RECT 0.04 0.452 0.122 0.47 ;
        RECT 0.04 0.61 0.122 0.628 ;
        RECT 0.04 0.992 0.122 1.01 ;
      LAYER M3 ;
        RECT 0.045 0.05 0.063 1.03 ;
      LAYER M1 ;
        RECT 0.099 0.164 0.117 0.236 ;
        RECT 0.072 0.07 0.117 0.106 ;
        RECT 0.099 0.034 0.117 0.106 ;
        RECT 0.072 0.164 0.117 0.2 ;
        RECT 0.072 0.07 0.09 0.2 ;
        RECT 0.099 0.434 0.117 0.506 ;
        RECT 0.072 0.34 0.117 0.376 ;
        RECT 0.099 0.304 0.117 0.376 ;
        RECT 0.072 0.434 0.117 0.47 ;
        RECT 0.072 0.34 0.09 0.47 ;
        RECT 0.099 0.704 0.117 0.776 ;
        RECT 0.072 0.61 0.117 0.646 ;
        RECT 0.099 0.574 0.117 0.646 ;
        RECT 0.072 0.704 0.117 0.74 ;
        RECT 0.072 0.61 0.09 0.74 ;
        RECT 0.099 0.974 0.117 1.046 ;
        RECT 0.072 0.88 0.117 0.916 ;
        RECT 0.099 0.844 0.117 0.916 ;
        RECT 0.072 0.974 0.117 1.01 ;
        RECT 0.072 0.88 0.09 1.01 ;
      LAYER V2 ;
        RECT 0.045 0.992 0.063 1.01 ;
        RECT 0.045 0.61 0.063 0.628 ;
        RECT 0.045 0.452 0.063 0.47 ;
        RECT 0.045 0.07 0.063 0.088 ;
      LAYER V1 ;
        RECT 0.099 0.992 0.117 1.01 ;
        RECT 0.099 0.61 0.117 0.628 ;
        RECT 0.099 0.452 0.117 0.47 ;
        RECT 0.099 0.07 0.117 0.088 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 0.85 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.774 0.027 0.792 0.119 ;
      RECT 0.774 0.027 0.954 0.045 ;
      RECT 0.774 0.495 0.954 0.513 ;
      RECT 0.936 0.297 0.954 0.513 ;
      RECT 0.774 0.421 0.792 0.513 ;
      RECT 0.85 0.297 0.954 0.315 ;
      RECT 0.85 0.765 0.954 0.783 ;
      RECT 0.936 0.567 0.954 0.783 ;
      RECT 0.774 0.567 0.792 0.659 ;
      RECT 0.774 0.567 0.954 0.585 ;
      RECT 0.774 1.035 0.954 1.053 ;
      RECT 0.936 0.837 0.954 1.053 ;
      RECT 0.774 0.961 0.792 1.053 ;
      RECT 0.85 0.837 0.954 0.855 ;
      RECT 0.688 0.224 0.738 0.242 ;
      RECT 0.72 0.027 0.738 0.242 ;
      RECT 0.72 0.153 0.9 0.171 ;
      RECT 0.882 0.117 0.9 0.171 ;
      RECT 0.828 0.117 0.846 0.171 ;
      RECT 0.634 0.027 0.738 0.045 ;
      RECT 0.634 0.495 0.738 0.513 ;
      RECT 0.72 0.298 0.738 0.513 ;
      RECT 0.882 0.369 0.9 0.423 ;
      RECT 0.828 0.369 0.846 0.423 ;
      RECT 0.72 0.369 0.9 0.387 ;
      RECT 0.688 0.298 0.738 0.316 ;
      RECT 0.688 0.764 0.738 0.782 ;
      RECT 0.72 0.567 0.738 0.782 ;
      RECT 0.72 0.693 0.9 0.711 ;
      RECT 0.882 0.657 0.9 0.711 ;
      RECT 0.828 0.657 0.846 0.711 ;
      RECT 0.634 0.567 0.738 0.585 ;
      RECT 0.634 1.035 0.738 1.053 ;
      RECT 0.72 0.838 0.738 1.053 ;
      RECT 0.882 0.909 0.9 0.963 ;
      RECT 0.828 0.909 0.846 0.963 ;
      RECT 0.72 0.909 0.9 0.927 ;
      RECT 0.688 0.838 0.738 0.856 ;
      RECT 0.576 0.225 0.63 0.243 ;
      RECT 0.612 0.081 0.63 0.243 ;
      RECT 0.496 0.081 0.63 0.099 ;
      RECT 0.585 0.045 0.603 0.099 ;
      RECT 0.585 0.441 0.603 0.495 ;
      RECT 0.496 0.441 0.63 0.459 ;
      RECT 0.612 0.297 0.63 0.459 ;
      RECT 0.576 0.297 0.63 0.315 ;
      RECT 0.576 0.765 0.63 0.783 ;
      RECT 0.612 0.621 0.63 0.783 ;
      RECT 0.496 0.621 0.63 0.639 ;
      RECT 0.585 0.585 0.603 0.639 ;
      RECT 0.585 0.981 0.603 1.035 ;
      RECT 0.496 0.981 0.63 0.999 ;
      RECT 0.612 0.837 0.63 0.999 ;
      RECT 0.576 0.837 0.63 0.855 ;
      RECT 0.364 0.225 0.468 0.243 ;
      RECT 0.45 0.027 0.468 0.243 ;
      RECT 0.45 0.122 0.576 0.14 ;
      RECT 0.418 0.027 0.468 0.045 ;
      RECT 0.418 0.495 0.468 0.513 ;
      RECT 0.45 0.297 0.468 0.513 ;
      RECT 0.45 0.4 0.576 0.418 ;
      RECT 0.364 0.297 0.468 0.315 ;
      RECT 0.364 0.765 0.468 0.783 ;
      RECT 0.45 0.567 0.468 0.783 ;
      RECT 0.45 0.662 0.576 0.68 ;
      RECT 0.418 0.567 0.468 0.585 ;
      RECT 0.418 1.035 0.468 1.053 ;
      RECT 0.45 0.837 0.468 1.053 ;
      RECT 0.45 0.94 0.576 0.958 ;
      RECT 0.364 0.837 0.468 0.855 ;
      RECT 0.315 0.126 0.333 0.203 ;
      RECT 0.315 0.126 0.367 0.144 ;
      RECT 0.315 0.396 0.367 0.414 ;
      RECT 0.315 0.337 0.333 0.414 ;
      RECT 0.315 0.666 0.333 0.743 ;
      RECT 0.315 0.666 0.367 0.684 ;
      RECT 0.315 0.936 0.367 0.954 ;
      RECT 0.315 0.877 0.333 0.954 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.148 0.495 0.198 0.513 ;
      RECT 0.18 0.297 0.198 0.513 ;
      RECT 0.148 0.297 0.198 0.315 ;
      RECT 0.148 0.765 0.198 0.783 ;
      RECT 0.18 0.567 0.198 0.783 ;
      RECT 0.148 0.567 0.198 0.585 ;
      RECT 0.148 1.035 0.198 1.053 ;
      RECT 0.18 0.837 0.198 1.053 ;
      RECT 0.148 0.837 0.198 0.855 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.144 0.047 0.162 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 0.009 0.495 0.068 0.513 ;
      RECT 0.009 0.297 0.027 0.513 ;
      RECT 0.009 0.378 0.047 0.396 ;
      RECT 0.009 0.297 0.068 0.315 ;
      RECT 0.009 0.765 0.068 0.783 ;
      RECT 0.009 0.567 0.027 0.783 ;
      RECT 0.009 0.684 0.047 0.702 ;
      RECT 0.009 0.567 0.068 0.585 ;
      RECT 0.009 1.035 0.068 1.053 ;
      RECT 0.009 0.837 0.027 1.053 ;
      RECT 0.009 0.918 0.047 0.936 ;
      RECT 0.009 0.837 0.068 0.855 ;
      RECT 0.99 0.09 1.008 0.167 ;
      RECT 0.99 0.373 1.008 0.45 ;
      RECT 0.99 0.63 1.008 0.707 ;
      RECT 0.99 0.913 1.008 0.99 ;
      RECT 0.666 0.101 0.684 0.167 ;
      RECT 0.666 0.373 0.684 0.439 ;
      RECT 0.666 0.641 0.684 0.707 ;
      RECT 0.666 0.913 0.684 0.979 ;
      RECT 0.504 0.165 0.522 0.203 ;
      RECT 0.504 0.337 0.522 0.375 ;
      RECT 0.504 0.705 0.522 0.743 ;
      RECT 0.504 0.877 0.522 0.915 ;
      RECT 0.396 0.106 0.414 0.167 ;
      RECT 0.396 0.373 0.414 0.434 ;
      RECT 0.396 0.646 0.414 0.707 ;
      RECT 0.396 0.913 0.414 0.974 ;
      RECT 0.142 0.106 0.16 0.167 ;
      RECT 0.142 0.373 0.16 0.434 ;
      RECT 0.142 0.646 0.16 0.707 ;
      RECT 0.142 0.913 0.16 0.974 ;
    LAYER M2 ;
      RECT 0.877 0.144 1.013 0.162 ;
      RECT 0.877 0.378 1.013 0.396 ;
      RECT 0.877 0.684 1.013 0.702 ;
      RECT 0.877 0.918 1.013 0.936 ;
      RECT 0.019 0.144 0.689 0.162 ;
      RECT 0.019 0.378 0.689 0.396 ;
      RECT 0.019 0.684 0.689 0.702 ;
      RECT 0.019 0.918 0.689 0.936 ;
      RECT 0.175 0.18 0.527 0.198 ;
      RECT 0.175 0.342 0.527 0.36 ;
      RECT 0.175 0.72 0.527 0.738 ;
      RECT 0.175 0.882 0.527 0.9 ;
    LAYER V1 ;
      RECT 0.99 0.144 1.008 0.162 ;
      RECT 0.99 0.378 1.008 0.396 ;
      RECT 0.99 0.684 1.008 0.702 ;
      RECT 0.99 0.918 1.008 0.936 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.882 0.378 0.9 0.396 ;
      RECT 0.882 0.684 0.9 0.702 ;
      RECT 0.882 0.918 0.9 0.936 ;
      RECT 0.666 0.144 0.684 0.162 ;
      RECT 0.666 0.378 0.684 0.396 ;
      RECT 0.666 0.684 0.684 0.702 ;
      RECT 0.666 0.918 0.684 0.936 ;
      RECT 0.504 0.18 0.522 0.198 ;
      RECT 0.504 0.342 0.522 0.36 ;
      RECT 0.504 0.72 0.522 0.738 ;
      RECT 0.504 0.882 0.522 0.9 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.396 0.378 0.414 0.396 ;
      RECT 0.396 0.684 0.414 0.702 ;
      RECT 0.396 0.918 0.414 0.936 ;
      RECT 0.315 0.18 0.333 0.198 ;
      RECT 0.315 0.342 0.333 0.36 ;
      RECT 0.315 0.72 0.333 0.738 ;
      RECT 0.315 0.882 0.333 0.9 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.18 0.342 0.198 0.36 ;
      RECT 0.18 0.72 0.198 0.738 ;
      RECT 0.18 0.882 0.198 0.9 ;
      RECT 0.142 0.144 0.16 0.162 ;
      RECT 0.142 0.378 0.16 0.396 ;
      RECT 0.142 0.684 0.16 0.702 ;
      RECT 0.142 0.918 0.16 0.936 ;
      RECT 0.024 0.144 0.042 0.162 ;
      RECT 0.024 0.378 0.042 0.396 ;
      RECT 0.024 0.684 0.042 0.702 ;
      RECT 0.024 0.918 0.042 0.936 ;
  END
END DFFHQNV4Xx2_ASAP7_75t_L

MACRO DFFHQNV4Xx2_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNV4Xx2_ASAP7_75t_R 0 0 ;
  SIZE 1.134 BY 1.08 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.126 0.29 0.144 ;
        RECT 0.234 0.225 0.271 0.243 ;
        RECT 0.234 0.027 0.271 0.045 ;
        RECT 0.234 0.027 0.252 0.243 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.396 0.29 0.414 ;
        RECT 0.234 0.495 0.271 0.513 ;
        RECT 0.234 0.297 0.271 0.315 ;
        RECT 0.234 0.297 0.252 0.513 ;
    END
  END D1
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.666 0.29 0.684 ;
        RECT 0.234 0.765 0.271 0.783 ;
        RECT 0.234 0.567 0.271 0.585 ;
        RECT 0.234 0.567 0.252 0.783 ;
    END
  END D2
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.936 0.29 0.954 ;
        RECT 0.234 1.035 0.271 1.053 ;
        RECT 0.234 0.837 0.271 0.855 ;
        RECT 0.234 0.837 0.252 1.053 ;
    END
  END D3
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.216 1.117 0.234 ;
        RECT 1.099 0.036 1.117 0.234 ;
        RECT 1.012 0.036 1.117 0.054 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.486 1.117 0.504 ;
        RECT 1.099 0.306 1.117 0.504 ;
        RECT 1.012 0.306 1.117 0.324 ;
    END
  END QN1
  PIN QN2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.756 1.117 0.774 ;
        RECT 1.099 0.576 1.117 0.774 ;
        RECT 1.012 0.576 1.117 0.594 ;
    END
  END QN2
  PIN QN3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 1.026 1.117 1.044 ;
        RECT 1.099 0.846 1.117 1.044 ;
        RECT 1.012 0.846 1.117 0.864 ;
    END
  END QN3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.134 0.279 ;
        RECT 0 0.801 1.134 0.819 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.134 0.009 ;
        RECT 0 0.531 1.134 0.549 ;
        RECT 0 1.071 1.134 1.089 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 0.04 0.07 0.122 0.088 ;
        RECT 0.04 0.452 0.122 0.47 ;
        RECT 0.04 0.61 0.122 0.628 ;
        RECT 0.04 0.992 0.122 1.01 ;
      LAYER M3 ;
        RECT 0.045 0.05 0.063 1.03 ;
      LAYER M1 ;
        RECT 0.099 0.164 0.117 0.236 ;
        RECT 0.072 0.07 0.117 0.106 ;
        RECT 0.099 0.034 0.117 0.106 ;
        RECT 0.072 0.164 0.117 0.2 ;
        RECT 0.072 0.07 0.09 0.2 ;
        RECT 0.099 0.434 0.117 0.506 ;
        RECT 0.072 0.34 0.117 0.376 ;
        RECT 0.099 0.304 0.117 0.376 ;
        RECT 0.072 0.434 0.117 0.47 ;
        RECT 0.072 0.34 0.09 0.47 ;
        RECT 0.099 0.704 0.117 0.776 ;
        RECT 0.072 0.61 0.117 0.646 ;
        RECT 0.099 0.574 0.117 0.646 ;
        RECT 0.072 0.704 0.117 0.74 ;
        RECT 0.072 0.61 0.09 0.74 ;
        RECT 0.099 0.974 0.117 1.046 ;
        RECT 0.072 0.88 0.117 0.916 ;
        RECT 0.099 0.844 0.117 0.916 ;
        RECT 0.072 0.974 0.117 1.01 ;
        RECT 0.072 0.88 0.09 1.01 ;
      LAYER V2 ;
        RECT 0.045 0.992 0.063 1.01 ;
        RECT 0.045 0.61 0.063 0.628 ;
        RECT 0.045 0.452 0.063 0.47 ;
        RECT 0.045 0.07 0.063 0.088 ;
      LAYER V1 ;
        RECT 0.099 0.992 0.117 1.01 ;
        RECT 0.099 0.61 0.117 0.628 ;
        RECT 0.099 0.452 0.117 0.47 ;
        RECT 0.099 0.07 0.117 0.088 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 0.85 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.774 0.027 0.792 0.119 ;
      RECT 0.774 0.027 0.954 0.045 ;
      RECT 0.774 0.495 0.954 0.513 ;
      RECT 0.936 0.297 0.954 0.513 ;
      RECT 0.774 0.421 0.792 0.513 ;
      RECT 0.85 0.297 0.954 0.315 ;
      RECT 0.85 0.765 0.954 0.783 ;
      RECT 0.936 0.567 0.954 0.783 ;
      RECT 0.774 0.567 0.792 0.659 ;
      RECT 0.774 0.567 0.954 0.585 ;
      RECT 0.774 1.035 0.954 1.053 ;
      RECT 0.936 0.837 0.954 1.053 ;
      RECT 0.774 0.961 0.792 1.053 ;
      RECT 0.85 0.837 0.954 0.855 ;
      RECT 0.688 0.224 0.738 0.242 ;
      RECT 0.72 0.027 0.738 0.242 ;
      RECT 0.72 0.153 0.9 0.171 ;
      RECT 0.882 0.117 0.9 0.171 ;
      RECT 0.828 0.117 0.846 0.171 ;
      RECT 0.634 0.027 0.738 0.045 ;
      RECT 0.634 0.495 0.738 0.513 ;
      RECT 0.72 0.298 0.738 0.513 ;
      RECT 0.882 0.369 0.9 0.423 ;
      RECT 0.828 0.369 0.846 0.423 ;
      RECT 0.72 0.369 0.9 0.387 ;
      RECT 0.688 0.298 0.738 0.316 ;
      RECT 0.688 0.764 0.738 0.782 ;
      RECT 0.72 0.567 0.738 0.782 ;
      RECT 0.72 0.693 0.9 0.711 ;
      RECT 0.882 0.657 0.9 0.711 ;
      RECT 0.828 0.657 0.846 0.711 ;
      RECT 0.634 0.567 0.738 0.585 ;
      RECT 0.634 1.035 0.738 1.053 ;
      RECT 0.72 0.838 0.738 1.053 ;
      RECT 0.882 0.909 0.9 0.963 ;
      RECT 0.828 0.909 0.846 0.963 ;
      RECT 0.72 0.909 0.9 0.927 ;
      RECT 0.688 0.838 0.738 0.856 ;
      RECT 0.576 0.225 0.63 0.243 ;
      RECT 0.612 0.081 0.63 0.243 ;
      RECT 0.496 0.081 0.63 0.099 ;
      RECT 0.585 0.045 0.603 0.099 ;
      RECT 0.585 0.441 0.603 0.495 ;
      RECT 0.496 0.441 0.63 0.459 ;
      RECT 0.612 0.297 0.63 0.459 ;
      RECT 0.576 0.297 0.63 0.315 ;
      RECT 0.576 0.765 0.63 0.783 ;
      RECT 0.612 0.621 0.63 0.783 ;
      RECT 0.496 0.621 0.63 0.639 ;
      RECT 0.585 0.585 0.603 0.639 ;
      RECT 0.585 0.981 0.603 1.035 ;
      RECT 0.496 0.981 0.63 0.999 ;
      RECT 0.612 0.837 0.63 0.999 ;
      RECT 0.576 0.837 0.63 0.855 ;
      RECT 0.364 0.225 0.468 0.243 ;
      RECT 0.45 0.027 0.468 0.243 ;
      RECT 0.45 0.122 0.576 0.14 ;
      RECT 0.418 0.027 0.468 0.045 ;
      RECT 0.418 0.495 0.468 0.513 ;
      RECT 0.45 0.297 0.468 0.513 ;
      RECT 0.45 0.4 0.576 0.418 ;
      RECT 0.364 0.297 0.468 0.315 ;
      RECT 0.364 0.765 0.468 0.783 ;
      RECT 0.45 0.567 0.468 0.783 ;
      RECT 0.45 0.662 0.576 0.68 ;
      RECT 0.418 0.567 0.468 0.585 ;
      RECT 0.418 1.035 0.468 1.053 ;
      RECT 0.45 0.837 0.468 1.053 ;
      RECT 0.45 0.94 0.576 0.958 ;
      RECT 0.364 0.837 0.468 0.855 ;
      RECT 0.315 0.126 0.333 0.203 ;
      RECT 0.315 0.126 0.367 0.144 ;
      RECT 0.315 0.396 0.367 0.414 ;
      RECT 0.315 0.337 0.333 0.414 ;
      RECT 0.315 0.666 0.333 0.743 ;
      RECT 0.315 0.666 0.367 0.684 ;
      RECT 0.315 0.936 0.367 0.954 ;
      RECT 0.315 0.877 0.333 0.954 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.148 0.495 0.198 0.513 ;
      RECT 0.18 0.297 0.198 0.513 ;
      RECT 0.148 0.297 0.198 0.315 ;
      RECT 0.148 0.765 0.198 0.783 ;
      RECT 0.18 0.567 0.198 0.783 ;
      RECT 0.148 0.567 0.198 0.585 ;
      RECT 0.148 1.035 0.198 1.053 ;
      RECT 0.18 0.837 0.198 1.053 ;
      RECT 0.148 0.837 0.198 0.855 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.144 0.047 0.162 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 0.009 0.495 0.068 0.513 ;
      RECT 0.009 0.297 0.027 0.513 ;
      RECT 0.009 0.378 0.047 0.396 ;
      RECT 0.009 0.297 0.068 0.315 ;
      RECT 0.009 0.765 0.068 0.783 ;
      RECT 0.009 0.567 0.027 0.783 ;
      RECT 0.009 0.684 0.047 0.702 ;
      RECT 0.009 0.567 0.068 0.585 ;
      RECT 0.009 1.035 0.068 1.053 ;
      RECT 0.009 0.837 0.027 1.053 ;
      RECT 0.009 0.918 0.047 0.936 ;
      RECT 0.009 0.837 0.068 0.855 ;
      RECT 0.99 0.09 1.008 0.167 ;
      RECT 0.99 0.373 1.008 0.45 ;
      RECT 0.99 0.63 1.008 0.707 ;
      RECT 0.99 0.913 1.008 0.99 ;
      RECT 0.666 0.101 0.684 0.167 ;
      RECT 0.666 0.373 0.684 0.439 ;
      RECT 0.666 0.641 0.684 0.707 ;
      RECT 0.666 0.913 0.684 0.979 ;
      RECT 0.504 0.165 0.522 0.203 ;
      RECT 0.504 0.337 0.522 0.375 ;
      RECT 0.504 0.705 0.522 0.743 ;
      RECT 0.504 0.877 0.522 0.915 ;
      RECT 0.396 0.106 0.414 0.167 ;
      RECT 0.396 0.373 0.414 0.434 ;
      RECT 0.396 0.646 0.414 0.707 ;
      RECT 0.396 0.913 0.414 0.974 ;
      RECT 0.142 0.106 0.16 0.167 ;
      RECT 0.142 0.373 0.16 0.434 ;
      RECT 0.142 0.646 0.16 0.707 ;
      RECT 0.142 0.913 0.16 0.974 ;
    LAYER M2 ;
      RECT 0.877 0.144 1.013 0.162 ;
      RECT 0.877 0.378 1.013 0.396 ;
      RECT 0.877 0.684 1.013 0.702 ;
      RECT 0.877 0.918 1.013 0.936 ;
      RECT 0.019 0.144 0.689 0.162 ;
      RECT 0.019 0.378 0.689 0.396 ;
      RECT 0.019 0.684 0.689 0.702 ;
      RECT 0.019 0.918 0.689 0.936 ;
      RECT 0.175 0.18 0.527 0.198 ;
      RECT 0.175 0.342 0.527 0.36 ;
      RECT 0.175 0.72 0.527 0.738 ;
      RECT 0.175 0.882 0.527 0.9 ;
    LAYER V1 ;
      RECT 0.99 0.144 1.008 0.162 ;
      RECT 0.99 0.378 1.008 0.396 ;
      RECT 0.99 0.684 1.008 0.702 ;
      RECT 0.99 0.918 1.008 0.936 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.882 0.378 0.9 0.396 ;
      RECT 0.882 0.684 0.9 0.702 ;
      RECT 0.882 0.918 0.9 0.936 ;
      RECT 0.666 0.144 0.684 0.162 ;
      RECT 0.666 0.378 0.684 0.396 ;
      RECT 0.666 0.684 0.684 0.702 ;
      RECT 0.666 0.918 0.684 0.936 ;
      RECT 0.504 0.18 0.522 0.198 ;
      RECT 0.504 0.342 0.522 0.36 ;
      RECT 0.504 0.72 0.522 0.738 ;
      RECT 0.504 0.882 0.522 0.9 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.396 0.378 0.414 0.396 ;
      RECT 0.396 0.684 0.414 0.702 ;
      RECT 0.396 0.918 0.414 0.936 ;
      RECT 0.315 0.18 0.333 0.198 ;
      RECT 0.315 0.342 0.333 0.36 ;
      RECT 0.315 0.72 0.333 0.738 ;
      RECT 0.315 0.882 0.333 0.9 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.18 0.342 0.198 0.36 ;
      RECT 0.18 0.72 0.198 0.738 ;
      RECT 0.18 0.882 0.198 0.9 ;
      RECT 0.142 0.144 0.16 0.162 ;
      RECT 0.142 0.378 0.16 0.396 ;
      RECT 0.142 0.684 0.16 0.702 ;
      RECT 0.142 0.918 0.16 0.936 ;
      RECT 0.024 0.144 0.042 0.162 ;
      RECT 0.024 0.378 0.042 0.396 ;
      RECT 0.024 0.684 0.042 0.702 ;
      RECT 0.024 0.918 0.042 0.936 ;
  END
END DFFHQNV4Xx2_ASAP7_75t_R

MACRO DFFHQNV4Xx2_ASAP7_75t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNV4Xx2_ASAP7_75t_SL 0 0 ;
  SIZE 1.134 BY 1.08 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.126 0.29 0.144 ;
        RECT 0.234 0.225 0.271 0.243 ;
        RECT 0.234 0.027 0.271 0.045 ;
        RECT 0.234 0.027 0.252 0.243 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.396 0.29 0.414 ;
        RECT 0.234 0.495 0.271 0.513 ;
        RECT 0.234 0.297 0.271 0.315 ;
        RECT 0.234 0.297 0.252 0.513 ;
    END
  END D1
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.666 0.29 0.684 ;
        RECT 0.234 0.765 0.271 0.783 ;
        RECT 0.234 0.567 0.271 0.585 ;
        RECT 0.234 0.567 0.252 0.783 ;
    END
  END D2
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.936 0.29 0.954 ;
        RECT 0.234 1.035 0.271 1.053 ;
        RECT 0.234 0.837 0.271 0.855 ;
        RECT 0.234 0.837 0.252 1.053 ;
    END
  END D3
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.216 1.117 0.234 ;
        RECT 1.099 0.036 1.117 0.234 ;
        RECT 1.012 0.036 1.117 0.054 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.486 1.117 0.504 ;
        RECT 1.099 0.306 1.117 0.504 ;
        RECT 1.012 0.306 1.117 0.324 ;
    END
  END QN1
  PIN QN2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.756 1.117 0.774 ;
        RECT 1.099 0.576 1.117 0.774 ;
        RECT 1.012 0.576 1.117 0.594 ;
    END
  END QN2
  PIN QN3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 1.026 1.117 1.044 ;
        RECT 1.099 0.846 1.117 1.044 ;
        RECT 1.012 0.846 1.117 0.864 ;
    END
  END QN3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.134 0.279 ;
        RECT 0 0.801 1.134 0.819 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.134 0.009 ;
        RECT 0 0.531 1.134 0.549 ;
        RECT 0 1.071 1.134 1.089 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 0.04 0.07 0.122 0.088 ;
        RECT 0.04 0.452 0.122 0.47 ;
        RECT 0.04 0.61 0.122 0.628 ;
        RECT 0.04 0.992 0.122 1.01 ;
      LAYER M3 ;
        RECT 0.045 0.05 0.063 1.03 ;
      LAYER M1 ;
        RECT 0.099 0.164 0.117 0.236 ;
        RECT 0.072 0.07 0.117 0.106 ;
        RECT 0.099 0.034 0.117 0.106 ;
        RECT 0.072 0.164 0.117 0.2 ;
        RECT 0.072 0.07 0.09 0.2 ;
        RECT 0.099 0.434 0.117 0.506 ;
        RECT 0.072 0.34 0.117 0.376 ;
        RECT 0.099 0.304 0.117 0.376 ;
        RECT 0.072 0.434 0.117 0.47 ;
        RECT 0.072 0.34 0.09 0.47 ;
        RECT 0.099 0.704 0.117 0.776 ;
        RECT 0.072 0.61 0.117 0.646 ;
        RECT 0.099 0.574 0.117 0.646 ;
        RECT 0.072 0.704 0.117 0.74 ;
        RECT 0.072 0.61 0.09 0.74 ;
        RECT 0.099 0.974 0.117 1.046 ;
        RECT 0.072 0.88 0.117 0.916 ;
        RECT 0.099 0.844 0.117 0.916 ;
        RECT 0.072 0.974 0.117 1.01 ;
        RECT 0.072 0.88 0.09 1.01 ;
      LAYER V2 ;
        RECT 0.045 0.992 0.063 1.01 ;
        RECT 0.045 0.61 0.063 0.628 ;
        RECT 0.045 0.452 0.063 0.47 ;
        RECT 0.045 0.07 0.063 0.088 ;
      LAYER V1 ;
        RECT 0.099 0.992 0.117 1.01 ;
        RECT 0.099 0.61 0.117 0.628 ;
        RECT 0.099 0.452 0.117 0.47 ;
        RECT 0.099 0.07 0.117 0.088 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 0.85 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.774 0.027 0.792 0.119 ;
      RECT 0.774 0.027 0.954 0.045 ;
      RECT 0.774 0.495 0.954 0.513 ;
      RECT 0.936 0.297 0.954 0.513 ;
      RECT 0.774 0.421 0.792 0.513 ;
      RECT 0.85 0.297 0.954 0.315 ;
      RECT 0.85 0.765 0.954 0.783 ;
      RECT 0.936 0.567 0.954 0.783 ;
      RECT 0.774 0.567 0.792 0.659 ;
      RECT 0.774 0.567 0.954 0.585 ;
      RECT 0.774 1.035 0.954 1.053 ;
      RECT 0.936 0.837 0.954 1.053 ;
      RECT 0.774 0.961 0.792 1.053 ;
      RECT 0.85 0.837 0.954 0.855 ;
      RECT 0.688 0.224 0.738 0.242 ;
      RECT 0.72 0.027 0.738 0.242 ;
      RECT 0.72 0.153 0.9 0.171 ;
      RECT 0.882 0.117 0.9 0.171 ;
      RECT 0.828 0.117 0.846 0.171 ;
      RECT 0.634 0.027 0.738 0.045 ;
      RECT 0.634 0.495 0.738 0.513 ;
      RECT 0.72 0.298 0.738 0.513 ;
      RECT 0.882 0.369 0.9 0.423 ;
      RECT 0.828 0.369 0.846 0.423 ;
      RECT 0.72 0.369 0.9 0.387 ;
      RECT 0.688 0.298 0.738 0.316 ;
      RECT 0.688 0.764 0.738 0.782 ;
      RECT 0.72 0.567 0.738 0.782 ;
      RECT 0.72 0.693 0.9 0.711 ;
      RECT 0.882 0.657 0.9 0.711 ;
      RECT 0.828 0.657 0.846 0.711 ;
      RECT 0.634 0.567 0.738 0.585 ;
      RECT 0.634 1.035 0.738 1.053 ;
      RECT 0.72 0.838 0.738 1.053 ;
      RECT 0.882 0.909 0.9 0.963 ;
      RECT 0.828 0.909 0.846 0.963 ;
      RECT 0.72 0.909 0.9 0.927 ;
      RECT 0.688 0.838 0.738 0.856 ;
      RECT 0.576 0.225 0.63 0.243 ;
      RECT 0.612 0.081 0.63 0.243 ;
      RECT 0.496 0.081 0.63 0.099 ;
      RECT 0.585 0.045 0.603 0.099 ;
      RECT 0.585 0.441 0.603 0.495 ;
      RECT 0.496 0.441 0.63 0.459 ;
      RECT 0.612 0.297 0.63 0.459 ;
      RECT 0.576 0.297 0.63 0.315 ;
      RECT 0.576 0.765 0.63 0.783 ;
      RECT 0.612 0.621 0.63 0.783 ;
      RECT 0.496 0.621 0.63 0.639 ;
      RECT 0.585 0.585 0.603 0.639 ;
      RECT 0.585 0.981 0.603 1.035 ;
      RECT 0.496 0.981 0.63 0.999 ;
      RECT 0.612 0.837 0.63 0.999 ;
      RECT 0.576 0.837 0.63 0.855 ;
      RECT 0.364 0.225 0.468 0.243 ;
      RECT 0.45 0.027 0.468 0.243 ;
      RECT 0.45 0.122 0.576 0.14 ;
      RECT 0.418 0.027 0.468 0.045 ;
      RECT 0.418 0.495 0.468 0.513 ;
      RECT 0.45 0.297 0.468 0.513 ;
      RECT 0.45 0.4 0.576 0.418 ;
      RECT 0.364 0.297 0.468 0.315 ;
      RECT 0.364 0.765 0.468 0.783 ;
      RECT 0.45 0.567 0.468 0.783 ;
      RECT 0.45 0.662 0.576 0.68 ;
      RECT 0.418 0.567 0.468 0.585 ;
      RECT 0.418 1.035 0.468 1.053 ;
      RECT 0.45 0.837 0.468 1.053 ;
      RECT 0.45 0.94 0.576 0.958 ;
      RECT 0.364 0.837 0.468 0.855 ;
      RECT 0.315 0.126 0.333 0.203 ;
      RECT 0.315 0.126 0.367 0.144 ;
      RECT 0.315 0.396 0.367 0.414 ;
      RECT 0.315 0.337 0.333 0.414 ;
      RECT 0.315 0.666 0.333 0.743 ;
      RECT 0.315 0.666 0.367 0.684 ;
      RECT 0.315 0.936 0.367 0.954 ;
      RECT 0.315 0.877 0.333 0.954 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.148 0.495 0.198 0.513 ;
      RECT 0.18 0.297 0.198 0.513 ;
      RECT 0.148 0.297 0.198 0.315 ;
      RECT 0.148 0.765 0.198 0.783 ;
      RECT 0.18 0.567 0.198 0.783 ;
      RECT 0.148 0.567 0.198 0.585 ;
      RECT 0.148 1.035 0.198 1.053 ;
      RECT 0.18 0.837 0.198 1.053 ;
      RECT 0.148 0.837 0.198 0.855 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.144 0.047 0.162 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 0.009 0.495 0.068 0.513 ;
      RECT 0.009 0.297 0.027 0.513 ;
      RECT 0.009 0.378 0.047 0.396 ;
      RECT 0.009 0.297 0.068 0.315 ;
      RECT 0.009 0.765 0.068 0.783 ;
      RECT 0.009 0.567 0.027 0.783 ;
      RECT 0.009 0.684 0.047 0.702 ;
      RECT 0.009 0.567 0.068 0.585 ;
      RECT 0.009 1.035 0.068 1.053 ;
      RECT 0.009 0.837 0.027 1.053 ;
      RECT 0.009 0.918 0.047 0.936 ;
      RECT 0.009 0.837 0.068 0.855 ;
      RECT 0.99 0.09 1.008 0.167 ;
      RECT 0.99 0.373 1.008 0.45 ;
      RECT 0.99 0.63 1.008 0.707 ;
      RECT 0.99 0.913 1.008 0.99 ;
      RECT 0.666 0.101 0.684 0.167 ;
      RECT 0.666 0.373 0.684 0.439 ;
      RECT 0.666 0.641 0.684 0.707 ;
      RECT 0.666 0.913 0.684 0.979 ;
      RECT 0.504 0.165 0.522 0.203 ;
      RECT 0.504 0.337 0.522 0.375 ;
      RECT 0.504 0.705 0.522 0.743 ;
      RECT 0.504 0.877 0.522 0.915 ;
      RECT 0.396 0.106 0.414 0.167 ;
      RECT 0.396 0.373 0.414 0.434 ;
      RECT 0.396 0.646 0.414 0.707 ;
      RECT 0.396 0.913 0.414 0.974 ;
      RECT 0.142 0.106 0.16 0.167 ;
      RECT 0.142 0.373 0.16 0.434 ;
      RECT 0.142 0.646 0.16 0.707 ;
      RECT 0.142 0.913 0.16 0.974 ;
    LAYER M2 ;
      RECT 0.877 0.144 1.013 0.162 ;
      RECT 0.877 0.378 1.013 0.396 ;
      RECT 0.877 0.684 1.013 0.702 ;
      RECT 0.877 0.918 1.013 0.936 ;
      RECT 0.019 0.144 0.689 0.162 ;
      RECT 0.019 0.378 0.689 0.396 ;
      RECT 0.019 0.684 0.689 0.702 ;
      RECT 0.019 0.918 0.689 0.936 ;
      RECT 0.175 0.18 0.527 0.198 ;
      RECT 0.175 0.342 0.527 0.36 ;
      RECT 0.175 0.72 0.527 0.738 ;
      RECT 0.175 0.882 0.527 0.9 ;
    LAYER V1 ;
      RECT 0.99 0.144 1.008 0.162 ;
      RECT 0.99 0.378 1.008 0.396 ;
      RECT 0.99 0.684 1.008 0.702 ;
      RECT 0.99 0.918 1.008 0.936 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.882 0.378 0.9 0.396 ;
      RECT 0.882 0.684 0.9 0.702 ;
      RECT 0.882 0.918 0.9 0.936 ;
      RECT 0.666 0.144 0.684 0.162 ;
      RECT 0.666 0.378 0.684 0.396 ;
      RECT 0.666 0.684 0.684 0.702 ;
      RECT 0.666 0.918 0.684 0.936 ;
      RECT 0.504 0.18 0.522 0.198 ;
      RECT 0.504 0.342 0.522 0.36 ;
      RECT 0.504 0.72 0.522 0.738 ;
      RECT 0.504 0.882 0.522 0.9 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.396 0.378 0.414 0.396 ;
      RECT 0.396 0.684 0.414 0.702 ;
      RECT 0.396 0.918 0.414 0.936 ;
      RECT 0.315 0.18 0.333 0.198 ;
      RECT 0.315 0.342 0.333 0.36 ;
      RECT 0.315 0.72 0.333 0.738 ;
      RECT 0.315 0.882 0.333 0.9 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.18 0.342 0.198 0.36 ;
      RECT 0.18 0.72 0.198 0.738 ;
      RECT 0.18 0.882 0.198 0.9 ;
      RECT 0.142 0.144 0.16 0.162 ;
      RECT 0.142 0.378 0.16 0.396 ;
      RECT 0.142 0.684 0.16 0.702 ;
      RECT 0.142 0.918 0.16 0.936 ;
      RECT 0.024 0.144 0.042 0.162 ;
      RECT 0.024 0.378 0.042 0.396 ;
      RECT 0.024 0.684 0.042 0.702 ;
      RECT 0.024 0.918 0.042 0.936 ;
  END
END DFFHQNV4Xx2_ASAP7_75t_SL

MACRO DFFHQNV4Xx3_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNV4Xx3_ASAP7_75t_L 0 0 ;
  SIZE 1.188 BY 1.08 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.126 0.29 0.144 ;
        RECT 0.234 0.225 0.271 0.243 ;
        RECT 0.234 0.027 0.271 0.045 ;
        RECT 0.234 0.027 0.252 0.243 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.396 0.29 0.414 ;
        RECT 0.234 0.495 0.271 0.513 ;
        RECT 0.234 0.297 0.271 0.315 ;
        RECT 0.234 0.297 0.252 0.513 ;
    END
  END D1
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.666 0.29 0.684 ;
        RECT 0.234 0.765 0.271 0.783 ;
        RECT 0.234 0.567 0.271 0.585 ;
        RECT 0.234 0.567 0.252 0.783 ;
    END
  END D2
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.936 0.29 0.954 ;
        RECT 0.234 1.035 0.271 1.053 ;
        RECT 0.234 0.837 0.271 0.855 ;
        RECT 0.234 0.837 0.252 1.053 ;
    END
  END D3
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.225 1.171 0.243 ;
        RECT 1.153 0.027 1.171 0.243 ;
        RECT 1.012 0.027 1.171 0.045 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.495 1.171 0.513 ;
        RECT 1.153 0.297 1.171 0.513 ;
        RECT 1.012 0.297 1.171 0.315 ;
    END
  END QN1
  PIN QN2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.765 1.171 0.783 ;
        RECT 1.153 0.567 1.171 0.783 ;
        RECT 1.012 0.567 1.171 0.585 ;
    END
  END QN2
  PIN QN3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 1.035 1.171 1.053 ;
        RECT 1.153 0.837 1.171 1.053 ;
        RECT 1.012 0.837 1.171 0.855 ;
    END
  END QN3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.188 0.279 ;
        RECT 0 0.801 1.188 0.819 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.188 0.009 ;
        RECT 0 0.531 1.188 0.549 ;
        RECT 0 1.071 1.188 1.089 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 0.04 0.07 0.122 0.088 ;
        RECT 0.04 0.452 0.122 0.47 ;
        RECT 0.04 0.61 0.122 0.628 ;
        RECT 0.04 0.992 0.122 1.01 ;
      LAYER M3 ;
        RECT 0.045 0.05 0.063 1.03 ;
      LAYER M1 ;
        RECT 0.099 0.164 0.117 0.236 ;
        RECT 0.072 0.07 0.117 0.106 ;
        RECT 0.099 0.034 0.117 0.106 ;
        RECT 0.072 0.164 0.117 0.2 ;
        RECT 0.072 0.07 0.09 0.2 ;
        RECT 0.099 0.434 0.117 0.506 ;
        RECT 0.072 0.34 0.117 0.376 ;
        RECT 0.099 0.304 0.117 0.376 ;
        RECT 0.072 0.434 0.117 0.47 ;
        RECT 0.072 0.34 0.09 0.47 ;
        RECT 0.099 0.704 0.117 0.776 ;
        RECT 0.072 0.61 0.117 0.646 ;
        RECT 0.099 0.574 0.117 0.646 ;
        RECT 0.072 0.704 0.117 0.74 ;
        RECT 0.072 0.61 0.09 0.74 ;
        RECT 0.099 0.974 0.117 1.046 ;
        RECT 0.072 0.88 0.117 0.916 ;
        RECT 0.099 0.844 0.117 0.916 ;
        RECT 0.072 0.974 0.117 1.01 ;
        RECT 0.072 0.88 0.09 1.01 ;
      LAYER V2 ;
        RECT 0.045 0.992 0.063 1.01 ;
        RECT 0.045 0.61 0.063 0.628 ;
        RECT 0.045 0.452 0.063 0.47 ;
        RECT 0.045 0.07 0.063 0.088 ;
      LAYER V1 ;
        RECT 0.099 0.992 0.117 1.01 ;
        RECT 0.099 0.61 0.117 0.628 ;
        RECT 0.099 0.452 0.117 0.47 ;
        RECT 0.099 0.07 0.117 0.088 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 0.85 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.774 0.027 0.792 0.119 ;
      RECT 0.774 0.027 0.954 0.045 ;
      RECT 0.774 0.495 0.954 0.513 ;
      RECT 0.936 0.297 0.954 0.513 ;
      RECT 0.774 0.421 0.792 0.513 ;
      RECT 0.85 0.297 0.954 0.315 ;
      RECT 0.85 0.765 0.954 0.783 ;
      RECT 0.936 0.567 0.954 0.783 ;
      RECT 0.774 0.567 0.792 0.659 ;
      RECT 0.774 0.567 0.954 0.585 ;
      RECT 0.774 1.035 0.954 1.053 ;
      RECT 0.936 0.837 0.954 1.053 ;
      RECT 0.774 0.961 0.792 1.053 ;
      RECT 0.85 0.837 0.954 0.855 ;
      RECT 0.688 0.224 0.738 0.242 ;
      RECT 0.72 0.027 0.738 0.242 ;
      RECT 0.72 0.153 0.9 0.171 ;
      RECT 0.882 0.117 0.9 0.171 ;
      RECT 0.828 0.117 0.846 0.171 ;
      RECT 0.634 0.027 0.738 0.045 ;
      RECT 0.634 0.495 0.738 0.513 ;
      RECT 0.72 0.298 0.738 0.513 ;
      RECT 0.882 0.369 0.9 0.423 ;
      RECT 0.828 0.369 0.846 0.423 ;
      RECT 0.72 0.369 0.9 0.387 ;
      RECT 0.688 0.298 0.738 0.316 ;
      RECT 0.688 0.764 0.738 0.782 ;
      RECT 0.72 0.567 0.738 0.782 ;
      RECT 0.72 0.693 0.9 0.711 ;
      RECT 0.882 0.657 0.9 0.711 ;
      RECT 0.828 0.657 0.846 0.711 ;
      RECT 0.634 0.567 0.738 0.585 ;
      RECT 0.634 1.035 0.738 1.053 ;
      RECT 0.72 0.838 0.738 1.053 ;
      RECT 0.882 0.909 0.9 0.963 ;
      RECT 0.828 0.909 0.846 0.963 ;
      RECT 0.72 0.909 0.9 0.927 ;
      RECT 0.688 0.838 0.738 0.856 ;
      RECT 0.576 0.225 0.63 0.243 ;
      RECT 0.612 0.081 0.63 0.243 ;
      RECT 0.496 0.081 0.63 0.099 ;
      RECT 0.585 0.045 0.603 0.099 ;
      RECT 0.585 0.441 0.603 0.495 ;
      RECT 0.496 0.441 0.63 0.459 ;
      RECT 0.612 0.297 0.63 0.459 ;
      RECT 0.576 0.297 0.63 0.315 ;
      RECT 0.576 0.765 0.63 0.783 ;
      RECT 0.612 0.621 0.63 0.783 ;
      RECT 0.496 0.621 0.63 0.639 ;
      RECT 0.585 0.585 0.603 0.639 ;
      RECT 0.585 0.981 0.603 1.035 ;
      RECT 0.496 0.981 0.63 0.999 ;
      RECT 0.612 0.837 0.63 0.999 ;
      RECT 0.576 0.837 0.63 0.855 ;
      RECT 0.364 0.225 0.468 0.243 ;
      RECT 0.45 0.027 0.468 0.243 ;
      RECT 0.45 0.122 0.576 0.14 ;
      RECT 0.418 0.027 0.468 0.045 ;
      RECT 0.418 0.495 0.468 0.513 ;
      RECT 0.45 0.297 0.468 0.513 ;
      RECT 0.45 0.4 0.576 0.418 ;
      RECT 0.364 0.297 0.468 0.315 ;
      RECT 0.364 0.765 0.468 0.783 ;
      RECT 0.45 0.567 0.468 0.783 ;
      RECT 0.45 0.662 0.576 0.68 ;
      RECT 0.418 0.567 0.468 0.585 ;
      RECT 0.418 1.035 0.468 1.053 ;
      RECT 0.45 0.837 0.468 1.053 ;
      RECT 0.45 0.94 0.576 0.958 ;
      RECT 0.364 0.837 0.468 0.855 ;
      RECT 0.315 0.126 0.333 0.203 ;
      RECT 0.315 0.126 0.367 0.144 ;
      RECT 0.315 0.396 0.367 0.414 ;
      RECT 0.315 0.337 0.333 0.414 ;
      RECT 0.315 0.666 0.333 0.743 ;
      RECT 0.315 0.666 0.367 0.684 ;
      RECT 0.315 0.936 0.367 0.954 ;
      RECT 0.315 0.877 0.333 0.954 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.148 0.495 0.198 0.513 ;
      RECT 0.18 0.297 0.198 0.513 ;
      RECT 0.148 0.297 0.198 0.315 ;
      RECT 0.148 0.765 0.198 0.783 ;
      RECT 0.18 0.567 0.198 0.783 ;
      RECT 0.148 0.567 0.198 0.585 ;
      RECT 0.148 1.035 0.198 1.053 ;
      RECT 0.18 0.837 0.198 1.053 ;
      RECT 0.148 0.837 0.198 0.855 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.144 0.047 0.162 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 0.009 0.495 0.068 0.513 ;
      RECT 0.009 0.297 0.027 0.513 ;
      RECT 0.009 0.378 0.047 0.396 ;
      RECT 0.009 0.297 0.068 0.315 ;
      RECT 0.009 0.765 0.068 0.783 ;
      RECT 0.009 0.567 0.027 0.783 ;
      RECT 0.009 0.684 0.047 0.702 ;
      RECT 0.009 0.567 0.068 0.585 ;
      RECT 0.009 1.035 0.068 1.053 ;
      RECT 0.009 0.837 0.027 1.053 ;
      RECT 0.009 0.918 0.047 0.936 ;
      RECT 0.009 0.837 0.068 0.855 ;
      RECT 0.99 0.122 1.008 0.167 ;
      RECT 0.99 0.373 1.008 0.418 ;
      RECT 0.99 0.662 1.008 0.707 ;
      RECT 0.99 0.913 1.008 0.958 ;
      RECT 0.666 0.101 0.684 0.167 ;
      RECT 0.666 0.373 0.684 0.439 ;
      RECT 0.666 0.641 0.684 0.707 ;
      RECT 0.666 0.913 0.684 0.979 ;
      RECT 0.504 0.165 0.522 0.203 ;
      RECT 0.504 0.337 0.522 0.375 ;
      RECT 0.504 0.705 0.522 0.743 ;
      RECT 0.504 0.877 0.522 0.915 ;
      RECT 0.396 0.106 0.414 0.167 ;
      RECT 0.396 0.373 0.414 0.434 ;
      RECT 0.396 0.646 0.414 0.707 ;
      RECT 0.396 0.913 0.414 0.974 ;
      RECT 0.142 0.106 0.16 0.167 ;
      RECT 0.142 0.373 0.16 0.434 ;
      RECT 0.142 0.646 0.16 0.707 ;
      RECT 0.142 0.913 0.16 0.974 ;
    LAYER M2 ;
      RECT 0.877 0.144 1.013 0.162 ;
      RECT 0.877 0.378 1.013 0.396 ;
      RECT 0.877 0.684 1.013 0.702 ;
      RECT 0.877 0.918 1.013 0.936 ;
      RECT 0.019 0.144 0.689 0.162 ;
      RECT 0.019 0.378 0.689 0.396 ;
      RECT 0.019 0.684 0.689 0.702 ;
      RECT 0.019 0.918 0.689 0.936 ;
      RECT 0.175 0.18 0.527 0.198 ;
      RECT 0.175 0.342 0.527 0.36 ;
      RECT 0.175 0.72 0.527 0.738 ;
      RECT 0.175 0.882 0.527 0.9 ;
    LAYER V1 ;
      RECT 0.99 0.144 1.008 0.162 ;
      RECT 0.99 0.378 1.008 0.396 ;
      RECT 0.99 0.684 1.008 0.702 ;
      RECT 0.99 0.918 1.008 0.936 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.882 0.378 0.9 0.396 ;
      RECT 0.882 0.684 0.9 0.702 ;
      RECT 0.882 0.918 0.9 0.936 ;
      RECT 0.666 0.144 0.684 0.162 ;
      RECT 0.666 0.378 0.684 0.396 ;
      RECT 0.666 0.684 0.684 0.702 ;
      RECT 0.666 0.918 0.684 0.936 ;
      RECT 0.504 0.18 0.522 0.198 ;
      RECT 0.504 0.342 0.522 0.36 ;
      RECT 0.504 0.72 0.522 0.738 ;
      RECT 0.504 0.882 0.522 0.9 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.396 0.378 0.414 0.396 ;
      RECT 0.396 0.684 0.414 0.702 ;
      RECT 0.396 0.918 0.414 0.936 ;
      RECT 0.315 0.18 0.333 0.198 ;
      RECT 0.315 0.342 0.333 0.36 ;
      RECT 0.315 0.72 0.333 0.738 ;
      RECT 0.315 0.882 0.333 0.9 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.18 0.342 0.198 0.36 ;
      RECT 0.18 0.72 0.198 0.738 ;
      RECT 0.18 0.882 0.198 0.9 ;
      RECT 0.142 0.144 0.16 0.162 ;
      RECT 0.142 0.378 0.16 0.396 ;
      RECT 0.142 0.684 0.16 0.702 ;
      RECT 0.142 0.918 0.16 0.936 ;
      RECT 0.024 0.144 0.042 0.162 ;
      RECT 0.024 0.378 0.042 0.396 ;
      RECT 0.024 0.684 0.042 0.702 ;
      RECT 0.024 0.918 0.042 0.936 ;
  END
END DFFHQNV4Xx3_ASAP7_75t_L

MACRO DFFHQNV4Xx3_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNV4Xx3_ASAP7_75t_R 0 0 ;
  SIZE 1.188 BY 1.08 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.126 0.29 0.144 ;
        RECT 0.234 0.225 0.271 0.243 ;
        RECT 0.234 0.027 0.271 0.045 ;
        RECT 0.234 0.027 0.252 0.243 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.396 0.29 0.414 ;
        RECT 0.234 0.495 0.271 0.513 ;
        RECT 0.234 0.297 0.271 0.315 ;
        RECT 0.234 0.297 0.252 0.513 ;
    END
  END D1
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.666 0.29 0.684 ;
        RECT 0.234 0.765 0.271 0.783 ;
        RECT 0.234 0.567 0.271 0.585 ;
        RECT 0.234 0.567 0.252 0.783 ;
    END
  END D2
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.936 0.29 0.954 ;
        RECT 0.234 1.035 0.271 1.053 ;
        RECT 0.234 0.837 0.271 0.855 ;
        RECT 0.234 0.837 0.252 1.053 ;
    END
  END D3
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.225 1.171 0.243 ;
        RECT 1.153 0.027 1.171 0.243 ;
        RECT 1.012 0.027 1.171 0.045 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.495 1.171 0.513 ;
        RECT 1.153 0.297 1.171 0.513 ;
        RECT 1.012 0.297 1.171 0.315 ;
    END
  END QN1
  PIN QN2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.765 1.171 0.783 ;
        RECT 1.153 0.567 1.171 0.783 ;
        RECT 1.012 0.567 1.171 0.585 ;
    END
  END QN2
  PIN QN3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 1.035 1.171 1.053 ;
        RECT 1.153 0.837 1.171 1.053 ;
        RECT 1.012 0.837 1.171 0.855 ;
    END
  END QN3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.188 0.279 ;
        RECT 0 0.801 1.188 0.819 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.188 0.009 ;
        RECT 0 0.531 1.188 0.549 ;
        RECT 0 1.071 1.188 1.089 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 0.04 0.07 0.122 0.088 ;
        RECT 0.04 0.452 0.122 0.47 ;
        RECT 0.04 0.61 0.122 0.628 ;
        RECT 0.04 0.992 0.122 1.01 ;
      LAYER M3 ;
        RECT 0.045 0.05 0.063 1.03 ;
      LAYER M1 ;
        RECT 0.099 0.164 0.117 0.236 ;
        RECT 0.072 0.07 0.117 0.106 ;
        RECT 0.099 0.034 0.117 0.106 ;
        RECT 0.072 0.164 0.117 0.2 ;
        RECT 0.072 0.07 0.09 0.2 ;
        RECT 0.099 0.434 0.117 0.506 ;
        RECT 0.072 0.34 0.117 0.376 ;
        RECT 0.099 0.304 0.117 0.376 ;
        RECT 0.072 0.434 0.117 0.47 ;
        RECT 0.072 0.34 0.09 0.47 ;
        RECT 0.099 0.704 0.117 0.776 ;
        RECT 0.072 0.61 0.117 0.646 ;
        RECT 0.099 0.574 0.117 0.646 ;
        RECT 0.072 0.704 0.117 0.74 ;
        RECT 0.072 0.61 0.09 0.74 ;
        RECT 0.099 0.974 0.117 1.046 ;
        RECT 0.072 0.88 0.117 0.916 ;
        RECT 0.099 0.844 0.117 0.916 ;
        RECT 0.072 0.974 0.117 1.01 ;
        RECT 0.072 0.88 0.09 1.01 ;
      LAYER V2 ;
        RECT 0.045 0.992 0.063 1.01 ;
        RECT 0.045 0.61 0.063 0.628 ;
        RECT 0.045 0.452 0.063 0.47 ;
        RECT 0.045 0.07 0.063 0.088 ;
      LAYER V1 ;
        RECT 0.099 0.992 0.117 1.01 ;
        RECT 0.099 0.61 0.117 0.628 ;
        RECT 0.099 0.452 0.117 0.47 ;
        RECT 0.099 0.07 0.117 0.088 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 0.85 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.774 0.027 0.792 0.119 ;
      RECT 0.774 0.027 0.954 0.045 ;
      RECT 0.774 0.495 0.954 0.513 ;
      RECT 0.936 0.297 0.954 0.513 ;
      RECT 0.774 0.421 0.792 0.513 ;
      RECT 0.85 0.297 0.954 0.315 ;
      RECT 0.85 0.765 0.954 0.783 ;
      RECT 0.936 0.567 0.954 0.783 ;
      RECT 0.774 0.567 0.792 0.659 ;
      RECT 0.774 0.567 0.954 0.585 ;
      RECT 0.774 1.035 0.954 1.053 ;
      RECT 0.936 0.837 0.954 1.053 ;
      RECT 0.774 0.961 0.792 1.053 ;
      RECT 0.85 0.837 0.954 0.855 ;
      RECT 0.688 0.224 0.738 0.242 ;
      RECT 0.72 0.027 0.738 0.242 ;
      RECT 0.72 0.153 0.9 0.171 ;
      RECT 0.882 0.117 0.9 0.171 ;
      RECT 0.828 0.117 0.846 0.171 ;
      RECT 0.634 0.027 0.738 0.045 ;
      RECT 0.634 0.495 0.738 0.513 ;
      RECT 0.72 0.298 0.738 0.513 ;
      RECT 0.882 0.369 0.9 0.423 ;
      RECT 0.828 0.369 0.846 0.423 ;
      RECT 0.72 0.369 0.9 0.387 ;
      RECT 0.688 0.298 0.738 0.316 ;
      RECT 0.688 0.764 0.738 0.782 ;
      RECT 0.72 0.567 0.738 0.782 ;
      RECT 0.72 0.693 0.9 0.711 ;
      RECT 0.882 0.657 0.9 0.711 ;
      RECT 0.828 0.657 0.846 0.711 ;
      RECT 0.634 0.567 0.738 0.585 ;
      RECT 0.634 1.035 0.738 1.053 ;
      RECT 0.72 0.838 0.738 1.053 ;
      RECT 0.882 0.909 0.9 0.963 ;
      RECT 0.828 0.909 0.846 0.963 ;
      RECT 0.72 0.909 0.9 0.927 ;
      RECT 0.688 0.838 0.738 0.856 ;
      RECT 0.576 0.225 0.63 0.243 ;
      RECT 0.612 0.081 0.63 0.243 ;
      RECT 0.496 0.081 0.63 0.099 ;
      RECT 0.585 0.045 0.603 0.099 ;
      RECT 0.585 0.441 0.603 0.495 ;
      RECT 0.496 0.441 0.63 0.459 ;
      RECT 0.612 0.297 0.63 0.459 ;
      RECT 0.576 0.297 0.63 0.315 ;
      RECT 0.576 0.765 0.63 0.783 ;
      RECT 0.612 0.621 0.63 0.783 ;
      RECT 0.496 0.621 0.63 0.639 ;
      RECT 0.585 0.585 0.603 0.639 ;
      RECT 0.585 0.981 0.603 1.035 ;
      RECT 0.496 0.981 0.63 0.999 ;
      RECT 0.612 0.837 0.63 0.999 ;
      RECT 0.576 0.837 0.63 0.855 ;
      RECT 0.364 0.225 0.468 0.243 ;
      RECT 0.45 0.027 0.468 0.243 ;
      RECT 0.45 0.122 0.576 0.14 ;
      RECT 0.418 0.027 0.468 0.045 ;
      RECT 0.418 0.495 0.468 0.513 ;
      RECT 0.45 0.297 0.468 0.513 ;
      RECT 0.45 0.4 0.576 0.418 ;
      RECT 0.364 0.297 0.468 0.315 ;
      RECT 0.364 0.765 0.468 0.783 ;
      RECT 0.45 0.567 0.468 0.783 ;
      RECT 0.45 0.662 0.576 0.68 ;
      RECT 0.418 0.567 0.468 0.585 ;
      RECT 0.418 1.035 0.468 1.053 ;
      RECT 0.45 0.837 0.468 1.053 ;
      RECT 0.45 0.94 0.576 0.958 ;
      RECT 0.364 0.837 0.468 0.855 ;
      RECT 0.315 0.126 0.333 0.203 ;
      RECT 0.315 0.126 0.367 0.144 ;
      RECT 0.315 0.396 0.367 0.414 ;
      RECT 0.315 0.337 0.333 0.414 ;
      RECT 0.315 0.666 0.333 0.743 ;
      RECT 0.315 0.666 0.367 0.684 ;
      RECT 0.315 0.936 0.367 0.954 ;
      RECT 0.315 0.877 0.333 0.954 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.148 0.495 0.198 0.513 ;
      RECT 0.18 0.297 0.198 0.513 ;
      RECT 0.148 0.297 0.198 0.315 ;
      RECT 0.148 0.765 0.198 0.783 ;
      RECT 0.18 0.567 0.198 0.783 ;
      RECT 0.148 0.567 0.198 0.585 ;
      RECT 0.148 1.035 0.198 1.053 ;
      RECT 0.18 0.837 0.198 1.053 ;
      RECT 0.148 0.837 0.198 0.855 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.144 0.047 0.162 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 0.009 0.495 0.068 0.513 ;
      RECT 0.009 0.297 0.027 0.513 ;
      RECT 0.009 0.378 0.047 0.396 ;
      RECT 0.009 0.297 0.068 0.315 ;
      RECT 0.009 0.765 0.068 0.783 ;
      RECT 0.009 0.567 0.027 0.783 ;
      RECT 0.009 0.684 0.047 0.702 ;
      RECT 0.009 0.567 0.068 0.585 ;
      RECT 0.009 1.035 0.068 1.053 ;
      RECT 0.009 0.837 0.027 1.053 ;
      RECT 0.009 0.918 0.047 0.936 ;
      RECT 0.009 0.837 0.068 0.855 ;
      RECT 0.99 0.122 1.008 0.167 ;
      RECT 0.99 0.373 1.008 0.418 ;
      RECT 0.99 0.662 1.008 0.707 ;
      RECT 0.99 0.913 1.008 0.958 ;
      RECT 0.666 0.101 0.684 0.167 ;
      RECT 0.666 0.373 0.684 0.439 ;
      RECT 0.666 0.641 0.684 0.707 ;
      RECT 0.666 0.913 0.684 0.979 ;
      RECT 0.504 0.165 0.522 0.203 ;
      RECT 0.504 0.337 0.522 0.375 ;
      RECT 0.504 0.705 0.522 0.743 ;
      RECT 0.504 0.877 0.522 0.915 ;
      RECT 0.396 0.106 0.414 0.167 ;
      RECT 0.396 0.373 0.414 0.434 ;
      RECT 0.396 0.646 0.414 0.707 ;
      RECT 0.396 0.913 0.414 0.974 ;
      RECT 0.142 0.106 0.16 0.167 ;
      RECT 0.142 0.373 0.16 0.434 ;
      RECT 0.142 0.646 0.16 0.707 ;
      RECT 0.142 0.913 0.16 0.974 ;
    LAYER M2 ;
      RECT 0.877 0.144 1.013 0.162 ;
      RECT 0.877 0.378 1.013 0.396 ;
      RECT 0.877 0.684 1.013 0.702 ;
      RECT 0.877 0.918 1.013 0.936 ;
      RECT 0.019 0.144 0.689 0.162 ;
      RECT 0.019 0.378 0.689 0.396 ;
      RECT 0.019 0.684 0.689 0.702 ;
      RECT 0.019 0.918 0.689 0.936 ;
      RECT 0.175 0.18 0.527 0.198 ;
      RECT 0.175 0.342 0.527 0.36 ;
      RECT 0.175 0.72 0.527 0.738 ;
      RECT 0.175 0.882 0.527 0.9 ;
    LAYER V1 ;
      RECT 0.99 0.144 1.008 0.162 ;
      RECT 0.99 0.378 1.008 0.396 ;
      RECT 0.99 0.684 1.008 0.702 ;
      RECT 0.99 0.918 1.008 0.936 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.882 0.378 0.9 0.396 ;
      RECT 0.882 0.684 0.9 0.702 ;
      RECT 0.882 0.918 0.9 0.936 ;
      RECT 0.666 0.144 0.684 0.162 ;
      RECT 0.666 0.378 0.684 0.396 ;
      RECT 0.666 0.684 0.684 0.702 ;
      RECT 0.666 0.918 0.684 0.936 ;
      RECT 0.504 0.18 0.522 0.198 ;
      RECT 0.504 0.342 0.522 0.36 ;
      RECT 0.504 0.72 0.522 0.738 ;
      RECT 0.504 0.882 0.522 0.9 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.396 0.378 0.414 0.396 ;
      RECT 0.396 0.684 0.414 0.702 ;
      RECT 0.396 0.918 0.414 0.936 ;
      RECT 0.315 0.18 0.333 0.198 ;
      RECT 0.315 0.342 0.333 0.36 ;
      RECT 0.315 0.72 0.333 0.738 ;
      RECT 0.315 0.882 0.333 0.9 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.18 0.342 0.198 0.36 ;
      RECT 0.18 0.72 0.198 0.738 ;
      RECT 0.18 0.882 0.198 0.9 ;
      RECT 0.142 0.144 0.16 0.162 ;
      RECT 0.142 0.378 0.16 0.396 ;
      RECT 0.142 0.684 0.16 0.702 ;
      RECT 0.142 0.918 0.16 0.936 ;
      RECT 0.024 0.144 0.042 0.162 ;
      RECT 0.024 0.378 0.042 0.396 ;
      RECT 0.024 0.684 0.042 0.702 ;
      RECT 0.024 0.918 0.042 0.936 ;
  END
END DFFHQNV4Xx3_ASAP7_75t_R

MACRO DFFHQNV4Xx3_ASAP7_75t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNV4Xx3_ASAP7_75t_SL 0 0 ;
  SIZE 1.188 BY 1.08 ;
  SYMMETRY X Y ;
  SITE asap7sc7p5t ;
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.126 0.29 0.144 ;
        RECT 0.234 0.225 0.271 0.243 ;
        RECT 0.234 0.027 0.271 0.045 ;
        RECT 0.234 0.027 0.252 0.243 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.396 0.29 0.414 ;
        RECT 0.234 0.495 0.271 0.513 ;
        RECT 0.234 0.297 0.271 0.315 ;
        RECT 0.234 0.297 0.252 0.513 ;
    END
  END D1
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.666 0.29 0.684 ;
        RECT 0.234 0.765 0.271 0.783 ;
        RECT 0.234 0.567 0.271 0.585 ;
        RECT 0.234 0.567 0.252 0.783 ;
    END
  END D2
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.936 0.29 0.954 ;
        RECT 0.234 1.035 0.271 1.053 ;
        RECT 0.234 0.837 0.271 0.855 ;
        RECT 0.234 0.837 0.252 1.053 ;
    END
  END D3
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.225 1.171 0.243 ;
        RECT 1.153 0.027 1.171 0.243 ;
        RECT 1.012 0.027 1.171 0.045 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.495 1.171 0.513 ;
        RECT 1.153 0.297 1.171 0.513 ;
        RECT 1.012 0.297 1.171 0.315 ;
    END
  END QN1
  PIN QN2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 0.765 1.171 0.783 ;
        RECT 1.153 0.567 1.171 0.783 ;
        RECT 1.012 0.567 1.171 0.585 ;
    END
  END QN2
  PIN QN3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.012 1.035 1.171 1.053 ;
        RECT 1.153 0.837 1.171 1.053 ;
        RECT 1.012 0.837 1.171 0.855 ;
    END
  END QN3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.188 0.279 ;
        RECT 0 0.801 1.188 0.819 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.188 0.009 ;
        RECT 0 0.531 1.188 0.549 ;
        RECT 0 1.071 1.188 1.089 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 0.04 0.07 0.122 0.088 ;
        RECT 0.04 0.452 0.122 0.47 ;
        RECT 0.04 0.61 0.122 0.628 ;
        RECT 0.04 0.992 0.122 1.01 ;
      LAYER M3 ;
        RECT 0.045 0.05 0.063 1.03 ;
      LAYER M1 ;
        RECT 0.099 0.164 0.117 0.236 ;
        RECT 0.072 0.07 0.117 0.106 ;
        RECT 0.099 0.034 0.117 0.106 ;
        RECT 0.072 0.164 0.117 0.2 ;
        RECT 0.072 0.07 0.09 0.2 ;
        RECT 0.099 0.434 0.117 0.506 ;
        RECT 0.072 0.34 0.117 0.376 ;
        RECT 0.099 0.304 0.117 0.376 ;
        RECT 0.072 0.434 0.117 0.47 ;
        RECT 0.072 0.34 0.09 0.47 ;
        RECT 0.099 0.704 0.117 0.776 ;
        RECT 0.072 0.61 0.117 0.646 ;
        RECT 0.099 0.574 0.117 0.646 ;
        RECT 0.072 0.704 0.117 0.74 ;
        RECT 0.072 0.61 0.09 0.74 ;
        RECT 0.099 0.974 0.117 1.046 ;
        RECT 0.072 0.88 0.117 0.916 ;
        RECT 0.099 0.844 0.117 0.916 ;
        RECT 0.072 0.974 0.117 1.01 ;
        RECT 0.072 0.88 0.09 1.01 ;
      LAYER V2 ;
        RECT 0.045 0.992 0.063 1.01 ;
        RECT 0.045 0.61 0.063 0.628 ;
        RECT 0.045 0.452 0.063 0.47 ;
        RECT 0.045 0.07 0.063 0.088 ;
      LAYER V1 ;
        RECT 0.099 0.992 0.117 1.01 ;
        RECT 0.099 0.61 0.117 0.628 ;
        RECT 0.099 0.452 0.117 0.47 ;
        RECT 0.099 0.07 0.117 0.088 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 0.85 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.774 0.027 0.792 0.119 ;
      RECT 0.774 0.027 0.954 0.045 ;
      RECT 0.774 0.495 0.954 0.513 ;
      RECT 0.936 0.297 0.954 0.513 ;
      RECT 0.774 0.421 0.792 0.513 ;
      RECT 0.85 0.297 0.954 0.315 ;
      RECT 0.85 0.765 0.954 0.783 ;
      RECT 0.936 0.567 0.954 0.783 ;
      RECT 0.774 0.567 0.792 0.659 ;
      RECT 0.774 0.567 0.954 0.585 ;
      RECT 0.774 1.035 0.954 1.053 ;
      RECT 0.936 0.837 0.954 1.053 ;
      RECT 0.774 0.961 0.792 1.053 ;
      RECT 0.85 0.837 0.954 0.855 ;
      RECT 0.688 0.224 0.738 0.242 ;
      RECT 0.72 0.027 0.738 0.242 ;
      RECT 0.72 0.153 0.9 0.171 ;
      RECT 0.882 0.117 0.9 0.171 ;
      RECT 0.828 0.117 0.846 0.171 ;
      RECT 0.634 0.027 0.738 0.045 ;
      RECT 0.634 0.495 0.738 0.513 ;
      RECT 0.72 0.298 0.738 0.513 ;
      RECT 0.882 0.369 0.9 0.423 ;
      RECT 0.828 0.369 0.846 0.423 ;
      RECT 0.72 0.369 0.9 0.387 ;
      RECT 0.688 0.298 0.738 0.316 ;
      RECT 0.688 0.764 0.738 0.782 ;
      RECT 0.72 0.567 0.738 0.782 ;
      RECT 0.72 0.693 0.9 0.711 ;
      RECT 0.882 0.657 0.9 0.711 ;
      RECT 0.828 0.657 0.846 0.711 ;
      RECT 0.634 0.567 0.738 0.585 ;
      RECT 0.634 1.035 0.738 1.053 ;
      RECT 0.72 0.838 0.738 1.053 ;
      RECT 0.882 0.909 0.9 0.963 ;
      RECT 0.828 0.909 0.846 0.963 ;
      RECT 0.72 0.909 0.9 0.927 ;
      RECT 0.688 0.838 0.738 0.856 ;
      RECT 0.576 0.225 0.63 0.243 ;
      RECT 0.612 0.081 0.63 0.243 ;
      RECT 0.496 0.081 0.63 0.099 ;
      RECT 0.585 0.045 0.603 0.099 ;
      RECT 0.585 0.441 0.603 0.495 ;
      RECT 0.496 0.441 0.63 0.459 ;
      RECT 0.612 0.297 0.63 0.459 ;
      RECT 0.576 0.297 0.63 0.315 ;
      RECT 0.576 0.765 0.63 0.783 ;
      RECT 0.612 0.621 0.63 0.783 ;
      RECT 0.496 0.621 0.63 0.639 ;
      RECT 0.585 0.585 0.603 0.639 ;
      RECT 0.585 0.981 0.603 1.035 ;
      RECT 0.496 0.981 0.63 0.999 ;
      RECT 0.612 0.837 0.63 0.999 ;
      RECT 0.576 0.837 0.63 0.855 ;
      RECT 0.364 0.225 0.468 0.243 ;
      RECT 0.45 0.027 0.468 0.243 ;
      RECT 0.45 0.122 0.576 0.14 ;
      RECT 0.418 0.027 0.468 0.045 ;
      RECT 0.418 0.495 0.468 0.513 ;
      RECT 0.45 0.297 0.468 0.513 ;
      RECT 0.45 0.4 0.576 0.418 ;
      RECT 0.364 0.297 0.468 0.315 ;
      RECT 0.364 0.765 0.468 0.783 ;
      RECT 0.45 0.567 0.468 0.783 ;
      RECT 0.45 0.662 0.576 0.68 ;
      RECT 0.418 0.567 0.468 0.585 ;
      RECT 0.418 1.035 0.468 1.053 ;
      RECT 0.45 0.837 0.468 1.053 ;
      RECT 0.45 0.94 0.576 0.958 ;
      RECT 0.364 0.837 0.468 0.855 ;
      RECT 0.315 0.126 0.333 0.203 ;
      RECT 0.315 0.126 0.367 0.144 ;
      RECT 0.315 0.396 0.367 0.414 ;
      RECT 0.315 0.337 0.333 0.414 ;
      RECT 0.315 0.666 0.333 0.743 ;
      RECT 0.315 0.666 0.367 0.684 ;
      RECT 0.315 0.936 0.367 0.954 ;
      RECT 0.315 0.877 0.333 0.954 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.148 0.495 0.198 0.513 ;
      RECT 0.18 0.297 0.198 0.513 ;
      RECT 0.148 0.297 0.198 0.315 ;
      RECT 0.148 0.765 0.198 0.783 ;
      RECT 0.18 0.567 0.198 0.783 ;
      RECT 0.148 0.567 0.198 0.585 ;
      RECT 0.148 1.035 0.198 1.053 ;
      RECT 0.18 0.837 0.198 1.053 ;
      RECT 0.148 0.837 0.198 0.855 ;
      RECT 0.009 0.225 0.068 0.243 ;
      RECT 0.009 0.027 0.027 0.243 ;
      RECT 0.009 0.144 0.047 0.162 ;
      RECT 0.009 0.027 0.068 0.045 ;
      RECT 0.009 0.495 0.068 0.513 ;
      RECT 0.009 0.297 0.027 0.513 ;
      RECT 0.009 0.378 0.047 0.396 ;
      RECT 0.009 0.297 0.068 0.315 ;
      RECT 0.009 0.765 0.068 0.783 ;
      RECT 0.009 0.567 0.027 0.783 ;
      RECT 0.009 0.684 0.047 0.702 ;
      RECT 0.009 0.567 0.068 0.585 ;
      RECT 0.009 1.035 0.068 1.053 ;
      RECT 0.009 0.837 0.027 1.053 ;
      RECT 0.009 0.918 0.047 0.936 ;
      RECT 0.009 0.837 0.068 0.855 ;
      RECT 0.99 0.122 1.008 0.167 ;
      RECT 0.99 0.373 1.008 0.418 ;
      RECT 0.99 0.662 1.008 0.707 ;
      RECT 0.99 0.913 1.008 0.958 ;
      RECT 0.666 0.101 0.684 0.167 ;
      RECT 0.666 0.373 0.684 0.439 ;
      RECT 0.666 0.641 0.684 0.707 ;
      RECT 0.666 0.913 0.684 0.979 ;
      RECT 0.504 0.165 0.522 0.203 ;
      RECT 0.504 0.337 0.522 0.375 ;
      RECT 0.504 0.705 0.522 0.743 ;
      RECT 0.504 0.877 0.522 0.915 ;
      RECT 0.396 0.106 0.414 0.167 ;
      RECT 0.396 0.373 0.414 0.434 ;
      RECT 0.396 0.646 0.414 0.707 ;
      RECT 0.396 0.913 0.414 0.974 ;
      RECT 0.142 0.106 0.16 0.167 ;
      RECT 0.142 0.373 0.16 0.434 ;
      RECT 0.142 0.646 0.16 0.707 ;
      RECT 0.142 0.913 0.16 0.974 ;
    LAYER M2 ;
      RECT 0.877 0.144 1.013 0.162 ;
      RECT 0.877 0.378 1.013 0.396 ;
      RECT 0.877 0.684 1.013 0.702 ;
      RECT 0.877 0.918 1.013 0.936 ;
      RECT 0.019 0.144 0.689 0.162 ;
      RECT 0.019 0.378 0.689 0.396 ;
      RECT 0.019 0.684 0.689 0.702 ;
      RECT 0.019 0.918 0.689 0.936 ;
      RECT 0.175 0.18 0.527 0.198 ;
      RECT 0.175 0.342 0.527 0.36 ;
      RECT 0.175 0.72 0.527 0.738 ;
      RECT 0.175 0.882 0.527 0.9 ;
    LAYER V1 ;
      RECT 0.99 0.144 1.008 0.162 ;
      RECT 0.99 0.378 1.008 0.396 ;
      RECT 0.99 0.684 1.008 0.702 ;
      RECT 0.99 0.918 1.008 0.936 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.882 0.378 0.9 0.396 ;
      RECT 0.882 0.684 0.9 0.702 ;
      RECT 0.882 0.918 0.9 0.936 ;
      RECT 0.666 0.144 0.684 0.162 ;
      RECT 0.666 0.378 0.684 0.396 ;
      RECT 0.666 0.684 0.684 0.702 ;
      RECT 0.666 0.918 0.684 0.936 ;
      RECT 0.504 0.18 0.522 0.198 ;
      RECT 0.504 0.342 0.522 0.36 ;
      RECT 0.504 0.72 0.522 0.738 ;
      RECT 0.504 0.882 0.522 0.9 ;
      RECT 0.396 0.144 0.414 0.162 ;
      RECT 0.396 0.378 0.414 0.396 ;
      RECT 0.396 0.684 0.414 0.702 ;
      RECT 0.396 0.918 0.414 0.936 ;
      RECT 0.315 0.18 0.333 0.198 ;
      RECT 0.315 0.342 0.333 0.36 ;
      RECT 0.315 0.72 0.333 0.738 ;
      RECT 0.315 0.882 0.333 0.9 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.18 0.342 0.198 0.36 ;
      RECT 0.18 0.72 0.198 0.738 ;
      RECT 0.18 0.882 0.198 0.9 ;
      RECT 0.142 0.144 0.16 0.162 ;
      RECT 0.142 0.378 0.16 0.396 ;
      RECT 0.142 0.684 0.16 0.702 ;
      RECT 0.142 0.918 0.16 0.936 ;
      RECT 0.024 0.144 0.042 0.162 ;
      RECT 0.024 0.378 0.042 0.396 ;
      RECT 0.024 0.684 0.042 0.702 ;
      RECT 0.024 0.918 0.042 0.936 ;
  END
END DFFHQNV4Xx3_ASAP7_75t_SL

END LIBRARY
