(* blackbox *)
module fakeram7_64x25 (
   output reg [24:0] rd_out,
   input [5:0] addr_in,
   input we_in,
   input [24:0] wd_in,
   input clk,
   input ce_in
);
endmodule
