(* blackbox *) module O2A1O1Ixp33_ASAP7_75t_SL (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module O2A1O1Ixp5_ASAP7_75t_SL (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module OA211x2_ASAP7_75t_SL (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module OA21x2_ASAP7_75t_SL (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module OA221x2_ASAP7_75t_SL (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module OA222x2_ASAP7_75t_SL (Y, A1, A2, B1, B2, C1, C2);
	output Y;
	input A1, A2, B1, B2, C1, C2;
endmodule
(* blackbox *) module OA22x2_ASAP7_75t_SL (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module OA31x2_ASAP7_75t_SL (Y, A1, A2, A3, B1);
	output Y;
	input A1, A2, A3, B1;
endmodule
(* blackbox *) module OA331x1_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1;
endmodule
(* blackbox *) module OA331x2_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1;
endmodule
(* blackbox *) module OA332x1_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module OA332x2_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module OA333x1_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module OA333x2_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module OA33x2_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3);
	output Y;
	input A1, A2, A3, B1, B2, B3;
endmodule
(* blackbox *) module OAI211xp5_ASAP7_75t_SL (Y, A1, A2, B, C);
	output Y;
	input A1, A2, B, C;
endmodule
(* blackbox *) module OAI21x1_ASAP7_75t_SL (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module OAI21xp33_ASAP7_75t_SL (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module OAI21xp5_ASAP7_75t_SL (Y, A1, A2, B);
	output Y;
	input A1, A2, B;
endmodule
(* blackbox *) module OAI221xp5_ASAP7_75t_SL (Y, A1, A2, B1, B2, C);
	output Y;
	input A1, A2, B1, B2, C;
endmodule
(* blackbox *) module OAI222xp33_ASAP7_75t_SL (Y, A1, A2, B1, B2, C1, C2);
	output Y;
	input A1, A2, B1, B2, C1, C2;
endmodule
(* blackbox *) module OAI22x1_ASAP7_75t_SL (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module OAI22xp33_ASAP7_75t_SL (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module OAI22xp5_ASAP7_75t_SL (Y, A1, A2, B1, B2);
	output Y;
	input A1, A2, B1, B2;
endmodule
(* blackbox *) module OAI311xp33_ASAP7_75t_SL (Y, A1, A2, A3, B1, C1);
	output Y;
	input A1, A2, A3, B1, C1;
endmodule
(* blackbox *) module OAI31xp33_ASAP7_75t_SL (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module OAI31xp67_ASAP7_75t_SL (Y, A1, A2, A3, B);
	output Y;
	input A1, A2, A3, B;
endmodule
(* blackbox *) module OAI321xp33_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, C);
	output Y;
	input A1, A2, A3, B1, B2, C;
endmodule
(* blackbox *) module OAI322xp33_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, C1, C2;
endmodule
(* blackbox *) module OAI32xp33_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2);
	output Y;
	input A1, A2, A3, B1, B2;
endmodule
(* blackbox *) module OAI331xp33_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1;
endmodule
(* blackbox *) module OAI332xp33_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1, C2);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2;
endmodule
(* blackbox *) module OAI333xp33_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3, C1, C2, C3);
	output Y;
	input A1, A2, A3, B1, B2, B3, C1, C2, C3;
endmodule
(* blackbox *) module OAI33xp33_ASAP7_75t_SL (Y, A1, A2, A3, B1, B2, B3);
	output Y;
	input A1, A2, A3, B1, B2, B3;
endmodule
