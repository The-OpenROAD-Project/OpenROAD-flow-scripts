module MockArray(
  input         clock,
  input         reset,
  input  [63:0] io_insHorizontal_0_0,
  input  [63:0] io_insHorizontal_0_1,
  input  [63:0] io_insHorizontal_0_2,
  input  [63:0] io_insHorizontal_0_3,
  input  [63:0] io_insHorizontal_0_4,
  input  [63:0] io_insHorizontal_0_5,
  input  [63:0] io_insHorizontal_0_6,
  input  [63:0] io_insHorizontal_0_7,
  input  [63:0] io_insHorizontal_0_8,
  input  [63:0] io_insHorizontal_0_9,
  input  [63:0] io_insHorizontal_0_10,
  input  [63:0] io_insHorizontal_0_11,
  input  [63:0] io_insHorizontal_0_12,
  input  [63:0] io_insHorizontal_0_13,
  input  [63:0] io_insHorizontal_0_14,
  input  [63:0] io_insHorizontal_0_15,
  input  [63:0] io_insHorizontal_1_0,
  input  [63:0] io_insHorizontal_1_1,
  input  [63:0] io_insHorizontal_1_2,
  input  [63:0] io_insHorizontal_1_3,
  input  [63:0] io_insHorizontal_1_4,
  input  [63:0] io_insHorizontal_1_5,
  input  [63:0] io_insHorizontal_1_6,
  input  [63:0] io_insHorizontal_1_7,
  input  [63:0] io_insHorizontal_1_8,
  input  [63:0] io_insHorizontal_1_9,
  input  [63:0] io_insHorizontal_1_10,
  input  [63:0] io_insHorizontal_1_11,
  input  [63:0] io_insHorizontal_1_12,
  input  [63:0] io_insHorizontal_1_13,
  input  [63:0] io_insHorizontal_1_14,
  input  [63:0] io_insHorizontal_1_15,
  output [63:0] io_outsHorizontal_0_0,
  output [63:0] io_outsHorizontal_0_1,
  output [63:0] io_outsHorizontal_0_2,
  output [63:0] io_outsHorizontal_0_3,
  output [63:0] io_outsHorizontal_0_4,
  output [63:0] io_outsHorizontal_0_5,
  output [63:0] io_outsHorizontal_0_6,
  output [63:0] io_outsHorizontal_0_7,
  output [63:0] io_outsHorizontal_0_8,
  output [63:0] io_outsHorizontal_0_9,
  output [63:0] io_outsHorizontal_0_10,
  output [63:0] io_outsHorizontal_0_11,
  output [63:0] io_outsHorizontal_0_12,
  output [63:0] io_outsHorizontal_0_13,
  output [63:0] io_outsHorizontal_0_14,
  output [63:0] io_outsHorizontal_0_15,
  output [63:0] io_outsHorizontal_1_0,
  output [63:0] io_outsHorizontal_1_1,
  output [63:0] io_outsHorizontal_1_2,
  output [63:0] io_outsHorizontal_1_3,
  output [63:0] io_outsHorizontal_1_4,
  output [63:0] io_outsHorizontal_1_5,
  output [63:0] io_outsHorizontal_1_6,
  output [63:0] io_outsHorizontal_1_7,
  output [63:0] io_outsHorizontal_1_8,
  output [63:0] io_outsHorizontal_1_9,
  output [63:0] io_outsHorizontal_1_10,
  output [63:0] io_outsHorizontal_1_11,
  output [63:0] io_outsHorizontal_1_12,
  output [63:0] io_outsHorizontal_1_13,
  output [63:0] io_outsHorizontal_1_14,
  output [63:0] io_outsHorizontal_1_15,
  input  [63:0] io_insVertical_0_0,
  input  [63:0] io_insVertical_0_1,
  input  [63:0] io_insVertical_0_2,
  input  [63:0] io_insVertical_0_3,
  input  [63:0] io_insVertical_0_4,
  input  [63:0] io_insVertical_0_5,
  input  [63:0] io_insVertical_0_6,
  input  [63:0] io_insVertical_0_7,
  input  [63:0] io_insVertical_1_0,
  input  [63:0] io_insVertical_1_1,
  input  [63:0] io_insVertical_1_2,
  input  [63:0] io_insVertical_1_3,
  input  [63:0] io_insVertical_1_4,
  input  [63:0] io_insVertical_1_5,
  input  [63:0] io_insVertical_1_6,
  input  [63:0] io_insVertical_1_7,
  output [63:0] io_outsVertical_0_0,
  output [63:0] io_outsVertical_0_1,
  output [63:0] io_outsVertical_0_2,
  output [63:0] io_outsVertical_0_3,
  output [63:0] io_outsVertical_0_4,
  output [63:0] io_outsVertical_0_5,
  output [63:0] io_outsVertical_0_6,
  output [63:0] io_outsVertical_0_7,
  output [63:0] io_outsVertical_1_0,
  output [63:0] io_outsVertical_1_1,
  output [63:0] io_outsVertical_1_2,
  output [63:0] io_outsVertical_1_3,
  output [63:0] io_outsVertical_1_4,
  output [63:0] io_outsVertical_1_5,
  output [63:0] io_outsVertical_1_6,
  output [63:0] io_outsVertical_1_7,
  output        io_lsbs_0,
  output        io_lsbs_1,
  output        io_lsbs_2,
  output        io_lsbs_3,
  output        io_lsbs_4,
  output        io_lsbs_5,
  output        io_lsbs_6,
  output        io_lsbs_7,
  output        io_lsbs_8,
  output        io_lsbs_9,
  output        io_lsbs_10,
  output        io_lsbs_11,
  output        io_lsbs_12,
  output        io_lsbs_13,
  output        io_lsbs_14,
  output        io_lsbs_15,
  output        io_lsbs_16,
  output        io_lsbs_17,
  output        io_lsbs_18,
  output        io_lsbs_19,
  output        io_lsbs_20,
  output        io_lsbs_21,
  output        io_lsbs_22,
  output        io_lsbs_23,
  output        io_lsbs_24,
  output        io_lsbs_25,
  output        io_lsbs_26,
  output        io_lsbs_27,
  output        io_lsbs_28,
  output        io_lsbs_29,
  output        io_lsbs_30,
  output        io_lsbs_31,
  output        io_lsbs_32,
  output        io_lsbs_33,
  output        io_lsbs_34,
  output        io_lsbs_35,
  output        io_lsbs_36,
  output        io_lsbs_37,
  output        io_lsbs_38,
  output        io_lsbs_39,
  output        io_lsbs_40,
  output        io_lsbs_41,
  output        io_lsbs_42,
  output        io_lsbs_43,
  output        io_lsbs_44,
  output        io_lsbs_45,
  output        io_lsbs_46,
  output        io_lsbs_47,
  output        io_lsbs_48,
  output        io_lsbs_49,
  output        io_lsbs_50,
  output        io_lsbs_51,
  output        io_lsbs_52,
  output        io_lsbs_53,
  output        io_lsbs_54,
  output        io_lsbs_55,
  output        io_lsbs_56,
  output        io_lsbs_57,
  output        io_lsbs_58,
  output        io_lsbs_59,
  output        io_lsbs_60,
  output        io_lsbs_61,
  output        io_lsbs_62,
  output        io_lsbs_63,
  output        io_lsbs_64,
  output        io_lsbs_65,
  output        io_lsbs_66,
  output        io_lsbs_67,
  output        io_lsbs_68,
  output        io_lsbs_69,
  output        io_lsbs_70,
  output        io_lsbs_71,
  output        io_lsbs_72,
  output        io_lsbs_73,
  output        io_lsbs_74,
  output        io_lsbs_75,
  output        io_lsbs_76,
  output        io_lsbs_77,
  output        io_lsbs_78,
  output        io_lsbs_79,
  output        io_lsbs_80,
  output        io_lsbs_81,
  output        io_lsbs_82,
  output        io_lsbs_83,
  output        io_lsbs_84,
  output        io_lsbs_85,
  output        io_lsbs_86,
  output        io_lsbs_87,
  output        io_lsbs_88,
  output        io_lsbs_89,
  output        io_lsbs_90,
  output        io_lsbs_91,
  output        io_lsbs_92,
  output        io_lsbs_93,
  output        io_lsbs_94,
  output        io_lsbs_95,
  output        io_lsbs_96,
  output        io_lsbs_97,
  output        io_lsbs_98,
  output        io_lsbs_99,
  output        io_lsbs_100,
  output        io_lsbs_101,
  output        io_lsbs_102,
  output        io_lsbs_103,
  output        io_lsbs_104,
  output        io_lsbs_105,
  output        io_lsbs_106,
  output        io_lsbs_107,
  output        io_lsbs_108,
  output        io_lsbs_109,
  output        io_lsbs_110,
  output        io_lsbs_111,
  output        io_lsbs_112,
  output        io_lsbs_113,
  output        io_lsbs_114,
  output        io_lsbs_115,
  output        io_lsbs_116,
  output        io_lsbs_117,
  output        io_lsbs_118,
  output        io_lsbs_119,
  output        io_lsbs_120,
  output        io_lsbs_121,
  output        io_lsbs_122,
  output        io_lsbs_123,
  output        io_lsbs_124,
  output        io_lsbs_125,
  output        io_lsbs_126,
  output        io_lsbs_127
);
  wire  ces_0_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_15_io_outs_3; // @[MockArray.scala 36:52]
  Element ces_0_0 ( // @[MockArray.scala 36:52]
    .clock(ces_0_0_clock),
    .io_ins_0(ces_0_0_io_ins_0),
    .io_ins_1(ces_0_0_io_ins_1),
    .io_ins_2(ces_0_0_io_ins_2),
    .io_ins_3(ces_0_0_io_ins_3),
    .io_outs_0(ces_0_0_io_outs_0),
    .io_outs_1(ces_0_0_io_outs_1),
    .io_outs_2(ces_0_0_io_outs_2),
    .io_outs_3(ces_0_0_io_outs_3)
  );
  Element ces_0_1 ( // @[MockArray.scala 36:52]
    .clock(ces_0_1_clock),
    .io_ins_0(ces_0_1_io_ins_0),
    .io_ins_1(ces_0_1_io_ins_1),
    .io_ins_2(ces_0_1_io_ins_2),
    .io_ins_3(ces_0_1_io_ins_3),
    .io_outs_0(ces_0_1_io_outs_0),
    .io_outs_1(ces_0_1_io_outs_1),
    .io_outs_2(ces_0_1_io_outs_2),
    .io_outs_3(ces_0_1_io_outs_3)
  );
  Element ces_0_2 ( // @[MockArray.scala 36:52]
    .clock(ces_0_2_clock),
    .io_ins_0(ces_0_2_io_ins_0),
    .io_ins_1(ces_0_2_io_ins_1),
    .io_ins_2(ces_0_2_io_ins_2),
    .io_ins_3(ces_0_2_io_ins_3),
    .io_outs_0(ces_0_2_io_outs_0),
    .io_outs_1(ces_0_2_io_outs_1),
    .io_outs_2(ces_0_2_io_outs_2),
    .io_outs_3(ces_0_2_io_outs_3)
  );
  Element ces_0_3 ( // @[MockArray.scala 36:52]
    .clock(ces_0_3_clock),
    .io_ins_0(ces_0_3_io_ins_0),
    .io_ins_1(ces_0_3_io_ins_1),
    .io_ins_2(ces_0_3_io_ins_2),
    .io_ins_3(ces_0_3_io_ins_3),
    .io_outs_0(ces_0_3_io_outs_0),
    .io_outs_1(ces_0_3_io_outs_1),
    .io_outs_2(ces_0_3_io_outs_2),
    .io_outs_3(ces_0_3_io_outs_3)
  );
  Element ces_0_4 ( // @[MockArray.scala 36:52]
    .clock(ces_0_4_clock),
    .io_ins_0(ces_0_4_io_ins_0),
    .io_ins_1(ces_0_4_io_ins_1),
    .io_ins_2(ces_0_4_io_ins_2),
    .io_ins_3(ces_0_4_io_ins_3),
    .io_outs_0(ces_0_4_io_outs_0),
    .io_outs_1(ces_0_4_io_outs_1),
    .io_outs_2(ces_0_4_io_outs_2),
    .io_outs_3(ces_0_4_io_outs_3)
  );
  Element ces_0_5 ( // @[MockArray.scala 36:52]
    .clock(ces_0_5_clock),
    .io_ins_0(ces_0_5_io_ins_0),
    .io_ins_1(ces_0_5_io_ins_1),
    .io_ins_2(ces_0_5_io_ins_2),
    .io_ins_3(ces_0_5_io_ins_3),
    .io_outs_0(ces_0_5_io_outs_0),
    .io_outs_1(ces_0_5_io_outs_1),
    .io_outs_2(ces_0_5_io_outs_2),
    .io_outs_3(ces_0_5_io_outs_3)
  );
  Element ces_0_6 ( // @[MockArray.scala 36:52]
    .clock(ces_0_6_clock),
    .io_ins_0(ces_0_6_io_ins_0),
    .io_ins_1(ces_0_6_io_ins_1),
    .io_ins_2(ces_0_6_io_ins_2),
    .io_ins_3(ces_0_6_io_ins_3),
    .io_outs_0(ces_0_6_io_outs_0),
    .io_outs_1(ces_0_6_io_outs_1),
    .io_outs_2(ces_0_6_io_outs_2),
    .io_outs_3(ces_0_6_io_outs_3)
  );
  Element ces_0_7 ( // @[MockArray.scala 36:52]
    .clock(ces_0_7_clock),
    .io_ins_0(ces_0_7_io_ins_0),
    .io_ins_1(ces_0_7_io_ins_1),
    .io_ins_2(ces_0_7_io_ins_2),
    .io_ins_3(ces_0_7_io_ins_3),
    .io_outs_0(ces_0_7_io_outs_0),
    .io_outs_1(ces_0_7_io_outs_1),
    .io_outs_2(ces_0_7_io_outs_2),
    .io_outs_3(ces_0_7_io_outs_3)
  );
  Element ces_0_8 ( // @[MockArray.scala 36:52]
    .clock(ces_0_8_clock),
    .io_ins_0(ces_0_8_io_ins_0),
    .io_ins_1(ces_0_8_io_ins_1),
    .io_ins_2(ces_0_8_io_ins_2),
    .io_ins_3(ces_0_8_io_ins_3),
    .io_outs_0(ces_0_8_io_outs_0),
    .io_outs_1(ces_0_8_io_outs_1),
    .io_outs_2(ces_0_8_io_outs_2),
    .io_outs_3(ces_0_8_io_outs_3)
  );
  Element ces_0_9 ( // @[MockArray.scala 36:52]
    .clock(ces_0_9_clock),
    .io_ins_0(ces_0_9_io_ins_0),
    .io_ins_1(ces_0_9_io_ins_1),
    .io_ins_2(ces_0_9_io_ins_2),
    .io_ins_3(ces_0_9_io_ins_3),
    .io_outs_0(ces_0_9_io_outs_0),
    .io_outs_1(ces_0_9_io_outs_1),
    .io_outs_2(ces_0_9_io_outs_2),
    .io_outs_3(ces_0_9_io_outs_3)
  );
  Element ces_0_10 ( // @[MockArray.scala 36:52]
    .clock(ces_0_10_clock),
    .io_ins_0(ces_0_10_io_ins_0),
    .io_ins_1(ces_0_10_io_ins_1),
    .io_ins_2(ces_0_10_io_ins_2),
    .io_ins_3(ces_0_10_io_ins_3),
    .io_outs_0(ces_0_10_io_outs_0),
    .io_outs_1(ces_0_10_io_outs_1),
    .io_outs_2(ces_0_10_io_outs_2),
    .io_outs_3(ces_0_10_io_outs_3)
  );
  Element ces_0_11 ( // @[MockArray.scala 36:52]
    .clock(ces_0_11_clock),
    .io_ins_0(ces_0_11_io_ins_0),
    .io_ins_1(ces_0_11_io_ins_1),
    .io_ins_2(ces_0_11_io_ins_2),
    .io_ins_3(ces_0_11_io_ins_3),
    .io_outs_0(ces_0_11_io_outs_0),
    .io_outs_1(ces_0_11_io_outs_1),
    .io_outs_2(ces_0_11_io_outs_2),
    .io_outs_3(ces_0_11_io_outs_3)
  );
  Element ces_0_12 ( // @[MockArray.scala 36:52]
    .clock(ces_0_12_clock),
    .io_ins_0(ces_0_12_io_ins_0),
    .io_ins_1(ces_0_12_io_ins_1),
    .io_ins_2(ces_0_12_io_ins_2),
    .io_ins_3(ces_0_12_io_ins_3),
    .io_outs_0(ces_0_12_io_outs_0),
    .io_outs_1(ces_0_12_io_outs_1),
    .io_outs_2(ces_0_12_io_outs_2),
    .io_outs_3(ces_0_12_io_outs_3)
  );
  Element ces_0_13 ( // @[MockArray.scala 36:52]
    .clock(ces_0_13_clock),
    .io_ins_0(ces_0_13_io_ins_0),
    .io_ins_1(ces_0_13_io_ins_1),
    .io_ins_2(ces_0_13_io_ins_2),
    .io_ins_3(ces_0_13_io_ins_3),
    .io_outs_0(ces_0_13_io_outs_0),
    .io_outs_1(ces_0_13_io_outs_1),
    .io_outs_2(ces_0_13_io_outs_2),
    .io_outs_3(ces_0_13_io_outs_3)
  );
  Element ces_0_14 ( // @[MockArray.scala 36:52]
    .clock(ces_0_14_clock),
    .io_ins_0(ces_0_14_io_ins_0),
    .io_ins_1(ces_0_14_io_ins_1),
    .io_ins_2(ces_0_14_io_ins_2),
    .io_ins_3(ces_0_14_io_ins_3),
    .io_outs_0(ces_0_14_io_outs_0),
    .io_outs_1(ces_0_14_io_outs_1),
    .io_outs_2(ces_0_14_io_outs_2),
    .io_outs_3(ces_0_14_io_outs_3)
  );
  Element ces_0_15 ( // @[MockArray.scala 36:52]
    .clock(ces_0_15_clock),
    .io_ins_0(ces_0_15_io_ins_0),
    .io_ins_1(ces_0_15_io_ins_1),
    .io_ins_2(ces_0_15_io_ins_2),
    .io_ins_3(ces_0_15_io_ins_3),
    .io_outs_0(ces_0_15_io_outs_0),
    .io_outs_1(ces_0_15_io_outs_1),
    .io_outs_2(ces_0_15_io_outs_2),
    .io_outs_3(ces_0_15_io_outs_3)
  );
  Element ces_1_0 ( // @[MockArray.scala 36:52]
    .clock(ces_1_0_clock),
    .io_ins_0(ces_1_0_io_ins_0),
    .io_ins_1(ces_1_0_io_ins_1),
    .io_ins_2(ces_1_0_io_ins_2),
    .io_ins_3(ces_1_0_io_ins_3),
    .io_outs_0(ces_1_0_io_outs_0),
    .io_outs_1(ces_1_0_io_outs_1),
    .io_outs_2(ces_1_0_io_outs_2),
    .io_outs_3(ces_1_0_io_outs_3)
  );
  Element ces_1_1 ( // @[MockArray.scala 36:52]
    .clock(ces_1_1_clock),
    .io_ins_0(ces_1_1_io_ins_0),
    .io_ins_1(ces_1_1_io_ins_1),
    .io_ins_2(ces_1_1_io_ins_2),
    .io_ins_3(ces_1_1_io_ins_3),
    .io_outs_0(ces_1_1_io_outs_0),
    .io_outs_1(ces_1_1_io_outs_1),
    .io_outs_2(ces_1_1_io_outs_2),
    .io_outs_3(ces_1_1_io_outs_3)
  );
  Element ces_1_2 ( // @[MockArray.scala 36:52]
    .clock(ces_1_2_clock),
    .io_ins_0(ces_1_2_io_ins_0),
    .io_ins_1(ces_1_2_io_ins_1),
    .io_ins_2(ces_1_2_io_ins_2),
    .io_ins_3(ces_1_2_io_ins_3),
    .io_outs_0(ces_1_2_io_outs_0),
    .io_outs_1(ces_1_2_io_outs_1),
    .io_outs_2(ces_1_2_io_outs_2),
    .io_outs_3(ces_1_2_io_outs_3)
  );
  Element ces_1_3 ( // @[MockArray.scala 36:52]
    .clock(ces_1_3_clock),
    .io_ins_0(ces_1_3_io_ins_0),
    .io_ins_1(ces_1_3_io_ins_1),
    .io_ins_2(ces_1_3_io_ins_2),
    .io_ins_3(ces_1_3_io_ins_3),
    .io_outs_0(ces_1_3_io_outs_0),
    .io_outs_1(ces_1_3_io_outs_1),
    .io_outs_2(ces_1_3_io_outs_2),
    .io_outs_3(ces_1_3_io_outs_3)
  );
  Element ces_1_4 ( // @[MockArray.scala 36:52]
    .clock(ces_1_4_clock),
    .io_ins_0(ces_1_4_io_ins_0),
    .io_ins_1(ces_1_4_io_ins_1),
    .io_ins_2(ces_1_4_io_ins_2),
    .io_ins_3(ces_1_4_io_ins_3),
    .io_outs_0(ces_1_4_io_outs_0),
    .io_outs_1(ces_1_4_io_outs_1),
    .io_outs_2(ces_1_4_io_outs_2),
    .io_outs_3(ces_1_4_io_outs_3)
  );
  Element ces_1_5 ( // @[MockArray.scala 36:52]
    .clock(ces_1_5_clock),
    .io_ins_0(ces_1_5_io_ins_0),
    .io_ins_1(ces_1_5_io_ins_1),
    .io_ins_2(ces_1_5_io_ins_2),
    .io_ins_3(ces_1_5_io_ins_3),
    .io_outs_0(ces_1_5_io_outs_0),
    .io_outs_1(ces_1_5_io_outs_1),
    .io_outs_2(ces_1_5_io_outs_2),
    .io_outs_3(ces_1_5_io_outs_3)
  );
  Element ces_1_6 ( // @[MockArray.scala 36:52]
    .clock(ces_1_6_clock),
    .io_ins_0(ces_1_6_io_ins_0),
    .io_ins_1(ces_1_6_io_ins_1),
    .io_ins_2(ces_1_6_io_ins_2),
    .io_ins_3(ces_1_6_io_ins_3),
    .io_outs_0(ces_1_6_io_outs_0),
    .io_outs_1(ces_1_6_io_outs_1),
    .io_outs_2(ces_1_6_io_outs_2),
    .io_outs_3(ces_1_6_io_outs_3)
  );
  Element ces_1_7 ( // @[MockArray.scala 36:52]
    .clock(ces_1_7_clock),
    .io_ins_0(ces_1_7_io_ins_0),
    .io_ins_1(ces_1_7_io_ins_1),
    .io_ins_2(ces_1_7_io_ins_2),
    .io_ins_3(ces_1_7_io_ins_3),
    .io_outs_0(ces_1_7_io_outs_0),
    .io_outs_1(ces_1_7_io_outs_1),
    .io_outs_2(ces_1_7_io_outs_2),
    .io_outs_3(ces_1_7_io_outs_3)
  );
  Element ces_1_8 ( // @[MockArray.scala 36:52]
    .clock(ces_1_8_clock),
    .io_ins_0(ces_1_8_io_ins_0),
    .io_ins_1(ces_1_8_io_ins_1),
    .io_ins_2(ces_1_8_io_ins_2),
    .io_ins_3(ces_1_8_io_ins_3),
    .io_outs_0(ces_1_8_io_outs_0),
    .io_outs_1(ces_1_8_io_outs_1),
    .io_outs_2(ces_1_8_io_outs_2),
    .io_outs_3(ces_1_8_io_outs_3)
  );
  Element ces_1_9 ( // @[MockArray.scala 36:52]
    .clock(ces_1_9_clock),
    .io_ins_0(ces_1_9_io_ins_0),
    .io_ins_1(ces_1_9_io_ins_1),
    .io_ins_2(ces_1_9_io_ins_2),
    .io_ins_3(ces_1_9_io_ins_3),
    .io_outs_0(ces_1_9_io_outs_0),
    .io_outs_1(ces_1_9_io_outs_1),
    .io_outs_2(ces_1_9_io_outs_2),
    .io_outs_3(ces_1_9_io_outs_3)
  );
  Element ces_1_10 ( // @[MockArray.scala 36:52]
    .clock(ces_1_10_clock),
    .io_ins_0(ces_1_10_io_ins_0),
    .io_ins_1(ces_1_10_io_ins_1),
    .io_ins_2(ces_1_10_io_ins_2),
    .io_ins_3(ces_1_10_io_ins_3),
    .io_outs_0(ces_1_10_io_outs_0),
    .io_outs_1(ces_1_10_io_outs_1),
    .io_outs_2(ces_1_10_io_outs_2),
    .io_outs_3(ces_1_10_io_outs_3)
  );
  Element ces_1_11 ( // @[MockArray.scala 36:52]
    .clock(ces_1_11_clock),
    .io_ins_0(ces_1_11_io_ins_0),
    .io_ins_1(ces_1_11_io_ins_1),
    .io_ins_2(ces_1_11_io_ins_2),
    .io_ins_3(ces_1_11_io_ins_3),
    .io_outs_0(ces_1_11_io_outs_0),
    .io_outs_1(ces_1_11_io_outs_1),
    .io_outs_2(ces_1_11_io_outs_2),
    .io_outs_3(ces_1_11_io_outs_3)
  );
  Element ces_1_12 ( // @[MockArray.scala 36:52]
    .clock(ces_1_12_clock),
    .io_ins_0(ces_1_12_io_ins_0),
    .io_ins_1(ces_1_12_io_ins_1),
    .io_ins_2(ces_1_12_io_ins_2),
    .io_ins_3(ces_1_12_io_ins_3),
    .io_outs_0(ces_1_12_io_outs_0),
    .io_outs_1(ces_1_12_io_outs_1),
    .io_outs_2(ces_1_12_io_outs_2),
    .io_outs_3(ces_1_12_io_outs_3)
  );
  Element ces_1_13 ( // @[MockArray.scala 36:52]
    .clock(ces_1_13_clock),
    .io_ins_0(ces_1_13_io_ins_0),
    .io_ins_1(ces_1_13_io_ins_1),
    .io_ins_2(ces_1_13_io_ins_2),
    .io_ins_3(ces_1_13_io_ins_3),
    .io_outs_0(ces_1_13_io_outs_0),
    .io_outs_1(ces_1_13_io_outs_1),
    .io_outs_2(ces_1_13_io_outs_2),
    .io_outs_3(ces_1_13_io_outs_3)
  );
  Element ces_1_14 ( // @[MockArray.scala 36:52]
    .clock(ces_1_14_clock),
    .io_ins_0(ces_1_14_io_ins_0),
    .io_ins_1(ces_1_14_io_ins_1),
    .io_ins_2(ces_1_14_io_ins_2),
    .io_ins_3(ces_1_14_io_ins_3),
    .io_outs_0(ces_1_14_io_outs_0),
    .io_outs_1(ces_1_14_io_outs_1),
    .io_outs_2(ces_1_14_io_outs_2),
    .io_outs_3(ces_1_14_io_outs_3)
  );
  Element ces_1_15 ( // @[MockArray.scala 36:52]
    .clock(ces_1_15_clock),
    .io_ins_0(ces_1_15_io_ins_0),
    .io_ins_1(ces_1_15_io_ins_1),
    .io_ins_2(ces_1_15_io_ins_2),
    .io_ins_3(ces_1_15_io_ins_3),
    .io_outs_0(ces_1_15_io_outs_0),
    .io_outs_1(ces_1_15_io_outs_1),
    .io_outs_2(ces_1_15_io_outs_2),
    .io_outs_3(ces_1_15_io_outs_3)
  );
  Element ces_2_0 ( // @[MockArray.scala 36:52]
    .clock(ces_2_0_clock),
    .io_ins_0(ces_2_0_io_ins_0),
    .io_ins_1(ces_2_0_io_ins_1),
    .io_ins_2(ces_2_0_io_ins_2),
    .io_ins_3(ces_2_0_io_ins_3),
    .io_outs_0(ces_2_0_io_outs_0),
    .io_outs_1(ces_2_0_io_outs_1),
    .io_outs_2(ces_2_0_io_outs_2),
    .io_outs_3(ces_2_0_io_outs_3)
  );
  Element ces_2_1 ( // @[MockArray.scala 36:52]
    .clock(ces_2_1_clock),
    .io_ins_0(ces_2_1_io_ins_0),
    .io_ins_1(ces_2_1_io_ins_1),
    .io_ins_2(ces_2_1_io_ins_2),
    .io_ins_3(ces_2_1_io_ins_3),
    .io_outs_0(ces_2_1_io_outs_0),
    .io_outs_1(ces_2_1_io_outs_1),
    .io_outs_2(ces_2_1_io_outs_2),
    .io_outs_3(ces_2_1_io_outs_3)
  );
  Element ces_2_2 ( // @[MockArray.scala 36:52]
    .clock(ces_2_2_clock),
    .io_ins_0(ces_2_2_io_ins_0),
    .io_ins_1(ces_2_2_io_ins_1),
    .io_ins_2(ces_2_2_io_ins_2),
    .io_ins_3(ces_2_2_io_ins_3),
    .io_outs_0(ces_2_2_io_outs_0),
    .io_outs_1(ces_2_2_io_outs_1),
    .io_outs_2(ces_2_2_io_outs_2),
    .io_outs_3(ces_2_2_io_outs_3)
  );
  Element ces_2_3 ( // @[MockArray.scala 36:52]
    .clock(ces_2_3_clock),
    .io_ins_0(ces_2_3_io_ins_0),
    .io_ins_1(ces_2_3_io_ins_1),
    .io_ins_2(ces_2_3_io_ins_2),
    .io_ins_3(ces_2_3_io_ins_3),
    .io_outs_0(ces_2_3_io_outs_0),
    .io_outs_1(ces_2_3_io_outs_1),
    .io_outs_2(ces_2_3_io_outs_2),
    .io_outs_3(ces_2_3_io_outs_3)
  );
  Element ces_2_4 ( // @[MockArray.scala 36:52]
    .clock(ces_2_4_clock),
    .io_ins_0(ces_2_4_io_ins_0),
    .io_ins_1(ces_2_4_io_ins_1),
    .io_ins_2(ces_2_4_io_ins_2),
    .io_ins_3(ces_2_4_io_ins_3),
    .io_outs_0(ces_2_4_io_outs_0),
    .io_outs_1(ces_2_4_io_outs_1),
    .io_outs_2(ces_2_4_io_outs_2),
    .io_outs_3(ces_2_4_io_outs_3)
  );
  Element ces_2_5 ( // @[MockArray.scala 36:52]
    .clock(ces_2_5_clock),
    .io_ins_0(ces_2_5_io_ins_0),
    .io_ins_1(ces_2_5_io_ins_1),
    .io_ins_2(ces_2_5_io_ins_2),
    .io_ins_3(ces_2_5_io_ins_3),
    .io_outs_0(ces_2_5_io_outs_0),
    .io_outs_1(ces_2_5_io_outs_1),
    .io_outs_2(ces_2_5_io_outs_2),
    .io_outs_3(ces_2_5_io_outs_3)
  );
  Element ces_2_6 ( // @[MockArray.scala 36:52]
    .clock(ces_2_6_clock),
    .io_ins_0(ces_2_6_io_ins_0),
    .io_ins_1(ces_2_6_io_ins_1),
    .io_ins_2(ces_2_6_io_ins_2),
    .io_ins_3(ces_2_6_io_ins_3),
    .io_outs_0(ces_2_6_io_outs_0),
    .io_outs_1(ces_2_6_io_outs_1),
    .io_outs_2(ces_2_6_io_outs_2),
    .io_outs_3(ces_2_6_io_outs_3)
  );
  Element ces_2_7 ( // @[MockArray.scala 36:52]
    .clock(ces_2_7_clock),
    .io_ins_0(ces_2_7_io_ins_0),
    .io_ins_1(ces_2_7_io_ins_1),
    .io_ins_2(ces_2_7_io_ins_2),
    .io_ins_3(ces_2_7_io_ins_3),
    .io_outs_0(ces_2_7_io_outs_0),
    .io_outs_1(ces_2_7_io_outs_1),
    .io_outs_2(ces_2_7_io_outs_2),
    .io_outs_3(ces_2_7_io_outs_3)
  );
  Element ces_2_8 ( // @[MockArray.scala 36:52]
    .clock(ces_2_8_clock),
    .io_ins_0(ces_2_8_io_ins_0),
    .io_ins_1(ces_2_8_io_ins_1),
    .io_ins_2(ces_2_8_io_ins_2),
    .io_ins_3(ces_2_8_io_ins_3),
    .io_outs_0(ces_2_8_io_outs_0),
    .io_outs_1(ces_2_8_io_outs_1),
    .io_outs_2(ces_2_8_io_outs_2),
    .io_outs_3(ces_2_8_io_outs_3)
  );
  Element ces_2_9 ( // @[MockArray.scala 36:52]
    .clock(ces_2_9_clock),
    .io_ins_0(ces_2_9_io_ins_0),
    .io_ins_1(ces_2_9_io_ins_1),
    .io_ins_2(ces_2_9_io_ins_2),
    .io_ins_3(ces_2_9_io_ins_3),
    .io_outs_0(ces_2_9_io_outs_0),
    .io_outs_1(ces_2_9_io_outs_1),
    .io_outs_2(ces_2_9_io_outs_2),
    .io_outs_3(ces_2_9_io_outs_3)
  );
  Element ces_2_10 ( // @[MockArray.scala 36:52]
    .clock(ces_2_10_clock),
    .io_ins_0(ces_2_10_io_ins_0),
    .io_ins_1(ces_2_10_io_ins_1),
    .io_ins_2(ces_2_10_io_ins_2),
    .io_ins_3(ces_2_10_io_ins_3),
    .io_outs_0(ces_2_10_io_outs_0),
    .io_outs_1(ces_2_10_io_outs_1),
    .io_outs_2(ces_2_10_io_outs_2),
    .io_outs_3(ces_2_10_io_outs_3)
  );
  Element ces_2_11 ( // @[MockArray.scala 36:52]
    .clock(ces_2_11_clock),
    .io_ins_0(ces_2_11_io_ins_0),
    .io_ins_1(ces_2_11_io_ins_1),
    .io_ins_2(ces_2_11_io_ins_2),
    .io_ins_3(ces_2_11_io_ins_3),
    .io_outs_0(ces_2_11_io_outs_0),
    .io_outs_1(ces_2_11_io_outs_1),
    .io_outs_2(ces_2_11_io_outs_2),
    .io_outs_3(ces_2_11_io_outs_3)
  );
  Element ces_2_12 ( // @[MockArray.scala 36:52]
    .clock(ces_2_12_clock),
    .io_ins_0(ces_2_12_io_ins_0),
    .io_ins_1(ces_2_12_io_ins_1),
    .io_ins_2(ces_2_12_io_ins_2),
    .io_ins_3(ces_2_12_io_ins_3),
    .io_outs_0(ces_2_12_io_outs_0),
    .io_outs_1(ces_2_12_io_outs_1),
    .io_outs_2(ces_2_12_io_outs_2),
    .io_outs_3(ces_2_12_io_outs_3)
  );
  Element ces_2_13 ( // @[MockArray.scala 36:52]
    .clock(ces_2_13_clock),
    .io_ins_0(ces_2_13_io_ins_0),
    .io_ins_1(ces_2_13_io_ins_1),
    .io_ins_2(ces_2_13_io_ins_2),
    .io_ins_3(ces_2_13_io_ins_3),
    .io_outs_0(ces_2_13_io_outs_0),
    .io_outs_1(ces_2_13_io_outs_1),
    .io_outs_2(ces_2_13_io_outs_2),
    .io_outs_3(ces_2_13_io_outs_3)
  );
  Element ces_2_14 ( // @[MockArray.scala 36:52]
    .clock(ces_2_14_clock),
    .io_ins_0(ces_2_14_io_ins_0),
    .io_ins_1(ces_2_14_io_ins_1),
    .io_ins_2(ces_2_14_io_ins_2),
    .io_ins_3(ces_2_14_io_ins_3),
    .io_outs_0(ces_2_14_io_outs_0),
    .io_outs_1(ces_2_14_io_outs_1),
    .io_outs_2(ces_2_14_io_outs_2),
    .io_outs_3(ces_2_14_io_outs_3)
  );
  Element ces_2_15 ( // @[MockArray.scala 36:52]
    .clock(ces_2_15_clock),
    .io_ins_0(ces_2_15_io_ins_0),
    .io_ins_1(ces_2_15_io_ins_1),
    .io_ins_2(ces_2_15_io_ins_2),
    .io_ins_3(ces_2_15_io_ins_3),
    .io_outs_0(ces_2_15_io_outs_0),
    .io_outs_1(ces_2_15_io_outs_1),
    .io_outs_2(ces_2_15_io_outs_2),
    .io_outs_3(ces_2_15_io_outs_3)
  );
  Element ces_3_0 ( // @[MockArray.scala 36:52]
    .clock(ces_3_0_clock),
    .io_ins_0(ces_3_0_io_ins_0),
    .io_ins_1(ces_3_0_io_ins_1),
    .io_ins_2(ces_3_0_io_ins_2),
    .io_ins_3(ces_3_0_io_ins_3),
    .io_outs_0(ces_3_0_io_outs_0),
    .io_outs_1(ces_3_0_io_outs_1),
    .io_outs_2(ces_3_0_io_outs_2),
    .io_outs_3(ces_3_0_io_outs_3)
  );
  Element ces_3_1 ( // @[MockArray.scala 36:52]
    .clock(ces_3_1_clock),
    .io_ins_0(ces_3_1_io_ins_0),
    .io_ins_1(ces_3_1_io_ins_1),
    .io_ins_2(ces_3_1_io_ins_2),
    .io_ins_3(ces_3_1_io_ins_3),
    .io_outs_0(ces_3_1_io_outs_0),
    .io_outs_1(ces_3_1_io_outs_1),
    .io_outs_2(ces_3_1_io_outs_2),
    .io_outs_3(ces_3_1_io_outs_3)
  );
  Element ces_3_2 ( // @[MockArray.scala 36:52]
    .clock(ces_3_2_clock),
    .io_ins_0(ces_3_2_io_ins_0),
    .io_ins_1(ces_3_2_io_ins_1),
    .io_ins_2(ces_3_2_io_ins_2),
    .io_ins_3(ces_3_2_io_ins_3),
    .io_outs_0(ces_3_2_io_outs_0),
    .io_outs_1(ces_3_2_io_outs_1),
    .io_outs_2(ces_3_2_io_outs_2),
    .io_outs_3(ces_3_2_io_outs_3)
  );
  Element ces_3_3 ( // @[MockArray.scala 36:52]
    .clock(ces_3_3_clock),
    .io_ins_0(ces_3_3_io_ins_0),
    .io_ins_1(ces_3_3_io_ins_1),
    .io_ins_2(ces_3_3_io_ins_2),
    .io_ins_3(ces_3_3_io_ins_3),
    .io_outs_0(ces_3_3_io_outs_0),
    .io_outs_1(ces_3_3_io_outs_1),
    .io_outs_2(ces_3_3_io_outs_2),
    .io_outs_3(ces_3_3_io_outs_3)
  );
  Element ces_3_4 ( // @[MockArray.scala 36:52]
    .clock(ces_3_4_clock),
    .io_ins_0(ces_3_4_io_ins_0),
    .io_ins_1(ces_3_4_io_ins_1),
    .io_ins_2(ces_3_4_io_ins_2),
    .io_ins_3(ces_3_4_io_ins_3),
    .io_outs_0(ces_3_4_io_outs_0),
    .io_outs_1(ces_3_4_io_outs_1),
    .io_outs_2(ces_3_4_io_outs_2),
    .io_outs_3(ces_3_4_io_outs_3)
  );
  Element ces_3_5 ( // @[MockArray.scala 36:52]
    .clock(ces_3_5_clock),
    .io_ins_0(ces_3_5_io_ins_0),
    .io_ins_1(ces_3_5_io_ins_1),
    .io_ins_2(ces_3_5_io_ins_2),
    .io_ins_3(ces_3_5_io_ins_3),
    .io_outs_0(ces_3_5_io_outs_0),
    .io_outs_1(ces_3_5_io_outs_1),
    .io_outs_2(ces_3_5_io_outs_2),
    .io_outs_3(ces_3_5_io_outs_3)
  );
  Element ces_3_6 ( // @[MockArray.scala 36:52]
    .clock(ces_3_6_clock),
    .io_ins_0(ces_3_6_io_ins_0),
    .io_ins_1(ces_3_6_io_ins_1),
    .io_ins_2(ces_3_6_io_ins_2),
    .io_ins_3(ces_3_6_io_ins_3),
    .io_outs_0(ces_3_6_io_outs_0),
    .io_outs_1(ces_3_6_io_outs_1),
    .io_outs_2(ces_3_6_io_outs_2),
    .io_outs_3(ces_3_6_io_outs_3)
  );
  Element ces_3_7 ( // @[MockArray.scala 36:52]
    .clock(ces_3_7_clock),
    .io_ins_0(ces_3_7_io_ins_0),
    .io_ins_1(ces_3_7_io_ins_1),
    .io_ins_2(ces_3_7_io_ins_2),
    .io_ins_3(ces_3_7_io_ins_3),
    .io_outs_0(ces_3_7_io_outs_0),
    .io_outs_1(ces_3_7_io_outs_1),
    .io_outs_2(ces_3_7_io_outs_2),
    .io_outs_3(ces_3_7_io_outs_3)
  );
  Element ces_3_8 ( // @[MockArray.scala 36:52]
    .clock(ces_3_8_clock),
    .io_ins_0(ces_3_8_io_ins_0),
    .io_ins_1(ces_3_8_io_ins_1),
    .io_ins_2(ces_3_8_io_ins_2),
    .io_ins_3(ces_3_8_io_ins_3),
    .io_outs_0(ces_3_8_io_outs_0),
    .io_outs_1(ces_3_8_io_outs_1),
    .io_outs_2(ces_3_8_io_outs_2),
    .io_outs_3(ces_3_8_io_outs_3)
  );
  Element ces_3_9 ( // @[MockArray.scala 36:52]
    .clock(ces_3_9_clock),
    .io_ins_0(ces_3_9_io_ins_0),
    .io_ins_1(ces_3_9_io_ins_1),
    .io_ins_2(ces_3_9_io_ins_2),
    .io_ins_3(ces_3_9_io_ins_3),
    .io_outs_0(ces_3_9_io_outs_0),
    .io_outs_1(ces_3_9_io_outs_1),
    .io_outs_2(ces_3_9_io_outs_2),
    .io_outs_3(ces_3_9_io_outs_3)
  );
  Element ces_3_10 ( // @[MockArray.scala 36:52]
    .clock(ces_3_10_clock),
    .io_ins_0(ces_3_10_io_ins_0),
    .io_ins_1(ces_3_10_io_ins_1),
    .io_ins_2(ces_3_10_io_ins_2),
    .io_ins_3(ces_3_10_io_ins_3),
    .io_outs_0(ces_3_10_io_outs_0),
    .io_outs_1(ces_3_10_io_outs_1),
    .io_outs_2(ces_3_10_io_outs_2),
    .io_outs_3(ces_3_10_io_outs_3)
  );
  Element ces_3_11 ( // @[MockArray.scala 36:52]
    .clock(ces_3_11_clock),
    .io_ins_0(ces_3_11_io_ins_0),
    .io_ins_1(ces_3_11_io_ins_1),
    .io_ins_2(ces_3_11_io_ins_2),
    .io_ins_3(ces_3_11_io_ins_3),
    .io_outs_0(ces_3_11_io_outs_0),
    .io_outs_1(ces_3_11_io_outs_1),
    .io_outs_2(ces_3_11_io_outs_2),
    .io_outs_3(ces_3_11_io_outs_3)
  );
  Element ces_3_12 ( // @[MockArray.scala 36:52]
    .clock(ces_3_12_clock),
    .io_ins_0(ces_3_12_io_ins_0),
    .io_ins_1(ces_3_12_io_ins_1),
    .io_ins_2(ces_3_12_io_ins_2),
    .io_ins_3(ces_3_12_io_ins_3),
    .io_outs_0(ces_3_12_io_outs_0),
    .io_outs_1(ces_3_12_io_outs_1),
    .io_outs_2(ces_3_12_io_outs_2),
    .io_outs_3(ces_3_12_io_outs_3)
  );
  Element ces_3_13 ( // @[MockArray.scala 36:52]
    .clock(ces_3_13_clock),
    .io_ins_0(ces_3_13_io_ins_0),
    .io_ins_1(ces_3_13_io_ins_1),
    .io_ins_2(ces_3_13_io_ins_2),
    .io_ins_3(ces_3_13_io_ins_3),
    .io_outs_0(ces_3_13_io_outs_0),
    .io_outs_1(ces_3_13_io_outs_1),
    .io_outs_2(ces_3_13_io_outs_2),
    .io_outs_3(ces_3_13_io_outs_3)
  );
  Element ces_3_14 ( // @[MockArray.scala 36:52]
    .clock(ces_3_14_clock),
    .io_ins_0(ces_3_14_io_ins_0),
    .io_ins_1(ces_3_14_io_ins_1),
    .io_ins_2(ces_3_14_io_ins_2),
    .io_ins_3(ces_3_14_io_ins_3),
    .io_outs_0(ces_3_14_io_outs_0),
    .io_outs_1(ces_3_14_io_outs_1),
    .io_outs_2(ces_3_14_io_outs_2),
    .io_outs_3(ces_3_14_io_outs_3)
  );
  Element ces_3_15 ( // @[MockArray.scala 36:52]
    .clock(ces_3_15_clock),
    .io_ins_0(ces_3_15_io_ins_0),
    .io_ins_1(ces_3_15_io_ins_1),
    .io_ins_2(ces_3_15_io_ins_2),
    .io_ins_3(ces_3_15_io_ins_3),
    .io_outs_0(ces_3_15_io_outs_0),
    .io_outs_1(ces_3_15_io_outs_1),
    .io_outs_2(ces_3_15_io_outs_2),
    .io_outs_3(ces_3_15_io_outs_3)
  );
  Element ces_4_0 ( // @[MockArray.scala 36:52]
    .clock(ces_4_0_clock),
    .io_ins_0(ces_4_0_io_ins_0),
    .io_ins_1(ces_4_0_io_ins_1),
    .io_ins_2(ces_4_0_io_ins_2),
    .io_ins_3(ces_4_0_io_ins_3),
    .io_outs_0(ces_4_0_io_outs_0),
    .io_outs_1(ces_4_0_io_outs_1),
    .io_outs_2(ces_4_0_io_outs_2),
    .io_outs_3(ces_4_0_io_outs_3)
  );
  Element ces_4_1 ( // @[MockArray.scala 36:52]
    .clock(ces_4_1_clock),
    .io_ins_0(ces_4_1_io_ins_0),
    .io_ins_1(ces_4_1_io_ins_1),
    .io_ins_2(ces_4_1_io_ins_2),
    .io_ins_3(ces_4_1_io_ins_3),
    .io_outs_0(ces_4_1_io_outs_0),
    .io_outs_1(ces_4_1_io_outs_1),
    .io_outs_2(ces_4_1_io_outs_2),
    .io_outs_3(ces_4_1_io_outs_3)
  );
  Element ces_4_2 ( // @[MockArray.scala 36:52]
    .clock(ces_4_2_clock),
    .io_ins_0(ces_4_2_io_ins_0),
    .io_ins_1(ces_4_2_io_ins_1),
    .io_ins_2(ces_4_2_io_ins_2),
    .io_ins_3(ces_4_2_io_ins_3),
    .io_outs_0(ces_4_2_io_outs_0),
    .io_outs_1(ces_4_2_io_outs_1),
    .io_outs_2(ces_4_2_io_outs_2),
    .io_outs_3(ces_4_2_io_outs_3)
  );
  Element ces_4_3 ( // @[MockArray.scala 36:52]
    .clock(ces_4_3_clock),
    .io_ins_0(ces_4_3_io_ins_0),
    .io_ins_1(ces_4_3_io_ins_1),
    .io_ins_2(ces_4_3_io_ins_2),
    .io_ins_3(ces_4_3_io_ins_3),
    .io_outs_0(ces_4_3_io_outs_0),
    .io_outs_1(ces_4_3_io_outs_1),
    .io_outs_2(ces_4_3_io_outs_2),
    .io_outs_3(ces_4_3_io_outs_3)
  );
  Element ces_4_4 ( // @[MockArray.scala 36:52]
    .clock(ces_4_4_clock),
    .io_ins_0(ces_4_4_io_ins_0),
    .io_ins_1(ces_4_4_io_ins_1),
    .io_ins_2(ces_4_4_io_ins_2),
    .io_ins_3(ces_4_4_io_ins_3),
    .io_outs_0(ces_4_4_io_outs_0),
    .io_outs_1(ces_4_4_io_outs_1),
    .io_outs_2(ces_4_4_io_outs_2),
    .io_outs_3(ces_4_4_io_outs_3)
  );
  Element ces_4_5 ( // @[MockArray.scala 36:52]
    .clock(ces_4_5_clock),
    .io_ins_0(ces_4_5_io_ins_0),
    .io_ins_1(ces_4_5_io_ins_1),
    .io_ins_2(ces_4_5_io_ins_2),
    .io_ins_3(ces_4_5_io_ins_3),
    .io_outs_0(ces_4_5_io_outs_0),
    .io_outs_1(ces_4_5_io_outs_1),
    .io_outs_2(ces_4_5_io_outs_2),
    .io_outs_3(ces_4_5_io_outs_3)
  );
  Element ces_4_6 ( // @[MockArray.scala 36:52]
    .clock(ces_4_6_clock),
    .io_ins_0(ces_4_6_io_ins_0),
    .io_ins_1(ces_4_6_io_ins_1),
    .io_ins_2(ces_4_6_io_ins_2),
    .io_ins_3(ces_4_6_io_ins_3),
    .io_outs_0(ces_4_6_io_outs_0),
    .io_outs_1(ces_4_6_io_outs_1),
    .io_outs_2(ces_4_6_io_outs_2),
    .io_outs_3(ces_4_6_io_outs_3)
  );
  Element ces_4_7 ( // @[MockArray.scala 36:52]
    .clock(ces_4_7_clock),
    .io_ins_0(ces_4_7_io_ins_0),
    .io_ins_1(ces_4_7_io_ins_1),
    .io_ins_2(ces_4_7_io_ins_2),
    .io_ins_3(ces_4_7_io_ins_3),
    .io_outs_0(ces_4_7_io_outs_0),
    .io_outs_1(ces_4_7_io_outs_1),
    .io_outs_2(ces_4_7_io_outs_2),
    .io_outs_3(ces_4_7_io_outs_3)
  );
  Element ces_4_8 ( // @[MockArray.scala 36:52]
    .clock(ces_4_8_clock),
    .io_ins_0(ces_4_8_io_ins_0),
    .io_ins_1(ces_4_8_io_ins_1),
    .io_ins_2(ces_4_8_io_ins_2),
    .io_ins_3(ces_4_8_io_ins_3),
    .io_outs_0(ces_4_8_io_outs_0),
    .io_outs_1(ces_4_8_io_outs_1),
    .io_outs_2(ces_4_8_io_outs_2),
    .io_outs_3(ces_4_8_io_outs_3)
  );
  Element ces_4_9 ( // @[MockArray.scala 36:52]
    .clock(ces_4_9_clock),
    .io_ins_0(ces_4_9_io_ins_0),
    .io_ins_1(ces_4_9_io_ins_1),
    .io_ins_2(ces_4_9_io_ins_2),
    .io_ins_3(ces_4_9_io_ins_3),
    .io_outs_0(ces_4_9_io_outs_0),
    .io_outs_1(ces_4_9_io_outs_1),
    .io_outs_2(ces_4_9_io_outs_2),
    .io_outs_3(ces_4_9_io_outs_3)
  );
  Element ces_4_10 ( // @[MockArray.scala 36:52]
    .clock(ces_4_10_clock),
    .io_ins_0(ces_4_10_io_ins_0),
    .io_ins_1(ces_4_10_io_ins_1),
    .io_ins_2(ces_4_10_io_ins_2),
    .io_ins_3(ces_4_10_io_ins_3),
    .io_outs_0(ces_4_10_io_outs_0),
    .io_outs_1(ces_4_10_io_outs_1),
    .io_outs_2(ces_4_10_io_outs_2),
    .io_outs_3(ces_4_10_io_outs_3)
  );
  Element ces_4_11 ( // @[MockArray.scala 36:52]
    .clock(ces_4_11_clock),
    .io_ins_0(ces_4_11_io_ins_0),
    .io_ins_1(ces_4_11_io_ins_1),
    .io_ins_2(ces_4_11_io_ins_2),
    .io_ins_3(ces_4_11_io_ins_3),
    .io_outs_0(ces_4_11_io_outs_0),
    .io_outs_1(ces_4_11_io_outs_1),
    .io_outs_2(ces_4_11_io_outs_2),
    .io_outs_3(ces_4_11_io_outs_3)
  );
  Element ces_4_12 ( // @[MockArray.scala 36:52]
    .clock(ces_4_12_clock),
    .io_ins_0(ces_4_12_io_ins_0),
    .io_ins_1(ces_4_12_io_ins_1),
    .io_ins_2(ces_4_12_io_ins_2),
    .io_ins_3(ces_4_12_io_ins_3),
    .io_outs_0(ces_4_12_io_outs_0),
    .io_outs_1(ces_4_12_io_outs_1),
    .io_outs_2(ces_4_12_io_outs_2),
    .io_outs_3(ces_4_12_io_outs_3)
  );
  Element ces_4_13 ( // @[MockArray.scala 36:52]
    .clock(ces_4_13_clock),
    .io_ins_0(ces_4_13_io_ins_0),
    .io_ins_1(ces_4_13_io_ins_1),
    .io_ins_2(ces_4_13_io_ins_2),
    .io_ins_3(ces_4_13_io_ins_3),
    .io_outs_0(ces_4_13_io_outs_0),
    .io_outs_1(ces_4_13_io_outs_1),
    .io_outs_2(ces_4_13_io_outs_2),
    .io_outs_3(ces_4_13_io_outs_3)
  );
  Element ces_4_14 ( // @[MockArray.scala 36:52]
    .clock(ces_4_14_clock),
    .io_ins_0(ces_4_14_io_ins_0),
    .io_ins_1(ces_4_14_io_ins_1),
    .io_ins_2(ces_4_14_io_ins_2),
    .io_ins_3(ces_4_14_io_ins_3),
    .io_outs_0(ces_4_14_io_outs_0),
    .io_outs_1(ces_4_14_io_outs_1),
    .io_outs_2(ces_4_14_io_outs_2),
    .io_outs_3(ces_4_14_io_outs_3)
  );
  Element ces_4_15 ( // @[MockArray.scala 36:52]
    .clock(ces_4_15_clock),
    .io_ins_0(ces_4_15_io_ins_0),
    .io_ins_1(ces_4_15_io_ins_1),
    .io_ins_2(ces_4_15_io_ins_2),
    .io_ins_3(ces_4_15_io_ins_3),
    .io_outs_0(ces_4_15_io_outs_0),
    .io_outs_1(ces_4_15_io_outs_1),
    .io_outs_2(ces_4_15_io_outs_2),
    .io_outs_3(ces_4_15_io_outs_3)
  );
  Element ces_5_0 ( // @[MockArray.scala 36:52]
    .clock(ces_5_0_clock),
    .io_ins_0(ces_5_0_io_ins_0),
    .io_ins_1(ces_5_0_io_ins_1),
    .io_ins_2(ces_5_0_io_ins_2),
    .io_ins_3(ces_5_0_io_ins_3),
    .io_outs_0(ces_5_0_io_outs_0),
    .io_outs_1(ces_5_0_io_outs_1),
    .io_outs_2(ces_5_0_io_outs_2),
    .io_outs_3(ces_5_0_io_outs_3)
  );
  Element ces_5_1 ( // @[MockArray.scala 36:52]
    .clock(ces_5_1_clock),
    .io_ins_0(ces_5_1_io_ins_0),
    .io_ins_1(ces_5_1_io_ins_1),
    .io_ins_2(ces_5_1_io_ins_2),
    .io_ins_3(ces_5_1_io_ins_3),
    .io_outs_0(ces_5_1_io_outs_0),
    .io_outs_1(ces_5_1_io_outs_1),
    .io_outs_2(ces_5_1_io_outs_2),
    .io_outs_3(ces_5_1_io_outs_3)
  );
  Element ces_5_2 ( // @[MockArray.scala 36:52]
    .clock(ces_5_2_clock),
    .io_ins_0(ces_5_2_io_ins_0),
    .io_ins_1(ces_5_2_io_ins_1),
    .io_ins_2(ces_5_2_io_ins_2),
    .io_ins_3(ces_5_2_io_ins_3),
    .io_outs_0(ces_5_2_io_outs_0),
    .io_outs_1(ces_5_2_io_outs_1),
    .io_outs_2(ces_5_2_io_outs_2),
    .io_outs_3(ces_5_2_io_outs_3)
  );
  Element ces_5_3 ( // @[MockArray.scala 36:52]
    .clock(ces_5_3_clock),
    .io_ins_0(ces_5_3_io_ins_0),
    .io_ins_1(ces_5_3_io_ins_1),
    .io_ins_2(ces_5_3_io_ins_2),
    .io_ins_3(ces_5_3_io_ins_3),
    .io_outs_0(ces_5_3_io_outs_0),
    .io_outs_1(ces_5_3_io_outs_1),
    .io_outs_2(ces_5_3_io_outs_2),
    .io_outs_3(ces_5_3_io_outs_3)
  );
  Element ces_5_4 ( // @[MockArray.scala 36:52]
    .clock(ces_5_4_clock),
    .io_ins_0(ces_5_4_io_ins_0),
    .io_ins_1(ces_5_4_io_ins_1),
    .io_ins_2(ces_5_4_io_ins_2),
    .io_ins_3(ces_5_4_io_ins_3),
    .io_outs_0(ces_5_4_io_outs_0),
    .io_outs_1(ces_5_4_io_outs_1),
    .io_outs_2(ces_5_4_io_outs_2),
    .io_outs_3(ces_5_4_io_outs_3)
  );
  Element ces_5_5 ( // @[MockArray.scala 36:52]
    .clock(ces_5_5_clock),
    .io_ins_0(ces_5_5_io_ins_0),
    .io_ins_1(ces_5_5_io_ins_1),
    .io_ins_2(ces_5_5_io_ins_2),
    .io_ins_3(ces_5_5_io_ins_3),
    .io_outs_0(ces_5_5_io_outs_0),
    .io_outs_1(ces_5_5_io_outs_1),
    .io_outs_2(ces_5_5_io_outs_2),
    .io_outs_3(ces_5_5_io_outs_3)
  );
  Element ces_5_6 ( // @[MockArray.scala 36:52]
    .clock(ces_5_6_clock),
    .io_ins_0(ces_5_6_io_ins_0),
    .io_ins_1(ces_5_6_io_ins_1),
    .io_ins_2(ces_5_6_io_ins_2),
    .io_ins_3(ces_5_6_io_ins_3),
    .io_outs_0(ces_5_6_io_outs_0),
    .io_outs_1(ces_5_6_io_outs_1),
    .io_outs_2(ces_5_6_io_outs_2),
    .io_outs_3(ces_5_6_io_outs_3)
  );
  Element ces_5_7 ( // @[MockArray.scala 36:52]
    .clock(ces_5_7_clock),
    .io_ins_0(ces_5_7_io_ins_0),
    .io_ins_1(ces_5_7_io_ins_1),
    .io_ins_2(ces_5_7_io_ins_2),
    .io_ins_3(ces_5_7_io_ins_3),
    .io_outs_0(ces_5_7_io_outs_0),
    .io_outs_1(ces_5_7_io_outs_1),
    .io_outs_2(ces_5_7_io_outs_2),
    .io_outs_3(ces_5_7_io_outs_3)
  );
  Element ces_5_8 ( // @[MockArray.scala 36:52]
    .clock(ces_5_8_clock),
    .io_ins_0(ces_5_8_io_ins_0),
    .io_ins_1(ces_5_8_io_ins_1),
    .io_ins_2(ces_5_8_io_ins_2),
    .io_ins_3(ces_5_8_io_ins_3),
    .io_outs_0(ces_5_8_io_outs_0),
    .io_outs_1(ces_5_8_io_outs_1),
    .io_outs_2(ces_5_8_io_outs_2),
    .io_outs_3(ces_5_8_io_outs_3)
  );
  Element ces_5_9 ( // @[MockArray.scala 36:52]
    .clock(ces_5_9_clock),
    .io_ins_0(ces_5_9_io_ins_0),
    .io_ins_1(ces_5_9_io_ins_1),
    .io_ins_2(ces_5_9_io_ins_2),
    .io_ins_3(ces_5_9_io_ins_3),
    .io_outs_0(ces_5_9_io_outs_0),
    .io_outs_1(ces_5_9_io_outs_1),
    .io_outs_2(ces_5_9_io_outs_2),
    .io_outs_3(ces_5_9_io_outs_3)
  );
  Element ces_5_10 ( // @[MockArray.scala 36:52]
    .clock(ces_5_10_clock),
    .io_ins_0(ces_5_10_io_ins_0),
    .io_ins_1(ces_5_10_io_ins_1),
    .io_ins_2(ces_5_10_io_ins_2),
    .io_ins_3(ces_5_10_io_ins_3),
    .io_outs_0(ces_5_10_io_outs_0),
    .io_outs_1(ces_5_10_io_outs_1),
    .io_outs_2(ces_5_10_io_outs_2),
    .io_outs_3(ces_5_10_io_outs_3)
  );
  Element ces_5_11 ( // @[MockArray.scala 36:52]
    .clock(ces_5_11_clock),
    .io_ins_0(ces_5_11_io_ins_0),
    .io_ins_1(ces_5_11_io_ins_1),
    .io_ins_2(ces_5_11_io_ins_2),
    .io_ins_3(ces_5_11_io_ins_3),
    .io_outs_0(ces_5_11_io_outs_0),
    .io_outs_1(ces_5_11_io_outs_1),
    .io_outs_2(ces_5_11_io_outs_2),
    .io_outs_3(ces_5_11_io_outs_3)
  );
  Element ces_5_12 ( // @[MockArray.scala 36:52]
    .clock(ces_5_12_clock),
    .io_ins_0(ces_5_12_io_ins_0),
    .io_ins_1(ces_5_12_io_ins_1),
    .io_ins_2(ces_5_12_io_ins_2),
    .io_ins_3(ces_5_12_io_ins_3),
    .io_outs_0(ces_5_12_io_outs_0),
    .io_outs_1(ces_5_12_io_outs_1),
    .io_outs_2(ces_5_12_io_outs_2),
    .io_outs_3(ces_5_12_io_outs_3)
  );
  Element ces_5_13 ( // @[MockArray.scala 36:52]
    .clock(ces_5_13_clock),
    .io_ins_0(ces_5_13_io_ins_0),
    .io_ins_1(ces_5_13_io_ins_1),
    .io_ins_2(ces_5_13_io_ins_2),
    .io_ins_3(ces_5_13_io_ins_3),
    .io_outs_0(ces_5_13_io_outs_0),
    .io_outs_1(ces_5_13_io_outs_1),
    .io_outs_2(ces_5_13_io_outs_2),
    .io_outs_3(ces_5_13_io_outs_3)
  );
  Element ces_5_14 ( // @[MockArray.scala 36:52]
    .clock(ces_5_14_clock),
    .io_ins_0(ces_5_14_io_ins_0),
    .io_ins_1(ces_5_14_io_ins_1),
    .io_ins_2(ces_5_14_io_ins_2),
    .io_ins_3(ces_5_14_io_ins_3),
    .io_outs_0(ces_5_14_io_outs_0),
    .io_outs_1(ces_5_14_io_outs_1),
    .io_outs_2(ces_5_14_io_outs_2),
    .io_outs_3(ces_5_14_io_outs_3)
  );
  Element ces_5_15 ( // @[MockArray.scala 36:52]
    .clock(ces_5_15_clock),
    .io_ins_0(ces_5_15_io_ins_0),
    .io_ins_1(ces_5_15_io_ins_1),
    .io_ins_2(ces_5_15_io_ins_2),
    .io_ins_3(ces_5_15_io_ins_3),
    .io_outs_0(ces_5_15_io_outs_0),
    .io_outs_1(ces_5_15_io_outs_1),
    .io_outs_2(ces_5_15_io_outs_2),
    .io_outs_3(ces_5_15_io_outs_3)
  );
  Element ces_6_0 ( // @[MockArray.scala 36:52]
    .clock(ces_6_0_clock),
    .io_ins_0(ces_6_0_io_ins_0),
    .io_ins_1(ces_6_0_io_ins_1),
    .io_ins_2(ces_6_0_io_ins_2),
    .io_ins_3(ces_6_0_io_ins_3),
    .io_outs_0(ces_6_0_io_outs_0),
    .io_outs_1(ces_6_0_io_outs_1),
    .io_outs_2(ces_6_0_io_outs_2),
    .io_outs_3(ces_6_0_io_outs_3)
  );
  Element ces_6_1 ( // @[MockArray.scala 36:52]
    .clock(ces_6_1_clock),
    .io_ins_0(ces_6_1_io_ins_0),
    .io_ins_1(ces_6_1_io_ins_1),
    .io_ins_2(ces_6_1_io_ins_2),
    .io_ins_3(ces_6_1_io_ins_3),
    .io_outs_0(ces_6_1_io_outs_0),
    .io_outs_1(ces_6_1_io_outs_1),
    .io_outs_2(ces_6_1_io_outs_2),
    .io_outs_3(ces_6_1_io_outs_3)
  );
  Element ces_6_2 ( // @[MockArray.scala 36:52]
    .clock(ces_6_2_clock),
    .io_ins_0(ces_6_2_io_ins_0),
    .io_ins_1(ces_6_2_io_ins_1),
    .io_ins_2(ces_6_2_io_ins_2),
    .io_ins_3(ces_6_2_io_ins_3),
    .io_outs_0(ces_6_2_io_outs_0),
    .io_outs_1(ces_6_2_io_outs_1),
    .io_outs_2(ces_6_2_io_outs_2),
    .io_outs_3(ces_6_2_io_outs_3)
  );
  Element ces_6_3 ( // @[MockArray.scala 36:52]
    .clock(ces_6_3_clock),
    .io_ins_0(ces_6_3_io_ins_0),
    .io_ins_1(ces_6_3_io_ins_1),
    .io_ins_2(ces_6_3_io_ins_2),
    .io_ins_3(ces_6_3_io_ins_3),
    .io_outs_0(ces_6_3_io_outs_0),
    .io_outs_1(ces_6_3_io_outs_1),
    .io_outs_2(ces_6_3_io_outs_2),
    .io_outs_3(ces_6_3_io_outs_3)
  );
  Element ces_6_4 ( // @[MockArray.scala 36:52]
    .clock(ces_6_4_clock),
    .io_ins_0(ces_6_4_io_ins_0),
    .io_ins_1(ces_6_4_io_ins_1),
    .io_ins_2(ces_6_4_io_ins_2),
    .io_ins_3(ces_6_4_io_ins_3),
    .io_outs_0(ces_6_4_io_outs_0),
    .io_outs_1(ces_6_4_io_outs_1),
    .io_outs_2(ces_6_4_io_outs_2),
    .io_outs_3(ces_6_4_io_outs_3)
  );
  Element ces_6_5 ( // @[MockArray.scala 36:52]
    .clock(ces_6_5_clock),
    .io_ins_0(ces_6_5_io_ins_0),
    .io_ins_1(ces_6_5_io_ins_1),
    .io_ins_2(ces_6_5_io_ins_2),
    .io_ins_3(ces_6_5_io_ins_3),
    .io_outs_0(ces_6_5_io_outs_0),
    .io_outs_1(ces_6_5_io_outs_1),
    .io_outs_2(ces_6_5_io_outs_2),
    .io_outs_3(ces_6_5_io_outs_3)
  );
  Element ces_6_6 ( // @[MockArray.scala 36:52]
    .clock(ces_6_6_clock),
    .io_ins_0(ces_6_6_io_ins_0),
    .io_ins_1(ces_6_6_io_ins_1),
    .io_ins_2(ces_6_6_io_ins_2),
    .io_ins_3(ces_6_6_io_ins_3),
    .io_outs_0(ces_6_6_io_outs_0),
    .io_outs_1(ces_6_6_io_outs_1),
    .io_outs_2(ces_6_6_io_outs_2),
    .io_outs_3(ces_6_6_io_outs_3)
  );
  Element ces_6_7 ( // @[MockArray.scala 36:52]
    .clock(ces_6_7_clock),
    .io_ins_0(ces_6_7_io_ins_0),
    .io_ins_1(ces_6_7_io_ins_1),
    .io_ins_2(ces_6_7_io_ins_2),
    .io_ins_3(ces_6_7_io_ins_3),
    .io_outs_0(ces_6_7_io_outs_0),
    .io_outs_1(ces_6_7_io_outs_1),
    .io_outs_2(ces_6_7_io_outs_2),
    .io_outs_3(ces_6_7_io_outs_3)
  );
  Element ces_6_8 ( // @[MockArray.scala 36:52]
    .clock(ces_6_8_clock),
    .io_ins_0(ces_6_8_io_ins_0),
    .io_ins_1(ces_6_8_io_ins_1),
    .io_ins_2(ces_6_8_io_ins_2),
    .io_ins_3(ces_6_8_io_ins_3),
    .io_outs_0(ces_6_8_io_outs_0),
    .io_outs_1(ces_6_8_io_outs_1),
    .io_outs_2(ces_6_8_io_outs_2),
    .io_outs_3(ces_6_8_io_outs_3)
  );
  Element ces_6_9 ( // @[MockArray.scala 36:52]
    .clock(ces_6_9_clock),
    .io_ins_0(ces_6_9_io_ins_0),
    .io_ins_1(ces_6_9_io_ins_1),
    .io_ins_2(ces_6_9_io_ins_2),
    .io_ins_3(ces_6_9_io_ins_3),
    .io_outs_0(ces_6_9_io_outs_0),
    .io_outs_1(ces_6_9_io_outs_1),
    .io_outs_2(ces_6_9_io_outs_2),
    .io_outs_3(ces_6_9_io_outs_3)
  );
  Element ces_6_10 ( // @[MockArray.scala 36:52]
    .clock(ces_6_10_clock),
    .io_ins_0(ces_6_10_io_ins_0),
    .io_ins_1(ces_6_10_io_ins_1),
    .io_ins_2(ces_6_10_io_ins_2),
    .io_ins_3(ces_6_10_io_ins_3),
    .io_outs_0(ces_6_10_io_outs_0),
    .io_outs_1(ces_6_10_io_outs_1),
    .io_outs_2(ces_6_10_io_outs_2),
    .io_outs_3(ces_6_10_io_outs_3)
  );
  Element ces_6_11 ( // @[MockArray.scala 36:52]
    .clock(ces_6_11_clock),
    .io_ins_0(ces_6_11_io_ins_0),
    .io_ins_1(ces_6_11_io_ins_1),
    .io_ins_2(ces_6_11_io_ins_2),
    .io_ins_3(ces_6_11_io_ins_3),
    .io_outs_0(ces_6_11_io_outs_0),
    .io_outs_1(ces_6_11_io_outs_1),
    .io_outs_2(ces_6_11_io_outs_2),
    .io_outs_3(ces_6_11_io_outs_3)
  );
  Element ces_6_12 ( // @[MockArray.scala 36:52]
    .clock(ces_6_12_clock),
    .io_ins_0(ces_6_12_io_ins_0),
    .io_ins_1(ces_6_12_io_ins_1),
    .io_ins_2(ces_6_12_io_ins_2),
    .io_ins_3(ces_6_12_io_ins_3),
    .io_outs_0(ces_6_12_io_outs_0),
    .io_outs_1(ces_6_12_io_outs_1),
    .io_outs_2(ces_6_12_io_outs_2),
    .io_outs_3(ces_6_12_io_outs_3)
  );
  Element ces_6_13 ( // @[MockArray.scala 36:52]
    .clock(ces_6_13_clock),
    .io_ins_0(ces_6_13_io_ins_0),
    .io_ins_1(ces_6_13_io_ins_1),
    .io_ins_2(ces_6_13_io_ins_2),
    .io_ins_3(ces_6_13_io_ins_3),
    .io_outs_0(ces_6_13_io_outs_0),
    .io_outs_1(ces_6_13_io_outs_1),
    .io_outs_2(ces_6_13_io_outs_2),
    .io_outs_3(ces_6_13_io_outs_3)
  );
  Element ces_6_14 ( // @[MockArray.scala 36:52]
    .clock(ces_6_14_clock),
    .io_ins_0(ces_6_14_io_ins_0),
    .io_ins_1(ces_6_14_io_ins_1),
    .io_ins_2(ces_6_14_io_ins_2),
    .io_ins_3(ces_6_14_io_ins_3),
    .io_outs_0(ces_6_14_io_outs_0),
    .io_outs_1(ces_6_14_io_outs_1),
    .io_outs_2(ces_6_14_io_outs_2),
    .io_outs_3(ces_6_14_io_outs_3)
  );
  Element ces_6_15 ( // @[MockArray.scala 36:52]
    .clock(ces_6_15_clock),
    .io_ins_0(ces_6_15_io_ins_0),
    .io_ins_1(ces_6_15_io_ins_1),
    .io_ins_2(ces_6_15_io_ins_2),
    .io_ins_3(ces_6_15_io_ins_3),
    .io_outs_0(ces_6_15_io_outs_0),
    .io_outs_1(ces_6_15_io_outs_1),
    .io_outs_2(ces_6_15_io_outs_2),
    .io_outs_3(ces_6_15_io_outs_3)
  );
  Element ces_7_0 ( // @[MockArray.scala 36:52]
    .clock(ces_7_0_clock),
    .io_ins_0(ces_7_0_io_ins_0),
    .io_ins_1(ces_7_0_io_ins_1),
    .io_ins_2(ces_7_0_io_ins_2),
    .io_ins_3(ces_7_0_io_ins_3),
    .io_outs_0(ces_7_0_io_outs_0),
    .io_outs_1(ces_7_0_io_outs_1),
    .io_outs_2(ces_7_0_io_outs_2),
    .io_outs_3(ces_7_0_io_outs_3)
  );
  Element ces_7_1 ( // @[MockArray.scala 36:52]
    .clock(ces_7_1_clock),
    .io_ins_0(ces_7_1_io_ins_0),
    .io_ins_1(ces_7_1_io_ins_1),
    .io_ins_2(ces_7_1_io_ins_2),
    .io_ins_3(ces_7_1_io_ins_3),
    .io_outs_0(ces_7_1_io_outs_0),
    .io_outs_1(ces_7_1_io_outs_1),
    .io_outs_2(ces_7_1_io_outs_2),
    .io_outs_3(ces_7_1_io_outs_3)
  );
  Element ces_7_2 ( // @[MockArray.scala 36:52]
    .clock(ces_7_2_clock),
    .io_ins_0(ces_7_2_io_ins_0),
    .io_ins_1(ces_7_2_io_ins_1),
    .io_ins_2(ces_7_2_io_ins_2),
    .io_ins_3(ces_7_2_io_ins_3),
    .io_outs_0(ces_7_2_io_outs_0),
    .io_outs_1(ces_7_2_io_outs_1),
    .io_outs_2(ces_7_2_io_outs_2),
    .io_outs_3(ces_7_2_io_outs_3)
  );
  Element ces_7_3 ( // @[MockArray.scala 36:52]
    .clock(ces_7_3_clock),
    .io_ins_0(ces_7_3_io_ins_0),
    .io_ins_1(ces_7_3_io_ins_1),
    .io_ins_2(ces_7_3_io_ins_2),
    .io_ins_3(ces_7_3_io_ins_3),
    .io_outs_0(ces_7_3_io_outs_0),
    .io_outs_1(ces_7_3_io_outs_1),
    .io_outs_2(ces_7_3_io_outs_2),
    .io_outs_3(ces_7_3_io_outs_3)
  );
  Element ces_7_4 ( // @[MockArray.scala 36:52]
    .clock(ces_7_4_clock),
    .io_ins_0(ces_7_4_io_ins_0),
    .io_ins_1(ces_7_4_io_ins_1),
    .io_ins_2(ces_7_4_io_ins_2),
    .io_ins_3(ces_7_4_io_ins_3),
    .io_outs_0(ces_7_4_io_outs_0),
    .io_outs_1(ces_7_4_io_outs_1),
    .io_outs_2(ces_7_4_io_outs_2),
    .io_outs_3(ces_7_4_io_outs_3)
  );
  Element ces_7_5 ( // @[MockArray.scala 36:52]
    .clock(ces_7_5_clock),
    .io_ins_0(ces_7_5_io_ins_0),
    .io_ins_1(ces_7_5_io_ins_1),
    .io_ins_2(ces_7_5_io_ins_2),
    .io_ins_3(ces_7_5_io_ins_3),
    .io_outs_0(ces_7_5_io_outs_0),
    .io_outs_1(ces_7_5_io_outs_1),
    .io_outs_2(ces_7_5_io_outs_2),
    .io_outs_3(ces_7_5_io_outs_3)
  );
  Element ces_7_6 ( // @[MockArray.scala 36:52]
    .clock(ces_7_6_clock),
    .io_ins_0(ces_7_6_io_ins_0),
    .io_ins_1(ces_7_6_io_ins_1),
    .io_ins_2(ces_7_6_io_ins_2),
    .io_ins_3(ces_7_6_io_ins_3),
    .io_outs_0(ces_7_6_io_outs_0),
    .io_outs_1(ces_7_6_io_outs_1),
    .io_outs_2(ces_7_6_io_outs_2),
    .io_outs_3(ces_7_6_io_outs_3)
  );
  Element ces_7_7 ( // @[MockArray.scala 36:52]
    .clock(ces_7_7_clock),
    .io_ins_0(ces_7_7_io_ins_0),
    .io_ins_1(ces_7_7_io_ins_1),
    .io_ins_2(ces_7_7_io_ins_2),
    .io_ins_3(ces_7_7_io_ins_3),
    .io_outs_0(ces_7_7_io_outs_0),
    .io_outs_1(ces_7_7_io_outs_1),
    .io_outs_2(ces_7_7_io_outs_2),
    .io_outs_3(ces_7_7_io_outs_3)
  );
  Element ces_7_8 ( // @[MockArray.scala 36:52]
    .clock(ces_7_8_clock),
    .io_ins_0(ces_7_8_io_ins_0),
    .io_ins_1(ces_7_8_io_ins_1),
    .io_ins_2(ces_7_8_io_ins_2),
    .io_ins_3(ces_7_8_io_ins_3),
    .io_outs_0(ces_7_8_io_outs_0),
    .io_outs_1(ces_7_8_io_outs_1),
    .io_outs_2(ces_7_8_io_outs_2),
    .io_outs_3(ces_7_8_io_outs_3)
  );
  Element ces_7_9 ( // @[MockArray.scala 36:52]
    .clock(ces_7_9_clock),
    .io_ins_0(ces_7_9_io_ins_0),
    .io_ins_1(ces_7_9_io_ins_1),
    .io_ins_2(ces_7_9_io_ins_2),
    .io_ins_3(ces_7_9_io_ins_3),
    .io_outs_0(ces_7_9_io_outs_0),
    .io_outs_1(ces_7_9_io_outs_1),
    .io_outs_2(ces_7_9_io_outs_2),
    .io_outs_3(ces_7_9_io_outs_3)
  );
  Element ces_7_10 ( // @[MockArray.scala 36:52]
    .clock(ces_7_10_clock),
    .io_ins_0(ces_7_10_io_ins_0),
    .io_ins_1(ces_7_10_io_ins_1),
    .io_ins_2(ces_7_10_io_ins_2),
    .io_ins_3(ces_7_10_io_ins_3),
    .io_outs_0(ces_7_10_io_outs_0),
    .io_outs_1(ces_7_10_io_outs_1),
    .io_outs_2(ces_7_10_io_outs_2),
    .io_outs_3(ces_7_10_io_outs_3)
  );
  Element ces_7_11 ( // @[MockArray.scala 36:52]
    .clock(ces_7_11_clock),
    .io_ins_0(ces_7_11_io_ins_0),
    .io_ins_1(ces_7_11_io_ins_1),
    .io_ins_2(ces_7_11_io_ins_2),
    .io_ins_3(ces_7_11_io_ins_3),
    .io_outs_0(ces_7_11_io_outs_0),
    .io_outs_1(ces_7_11_io_outs_1),
    .io_outs_2(ces_7_11_io_outs_2),
    .io_outs_3(ces_7_11_io_outs_3)
  );
  Element ces_7_12 ( // @[MockArray.scala 36:52]
    .clock(ces_7_12_clock),
    .io_ins_0(ces_7_12_io_ins_0),
    .io_ins_1(ces_7_12_io_ins_1),
    .io_ins_2(ces_7_12_io_ins_2),
    .io_ins_3(ces_7_12_io_ins_3),
    .io_outs_0(ces_7_12_io_outs_0),
    .io_outs_1(ces_7_12_io_outs_1),
    .io_outs_2(ces_7_12_io_outs_2),
    .io_outs_3(ces_7_12_io_outs_3)
  );
  Element ces_7_13 ( // @[MockArray.scala 36:52]
    .clock(ces_7_13_clock),
    .io_ins_0(ces_7_13_io_ins_0),
    .io_ins_1(ces_7_13_io_ins_1),
    .io_ins_2(ces_7_13_io_ins_2),
    .io_ins_3(ces_7_13_io_ins_3),
    .io_outs_0(ces_7_13_io_outs_0),
    .io_outs_1(ces_7_13_io_outs_1),
    .io_outs_2(ces_7_13_io_outs_2),
    .io_outs_3(ces_7_13_io_outs_3)
  );
  Element ces_7_14 ( // @[MockArray.scala 36:52]
    .clock(ces_7_14_clock),
    .io_ins_0(ces_7_14_io_ins_0),
    .io_ins_1(ces_7_14_io_ins_1),
    .io_ins_2(ces_7_14_io_ins_2),
    .io_ins_3(ces_7_14_io_ins_3),
    .io_outs_0(ces_7_14_io_outs_0),
    .io_outs_1(ces_7_14_io_outs_1),
    .io_outs_2(ces_7_14_io_outs_2),
    .io_outs_3(ces_7_14_io_outs_3)
  );
  Element ces_7_15 ( // @[MockArray.scala 36:52]
    .clock(ces_7_15_clock),
    .io_ins_0(ces_7_15_io_ins_0),
    .io_ins_1(ces_7_15_io_ins_1),
    .io_ins_2(ces_7_15_io_ins_2),
    .io_ins_3(ces_7_15_io_ins_3),
    .io_outs_0(ces_7_15_io_outs_0),
    .io_outs_1(ces_7_15_io_outs_1),
    .io_outs_2(ces_7_15_io_outs_2),
    .io_outs_3(ces_7_15_io_outs_3)
  );
  assign io_outsHorizontal_0_0 = ces_0_0_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_1 = ces_0_1_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_2 = ces_0_2_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_3 = ces_0_3_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_4 = ces_0_4_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_5 = ces_0_5_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_6 = ces_0_6_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_7 = ces_0_7_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_8 = ces_0_8_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_9 = ces_0_9_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_10 = ces_0_10_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_11 = ces_0_11_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_12 = ces_0_12_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_13 = ces_0_13_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_14 = ces_0_14_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_15 = ces_0_15_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_1_0 = ces_7_0_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_1 = ces_7_1_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_2 = ces_7_2_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_3 = ces_7_3_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_4 = ces_7_4_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_5 = ces_7_5_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_6 = ces_7_6_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_7 = ces_7_7_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_8 = ces_7_8_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_9 = ces_7_9_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_10 = ces_7_10_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_11 = ces_7_11_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_12 = ces_7_12_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_13 = ces_7_13_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_14 = ces_7_14_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_15 = ces_7_15_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_0 = ces_0_15_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_1 = ces_1_15_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_2 = ces_2_15_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_3 = ces_3_15_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_4 = ces_4_15_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_5 = ces_5_15_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_6 = ces_6_15_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_7 = ces_7_15_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_1_0 = ces_0_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_1 = ces_1_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_2 = ces_2_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_3 = ces_3_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_4 = ces_4_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_5 = ces_5_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_6 = ces_6_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_7 = ces_7_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_lsbs_0 = ces_0_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1 = ces_0_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_2 = ces_0_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_3 = ces_0_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_4 = ces_0_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_5 = ces_0_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_6 = ces_0_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_7 = ces_0_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_8 = ces_0_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_9 = ces_0_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_10 = ces_0_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_11 = ces_0_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_12 = ces_0_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_13 = ces_0_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_14 = ces_0_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_15 = ces_0_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_16 = ces_1_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_17 = ces_1_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_18 = ces_1_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_19 = ces_1_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_20 = ces_1_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_21 = ces_1_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_22 = ces_1_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_23 = ces_1_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_24 = ces_1_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_25 = ces_1_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_26 = ces_1_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_27 = ces_1_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_28 = ces_1_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_29 = ces_1_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_30 = ces_1_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_31 = ces_1_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_32 = ces_2_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_33 = ces_2_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_34 = ces_2_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_35 = ces_2_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_36 = ces_2_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_37 = ces_2_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_38 = ces_2_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_39 = ces_2_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_40 = ces_2_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_41 = ces_2_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_42 = ces_2_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_43 = ces_2_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_44 = ces_2_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_45 = ces_2_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_46 = ces_2_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_47 = ces_2_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_48 = ces_3_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_49 = ces_3_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_50 = ces_3_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_51 = ces_3_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_52 = ces_3_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_53 = ces_3_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_54 = ces_3_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_55 = ces_3_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_56 = ces_3_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_57 = ces_3_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_58 = ces_3_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_59 = ces_3_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_60 = ces_3_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_61 = ces_3_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_62 = ces_3_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_63 = ces_3_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_64 = ces_4_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_65 = ces_4_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_66 = ces_4_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_67 = ces_4_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_68 = ces_4_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_69 = ces_4_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_70 = ces_4_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_71 = ces_4_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_72 = ces_4_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_73 = ces_4_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_74 = ces_4_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_75 = ces_4_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_76 = ces_4_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_77 = ces_4_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_78 = ces_4_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_79 = ces_4_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_80 = ces_5_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_81 = ces_5_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_82 = ces_5_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_83 = ces_5_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_84 = ces_5_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_85 = ces_5_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_86 = ces_5_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_87 = ces_5_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_88 = ces_5_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_89 = ces_5_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_90 = ces_5_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_91 = ces_5_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_92 = ces_5_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_93 = ces_5_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_94 = ces_5_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_95 = ces_5_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_96 = ces_6_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_97 = ces_6_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_98 = ces_6_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_99 = ces_6_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_100 = ces_6_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_101 = ces_6_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_102 = ces_6_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_103 = ces_6_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_104 = ces_6_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_105 = ces_6_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_106 = ces_6_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_107 = ces_6_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_108 = ces_6_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_109 = ces_6_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_110 = ces_6_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_111 = ces_6_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_112 = ces_7_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_113 = ces_7_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_114 = ces_7_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_115 = ces_7_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_116 = ces_7_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_117 = ces_7_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_118 = ces_7_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_119 = ces_7_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_120 = ces_7_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_121 = ces_7_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_122 = ces_7_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_123 = ces_7_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_124 = ces_7_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_125 = ces_7_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_126 = ces_7_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_127 = ces_7_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign ces_0_0_clock = clock;
  assign ces_0_0_io_ins_0 = io_insHorizontal_0_0; // @[MockArray.scala 44:87]
  assign ces_0_0_io_ins_1 = ces_0_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_0_io_ins_2 = ces_1_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_0_io_ins_3 = io_insVertical_1_0; // @[MockArray.scala 47:87]
  assign ces_0_1_clock = clock;
  assign ces_0_1_io_ins_0 = io_insHorizontal_0_1; // @[MockArray.scala 44:87]
  assign ces_0_1_io_ins_1 = ces_0_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_1_io_ins_2 = ces_1_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_1_io_ins_3 = ces_0_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_2_clock = clock;
  assign ces_0_2_io_ins_0 = io_insHorizontal_0_2; // @[MockArray.scala 44:87]
  assign ces_0_2_io_ins_1 = ces_0_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_2_io_ins_2 = ces_1_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_2_io_ins_3 = ces_0_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_3_clock = clock;
  assign ces_0_3_io_ins_0 = io_insHorizontal_0_3; // @[MockArray.scala 44:87]
  assign ces_0_3_io_ins_1 = ces_0_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_3_io_ins_2 = ces_1_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_3_io_ins_3 = ces_0_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_4_clock = clock;
  assign ces_0_4_io_ins_0 = io_insHorizontal_0_4; // @[MockArray.scala 44:87]
  assign ces_0_4_io_ins_1 = ces_0_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_4_io_ins_2 = ces_1_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_4_io_ins_3 = ces_0_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_5_clock = clock;
  assign ces_0_5_io_ins_0 = io_insHorizontal_0_5; // @[MockArray.scala 44:87]
  assign ces_0_5_io_ins_1 = ces_0_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_5_io_ins_2 = ces_1_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_5_io_ins_3 = ces_0_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_6_clock = clock;
  assign ces_0_6_io_ins_0 = io_insHorizontal_0_6; // @[MockArray.scala 44:87]
  assign ces_0_6_io_ins_1 = ces_0_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_6_io_ins_2 = ces_1_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_6_io_ins_3 = ces_0_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_7_clock = clock;
  assign ces_0_7_io_ins_0 = io_insHorizontal_0_7; // @[MockArray.scala 44:87]
  assign ces_0_7_io_ins_1 = ces_0_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_7_io_ins_2 = ces_1_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_7_io_ins_3 = ces_0_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_8_clock = clock;
  assign ces_0_8_io_ins_0 = io_insHorizontal_0_8; // @[MockArray.scala 44:87]
  assign ces_0_8_io_ins_1 = ces_0_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_8_io_ins_2 = ces_1_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_8_io_ins_3 = ces_0_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_9_clock = clock;
  assign ces_0_9_io_ins_0 = io_insHorizontal_0_9; // @[MockArray.scala 44:87]
  assign ces_0_9_io_ins_1 = ces_0_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_9_io_ins_2 = ces_1_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_9_io_ins_3 = ces_0_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_10_clock = clock;
  assign ces_0_10_io_ins_0 = io_insHorizontal_0_10; // @[MockArray.scala 44:87]
  assign ces_0_10_io_ins_1 = ces_0_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_10_io_ins_2 = ces_1_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_10_io_ins_3 = ces_0_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_11_clock = clock;
  assign ces_0_11_io_ins_0 = io_insHorizontal_0_11; // @[MockArray.scala 44:87]
  assign ces_0_11_io_ins_1 = ces_0_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_11_io_ins_2 = ces_1_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_11_io_ins_3 = ces_0_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_12_clock = clock;
  assign ces_0_12_io_ins_0 = io_insHorizontal_0_12; // @[MockArray.scala 44:87]
  assign ces_0_12_io_ins_1 = ces_0_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_12_io_ins_2 = ces_1_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_12_io_ins_3 = ces_0_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_13_clock = clock;
  assign ces_0_13_io_ins_0 = io_insHorizontal_0_13; // @[MockArray.scala 44:87]
  assign ces_0_13_io_ins_1 = ces_0_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_13_io_ins_2 = ces_1_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_13_io_ins_3 = ces_0_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_14_clock = clock;
  assign ces_0_14_io_ins_0 = io_insHorizontal_0_14; // @[MockArray.scala 44:87]
  assign ces_0_14_io_ins_1 = ces_0_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_14_io_ins_2 = ces_1_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_14_io_ins_3 = ces_0_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_15_clock = clock;
  assign ces_0_15_io_ins_0 = io_insHorizontal_0_15; // @[MockArray.scala 44:87]
  assign ces_0_15_io_ins_1 = io_insVertical_0_0; // @[MockArray.scala 45:87]
  assign ces_0_15_io_ins_2 = ces_1_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_15_io_ins_3 = ces_0_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_0_clock = clock;
  assign ces_1_0_io_ins_0 = ces_0_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_0_io_ins_1 = ces_1_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_0_io_ins_2 = ces_2_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_0_io_ins_3 = io_insVertical_1_1; // @[MockArray.scala 47:87]
  assign ces_1_1_clock = clock;
  assign ces_1_1_io_ins_0 = ces_0_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_1_io_ins_1 = ces_1_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_1_io_ins_2 = ces_2_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_1_io_ins_3 = ces_1_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_2_clock = clock;
  assign ces_1_2_io_ins_0 = ces_0_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_2_io_ins_1 = ces_1_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_2_io_ins_2 = ces_2_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_2_io_ins_3 = ces_1_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_3_clock = clock;
  assign ces_1_3_io_ins_0 = ces_0_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_3_io_ins_1 = ces_1_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_3_io_ins_2 = ces_2_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_3_io_ins_3 = ces_1_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_4_clock = clock;
  assign ces_1_4_io_ins_0 = ces_0_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_4_io_ins_1 = ces_1_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_4_io_ins_2 = ces_2_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_4_io_ins_3 = ces_1_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_5_clock = clock;
  assign ces_1_5_io_ins_0 = ces_0_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_5_io_ins_1 = ces_1_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_5_io_ins_2 = ces_2_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_5_io_ins_3 = ces_1_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_6_clock = clock;
  assign ces_1_6_io_ins_0 = ces_0_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_6_io_ins_1 = ces_1_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_6_io_ins_2 = ces_2_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_6_io_ins_3 = ces_1_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_7_clock = clock;
  assign ces_1_7_io_ins_0 = ces_0_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_7_io_ins_1 = ces_1_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_7_io_ins_2 = ces_2_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_7_io_ins_3 = ces_1_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_8_clock = clock;
  assign ces_1_8_io_ins_0 = ces_0_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_8_io_ins_1 = ces_1_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_8_io_ins_2 = ces_2_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_8_io_ins_3 = ces_1_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_9_clock = clock;
  assign ces_1_9_io_ins_0 = ces_0_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_9_io_ins_1 = ces_1_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_9_io_ins_2 = ces_2_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_9_io_ins_3 = ces_1_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_10_clock = clock;
  assign ces_1_10_io_ins_0 = ces_0_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_10_io_ins_1 = ces_1_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_10_io_ins_2 = ces_2_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_10_io_ins_3 = ces_1_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_11_clock = clock;
  assign ces_1_11_io_ins_0 = ces_0_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_11_io_ins_1 = ces_1_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_11_io_ins_2 = ces_2_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_11_io_ins_3 = ces_1_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_12_clock = clock;
  assign ces_1_12_io_ins_0 = ces_0_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_12_io_ins_1 = ces_1_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_12_io_ins_2 = ces_2_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_12_io_ins_3 = ces_1_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_13_clock = clock;
  assign ces_1_13_io_ins_0 = ces_0_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_13_io_ins_1 = ces_1_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_13_io_ins_2 = ces_2_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_13_io_ins_3 = ces_1_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_14_clock = clock;
  assign ces_1_14_io_ins_0 = ces_0_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_14_io_ins_1 = ces_1_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_14_io_ins_2 = ces_2_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_14_io_ins_3 = ces_1_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_15_clock = clock;
  assign ces_1_15_io_ins_0 = ces_0_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_15_io_ins_1 = io_insVertical_0_1; // @[MockArray.scala 45:87]
  assign ces_1_15_io_ins_2 = ces_2_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_15_io_ins_3 = ces_1_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_0_clock = clock;
  assign ces_2_0_io_ins_0 = ces_1_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_0_io_ins_1 = ces_2_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_0_io_ins_2 = ces_3_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_0_io_ins_3 = io_insVertical_1_2; // @[MockArray.scala 47:87]
  assign ces_2_1_clock = clock;
  assign ces_2_1_io_ins_0 = ces_1_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_1_io_ins_1 = ces_2_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_1_io_ins_2 = ces_3_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_1_io_ins_3 = ces_2_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_2_clock = clock;
  assign ces_2_2_io_ins_0 = ces_1_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_2_io_ins_1 = ces_2_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_2_io_ins_2 = ces_3_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_2_io_ins_3 = ces_2_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_3_clock = clock;
  assign ces_2_3_io_ins_0 = ces_1_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_3_io_ins_1 = ces_2_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_3_io_ins_2 = ces_3_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_3_io_ins_3 = ces_2_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_4_clock = clock;
  assign ces_2_4_io_ins_0 = ces_1_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_4_io_ins_1 = ces_2_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_4_io_ins_2 = ces_3_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_4_io_ins_3 = ces_2_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_5_clock = clock;
  assign ces_2_5_io_ins_0 = ces_1_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_5_io_ins_1 = ces_2_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_5_io_ins_2 = ces_3_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_5_io_ins_3 = ces_2_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_6_clock = clock;
  assign ces_2_6_io_ins_0 = ces_1_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_6_io_ins_1 = ces_2_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_6_io_ins_2 = ces_3_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_6_io_ins_3 = ces_2_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_7_clock = clock;
  assign ces_2_7_io_ins_0 = ces_1_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_7_io_ins_1 = ces_2_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_7_io_ins_2 = ces_3_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_7_io_ins_3 = ces_2_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_8_clock = clock;
  assign ces_2_8_io_ins_0 = ces_1_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_8_io_ins_1 = ces_2_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_8_io_ins_2 = ces_3_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_8_io_ins_3 = ces_2_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_9_clock = clock;
  assign ces_2_9_io_ins_0 = ces_1_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_9_io_ins_1 = ces_2_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_9_io_ins_2 = ces_3_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_9_io_ins_3 = ces_2_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_10_clock = clock;
  assign ces_2_10_io_ins_0 = ces_1_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_10_io_ins_1 = ces_2_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_10_io_ins_2 = ces_3_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_10_io_ins_3 = ces_2_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_11_clock = clock;
  assign ces_2_11_io_ins_0 = ces_1_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_11_io_ins_1 = ces_2_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_11_io_ins_2 = ces_3_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_11_io_ins_3 = ces_2_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_12_clock = clock;
  assign ces_2_12_io_ins_0 = ces_1_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_12_io_ins_1 = ces_2_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_12_io_ins_2 = ces_3_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_12_io_ins_3 = ces_2_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_13_clock = clock;
  assign ces_2_13_io_ins_0 = ces_1_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_13_io_ins_1 = ces_2_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_13_io_ins_2 = ces_3_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_13_io_ins_3 = ces_2_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_14_clock = clock;
  assign ces_2_14_io_ins_0 = ces_1_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_14_io_ins_1 = ces_2_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_14_io_ins_2 = ces_3_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_14_io_ins_3 = ces_2_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_15_clock = clock;
  assign ces_2_15_io_ins_0 = ces_1_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_15_io_ins_1 = io_insVertical_0_2; // @[MockArray.scala 45:87]
  assign ces_2_15_io_ins_2 = ces_3_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_15_io_ins_3 = ces_2_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_0_clock = clock;
  assign ces_3_0_io_ins_0 = ces_2_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_0_io_ins_1 = ces_3_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_0_io_ins_2 = ces_4_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_0_io_ins_3 = io_insVertical_1_3; // @[MockArray.scala 47:87]
  assign ces_3_1_clock = clock;
  assign ces_3_1_io_ins_0 = ces_2_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_1_io_ins_1 = ces_3_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_1_io_ins_2 = ces_4_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_1_io_ins_3 = ces_3_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_2_clock = clock;
  assign ces_3_2_io_ins_0 = ces_2_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_2_io_ins_1 = ces_3_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_2_io_ins_2 = ces_4_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_2_io_ins_3 = ces_3_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_3_clock = clock;
  assign ces_3_3_io_ins_0 = ces_2_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_3_io_ins_1 = ces_3_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_3_io_ins_2 = ces_4_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_3_io_ins_3 = ces_3_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_4_clock = clock;
  assign ces_3_4_io_ins_0 = ces_2_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_4_io_ins_1 = ces_3_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_4_io_ins_2 = ces_4_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_4_io_ins_3 = ces_3_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_5_clock = clock;
  assign ces_3_5_io_ins_0 = ces_2_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_5_io_ins_1 = ces_3_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_5_io_ins_2 = ces_4_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_5_io_ins_3 = ces_3_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_6_clock = clock;
  assign ces_3_6_io_ins_0 = ces_2_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_6_io_ins_1 = ces_3_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_6_io_ins_2 = ces_4_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_6_io_ins_3 = ces_3_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_7_clock = clock;
  assign ces_3_7_io_ins_0 = ces_2_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_7_io_ins_1 = ces_3_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_7_io_ins_2 = ces_4_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_7_io_ins_3 = ces_3_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_8_clock = clock;
  assign ces_3_8_io_ins_0 = ces_2_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_8_io_ins_1 = ces_3_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_8_io_ins_2 = ces_4_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_8_io_ins_3 = ces_3_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_9_clock = clock;
  assign ces_3_9_io_ins_0 = ces_2_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_9_io_ins_1 = ces_3_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_9_io_ins_2 = ces_4_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_9_io_ins_3 = ces_3_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_10_clock = clock;
  assign ces_3_10_io_ins_0 = ces_2_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_10_io_ins_1 = ces_3_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_10_io_ins_2 = ces_4_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_10_io_ins_3 = ces_3_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_11_clock = clock;
  assign ces_3_11_io_ins_0 = ces_2_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_11_io_ins_1 = ces_3_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_11_io_ins_2 = ces_4_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_11_io_ins_3 = ces_3_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_12_clock = clock;
  assign ces_3_12_io_ins_0 = ces_2_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_12_io_ins_1 = ces_3_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_12_io_ins_2 = ces_4_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_12_io_ins_3 = ces_3_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_13_clock = clock;
  assign ces_3_13_io_ins_0 = ces_2_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_13_io_ins_1 = ces_3_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_13_io_ins_2 = ces_4_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_13_io_ins_3 = ces_3_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_14_clock = clock;
  assign ces_3_14_io_ins_0 = ces_2_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_14_io_ins_1 = ces_3_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_14_io_ins_2 = ces_4_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_14_io_ins_3 = ces_3_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_15_clock = clock;
  assign ces_3_15_io_ins_0 = ces_2_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_15_io_ins_1 = io_insVertical_0_3; // @[MockArray.scala 45:87]
  assign ces_3_15_io_ins_2 = ces_4_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_15_io_ins_3 = ces_3_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_0_clock = clock;
  assign ces_4_0_io_ins_0 = ces_3_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_0_io_ins_1 = ces_4_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_0_io_ins_2 = ces_5_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_0_io_ins_3 = io_insVertical_1_4; // @[MockArray.scala 47:87]
  assign ces_4_1_clock = clock;
  assign ces_4_1_io_ins_0 = ces_3_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_1_io_ins_1 = ces_4_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_1_io_ins_2 = ces_5_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_1_io_ins_3 = ces_4_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_2_clock = clock;
  assign ces_4_2_io_ins_0 = ces_3_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_2_io_ins_1 = ces_4_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_2_io_ins_2 = ces_5_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_2_io_ins_3 = ces_4_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_3_clock = clock;
  assign ces_4_3_io_ins_0 = ces_3_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_3_io_ins_1 = ces_4_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_3_io_ins_2 = ces_5_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_3_io_ins_3 = ces_4_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_4_clock = clock;
  assign ces_4_4_io_ins_0 = ces_3_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_4_io_ins_1 = ces_4_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_4_io_ins_2 = ces_5_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_4_io_ins_3 = ces_4_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_5_clock = clock;
  assign ces_4_5_io_ins_0 = ces_3_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_5_io_ins_1 = ces_4_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_5_io_ins_2 = ces_5_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_5_io_ins_3 = ces_4_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_6_clock = clock;
  assign ces_4_6_io_ins_0 = ces_3_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_6_io_ins_1 = ces_4_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_6_io_ins_2 = ces_5_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_6_io_ins_3 = ces_4_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_7_clock = clock;
  assign ces_4_7_io_ins_0 = ces_3_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_7_io_ins_1 = ces_4_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_7_io_ins_2 = ces_5_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_7_io_ins_3 = ces_4_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_8_clock = clock;
  assign ces_4_8_io_ins_0 = ces_3_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_8_io_ins_1 = ces_4_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_8_io_ins_2 = ces_5_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_8_io_ins_3 = ces_4_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_9_clock = clock;
  assign ces_4_9_io_ins_0 = ces_3_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_9_io_ins_1 = ces_4_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_9_io_ins_2 = ces_5_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_9_io_ins_3 = ces_4_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_10_clock = clock;
  assign ces_4_10_io_ins_0 = ces_3_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_10_io_ins_1 = ces_4_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_10_io_ins_2 = ces_5_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_10_io_ins_3 = ces_4_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_11_clock = clock;
  assign ces_4_11_io_ins_0 = ces_3_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_11_io_ins_1 = ces_4_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_11_io_ins_2 = ces_5_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_11_io_ins_3 = ces_4_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_12_clock = clock;
  assign ces_4_12_io_ins_0 = ces_3_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_12_io_ins_1 = ces_4_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_12_io_ins_2 = ces_5_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_12_io_ins_3 = ces_4_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_13_clock = clock;
  assign ces_4_13_io_ins_0 = ces_3_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_13_io_ins_1 = ces_4_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_13_io_ins_2 = ces_5_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_13_io_ins_3 = ces_4_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_14_clock = clock;
  assign ces_4_14_io_ins_0 = ces_3_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_14_io_ins_1 = ces_4_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_14_io_ins_2 = ces_5_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_14_io_ins_3 = ces_4_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_15_clock = clock;
  assign ces_4_15_io_ins_0 = ces_3_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_15_io_ins_1 = io_insVertical_0_4; // @[MockArray.scala 45:87]
  assign ces_4_15_io_ins_2 = ces_5_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_15_io_ins_3 = ces_4_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_0_clock = clock;
  assign ces_5_0_io_ins_0 = ces_4_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_0_io_ins_1 = ces_5_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_0_io_ins_2 = ces_6_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_0_io_ins_3 = io_insVertical_1_5; // @[MockArray.scala 47:87]
  assign ces_5_1_clock = clock;
  assign ces_5_1_io_ins_0 = ces_4_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_1_io_ins_1 = ces_5_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_1_io_ins_2 = ces_6_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_1_io_ins_3 = ces_5_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_2_clock = clock;
  assign ces_5_2_io_ins_0 = ces_4_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_2_io_ins_1 = ces_5_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_2_io_ins_2 = ces_6_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_2_io_ins_3 = ces_5_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_3_clock = clock;
  assign ces_5_3_io_ins_0 = ces_4_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_3_io_ins_1 = ces_5_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_3_io_ins_2 = ces_6_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_3_io_ins_3 = ces_5_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_4_clock = clock;
  assign ces_5_4_io_ins_0 = ces_4_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_4_io_ins_1 = ces_5_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_4_io_ins_2 = ces_6_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_4_io_ins_3 = ces_5_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_5_clock = clock;
  assign ces_5_5_io_ins_0 = ces_4_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_5_io_ins_1 = ces_5_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_5_io_ins_2 = ces_6_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_5_io_ins_3 = ces_5_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_6_clock = clock;
  assign ces_5_6_io_ins_0 = ces_4_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_6_io_ins_1 = ces_5_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_6_io_ins_2 = ces_6_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_6_io_ins_3 = ces_5_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_7_clock = clock;
  assign ces_5_7_io_ins_0 = ces_4_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_7_io_ins_1 = ces_5_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_7_io_ins_2 = ces_6_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_7_io_ins_3 = ces_5_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_8_clock = clock;
  assign ces_5_8_io_ins_0 = ces_4_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_8_io_ins_1 = ces_5_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_8_io_ins_2 = ces_6_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_8_io_ins_3 = ces_5_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_9_clock = clock;
  assign ces_5_9_io_ins_0 = ces_4_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_9_io_ins_1 = ces_5_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_9_io_ins_2 = ces_6_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_9_io_ins_3 = ces_5_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_10_clock = clock;
  assign ces_5_10_io_ins_0 = ces_4_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_10_io_ins_1 = ces_5_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_10_io_ins_2 = ces_6_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_10_io_ins_3 = ces_5_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_11_clock = clock;
  assign ces_5_11_io_ins_0 = ces_4_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_11_io_ins_1 = ces_5_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_11_io_ins_2 = ces_6_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_11_io_ins_3 = ces_5_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_12_clock = clock;
  assign ces_5_12_io_ins_0 = ces_4_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_12_io_ins_1 = ces_5_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_12_io_ins_2 = ces_6_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_12_io_ins_3 = ces_5_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_13_clock = clock;
  assign ces_5_13_io_ins_0 = ces_4_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_13_io_ins_1 = ces_5_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_13_io_ins_2 = ces_6_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_13_io_ins_3 = ces_5_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_14_clock = clock;
  assign ces_5_14_io_ins_0 = ces_4_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_14_io_ins_1 = ces_5_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_14_io_ins_2 = ces_6_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_14_io_ins_3 = ces_5_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_15_clock = clock;
  assign ces_5_15_io_ins_0 = ces_4_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_15_io_ins_1 = io_insVertical_0_5; // @[MockArray.scala 45:87]
  assign ces_5_15_io_ins_2 = ces_6_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_15_io_ins_3 = ces_5_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_0_clock = clock;
  assign ces_6_0_io_ins_0 = ces_5_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_0_io_ins_1 = ces_6_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_0_io_ins_2 = ces_7_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_0_io_ins_3 = io_insVertical_1_6; // @[MockArray.scala 47:87]
  assign ces_6_1_clock = clock;
  assign ces_6_1_io_ins_0 = ces_5_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_1_io_ins_1 = ces_6_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_1_io_ins_2 = ces_7_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_1_io_ins_3 = ces_6_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_2_clock = clock;
  assign ces_6_2_io_ins_0 = ces_5_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_2_io_ins_1 = ces_6_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_2_io_ins_2 = ces_7_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_2_io_ins_3 = ces_6_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_3_clock = clock;
  assign ces_6_3_io_ins_0 = ces_5_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_3_io_ins_1 = ces_6_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_3_io_ins_2 = ces_7_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_3_io_ins_3 = ces_6_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_4_clock = clock;
  assign ces_6_4_io_ins_0 = ces_5_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_4_io_ins_1 = ces_6_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_4_io_ins_2 = ces_7_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_4_io_ins_3 = ces_6_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_5_clock = clock;
  assign ces_6_5_io_ins_0 = ces_5_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_5_io_ins_1 = ces_6_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_5_io_ins_2 = ces_7_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_5_io_ins_3 = ces_6_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_6_clock = clock;
  assign ces_6_6_io_ins_0 = ces_5_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_6_io_ins_1 = ces_6_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_6_io_ins_2 = ces_7_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_6_io_ins_3 = ces_6_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_7_clock = clock;
  assign ces_6_7_io_ins_0 = ces_5_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_7_io_ins_1 = ces_6_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_7_io_ins_2 = ces_7_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_7_io_ins_3 = ces_6_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_8_clock = clock;
  assign ces_6_8_io_ins_0 = ces_5_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_8_io_ins_1 = ces_6_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_8_io_ins_2 = ces_7_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_8_io_ins_3 = ces_6_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_9_clock = clock;
  assign ces_6_9_io_ins_0 = ces_5_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_9_io_ins_1 = ces_6_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_9_io_ins_2 = ces_7_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_9_io_ins_3 = ces_6_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_10_clock = clock;
  assign ces_6_10_io_ins_0 = ces_5_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_10_io_ins_1 = ces_6_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_10_io_ins_2 = ces_7_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_10_io_ins_3 = ces_6_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_11_clock = clock;
  assign ces_6_11_io_ins_0 = ces_5_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_11_io_ins_1 = ces_6_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_11_io_ins_2 = ces_7_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_11_io_ins_3 = ces_6_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_12_clock = clock;
  assign ces_6_12_io_ins_0 = ces_5_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_12_io_ins_1 = ces_6_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_12_io_ins_2 = ces_7_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_12_io_ins_3 = ces_6_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_13_clock = clock;
  assign ces_6_13_io_ins_0 = ces_5_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_13_io_ins_1 = ces_6_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_13_io_ins_2 = ces_7_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_13_io_ins_3 = ces_6_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_14_clock = clock;
  assign ces_6_14_io_ins_0 = ces_5_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_14_io_ins_1 = ces_6_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_14_io_ins_2 = ces_7_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_14_io_ins_3 = ces_6_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_15_clock = clock;
  assign ces_6_15_io_ins_0 = ces_5_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_15_io_ins_1 = io_insVertical_0_6; // @[MockArray.scala 45:87]
  assign ces_6_15_io_ins_2 = ces_7_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_15_io_ins_3 = ces_6_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_0_clock = clock;
  assign ces_7_0_io_ins_0 = ces_6_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_0_io_ins_1 = ces_7_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_0_io_ins_2 = io_insHorizontal_1_0; // @[MockArray.scala 46:87]
  assign ces_7_0_io_ins_3 = io_insVertical_1_7; // @[MockArray.scala 47:87]
  assign ces_7_1_clock = clock;
  assign ces_7_1_io_ins_0 = ces_6_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_1_io_ins_1 = ces_7_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_1_io_ins_2 = io_insHorizontal_1_1; // @[MockArray.scala 46:87]
  assign ces_7_1_io_ins_3 = ces_7_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_2_clock = clock;
  assign ces_7_2_io_ins_0 = ces_6_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_2_io_ins_1 = ces_7_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_2_io_ins_2 = io_insHorizontal_1_2; // @[MockArray.scala 46:87]
  assign ces_7_2_io_ins_3 = ces_7_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_3_clock = clock;
  assign ces_7_3_io_ins_0 = ces_6_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_3_io_ins_1 = ces_7_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_3_io_ins_2 = io_insHorizontal_1_3; // @[MockArray.scala 46:87]
  assign ces_7_3_io_ins_3 = ces_7_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_4_clock = clock;
  assign ces_7_4_io_ins_0 = ces_6_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_4_io_ins_1 = ces_7_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_4_io_ins_2 = io_insHorizontal_1_4; // @[MockArray.scala 46:87]
  assign ces_7_4_io_ins_3 = ces_7_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_5_clock = clock;
  assign ces_7_5_io_ins_0 = ces_6_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_5_io_ins_1 = ces_7_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_5_io_ins_2 = io_insHorizontal_1_5; // @[MockArray.scala 46:87]
  assign ces_7_5_io_ins_3 = ces_7_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_6_clock = clock;
  assign ces_7_6_io_ins_0 = ces_6_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_6_io_ins_1 = ces_7_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_6_io_ins_2 = io_insHorizontal_1_6; // @[MockArray.scala 46:87]
  assign ces_7_6_io_ins_3 = ces_7_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_7_clock = clock;
  assign ces_7_7_io_ins_0 = ces_6_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_7_io_ins_1 = ces_7_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_7_io_ins_2 = io_insHorizontal_1_7; // @[MockArray.scala 46:87]
  assign ces_7_7_io_ins_3 = ces_7_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_8_clock = clock;
  assign ces_7_8_io_ins_0 = ces_6_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_8_io_ins_1 = ces_7_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_8_io_ins_2 = io_insHorizontal_1_8; // @[MockArray.scala 46:87]
  assign ces_7_8_io_ins_3 = ces_7_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_9_clock = clock;
  assign ces_7_9_io_ins_0 = ces_6_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_9_io_ins_1 = ces_7_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_9_io_ins_2 = io_insHorizontal_1_9; // @[MockArray.scala 46:87]
  assign ces_7_9_io_ins_3 = ces_7_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_10_clock = clock;
  assign ces_7_10_io_ins_0 = ces_6_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_10_io_ins_1 = ces_7_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_10_io_ins_2 = io_insHorizontal_1_10; // @[MockArray.scala 46:87]
  assign ces_7_10_io_ins_3 = ces_7_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_11_clock = clock;
  assign ces_7_11_io_ins_0 = ces_6_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_11_io_ins_1 = ces_7_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_11_io_ins_2 = io_insHorizontal_1_11; // @[MockArray.scala 46:87]
  assign ces_7_11_io_ins_3 = ces_7_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_12_clock = clock;
  assign ces_7_12_io_ins_0 = ces_6_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_12_io_ins_1 = ces_7_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_12_io_ins_2 = io_insHorizontal_1_12; // @[MockArray.scala 46:87]
  assign ces_7_12_io_ins_3 = ces_7_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_13_clock = clock;
  assign ces_7_13_io_ins_0 = ces_6_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_13_io_ins_1 = ces_7_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_13_io_ins_2 = io_insHorizontal_1_13; // @[MockArray.scala 46:87]
  assign ces_7_13_io_ins_3 = ces_7_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_14_clock = clock;
  assign ces_7_14_io_ins_0 = ces_6_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_14_io_ins_1 = ces_7_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_14_io_ins_2 = io_insHorizontal_1_14; // @[MockArray.scala 46:87]
  assign ces_7_14_io_ins_3 = ces_7_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_15_clock = clock;
  assign ces_7_15_io_ins_0 = ces_6_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_15_io_ins_1 = io_insVertical_0_7; // @[MockArray.scala 45:87]
  assign ces_7_15_io_ins_2 = io_insHorizontal_1_15; // @[MockArray.scala 46:87]
  assign ces_7_15_io_ins_3 = ces_7_14_io_outs_1; // @[MockArray.scala 63:19]
endmodule
