module MuxTest_width_256_inputs_4_outputs_16_pipeline_5( // @[:@3.2]
  input          clock, // @[:@4.4]
  input          reset, // @[:@5.4]
  input  [1:0]   io_selects_0_0, // @[:@6.4]
  input  [1:0]   io_selects_0_1, // @[:@6.4]
  input  [1:0]   io_selects_1_0, // @[:@6.4]
  input  [1:0]   io_selects_1_1, // @[:@6.4]
  input  [1:0]   io_selects_2_0, // @[:@6.4]
  input  [1:0]   io_selects_2_1, // @[:@6.4]
  input  [1:0]   io_selects_3_0, // @[:@6.4]
  input  [1:0]   io_selects_3_1, // @[:@6.4]
  input  [1:0]   io_selects_4_0, // @[:@6.4]
  input  [1:0]   io_selects_4_1, // @[:@6.4]
  input  [1:0]   io_selects_5_0, // @[:@6.4]
  input  [1:0]   io_selects_5_1, // @[:@6.4]
  input  [1:0]   io_selects_6_0, // @[:@6.4]
  input  [1:0]   io_selects_6_1, // @[:@6.4]
  input  [1:0]   io_selects_7_0, // @[:@6.4]
  input  [1:0]   io_selects_7_1, // @[:@6.4]
  input  [1:0]   io_selects_8_0, // @[:@6.4]
  input  [1:0]   io_selects_8_1, // @[:@6.4]
  input  [1:0]   io_selects_9_0, // @[:@6.4]
  input  [1:0]   io_selects_9_1, // @[:@6.4]
  input  [1:0]   io_selects_10_0, // @[:@6.4]
  input  [1:0]   io_selects_10_1, // @[:@6.4]
  input  [1:0]   io_selects_11_0, // @[:@6.4]
  input  [1:0]   io_selects_11_1, // @[:@6.4]
  input  [1:0]   io_selects_12_0, // @[:@6.4]
  input  [1:0]   io_selects_12_1, // @[:@6.4]
  input  [1:0]   io_selects_13_0, // @[:@6.4]
  input  [1:0]   io_selects_13_1, // @[:@6.4]
  input  [1:0]   io_selects_14_0, // @[:@6.4]
  input  [1:0]   io_selects_14_1, // @[:@6.4]
  input  [1:0]   io_selects_15_0, // @[:@6.4]
  input  [1:0]   io_selects_15_1, // @[:@6.4]
  input  [2:0]   io_operation_0, // @[:@6.4]
  input  [2:0]   io_operation_1, // @[:@6.4]
  input  [2:0]   io_operation_2, // @[:@6.4]
  input  [2:0]   io_operation_3, // @[:@6.4]
  input  [2:0]   io_operation_4, // @[:@6.4]
  input  [2:0]   io_operation_5, // @[:@6.4]
  input  [2:0]   io_operation_6, // @[:@6.4]
  input  [2:0]   io_operation_7, // @[:@6.4]
  input  [2:0]   io_operation_8, // @[:@6.4]
  input  [2:0]   io_operation_9, // @[:@6.4]
  input  [2:0]   io_operation_10, // @[:@6.4]
  input  [2:0]   io_operation_11, // @[:@6.4]
  input  [2:0]   io_operation_12, // @[:@6.4]
  input  [2:0]   io_operation_13, // @[:@6.4]
  input  [2:0]   io_operation_14, // @[:@6.4]
  input  [2:0]   io_operation_15, // @[:@6.4]
  input  [255:0] io_inputs_0, // @[:@6.4]
  input  [255:0] io_inputs_1, // @[:@6.4]
  input  [255:0] io_inputs_2, // @[:@6.4]
  input  [255:0] io_inputs_3, // @[:@6.4]
  output [255:0] io_outputs_0, // @[:@6.4]
  output [255:0] io_outputs_1, // @[:@6.4]
  output [255:0] io_outputs_2, // @[:@6.4]
  output [255:0] io_outputs_3, // @[:@6.4]
  output [255:0] io_outputs_4, // @[:@6.4]
  output [255:0] io_outputs_5, // @[:@6.4]
  output [255:0] io_outputs_6, // @[:@6.4]
  output [255:0] io_outputs_7, // @[:@6.4]
  output [255:0] io_outputs_8, // @[:@6.4]
  output [255:0] io_outputs_9, // @[:@6.4]
  output [255:0] io_outputs_10, // @[:@6.4]
  output [255:0] io_outputs_11, // @[:@6.4]
  output [255:0] io_outputs_12, // @[:@6.4]
  output [255:0] io_outputs_13, // @[:@6.4]
  output [255:0] io_outputs_14, // @[:@6.4]
  output [255:0] io_outputs_15 // @[:@6.4]
);
  wire [255:0] _GEN_1; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [255:0] _GEN_2; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [255:0] _GEN_3; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [255:0] _GEN_5; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [255:0] _GEN_6; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [255:0] _GEN_7; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [256:0] _T_698; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [255:0] _T_699; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@9.4]
  wire [511:0] _T_701; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@10.4]
  wire [255:0] _T_703; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@11.4]
  wire  _T_704; // @[Mux.scala 46:19:@12.4]
  wire [255:0] _T_705; // @[Mux.scala 46:16:@13.4]
  wire  _T_706; // @[Mux.scala 46:19:@14.4]
  wire [511:0] _T_707; // @[Mux.scala 46:16:@15.4]
  wire  _T_708; // @[Mux.scala 46:19:@16.4]
  wire [511:0] _T_709; // @[Mux.scala 46:16:@17.4]
  wire  _T_710; // @[Mux.scala 46:19:@18.4]
  wire [255:0] _GEN_9; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [255:0] _GEN_10; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [255:0] _GEN_11; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [255:0] _GEN_13; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [255:0] _GEN_14; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [255:0] _GEN_15; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [256:0] _T_715; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@20.4]
  wire [255:0] _T_716; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@21.4]
  wire [511:0] _T_718; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@22.4]
  wire [255:0] _T_720; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@23.4]
  wire  _T_721; // @[Mux.scala 46:19:@24.4]
  wire [255:0] _T_722; // @[Mux.scala 46:16:@25.4]
  wire  _T_723; // @[Mux.scala 46:19:@26.4]
  wire [511:0] _T_724; // @[Mux.scala 46:16:@27.4]
  wire  _T_725; // @[Mux.scala 46:19:@28.4]
  wire [511:0] _T_726; // @[Mux.scala 46:16:@29.4]
  wire  _T_727; // @[Mux.scala 46:19:@30.4]
  wire [255:0] _GEN_17; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [255:0] _GEN_18; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [255:0] _GEN_19; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [255:0] _GEN_21; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [255:0] _GEN_22; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [255:0] _GEN_23; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [256:0] _T_732; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@32.4]
  wire [255:0] _T_733; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@33.4]
  wire [511:0] _T_735; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@34.4]
  wire [255:0] _T_737; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@35.4]
  wire  _T_738; // @[Mux.scala 46:19:@36.4]
  wire [255:0] _T_739; // @[Mux.scala 46:16:@37.4]
  wire  _T_740; // @[Mux.scala 46:19:@38.4]
  wire [511:0] _T_741; // @[Mux.scala 46:16:@39.4]
  wire  _T_742; // @[Mux.scala 46:19:@40.4]
  wire [511:0] _T_743; // @[Mux.scala 46:16:@41.4]
  wire  _T_744; // @[Mux.scala 46:19:@42.4]
  wire [255:0] _GEN_25; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [255:0] _GEN_26; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [255:0] _GEN_27; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [255:0] _GEN_29; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [255:0] _GEN_30; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [255:0] _GEN_31; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [256:0] _T_749; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@44.4]
  wire [255:0] _T_750; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@45.4]
  wire [511:0] _T_752; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@46.4]
  wire [255:0] _T_754; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@47.4]
  wire  _T_755; // @[Mux.scala 46:19:@48.4]
  wire [255:0] _T_756; // @[Mux.scala 46:16:@49.4]
  wire  _T_757; // @[Mux.scala 46:19:@50.4]
  wire [511:0] _T_758; // @[Mux.scala 46:16:@51.4]
  wire  _T_759; // @[Mux.scala 46:19:@52.4]
  wire [511:0] _T_760; // @[Mux.scala 46:16:@53.4]
  wire  _T_761; // @[Mux.scala 46:19:@54.4]
  wire [255:0] _GEN_33; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [255:0] _GEN_34; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [255:0] _GEN_35; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [255:0] _GEN_37; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [255:0] _GEN_38; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [255:0] _GEN_39; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [256:0] _T_766; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@56.4]
  wire [255:0] _T_767; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@57.4]
  wire [511:0] _T_769; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@58.4]
  wire [255:0] _T_771; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@59.4]
  wire  _T_772; // @[Mux.scala 46:19:@60.4]
  wire [255:0] _T_773; // @[Mux.scala 46:16:@61.4]
  wire  _T_774; // @[Mux.scala 46:19:@62.4]
  wire [511:0] _T_775; // @[Mux.scala 46:16:@63.4]
  wire  _T_776; // @[Mux.scala 46:19:@64.4]
  wire [511:0] _T_777; // @[Mux.scala 46:16:@65.4]
  wire  _T_778; // @[Mux.scala 46:19:@66.4]
  wire [255:0] _GEN_41; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [255:0] _GEN_42; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [255:0] _GEN_43; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [255:0] _GEN_45; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [255:0] _GEN_46; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [255:0] _GEN_47; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [256:0] _T_783; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@68.4]
  wire [255:0] _T_784; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@69.4]
  wire [511:0] _T_786; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@70.4]
  wire [255:0] _T_788; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@71.4]
  wire  _T_789; // @[Mux.scala 46:19:@72.4]
  wire [255:0] _T_790; // @[Mux.scala 46:16:@73.4]
  wire  _T_791; // @[Mux.scala 46:19:@74.4]
  wire [511:0] _T_792; // @[Mux.scala 46:16:@75.4]
  wire  _T_793; // @[Mux.scala 46:19:@76.4]
  wire [511:0] _T_794; // @[Mux.scala 46:16:@77.4]
  wire  _T_795; // @[Mux.scala 46:19:@78.4]
  wire [255:0] _GEN_49; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [255:0] _GEN_50; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [255:0] _GEN_51; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [255:0] _GEN_53; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [255:0] _GEN_54; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [255:0] _GEN_55; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [256:0] _T_800; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@80.4]
  wire [255:0] _T_801; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@81.4]
  wire [511:0] _T_803; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@82.4]
  wire [255:0] _T_805; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@83.4]
  wire  _T_806; // @[Mux.scala 46:19:@84.4]
  wire [255:0] _T_807; // @[Mux.scala 46:16:@85.4]
  wire  _T_808; // @[Mux.scala 46:19:@86.4]
  wire [511:0] _T_809; // @[Mux.scala 46:16:@87.4]
  wire  _T_810; // @[Mux.scala 46:19:@88.4]
  wire [511:0] _T_811; // @[Mux.scala 46:16:@89.4]
  wire  _T_812; // @[Mux.scala 46:19:@90.4]
  wire [255:0] _GEN_57; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [255:0] _GEN_58; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [255:0] _GEN_59; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [255:0] _GEN_61; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [255:0] _GEN_62; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [255:0] _GEN_63; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [256:0] _T_817; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@92.4]
  wire [255:0] _T_818; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@93.4]
  wire [511:0] _T_820; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@94.4]
  wire [255:0] _T_822; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@95.4]
  wire  _T_823; // @[Mux.scala 46:19:@96.4]
  wire [255:0] _T_824; // @[Mux.scala 46:16:@97.4]
  wire  _T_825; // @[Mux.scala 46:19:@98.4]
  wire [511:0] _T_826; // @[Mux.scala 46:16:@99.4]
  wire  _T_827; // @[Mux.scala 46:19:@100.4]
  wire [511:0] _T_828; // @[Mux.scala 46:16:@101.4]
  wire  _T_829; // @[Mux.scala 46:19:@102.4]
  wire [255:0] _GEN_65; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [255:0] _GEN_66; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [255:0] _GEN_67; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [255:0] _GEN_69; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [255:0] _GEN_70; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [255:0] _GEN_71; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [256:0] _T_834; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@104.4]
  wire [255:0] _T_835; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@105.4]
  wire [511:0] _T_837; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@106.4]
  wire [255:0] _T_839; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@107.4]
  wire  _T_840; // @[Mux.scala 46:19:@108.4]
  wire [255:0] _T_841; // @[Mux.scala 46:16:@109.4]
  wire  _T_842; // @[Mux.scala 46:19:@110.4]
  wire [511:0] _T_843; // @[Mux.scala 46:16:@111.4]
  wire  _T_844; // @[Mux.scala 46:19:@112.4]
  wire [511:0] _T_845; // @[Mux.scala 46:16:@113.4]
  wire  _T_846; // @[Mux.scala 46:19:@114.4]
  wire [255:0] _GEN_73; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [255:0] _GEN_74; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [255:0] _GEN_75; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [255:0] _GEN_77; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [255:0] _GEN_78; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [255:0] _GEN_79; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [256:0] _T_851; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@116.4]
  wire [255:0] _T_852; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@117.4]
  wire [511:0] _T_854; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@118.4]
  wire [255:0] _T_856; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@119.4]
  wire  _T_857; // @[Mux.scala 46:19:@120.4]
  wire [255:0] _T_858; // @[Mux.scala 46:16:@121.4]
  wire  _T_859; // @[Mux.scala 46:19:@122.4]
  wire [511:0] _T_860; // @[Mux.scala 46:16:@123.4]
  wire  _T_861; // @[Mux.scala 46:19:@124.4]
  wire [511:0] _T_862; // @[Mux.scala 46:16:@125.4]
  wire  _T_863; // @[Mux.scala 46:19:@126.4]
  wire [255:0] _GEN_81; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [255:0] _GEN_82; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [255:0] _GEN_83; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [255:0] _GEN_85; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [255:0] _GEN_86; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [255:0] _GEN_87; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [256:0] _T_868; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@128.4]
  wire [255:0] _T_869; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@129.4]
  wire [511:0] _T_871; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@130.4]
  wire [255:0] _T_873; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@131.4]
  wire  _T_874; // @[Mux.scala 46:19:@132.4]
  wire [255:0] _T_875; // @[Mux.scala 46:16:@133.4]
  wire  _T_876; // @[Mux.scala 46:19:@134.4]
  wire [511:0] _T_877; // @[Mux.scala 46:16:@135.4]
  wire  _T_878; // @[Mux.scala 46:19:@136.4]
  wire [511:0] _T_879; // @[Mux.scala 46:16:@137.4]
  wire  _T_880; // @[Mux.scala 46:19:@138.4]
  wire [255:0] _GEN_89; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [255:0] _GEN_90; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [255:0] _GEN_91; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [255:0] _GEN_93; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [255:0] _GEN_94; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [255:0] _GEN_95; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [256:0] _T_885; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@140.4]
  wire [255:0] _T_886; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@141.4]
  wire [511:0] _T_888; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@142.4]
  wire [255:0] _T_890; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@143.4]
  wire  _T_891; // @[Mux.scala 46:19:@144.4]
  wire [255:0] _T_892; // @[Mux.scala 46:16:@145.4]
  wire  _T_893; // @[Mux.scala 46:19:@146.4]
  wire [511:0] _T_894; // @[Mux.scala 46:16:@147.4]
  wire  _T_895; // @[Mux.scala 46:19:@148.4]
  wire [511:0] _T_896; // @[Mux.scala 46:16:@149.4]
  wire  _T_897; // @[Mux.scala 46:19:@150.4]
  wire [255:0] _GEN_97; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [255:0] _GEN_98; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [255:0] _GEN_99; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [255:0] _GEN_101; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [255:0] _GEN_102; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [255:0] _GEN_103; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [256:0] _T_902; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@152.4]
  wire [255:0] _T_903; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@153.4]
  wire [511:0] _T_905; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@154.4]
  wire [255:0] _T_907; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@155.4]
  wire  _T_908; // @[Mux.scala 46:19:@156.4]
  wire [255:0] _T_909; // @[Mux.scala 46:16:@157.4]
  wire  _T_910; // @[Mux.scala 46:19:@158.4]
  wire [511:0] _T_911; // @[Mux.scala 46:16:@159.4]
  wire  _T_912; // @[Mux.scala 46:19:@160.4]
  wire [511:0] _T_913; // @[Mux.scala 46:16:@161.4]
  wire  _T_914; // @[Mux.scala 46:19:@162.4]
  wire [255:0] _GEN_105; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [255:0] _GEN_106; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [255:0] _GEN_107; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [255:0] _GEN_109; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [255:0] _GEN_110; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [255:0] _GEN_111; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [256:0] _T_919; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@164.4]
  wire [255:0] _T_920; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@165.4]
  wire [511:0] _T_922; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@166.4]
  wire [255:0] _T_924; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@167.4]
  wire  _T_925; // @[Mux.scala 46:19:@168.4]
  wire [255:0] _T_926; // @[Mux.scala 46:16:@169.4]
  wire  _T_927; // @[Mux.scala 46:19:@170.4]
  wire [511:0] _T_928; // @[Mux.scala 46:16:@171.4]
  wire  _T_929; // @[Mux.scala 46:19:@172.4]
  wire [511:0] _T_930; // @[Mux.scala 46:16:@173.4]
  wire  _T_931; // @[Mux.scala 46:19:@174.4]
  wire [255:0] _GEN_113; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [255:0] _GEN_114; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [255:0] _GEN_115; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [255:0] _GEN_117; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [255:0] _GEN_118; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [255:0] _GEN_119; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [256:0] _T_936; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@176.4]
  wire [255:0] _T_937; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@177.4]
  wire [511:0] _T_939; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@178.4]
  wire [255:0] _T_941; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@179.4]
  wire  _T_942; // @[Mux.scala 46:19:@180.4]
  wire [255:0] _T_943; // @[Mux.scala 46:16:@181.4]
  wire  _T_944; // @[Mux.scala 46:19:@182.4]
  wire [511:0] _T_945; // @[Mux.scala 46:16:@183.4]
  wire  _T_946; // @[Mux.scala 46:19:@184.4]
  wire [511:0] _T_947; // @[Mux.scala 46:16:@185.4]
  wire  _T_948; // @[Mux.scala 46:19:@186.4]
  wire [255:0] _GEN_121; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [255:0] _GEN_122; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [255:0] _GEN_123; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [255:0] _GEN_125; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [255:0] _GEN_126; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [255:0] _GEN_127; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [256:0] _T_953; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@188.4]
  wire [255:0] _T_954; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@189.4]
  wire [511:0] _T_956; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@190.4]
  wire [255:0] _T_958; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@191.4]
  wire  _T_959; // @[Mux.scala 46:19:@192.4]
  wire [255:0] _T_960; // @[Mux.scala 46:16:@193.4]
  wire  _T_961; // @[Mux.scala 46:19:@194.4]
  wire [511:0] _T_962; // @[Mux.scala 46:16:@195.4]
  wire  _T_963; // @[Mux.scala 46:19:@196.4]
  wire [511:0] _T_964; // @[Mux.scala 46:16:@197.4]
  wire  _T_965; // @[Mux.scala 46:19:@198.4]
  reg [511:0] _T_969; // @[Reg.scala 11:16:@200.4]
  reg [511:0] _RAND_0;
  reg [511:0] _T_971; // @[Reg.scala 11:16:@204.4]
  reg [511:0] _RAND_1;
  reg [511:0] _T_973; // @[Reg.scala 11:16:@208.4]
  reg [511:0] _RAND_2;
  reg [511:0] _T_975; // @[Reg.scala 11:16:@212.4]
  reg [511:0] _RAND_3;
  reg [511:0] _T_977; // @[Reg.scala 11:16:@216.4]
  reg [511:0] _RAND_4;
  reg [511:0] _T_980; // @[Reg.scala 11:16:@220.4]
  reg [511:0] _RAND_5;
  reg [511:0] _T_982; // @[Reg.scala 11:16:@224.4]
  reg [511:0] _RAND_6;
  reg [511:0] _T_984; // @[Reg.scala 11:16:@228.4]
  reg [511:0] _RAND_7;
  reg [511:0] _T_986; // @[Reg.scala 11:16:@232.4]
  reg [511:0] _RAND_8;
  reg [511:0] _T_988; // @[Reg.scala 11:16:@236.4]
  reg [511:0] _RAND_9;
  reg [511:0] _T_991; // @[Reg.scala 11:16:@240.4]
  reg [511:0] _RAND_10;
  reg [511:0] _T_993; // @[Reg.scala 11:16:@244.4]
  reg [511:0] _RAND_11;
  reg [511:0] _T_995; // @[Reg.scala 11:16:@248.4]
  reg [511:0] _RAND_12;
  reg [511:0] _T_997; // @[Reg.scala 11:16:@252.4]
  reg [511:0] _RAND_13;
  reg [511:0] _T_999; // @[Reg.scala 11:16:@256.4]
  reg [511:0] _RAND_14;
  reg [511:0] _T_1002; // @[Reg.scala 11:16:@260.4]
  reg [511:0] _RAND_15;
  reg [511:0] _T_1004; // @[Reg.scala 11:16:@264.4]
  reg [511:0] _RAND_16;
  reg [511:0] _T_1006; // @[Reg.scala 11:16:@268.4]
  reg [511:0] _RAND_17;
  reg [511:0] _T_1008; // @[Reg.scala 11:16:@272.4]
  reg [511:0] _RAND_18;
  reg [511:0] _T_1010; // @[Reg.scala 11:16:@276.4]
  reg [511:0] _RAND_19;
  reg [511:0] _T_1013; // @[Reg.scala 11:16:@280.4]
  reg [511:0] _RAND_20;
  reg [511:0] _T_1015; // @[Reg.scala 11:16:@284.4]
  reg [511:0] _RAND_21;
  reg [511:0] _T_1017; // @[Reg.scala 11:16:@288.4]
  reg [511:0] _RAND_22;
  reg [511:0] _T_1019; // @[Reg.scala 11:16:@292.4]
  reg [511:0] _RAND_23;
  reg [511:0] _T_1021; // @[Reg.scala 11:16:@296.4]
  reg [511:0] _RAND_24;
  reg [511:0] _T_1024; // @[Reg.scala 11:16:@300.4]
  reg [511:0] _RAND_25;
  reg [511:0] _T_1026; // @[Reg.scala 11:16:@304.4]
  reg [511:0] _RAND_26;
  reg [511:0] _T_1028; // @[Reg.scala 11:16:@308.4]
  reg [511:0] _RAND_27;
  reg [511:0] _T_1030; // @[Reg.scala 11:16:@312.4]
  reg [511:0] _RAND_28;
  reg [511:0] _T_1032; // @[Reg.scala 11:16:@316.4]
  reg [511:0] _RAND_29;
  reg [511:0] _T_1035; // @[Reg.scala 11:16:@320.4]
  reg [511:0] _RAND_30;
  reg [511:0] _T_1037; // @[Reg.scala 11:16:@324.4]
  reg [511:0] _RAND_31;
  reg [511:0] _T_1039; // @[Reg.scala 11:16:@328.4]
  reg [511:0] _RAND_32;
  reg [511:0] _T_1041; // @[Reg.scala 11:16:@332.4]
  reg [511:0] _RAND_33;
  reg [511:0] _T_1043; // @[Reg.scala 11:16:@336.4]
  reg [511:0] _RAND_34;
  reg [511:0] _T_1046; // @[Reg.scala 11:16:@340.4]
  reg [511:0] _RAND_35;
  reg [511:0] _T_1048; // @[Reg.scala 11:16:@344.4]
  reg [511:0] _RAND_36;
  reg [511:0] _T_1050; // @[Reg.scala 11:16:@348.4]
  reg [511:0] _RAND_37;
  reg [511:0] _T_1052; // @[Reg.scala 11:16:@352.4]
  reg [511:0] _RAND_38;
  reg [511:0] _T_1054; // @[Reg.scala 11:16:@356.4]
  reg [511:0] _RAND_39;
  reg [511:0] _T_1057; // @[Reg.scala 11:16:@360.4]
  reg [511:0] _RAND_40;
  reg [511:0] _T_1059; // @[Reg.scala 11:16:@364.4]
  reg [511:0] _RAND_41;
  reg [511:0] _T_1061; // @[Reg.scala 11:16:@368.4]
  reg [511:0] _RAND_42;
  reg [511:0] _T_1063; // @[Reg.scala 11:16:@372.4]
  reg [511:0] _RAND_43;
  reg [511:0] _T_1065; // @[Reg.scala 11:16:@376.4]
  reg [511:0] _RAND_44;
  reg [511:0] _T_1068; // @[Reg.scala 11:16:@380.4]
  reg [511:0] _RAND_45;
  reg [511:0] _T_1070; // @[Reg.scala 11:16:@384.4]
  reg [511:0] _RAND_46;
  reg [511:0] _T_1072; // @[Reg.scala 11:16:@388.4]
  reg [511:0] _RAND_47;
  reg [511:0] _T_1074; // @[Reg.scala 11:16:@392.4]
  reg [511:0] _RAND_48;
  reg [511:0] _T_1076; // @[Reg.scala 11:16:@396.4]
  reg [511:0] _RAND_49;
  reg [511:0] _T_1079; // @[Reg.scala 11:16:@400.4]
  reg [511:0] _RAND_50;
  reg [511:0] _T_1081; // @[Reg.scala 11:16:@404.4]
  reg [511:0] _RAND_51;
  reg [511:0] _T_1083; // @[Reg.scala 11:16:@408.4]
  reg [511:0] _RAND_52;
  reg [511:0] _T_1085; // @[Reg.scala 11:16:@412.4]
  reg [511:0] _RAND_53;
  reg [511:0] _T_1087; // @[Reg.scala 11:16:@416.4]
  reg [511:0] _RAND_54;
  reg [511:0] _T_1090; // @[Reg.scala 11:16:@420.4]
  reg [511:0] _RAND_55;
  reg [511:0] _T_1092; // @[Reg.scala 11:16:@424.4]
  reg [511:0] _RAND_56;
  reg [511:0] _T_1094; // @[Reg.scala 11:16:@428.4]
  reg [511:0] _RAND_57;
  reg [511:0] _T_1096; // @[Reg.scala 11:16:@432.4]
  reg [511:0] _RAND_58;
  reg [511:0] _T_1098; // @[Reg.scala 11:16:@436.4]
  reg [511:0] _RAND_59;
  reg [511:0] _T_1101; // @[Reg.scala 11:16:@440.4]
  reg [511:0] _RAND_60;
  reg [511:0] _T_1103; // @[Reg.scala 11:16:@444.4]
  reg [511:0] _RAND_61;
  reg [511:0] _T_1105; // @[Reg.scala 11:16:@448.4]
  reg [511:0] _RAND_62;
  reg [511:0] _T_1107; // @[Reg.scala 11:16:@452.4]
  reg [511:0] _RAND_63;
  reg [511:0] _T_1109; // @[Reg.scala 11:16:@456.4]
  reg [511:0] _RAND_64;
  reg [511:0] _T_1112; // @[Reg.scala 11:16:@460.4]
  reg [511:0] _RAND_65;
  reg [511:0] _T_1114; // @[Reg.scala 11:16:@464.4]
  reg [511:0] _RAND_66;
  reg [511:0] _T_1116; // @[Reg.scala 11:16:@468.4]
  reg [511:0] _RAND_67;
  reg [511:0] _T_1118; // @[Reg.scala 11:16:@472.4]
  reg [511:0] _RAND_68;
  reg [511:0] _T_1120; // @[Reg.scala 11:16:@476.4]
  reg [511:0] _RAND_69;
  reg [511:0] _T_1123; // @[Reg.scala 11:16:@480.4]
  reg [511:0] _RAND_70;
  reg [511:0] _T_1125; // @[Reg.scala 11:16:@484.4]
  reg [511:0] _RAND_71;
  reg [511:0] _T_1127; // @[Reg.scala 11:16:@488.4]
  reg [511:0] _RAND_72;
  reg [511:0] _T_1129; // @[Reg.scala 11:16:@492.4]
  reg [511:0] _RAND_73;
  reg [511:0] _T_1131; // @[Reg.scala 11:16:@496.4]
  reg [511:0] _RAND_74;
  reg [511:0] _T_1134; // @[Reg.scala 11:16:@500.4]
  reg [511:0] _RAND_75;
  reg [511:0] _T_1136; // @[Reg.scala 11:16:@504.4]
  reg [511:0] _RAND_76;
  reg [511:0] _T_1138; // @[Reg.scala 11:16:@508.4]
  reg [511:0] _RAND_77;
  reg [511:0] _T_1140; // @[Reg.scala 11:16:@512.4]
  reg [511:0] _RAND_78;
  reg [511:0] _T_1142; // @[Reg.scala 11:16:@516.4]
  reg [511:0] _RAND_79;
  assign _GEN_1 = 2'h1 == io_selects_0_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_2 = 2'h2 == io_selects_0_0 ? io_inputs_2 : _GEN_1; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_3 = 2'h3 == io_selects_0_0 ? io_inputs_3 : _GEN_2; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_5 = 2'h1 == io_selects_0_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_6 = 2'h2 == io_selects_0_1 ? io_inputs_2 : _GEN_5; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_7 = 2'h3 == io_selects_0_1 ? io_inputs_3 : _GEN_6; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _T_698 = _GEN_3 + _GEN_7; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _T_699 = _GEN_3 + _GEN_7; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@9.4]
  assign _T_701 = _GEN_3 * _GEN_7; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@10.4]
  assign _T_703 = _GEN_3 / _GEN_7; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@11.4]
  assign _T_704 = 3'h3 == io_operation_0; // @[Mux.scala 46:19:@12.4]
  assign _T_705 = _T_704 ? _T_703 : 256'h0; // @[Mux.scala 46:16:@13.4]
  assign _T_706 = 3'h2 == io_operation_0; // @[Mux.scala 46:19:@14.4]
  assign _T_707 = _T_706 ? _T_701 : {{256'd0}, _T_705}; // @[Mux.scala 46:16:@15.4]
  assign _T_708 = 3'h1 == io_operation_0; // @[Mux.scala 46:19:@16.4]
  assign _T_709 = _T_708 ? {{256'd0}, _T_699} : _T_707; // @[Mux.scala 46:16:@17.4]
  assign _T_710 = 3'h0 == io_operation_0; // @[Mux.scala 46:19:@18.4]
  assign _GEN_9 = 2'h1 == io_selects_1_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_10 = 2'h2 == io_selects_1_0 ? io_inputs_2 : _GEN_9; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_11 = 2'h3 == io_selects_1_0 ? io_inputs_3 : _GEN_10; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_13 = 2'h1 == io_selects_1_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_14 = 2'h2 == io_selects_1_1 ? io_inputs_2 : _GEN_13; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_15 = 2'h3 == io_selects_1_1 ? io_inputs_3 : _GEN_14; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _T_715 = _GEN_11 + _GEN_15; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@20.4]
  assign _T_716 = _GEN_11 + _GEN_15; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@21.4]
  assign _T_718 = _GEN_11 * _GEN_15; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@22.4]
  assign _T_720 = _GEN_11 / _GEN_15; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@23.4]
  assign _T_721 = 3'h3 == io_operation_1; // @[Mux.scala 46:19:@24.4]
  assign _T_722 = _T_721 ? _T_720 : 256'h0; // @[Mux.scala 46:16:@25.4]
  assign _T_723 = 3'h2 == io_operation_1; // @[Mux.scala 46:19:@26.4]
  assign _T_724 = _T_723 ? _T_718 : {{256'd0}, _T_722}; // @[Mux.scala 46:16:@27.4]
  assign _T_725 = 3'h1 == io_operation_1; // @[Mux.scala 46:19:@28.4]
  assign _T_726 = _T_725 ? {{256'd0}, _T_716} : _T_724; // @[Mux.scala 46:16:@29.4]
  assign _T_727 = 3'h0 == io_operation_1; // @[Mux.scala 46:19:@30.4]
  assign _GEN_17 = 2'h1 == io_selects_2_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_18 = 2'h2 == io_selects_2_0 ? io_inputs_2 : _GEN_17; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_19 = 2'h3 == io_selects_2_0 ? io_inputs_3 : _GEN_18; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_21 = 2'h1 == io_selects_2_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_22 = 2'h2 == io_selects_2_1 ? io_inputs_2 : _GEN_21; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_23 = 2'h3 == io_selects_2_1 ? io_inputs_3 : _GEN_22; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _T_732 = _GEN_19 + _GEN_23; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@32.4]
  assign _T_733 = _GEN_19 + _GEN_23; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@33.4]
  assign _T_735 = _GEN_19 * _GEN_23; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@34.4]
  assign _T_737 = _GEN_19 / _GEN_23; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@35.4]
  assign _T_738 = 3'h3 == io_operation_2; // @[Mux.scala 46:19:@36.4]
  assign _T_739 = _T_738 ? _T_737 : 256'h0; // @[Mux.scala 46:16:@37.4]
  assign _T_740 = 3'h2 == io_operation_2; // @[Mux.scala 46:19:@38.4]
  assign _T_741 = _T_740 ? _T_735 : {{256'd0}, _T_739}; // @[Mux.scala 46:16:@39.4]
  assign _T_742 = 3'h1 == io_operation_2; // @[Mux.scala 46:19:@40.4]
  assign _T_743 = _T_742 ? {{256'd0}, _T_733} : _T_741; // @[Mux.scala 46:16:@41.4]
  assign _T_744 = 3'h0 == io_operation_2; // @[Mux.scala 46:19:@42.4]
  assign _GEN_25 = 2'h1 == io_selects_3_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_26 = 2'h2 == io_selects_3_0 ? io_inputs_2 : _GEN_25; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_27 = 2'h3 == io_selects_3_0 ? io_inputs_3 : _GEN_26; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_29 = 2'h1 == io_selects_3_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_30 = 2'h2 == io_selects_3_1 ? io_inputs_2 : _GEN_29; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_31 = 2'h3 == io_selects_3_1 ? io_inputs_3 : _GEN_30; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _T_749 = _GEN_27 + _GEN_31; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@44.4]
  assign _T_750 = _GEN_27 + _GEN_31; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@45.4]
  assign _T_752 = _GEN_27 * _GEN_31; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@46.4]
  assign _T_754 = _GEN_27 / _GEN_31; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@47.4]
  assign _T_755 = 3'h3 == io_operation_3; // @[Mux.scala 46:19:@48.4]
  assign _T_756 = _T_755 ? _T_754 : 256'h0; // @[Mux.scala 46:16:@49.4]
  assign _T_757 = 3'h2 == io_operation_3; // @[Mux.scala 46:19:@50.4]
  assign _T_758 = _T_757 ? _T_752 : {{256'd0}, _T_756}; // @[Mux.scala 46:16:@51.4]
  assign _T_759 = 3'h1 == io_operation_3; // @[Mux.scala 46:19:@52.4]
  assign _T_760 = _T_759 ? {{256'd0}, _T_750} : _T_758; // @[Mux.scala 46:16:@53.4]
  assign _T_761 = 3'h0 == io_operation_3; // @[Mux.scala 46:19:@54.4]
  assign _GEN_33 = 2'h1 == io_selects_4_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_34 = 2'h2 == io_selects_4_0 ? io_inputs_2 : _GEN_33; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_35 = 2'h3 == io_selects_4_0 ? io_inputs_3 : _GEN_34; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_37 = 2'h1 == io_selects_4_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_38 = 2'h2 == io_selects_4_1 ? io_inputs_2 : _GEN_37; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_39 = 2'h3 == io_selects_4_1 ? io_inputs_3 : _GEN_38; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _T_766 = _GEN_35 + _GEN_39; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@56.4]
  assign _T_767 = _GEN_35 + _GEN_39; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@57.4]
  assign _T_769 = _GEN_35 * _GEN_39; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@58.4]
  assign _T_771 = _GEN_35 / _GEN_39; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@59.4]
  assign _T_772 = 3'h3 == io_operation_4; // @[Mux.scala 46:19:@60.4]
  assign _T_773 = _T_772 ? _T_771 : 256'h0; // @[Mux.scala 46:16:@61.4]
  assign _T_774 = 3'h2 == io_operation_4; // @[Mux.scala 46:19:@62.4]
  assign _T_775 = _T_774 ? _T_769 : {{256'd0}, _T_773}; // @[Mux.scala 46:16:@63.4]
  assign _T_776 = 3'h1 == io_operation_4; // @[Mux.scala 46:19:@64.4]
  assign _T_777 = _T_776 ? {{256'd0}, _T_767} : _T_775; // @[Mux.scala 46:16:@65.4]
  assign _T_778 = 3'h0 == io_operation_4; // @[Mux.scala 46:19:@66.4]
  assign _GEN_41 = 2'h1 == io_selects_5_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_42 = 2'h2 == io_selects_5_0 ? io_inputs_2 : _GEN_41; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_43 = 2'h3 == io_selects_5_0 ? io_inputs_3 : _GEN_42; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_45 = 2'h1 == io_selects_5_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_46 = 2'h2 == io_selects_5_1 ? io_inputs_2 : _GEN_45; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_47 = 2'h3 == io_selects_5_1 ? io_inputs_3 : _GEN_46; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _T_783 = _GEN_43 + _GEN_47; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@68.4]
  assign _T_784 = _GEN_43 + _GEN_47; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@69.4]
  assign _T_786 = _GEN_43 * _GEN_47; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@70.4]
  assign _T_788 = _GEN_43 / _GEN_47; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@71.4]
  assign _T_789 = 3'h3 == io_operation_5; // @[Mux.scala 46:19:@72.4]
  assign _T_790 = _T_789 ? _T_788 : 256'h0; // @[Mux.scala 46:16:@73.4]
  assign _T_791 = 3'h2 == io_operation_5; // @[Mux.scala 46:19:@74.4]
  assign _T_792 = _T_791 ? _T_786 : {{256'd0}, _T_790}; // @[Mux.scala 46:16:@75.4]
  assign _T_793 = 3'h1 == io_operation_5; // @[Mux.scala 46:19:@76.4]
  assign _T_794 = _T_793 ? {{256'd0}, _T_784} : _T_792; // @[Mux.scala 46:16:@77.4]
  assign _T_795 = 3'h0 == io_operation_5; // @[Mux.scala 46:19:@78.4]
  assign _GEN_49 = 2'h1 == io_selects_6_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_50 = 2'h2 == io_selects_6_0 ? io_inputs_2 : _GEN_49; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_51 = 2'h3 == io_selects_6_0 ? io_inputs_3 : _GEN_50; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_53 = 2'h1 == io_selects_6_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_54 = 2'h2 == io_selects_6_1 ? io_inputs_2 : _GEN_53; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_55 = 2'h3 == io_selects_6_1 ? io_inputs_3 : _GEN_54; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _T_800 = _GEN_51 + _GEN_55; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@80.4]
  assign _T_801 = _GEN_51 + _GEN_55; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@81.4]
  assign _T_803 = _GEN_51 * _GEN_55; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@82.4]
  assign _T_805 = _GEN_51 / _GEN_55; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@83.4]
  assign _T_806 = 3'h3 == io_operation_6; // @[Mux.scala 46:19:@84.4]
  assign _T_807 = _T_806 ? _T_805 : 256'h0; // @[Mux.scala 46:16:@85.4]
  assign _T_808 = 3'h2 == io_operation_6; // @[Mux.scala 46:19:@86.4]
  assign _T_809 = _T_808 ? _T_803 : {{256'd0}, _T_807}; // @[Mux.scala 46:16:@87.4]
  assign _T_810 = 3'h1 == io_operation_6; // @[Mux.scala 46:19:@88.4]
  assign _T_811 = _T_810 ? {{256'd0}, _T_801} : _T_809; // @[Mux.scala 46:16:@89.4]
  assign _T_812 = 3'h0 == io_operation_6; // @[Mux.scala 46:19:@90.4]
  assign _GEN_57 = 2'h1 == io_selects_7_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_58 = 2'h2 == io_selects_7_0 ? io_inputs_2 : _GEN_57; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_59 = 2'h3 == io_selects_7_0 ? io_inputs_3 : _GEN_58; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_61 = 2'h1 == io_selects_7_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_62 = 2'h2 == io_selects_7_1 ? io_inputs_2 : _GEN_61; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_63 = 2'h3 == io_selects_7_1 ? io_inputs_3 : _GEN_62; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _T_817 = _GEN_59 + _GEN_63; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@92.4]
  assign _T_818 = _GEN_59 + _GEN_63; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@93.4]
  assign _T_820 = _GEN_59 * _GEN_63; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@94.4]
  assign _T_822 = _GEN_59 / _GEN_63; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@95.4]
  assign _T_823 = 3'h3 == io_operation_7; // @[Mux.scala 46:19:@96.4]
  assign _T_824 = _T_823 ? _T_822 : 256'h0; // @[Mux.scala 46:16:@97.4]
  assign _T_825 = 3'h2 == io_operation_7; // @[Mux.scala 46:19:@98.4]
  assign _T_826 = _T_825 ? _T_820 : {{256'd0}, _T_824}; // @[Mux.scala 46:16:@99.4]
  assign _T_827 = 3'h1 == io_operation_7; // @[Mux.scala 46:19:@100.4]
  assign _T_828 = _T_827 ? {{256'd0}, _T_818} : _T_826; // @[Mux.scala 46:16:@101.4]
  assign _T_829 = 3'h0 == io_operation_7; // @[Mux.scala 46:19:@102.4]
  assign _GEN_65 = 2'h1 == io_selects_8_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_66 = 2'h2 == io_selects_8_0 ? io_inputs_2 : _GEN_65; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_67 = 2'h3 == io_selects_8_0 ? io_inputs_3 : _GEN_66; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_69 = 2'h1 == io_selects_8_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_70 = 2'h2 == io_selects_8_1 ? io_inputs_2 : _GEN_69; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _GEN_71 = 2'h3 == io_selects_8_1 ? io_inputs_3 : _GEN_70; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _T_834 = _GEN_67 + _GEN_71; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@104.4]
  assign _T_835 = _GEN_67 + _GEN_71; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@105.4]
  assign _T_837 = _GEN_67 * _GEN_71; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@106.4]
  assign _T_839 = _GEN_67 / _GEN_71; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@107.4]
  assign _T_840 = 3'h3 == io_operation_8; // @[Mux.scala 46:19:@108.4]
  assign _T_841 = _T_840 ? _T_839 : 256'h0; // @[Mux.scala 46:16:@109.4]
  assign _T_842 = 3'h2 == io_operation_8; // @[Mux.scala 46:19:@110.4]
  assign _T_843 = _T_842 ? _T_837 : {{256'd0}, _T_841}; // @[Mux.scala 46:16:@111.4]
  assign _T_844 = 3'h1 == io_operation_8; // @[Mux.scala 46:19:@112.4]
  assign _T_845 = _T_844 ? {{256'd0}, _T_835} : _T_843; // @[Mux.scala 46:16:@113.4]
  assign _T_846 = 3'h0 == io_operation_8; // @[Mux.scala 46:19:@114.4]
  assign _GEN_73 = 2'h1 == io_selects_9_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_74 = 2'h2 == io_selects_9_0 ? io_inputs_2 : _GEN_73; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_75 = 2'h3 == io_selects_9_0 ? io_inputs_3 : _GEN_74; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_77 = 2'h1 == io_selects_9_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_78 = 2'h2 == io_selects_9_1 ? io_inputs_2 : _GEN_77; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _GEN_79 = 2'h3 == io_selects_9_1 ? io_inputs_3 : _GEN_78; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _T_851 = _GEN_75 + _GEN_79; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@116.4]
  assign _T_852 = _GEN_75 + _GEN_79; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@117.4]
  assign _T_854 = _GEN_75 * _GEN_79; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@118.4]
  assign _T_856 = _GEN_75 / _GEN_79; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@119.4]
  assign _T_857 = 3'h3 == io_operation_9; // @[Mux.scala 46:19:@120.4]
  assign _T_858 = _T_857 ? _T_856 : 256'h0; // @[Mux.scala 46:16:@121.4]
  assign _T_859 = 3'h2 == io_operation_9; // @[Mux.scala 46:19:@122.4]
  assign _T_860 = _T_859 ? _T_854 : {{256'd0}, _T_858}; // @[Mux.scala 46:16:@123.4]
  assign _T_861 = 3'h1 == io_operation_9; // @[Mux.scala 46:19:@124.4]
  assign _T_862 = _T_861 ? {{256'd0}, _T_852} : _T_860; // @[Mux.scala 46:16:@125.4]
  assign _T_863 = 3'h0 == io_operation_9; // @[Mux.scala 46:19:@126.4]
  assign _GEN_81 = 2'h1 == io_selects_10_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_82 = 2'h2 == io_selects_10_0 ? io_inputs_2 : _GEN_81; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_83 = 2'h3 == io_selects_10_0 ? io_inputs_3 : _GEN_82; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_85 = 2'h1 == io_selects_10_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_86 = 2'h2 == io_selects_10_1 ? io_inputs_2 : _GEN_85; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _GEN_87 = 2'h3 == io_selects_10_1 ? io_inputs_3 : _GEN_86; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _T_868 = _GEN_83 + _GEN_87; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@128.4]
  assign _T_869 = _GEN_83 + _GEN_87; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@129.4]
  assign _T_871 = _GEN_83 * _GEN_87; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@130.4]
  assign _T_873 = _GEN_83 / _GEN_87; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@131.4]
  assign _T_874 = 3'h3 == io_operation_10; // @[Mux.scala 46:19:@132.4]
  assign _T_875 = _T_874 ? _T_873 : 256'h0; // @[Mux.scala 46:16:@133.4]
  assign _T_876 = 3'h2 == io_operation_10; // @[Mux.scala 46:19:@134.4]
  assign _T_877 = _T_876 ? _T_871 : {{256'd0}, _T_875}; // @[Mux.scala 46:16:@135.4]
  assign _T_878 = 3'h1 == io_operation_10; // @[Mux.scala 46:19:@136.4]
  assign _T_879 = _T_878 ? {{256'd0}, _T_869} : _T_877; // @[Mux.scala 46:16:@137.4]
  assign _T_880 = 3'h0 == io_operation_10; // @[Mux.scala 46:19:@138.4]
  assign _GEN_89 = 2'h1 == io_selects_11_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_90 = 2'h2 == io_selects_11_0 ? io_inputs_2 : _GEN_89; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_91 = 2'h3 == io_selects_11_0 ? io_inputs_3 : _GEN_90; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_93 = 2'h1 == io_selects_11_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_94 = 2'h2 == io_selects_11_1 ? io_inputs_2 : _GEN_93; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _GEN_95 = 2'h3 == io_selects_11_1 ? io_inputs_3 : _GEN_94; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _T_885 = _GEN_91 + _GEN_95; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@140.4]
  assign _T_886 = _GEN_91 + _GEN_95; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@141.4]
  assign _T_888 = _GEN_91 * _GEN_95; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@142.4]
  assign _T_890 = _GEN_91 / _GEN_95; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@143.4]
  assign _T_891 = 3'h3 == io_operation_11; // @[Mux.scala 46:19:@144.4]
  assign _T_892 = _T_891 ? _T_890 : 256'h0; // @[Mux.scala 46:16:@145.4]
  assign _T_893 = 3'h2 == io_operation_11; // @[Mux.scala 46:19:@146.4]
  assign _T_894 = _T_893 ? _T_888 : {{256'd0}, _T_892}; // @[Mux.scala 46:16:@147.4]
  assign _T_895 = 3'h1 == io_operation_11; // @[Mux.scala 46:19:@148.4]
  assign _T_896 = _T_895 ? {{256'd0}, _T_886} : _T_894; // @[Mux.scala 46:16:@149.4]
  assign _T_897 = 3'h0 == io_operation_11; // @[Mux.scala 46:19:@150.4]
  assign _GEN_97 = 2'h1 == io_selects_12_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_98 = 2'h2 == io_selects_12_0 ? io_inputs_2 : _GEN_97; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_99 = 2'h3 == io_selects_12_0 ? io_inputs_3 : _GEN_98; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_101 = 2'h1 == io_selects_12_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_102 = 2'h2 == io_selects_12_1 ? io_inputs_2 : _GEN_101; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _GEN_103 = 2'h3 == io_selects_12_1 ? io_inputs_3 : _GEN_102; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _T_902 = _GEN_99 + _GEN_103; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@152.4]
  assign _T_903 = _GEN_99 + _GEN_103; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@153.4]
  assign _T_905 = _GEN_99 * _GEN_103; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@154.4]
  assign _T_907 = _GEN_99 / _GEN_103; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@155.4]
  assign _T_908 = 3'h3 == io_operation_12; // @[Mux.scala 46:19:@156.4]
  assign _T_909 = _T_908 ? _T_907 : 256'h0; // @[Mux.scala 46:16:@157.4]
  assign _T_910 = 3'h2 == io_operation_12; // @[Mux.scala 46:19:@158.4]
  assign _T_911 = _T_910 ? _T_905 : {{256'd0}, _T_909}; // @[Mux.scala 46:16:@159.4]
  assign _T_912 = 3'h1 == io_operation_12; // @[Mux.scala 46:19:@160.4]
  assign _T_913 = _T_912 ? {{256'd0}, _T_903} : _T_911; // @[Mux.scala 46:16:@161.4]
  assign _T_914 = 3'h0 == io_operation_12; // @[Mux.scala 46:19:@162.4]
  assign _GEN_105 = 2'h1 == io_selects_13_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_106 = 2'h2 == io_selects_13_0 ? io_inputs_2 : _GEN_105; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_107 = 2'h3 == io_selects_13_0 ? io_inputs_3 : _GEN_106; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_109 = 2'h1 == io_selects_13_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_110 = 2'h2 == io_selects_13_1 ? io_inputs_2 : _GEN_109; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _GEN_111 = 2'h3 == io_selects_13_1 ? io_inputs_3 : _GEN_110; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _T_919 = _GEN_107 + _GEN_111; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@164.4]
  assign _T_920 = _GEN_107 + _GEN_111; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@165.4]
  assign _T_922 = _GEN_107 * _GEN_111; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@166.4]
  assign _T_924 = _GEN_107 / _GEN_111; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@167.4]
  assign _T_925 = 3'h3 == io_operation_13; // @[Mux.scala 46:19:@168.4]
  assign _T_926 = _T_925 ? _T_924 : 256'h0; // @[Mux.scala 46:16:@169.4]
  assign _T_927 = 3'h2 == io_operation_13; // @[Mux.scala 46:19:@170.4]
  assign _T_928 = _T_927 ? _T_922 : {{256'd0}, _T_926}; // @[Mux.scala 46:16:@171.4]
  assign _T_929 = 3'h1 == io_operation_13; // @[Mux.scala 46:19:@172.4]
  assign _T_930 = _T_929 ? {{256'd0}, _T_920} : _T_928; // @[Mux.scala 46:16:@173.4]
  assign _T_931 = 3'h0 == io_operation_13; // @[Mux.scala 46:19:@174.4]
  assign _GEN_113 = 2'h1 == io_selects_14_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_114 = 2'h2 == io_selects_14_0 ? io_inputs_2 : _GEN_113; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_115 = 2'h3 == io_selects_14_0 ? io_inputs_3 : _GEN_114; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_117 = 2'h1 == io_selects_14_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_118 = 2'h2 == io_selects_14_1 ? io_inputs_2 : _GEN_117; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _GEN_119 = 2'h3 == io_selects_14_1 ? io_inputs_3 : _GEN_118; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _T_936 = _GEN_115 + _GEN_119; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@176.4]
  assign _T_937 = _GEN_115 + _GEN_119; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@177.4]
  assign _T_939 = _GEN_115 * _GEN_119; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@178.4]
  assign _T_941 = _GEN_115 / _GEN_119; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@179.4]
  assign _T_942 = 3'h3 == io_operation_14; // @[Mux.scala 46:19:@180.4]
  assign _T_943 = _T_942 ? _T_941 : 256'h0; // @[Mux.scala 46:16:@181.4]
  assign _T_944 = 3'h2 == io_operation_14; // @[Mux.scala 46:19:@182.4]
  assign _T_945 = _T_944 ? _T_939 : {{256'd0}, _T_943}; // @[Mux.scala 46:16:@183.4]
  assign _T_946 = 3'h1 == io_operation_14; // @[Mux.scala 46:19:@184.4]
  assign _T_947 = _T_946 ? {{256'd0}, _T_937} : _T_945; // @[Mux.scala 46:16:@185.4]
  assign _T_948 = 3'h0 == io_operation_14; // @[Mux.scala 46:19:@186.4]
  assign _GEN_121 = 2'h1 == io_selects_15_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_122 = 2'h2 == io_selects_15_0 ? io_inputs_2 : _GEN_121; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_123 = 2'h3 == io_selects_15_0 ? io_inputs_3 : _GEN_122; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_125 = 2'h1 == io_selects_15_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_126 = 2'h2 == io_selects_15_1 ? io_inputs_2 : _GEN_125; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _GEN_127 = 2'h3 == io_selects_15_1 ? io_inputs_3 : _GEN_126; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _T_953 = _GEN_123 + _GEN_127; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@188.4]
  assign _T_954 = _GEN_123 + _GEN_127; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 32:53:@189.4]
  assign _T_956 = _GEN_123 * _GEN_127; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 33:58:@190.4]
  assign _T_958 = _GEN_123 / _GEN_127; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 34:56:@191.4]
  assign _T_959 = 3'h3 == io_operation_15; // @[Mux.scala 46:19:@192.4]
  assign _T_960 = _T_959 ? _T_958 : 256'h0; // @[Mux.scala 46:16:@193.4]
  assign _T_961 = 3'h2 == io_operation_15; // @[Mux.scala 46:19:@194.4]
  assign _T_962 = _T_961 ? _T_956 : {{256'd0}, _T_960}; // @[Mux.scala 46:16:@195.4]
  assign _T_963 = 3'h1 == io_operation_15; // @[Mux.scala 46:19:@196.4]
  assign _T_964 = _T_963 ? {{256'd0}, _T_954} : _T_962; // @[Mux.scala 46:16:@197.4]
  assign _T_965 = 3'h0 == io_operation_15; // @[Mux.scala 46:19:@198.4]
  assign io_outputs_0 = _T_977[255:0]; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 23:14:@520.4]
  assign io_outputs_1 = _T_988[255:0]; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 23:14:@521.4]
  assign io_outputs_2 = _T_999[255:0]; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 23:14:@522.4]
  assign io_outputs_3 = _T_1010[255:0]; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 23:14:@523.4]
  assign io_outputs_4 = _T_1021[255:0]; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 23:14:@524.4]
  assign io_outputs_5 = _T_1032[255:0]; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 23:14:@525.4]
  assign io_outputs_6 = _T_1043[255:0]; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 23:14:@526.4]
  assign io_outputs_7 = _T_1054[255:0]; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 23:14:@527.4]
  assign io_outputs_8 = _T_1065[255:0]; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 23:14:@528.4]
  assign io_outputs_9 = _T_1076[255:0]; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 23:14:@529.4]
  assign io_outputs_10 = _T_1087[255:0]; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 23:14:@530.4]
  assign io_outputs_11 = _T_1098[255:0]; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 23:14:@531.4]
  assign io_outputs_12 = _T_1109[255:0]; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 23:14:@532.4]
  assign io_outputs_13 = _T_1120[255:0]; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 23:14:@533.4]
  assign io_outputs_14 = _T_1131[255:0]; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 23:14:@534.4]
  assign io_outputs_15 = _T_1142[255:0]; // @[MuxTest_width_256_inputs_4_outputs_16_pipeline_5s.scala 23:14:@535.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {16{`RANDOM}};
  _T_969 = _RAND_0[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {16{`RANDOM}};
  _T_971 = _RAND_1[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {16{`RANDOM}};
  _T_973 = _RAND_2[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {16{`RANDOM}};
  _T_975 = _RAND_3[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {16{`RANDOM}};
  _T_977 = _RAND_4[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {16{`RANDOM}};
  _T_980 = _RAND_5[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {16{`RANDOM}};
  _T_982 = _RAND_6[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {16{`RANDOM}};
  _T_984 = _RAND_7[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {16{`RANDOM}};
  _T_986 = _RAND_8[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {16{`RANDOM}};
  _T_988 = _RAND_9[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {16{`RANDOM}};
  _T_991 = _RAND_10[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {16{`RANDOM}};
  _T_993 = _RAND_11[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {16{`RANDOM}};
  _T_995 = _RAND_12[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {16{`RANDOM}};
  _T_997 = _RAND_13[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {16{`RANDOM}};
  _T_999 = _RAND_14[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {16{`RANDOM}};
  _T_1002 = _RAND_15[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {16{`RANDOM}};
  _T_1004 = _RAND_16[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {16{`RANDOM}};
  _T_1006 = _RAND_17[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {16{`RANDOM}};
  _T_1008 = _RAND_18[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {16{`RANDOM}};
  _T_1010 = _RAND_19[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {16{`RANDOM}};
  _T_1013 = _RAND_20[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {16{`RANDOM}};
  _T_1015 = _RAND_21[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {16{`RANDOM}};
  _T_1017 = _RAND_22[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {16{`RANDOM}};
  _T_1019 = _RAND_23[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {16{`RANDOM}};
  _T_1021 = _RAND_24[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {16{`RANDOM}};
  _T_1024 = _RAND_25[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {16{`RANDOM}};
  _T_1026 = _RAND_26[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {16{`RANDOM}};
  _T_1028 = _RAND_27[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {16{`RANDOM}};
  _T_1030 = _RAND_28[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {16{`RANDOM}};
  _T_1032 = _RAND_29[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {16{`RANDOM}};
  _T_1035 = _RAND_30[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {16{`RANDOM}};
  _T_1037 = _RAND_31[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {16{`RANDOM}};
  _T_1039 = _RAND_32[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {16{`RANDOM}};
  _T_1041 = _RAND_33[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {16{`RANDOM}};
  _T_1043 = _RAND_34[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {16{`RANDOM}};
  _T_1046 = _RAND_35[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {16{`RANDOM}};
  _T_1048 = _RAND_36[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {16{`RANDOM}};
  _T_1050 = _RAND_37[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {16{`RANDOM}};
  _T_1052 = _RAND_38[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {16{`RANDOM}};
  _T_1054 = _RAND_39[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {16{`RANDOM}};
  _T_1057 = _RAND_40[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {16{`RANDOM}};
  _T_1059 = _RAND_41[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {16{`RANDOM}};
  _T_1061 = _RAND_42[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {16{`RANDOM}};
  _T_1063 = _RAND_43[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {16{`RANDOM}};
  _T_1065 = _RAND_44[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {16{`RANDOM}};
  _T_1068 = _RAND_45[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {16{`RANDOM}};
  _T_1070 = _RAND_46[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {16{`RANDOM}};
  _T_1072 = _RAND_47[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {16{`RANDOM}};
  _T_1074 = _RAND_48[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {16{`RANDOM}};
  _T_1076 = _RAND_49[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {16{`RANDOM}};
  _T_1079 = _RAND_50[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {16{`RANDOM}};
  _T_1081 = _RAND_51[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {16{`RANDOM}};
  _T_1083 = _RAND_52[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {16{`RANDOM}};
  _T_1085 = _RAND_53[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {16{`RANDOM}};
  _T_1087 = _RAND_54[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {16{`RANDOM}};
  _T_1090 = _RAND_55[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {16{`RANDOM}};
  _T_1092 = _RAND_56[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {16{`RANDOM}};
  _T_1094 = _RAND_57[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {16{`RANDOM}};
  _T_1096 = _RAND_58[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {16{`RANDOM}};
  _T_1098 = _RAND_59[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {16{`RANDOM}};
  _T_1101 = _RAND_60[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {16{`RANDOM}};
  _T_1103 = _RAND_61[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {16{`RANDOM}};
  _T_1105 = _RAND_62[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {16{`RANDOM}};
  _T_1107 = _RAND_63[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {16{`RANDOM}};
  _T_1109 = _RAND_64[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {16{`RANDOM}};
  _T_1112 = _RAND_65[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {16{`RANDOM}};
  _T_1114 = _RAND_66[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {16{`RANDOM}};
  _T_1116 = _RAND_67[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {16{`RANDOM}};
  _T_1118 = _RAND_68[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {16{`RANDOM}};
  _T_1120 = _RAND_69[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {16{`RANDOM}};
  _T_1123 = _RAND_70[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {16{`RANDOM}};
  _T_1125 = _RAND_71[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {16{`RANDOM}};
  _T_1127 = _RAND_72[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {16{`RANDOM}};
  _T_1129 = _RAND_73[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {16{`RANDOM}};
  _T_1131 = _RAND_74[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {16{`RANDOM}};
  _T_1134 = _RAND_75[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {16{`RANDOM}};
  _T_1136 = _RAND_76[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {16{`RANDOM}};
  _T_1138 = _RAND_77[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {16{`RANDOM}};
  _T_1140 = _RAND_78[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {16{`RANDOM}};
  _T_1142 = _RAND_79[511:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_710) begin
      _T_969 <= {{256'd0}, _GEN_3};
    end else begin
      _T_969 <= _T_709;
    end
    _T_971 <= _T_969;
    _T_973 <= _T_971;
    _T_975 <= _T_973;
    _T_977 <= _T_975;
    if (_T_727) begin
      _T_980 <= {{256'd0}, _GEN_11};
    end else begin
      _T_980 <= _T_726;
    end
    _T_982 <= _T_980;
    _T_984 <= _T_982;
    _T_986 <= _T_984;
    _T_988 <= _T_986;
    if (_T_744) begin
      _T_991 <= {{256'd0}, _GEN_19};
    end else begin
      _T_991 <= _T_743;
    end
    _T_993 <= _T_991;
    _T_995 <= _T_993;
    _T_997 <= _T_995;
    _T_999 <= _T_997;
    if (_T_761) begin
      _T_1002 <= {{256'd0}, _GEN_27};
    end else begin
      _T_1002 <= _T_760;
    end
    _T_1004 <= _T_1002;
    _T_1006 <= _T_1004;
    _T_1008 <= _T_1006;
    _T_1010 <= _T_1008;
    if (_T_778) begin
      _T_1013 <= {{256'd0}, _GEN_35};
    end else begin
      _T_1013 <= _T_777;
    end
    _T_1015 <= _T_1013;
    _T_1017 <= _T_1015;
    _T_1019 <= _T_1017;
    _T_1021 <= _T_1019;
    if (_T_795) begin
      _T_1024 <= {{256'd0}, _GEN_43};
    end else begin
      _T_1024 <= _T_794;
    end
    _T_1026 <= _T_1024;
    _T_1028 <= _T_1026;
    _T_1030 <= _T_1028;
    _T_1032 <= _T_1030;
    if (_T_812) begin
      _T_1035 <= {{256'd0}, _GEN_51};
    end else begin
      _T_1035 <= _T_811;
    end
    _T_1037 <= _T_1035;
    _T_1039 <= _T_1037;
    _T_1041 <= _T_1039;
    _T_1043 <= _T_1041;
    if (_T_829) begin
      _T_1046 <= {{256'd0}, _GEN_59};
    end else begin
      _T_1046 <= _T_828;
    end
    _T_1048 <= _T_1046;
    _T_1050 <= _T_1048;
    _T_1052 <= _T_1050;
    _T_1054 <= _T_1052;
    if (_T_846) begin
      _T_1057 <= {{256'd0}, _GEN_67};
    end else begin
      _T_1057 <= _T_845;
    end
    _T_1059 <= _T_1057;
    _T_1061 <= _T_1059;
    _T_1063 <= _T_1061;
    _T_1065 <= _T_1063;
    if (_T_863) begin
      _T_1068 <= {{256'd0}, _GEN_75};
    end else begin
      _T_1068 <= _T_862;
    end
    _T_1070 <= _T_1068;
    _T_1072 <= _T_1070;
    _T_1074 <= _T_1072;
    _T_1076 <= _T_1074;
    if (_T_880) begin
      _T_1079 <= {{256'd0}, _GEN_83};
    end else begin
      _T_1079 <= _T_879;
    end
    _T_1081 <= _T_1079;
    _T_1083 <= _T_1081;
    _T_1085 <= _T_1083;
    _T_1087 <= _T_1085;
    if (_T_897) begin
      _T_1090 <= {{256'd0}, _GEN_91};
    end else begin
      _T_1090 <= _T_896;
    end
    _T_1092 <= _T_1090;
    _T_1094 <= _T_1092;
    _T_1096 <= _T_1094;
    _T_1098 <= _T_1096;
    if (_T_914) begin
      _T_1101 <= {{256'd0}, _GEN_99};
    end else begin
      _T_1101 <= _T_913;
    end
    _T_1103 <= _T_1101;
    _T_1105 <= _T_1103;
    _T_1107 <= _T_1105;
    _T_1109 <= _T_1107;
    if (_T_931) begin
      _T_1112 <= {{256'd0}, _GEN_107};
    end else begin
      _T_1112 <= _T_930;
    end
    _T_1114 <= _T_1112;
    _T_1116 <= _T_1114;
    _T_1118 <= _T_1116;
    _T_1120 <= _T_1118;
    if (_T_948) begin
      _T_1123 <= {{256'd0}, _GEN_115};
    end else begin
      _T_1123 <= _T_947;
    end
    _T_1125 <= _T_1123;
    _T_1127 <= _T_1125;
    _T_1129 <= _T_1127;
    _T_1131 <= _T_1129;
    if (_T_965) begin
      _T_1134 <= {{256'd0}, _GEN_123};
    end else begin
      _T_1134 <= _T_964;
    end
    _T_1136 <= _T_1134;
    _T_1138 <= _T_1136;
    _T_1140 <= _T_1138;
    _T_1142 <= _T_1140;
  end
endmodule
