../../../../platforms/asap7/lef/fakeram7_2048x39.lef